module lenet5_layer_2(clk,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81);
   input clk;
   input signed [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117;
   output reg signed [9:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81;
   wire signed [5:0] neg1,neg2,neg3,neg4,neg5,neg6,neg7,neg8,neg9,neg10,neg11,neg12,neg13,neg14,neg15,neg16,neg17,neg18,neg19,neg20,neg21,neg22,neg23,neg24,neg25,neg26,neg27,neg28,neg29,neg30,neg31,neg32,neg33,neg34,neg35,neg36,neg37,neg38,neg39,neg40,neg41,neg42,neg43,neg44,neg45,neg46,neg47,neg48,neg49,neg50,neg51,neg52,neg53,neg54,neg55,neg56,neg57,neg58,neg59,neg60,neg61,neg62,neg63,neg64,neg65,neg66,neg67,neg68,neg69,neg70,neg71,neg72,neg73,neg74,neg75,neg76,neg77,neg78,neg79,neg80,neg81,neg82,neg83,neg84,neg85,neg86,neg87,neg88,neg89,neg90,neg91,neg92,neg93,neg94,neg95,neg96,neg97,neg98,neg99,neg100,neg101,neg102,neg103,neg104,neg105,neg106,neg107,neg108,neg109,neg110,neg111,neg112,neg113,neg114,neg115,neg116,neg117;

   //Bias value
   wire signed [9:0] b1 = $signed(10'h6);
   wire signed [9:0] b2 = $signed(10'h5);
   wire signed [9:0] b3 = $signed(10'h5);
   wire signed [9:0] b4 = $signed(10'h4);
   wire signed [9:0] b5 = $signed(10'h5);
   wire signed [9:0] b6 = $signed(10'h3);
   wire signed [9:0] b7 = $signed(10'h4);
   wire signed [9:0] b8 = $signed(10'h8);
   wire signed [9:0] b9 = $signed(10'h6);
   wire signed [9:0] b10 = $signed(10'h4);
   wire signed [9:0] b11 = $signed(10'h3);
   wire signed [9:0] b12 = $signed(10'h8);
   wire signed [9:0] b13 = $signed(10'h3);
   wire signed [9:0] b14 = $signed(10'h5);
   wire signed [9:0] b15 = $signed(10'h9);
   wire signed [9:0] b16 = $signed(10'h3FE);
   wire signed [9:0] b17 = $signed(10'h7);
   wire signed [9:0] b18 = $signed(10'h4);
   wire signed [9:0] b19 = $signed(10'h5);
   wire signed [9:0] b20 = $signed(10'h4);
   wire signed [9:0] b21 = $signed(10'h6);
   wire signed [9:0] b22 = $signed(10'h9);
   wire signed [9:0] b23 = $signed(10'h3);
   wire signed [9:0] b24 = $signed(10'h5);
   wire signed [9:0] b25 = $signed(10'h8);
   wire signed [9:0] b26 = $signed(10'h3FF);
   wire signed [9:0] b27 = $signed(10'h0);
   wire signed [9:0] b28 = $signed(10'h2);
   wire signed [9:0] b29 = $signed(10'h5);
   wire signed [9:0] b30 = $signed(10'h5);
   wire signed [9:0] b31 = $signed(10'h7);
   wire signed [9:0] b32 = $signed(10'h6);
   wire signed [9:0] b33 = $signed(10'h1);
   wire signed [9:0] b34 = $signed(10'h7);
   wire signed [9:0] b35 = $signed(10'h1);
   wire signed [9:0] b36 = $signed(10'h3);
   wire signed [9:0] b37 = $signed(10'h5);
   wire signed [9:0] b38 = $signed(10'h4);
   wire signed [9:0] b39 = $signed(10'h8);
   wire signed [9:0] b40 = $signed(10'h5);
   wire signed [9:0] b41 = $signed(10'h3);
   wire signed [9:0] b42 = $signed(10'h7);
   wire signed [9:0] b43 = $signed(10'h6);
   wire signed [9:0] b44 = $signed(10'h2);
   wire signed [9:0] b45 = $signed(10'h4);
   wire signed [9:0] b46 = $signed(10'h0);
   wire signed [9:0] b47 = $signed(10'h7);
   wire signed [9:0] b48 = $signed(10'h6);
   wire signed [9:0] b49 = $signed(10'hB);
   wire signed [9:0] b50 = $signed(10'h4);
   wire signed [9:0] b51 = $signed(10'h7);
   wire signed [9:0] b52 = $signed(10'h7);
   wire signed [9:0] b53 = $signed(10'h5);
   wire signed [9:0] b54 = $signed(10'h6);
   wire signed [9:0] b55 = $signed(10'hA);
   wire signed [9:0] b56 = $signed(10'h3);
   wire signed [9:0] b57 = $signed(10'h8);
   wire signed [9:0] b58 = $signed(10'h8);
   wire signed [9:0] b59 = $signed(10'h7);
   wire signed [9:0] b60 = $signed(10'h7);
   wire signed [9:0] b61 = $signed(10'h5);
   wire signed [9:0] b62 = $signed(10'h3);
   wire signed [9:0] b63 = $signed(10'h3);
   wire signed [9:0] b64 = $signed(10'h9);
   wire signed [9:0] b65 = $signed(10'h8);
   wire signed [9:0] b66 = $signed(10'h5);
   wire signed [9:0] b67 = $signed(10'h5);
   wire signed [9:0] b68 = $signed(10'h5);
   wire signed [9:0] b69 = $signed(10'h3);
   wire signed [9:0] b70 = $signed(10'h5);
   wire signed [9:0] b71 = $signed(10'h1);
   wire signed [9:0] b72 = $signed(10'h9);
   wire signed [9:0] b73 = $signed(10'h3);
   wire signed [9:0] b74 = $signed(10'h6);
   wire signed [9:0] b75 = $signed(10'h1);
   wire signed [9:0] b76 = $signed(10'h4);
   wire signed [9:0] b77 = $signed(10'h5);
   wire signed [9:0] b78 = $signed(10'h5);
   wire signed [9:0] b79 = $signed(10'h5);
   wire signed [9:0] b80 = $signed(10'h4);
   wire signed [9:0] b81 = $signed(10'h2);

   //Negation modules
   negate #(6) N1(in1,neg1);
   negate #(6) N2(in2,neg2);
   negate #(6) N3(in3,neg3);
   negate #(6) N4(in4,neg4);
   negate #(6) N5(in5,neg5);
   negate #(6) N6(in6,neg6);
   negate #(6) N7(in7,neg7);
   negate #(6) N8(in8,neg8);
   negate #(6) N9(in9,neg9);
   negate #(6) N10(in10,neg10);
   negate #(6) N11(in11,neg11);
   negate #(6) N12(in12,neg12);
   negate #(6) N13(in13,neg13);
   negate #(6) N14(in14,neg14);
   negate #(6) N15(in15,neg15);
   negate #(6) N16(in16,neg16);
   negate #(6) N17(in17,neg17);
   negate #(6) N18(in18,neg18);
   negate #(6) N19(in19,neg19);
   negate #(6) N20(in20,neg20);
   negate #(6) N21(in21,neg21);
   negate #(6) N22(in22,neg22);
   negate #(6) N23(in23,neg23);
   negate #(6) N24(in24,neg24);
   negate #(6) N25(in25,neg25);
   negate #(6) N26(in26,neg26);
   negate #(6) N27(in27,neg27);
   negate #(6) N28(in28,neg28);
   negate #(6) N29(in29,neg29);
   negate #(6) N30(in30,neg30);
   negate #(6) N31(in31,neg31);
   negate #(6) N32(in32,neg32);
   negate #(6) N33(in33,neg33);
   negate #(6) N34(in34,neg34);
   negate #(6) N35(in35,neg35);
   negate #(6) N36(in36,neg36);
   negate #(6) N37(in37,neg37);
   negate #(6) N38(in38,neg38);
   negate #(6) N39(in39,neg39);
   negate #(6) N40(in40,neg40);
   negate #(6) N41(in41,neg41);
   negate #(6) N42(in42,neg42);
   negate #(6) N43(in43,neg43);
   negate #(6) N44(in44,neg44);
   negate #(6) N45(in45,neg45);
   negate #(6) N46(in46,neg46);
   negate #(6) N47(in47,neg47);
   negate #(6) N48(in48,neg48);
   negate #(6) N49(in49,neg49);
   negate #(6) N50(in50,neg50);
   negate #(6) N51(in51,neg51);
   negate #(6) N52(in52,neg52);
   negate #(6) N53(in53,neg53);
   negate #(6) N54(in54,neg54);
   negate #(6) N55(in55,neg55);
   negate #(6) N56(in56,neg56);
   negate #(6) N57(in57,neg57);
   negate #(6) N58(in58,neg58);
   negate #(6) N59(in59,neg59);
   negate #(6) N60(in60,neg60);
   negate #(6) N61(in61,neg61);
   negate #(6) N62(in62,neg62);
   negate #(6) N63(in63,neg63);
   negate #(6) N64(in64,neg64);
   negate #(6) N65(in65,neg65);
   negate #(6) N66(in66,neg66);
   negate #(6) N67(in67,neg67);
   negate #(6) N68(in68,neg68);
   negate #(6) N69(in69,neg69);
   negate #(6) N70(in70,neg70);
   negate #(6) N71(in71,neg71);
   negate #(6) N72(in72,neg72);
   negate #(6) N73(in73,neg73);
   negate #(6) N74(in74,neg74);
   negate #(6) N75(in75,neg75);
   negate #(6) N76(in76,neg76);
   negate #(6) N77(in77,neg77);
   negate #(6) N78(in78,neg78);
   negate #(6) N79(in79,neg79);
   negate #(6) N80(in80,neg80);
   negate #(6) N81(in81,neg81);
   negate #(6) N82(in82,neg82);
   negate #(6) N83(in83,neg83);
   negate #(6) N84(in84,neg84);
   negate #(6) N85(in85,neg85);
   negate #(6) N86(in86,neg86);
   negate #(6) N87(in87,neg87);
   negate #(6) N88(in88,neg88);
   negate #(6) N89(in89,neg89);
   negate #(6) N90(in90,neg90);
   negate #(6) N91(in91,neg91);
   negate #(6) N92(in92,neg92);
   negate #(6) N93(in93,neg93);
   negate #(6) N94(in94,neg94);
   negate #(6) N95(in95,neg95);
   negate #(6) N96(in96,neg96);
   negate #(6) N97(in97,neg97);
   negate #(6) N98(in98,neg98);
   negate #(6) N99(in99,neg99);
   negate #(6) N100(in100,neg100);
   negate #(6) N101(in101,neg101);
   negate #(6) N102(in102,neg102);
   negate #(6) N103(in103,neg103);
   negate #(6) N104(in104,neg104);
   negate #(6) N105(in105,neg105);
   negate #(6) N106(in106,neg106);
   negate #(6) N107(in107,neg107);
   negate #(6) N108(in108,neg108);
   negate #(6) N109(in109,neg109);
   negate #(6) N110(in110,neg110);
   negate #(6) N111(in111,neg111);
   negate #(6) N112(in112,neg112);
   negate #(6) N113(in113,neg113);
   negate #(6) N114(in114,neg114);
   negate #(6) N115(in115,neg115);
   negate #(6) N116(in116,neg116);
   negate #(6) N117(in117,neg117);

   // m1_1 = W*in
   wire signed [9:0] m1_1;
   assign m1_1 =10'b0;

   // m1_2 = W*in
   wire signed [9:0] m1_2;
   assign m1_2 =10'b0;

   // m1_3 = W*in
   wire signed [9:0] m1_3;
   assign m1_3 =10'b0;

   // m1_4 = W*in
   wire signed [9:0] m1_4;
   assign m1_4 =10'b0;

   // m1_5 = W*in
   wire signed [9:0] m1_5;
   assign m1_5 =10'b0;

   // m1_6 = W*in
   wire signed [9:0] m1_6;
   assign m1_6 =10'b0;

   // m1_7 = W*in
   wire signed [9:0] m1_7;
   assign m1_7 =10'b0;

   // m1_8 = W*in
   wire signed [9:0] m1_8;
   assign m1_8 =10'b0;

   // m1_9 = W*in
   wire signed [9:0] m1_9;
   assign m1_9 =10'b0;

   // m1_10 = W*in
   wire signed [9:0] m1_10;
   assign m1_10 =10'b0;

   // m1_11 = W*in
   wire signed [9:0] m1_11;
   assign m1_11 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_12 = W*in
   wire signed [9:0] m1_12;
   assign m1_12 =10'b0;

   // m1_13 = W*in
   wire signed [9:0] m1_13;
   assign m1_13 =10'b0;

   // m1_14 = W*in
   wire signed [9:0] m1_14;
   assign m1_14 =10'b0;

   // m1_15 = W*in
   wire signed [9:0] m1_15;
   assign m1_15 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_16 = W*in
   wire signed [9:0] m1_16;
   assign m1_16 =10'b0;

   // m1_17 = W*in
   wire signed [9:0] m1_17;
   assign m1_17 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_18 = W*in
   wire signed [9:0] m1_18;
   assign m1_18 =10'b0;

   // m1_19 = W*in
   wire signed [9:0] m1_19;
   assign m1_19 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_20 = W*in
   wire signed [9:0] m1_20;
   assign m1_20 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_21 = W*in
   wire signed [9:0] m1_21;
   assign m1_21 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_22 = W*in
   wire signed [9:0] m1_22;
   assign m1_22 =10'b0;

   // m1_23 = W*in
   wire signed [9:0] m1_23;
   assign m1_23 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_24 = W*in
   wire signed [9:0] m1_24;
   assign m1_24 =10'b0;

   // m1_25 = W*in
   wire signed [9:0] m1_25;
   assign m1_25 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_26 = W*in
   wire signed [9:0] m1_26;
   assign m1_26 =10'b0;

   // m1_27 = W*in
   wire signed [9:0] m1_27;
   assign m1_27 =10'b0;

   // m1_28 = W*in
   wire signed [9:0] m1_28;
   assign m1_28 =10'b0;

   // m1_29 = W*in
   wire signed [9:0] m1_29;
   assign m1_29 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_30 = W*in
   wire signed [9:0] m1_30;
   assign m1_30 =10'b0;

   // m1_31 = W*in
   wire signed [9:0] m1_31;
   assign m1_31 =10'b0;

   // m1_32 = W*in
   wire signed [9:0] m1_32;
   assign m1_32 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_33 = W*in
   wire signed [9:0] m1_33;
   assign m1_33 =10'b0;

   // m1_34 = W*in
   wire signed [9:0] m1_34;
   assign m1_34 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_35 = W*in
   wire signed [9:0] m1_35;
   assign m1_35 =10'b0;

   // m1_36 = W*in
   wire signed [9:0] m1_36;
   assign m1_36 =10'b0;

   // m1_37 = W*in
   wire signed [9:0] m1_37;
   assign m1_37 =10'b0;

   // m1_38 = W*in
   wire signed [9:0] m1_38;
   assign m1_38 =10'b0;

   // m1_39 = W*in
   wire signed [9:0] m1_39;
   assign m1_39 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_40 = W*in
   wire signed [9:0] m1_40;
   assign m1_40 =10'b0;

   // m1_41 = W*in
   wire signed [9:0] m1_41;
   assign m1_41 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_42 = W*in
   wire signed [9:0] m1_42;
   assign m1_42 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_43 = W*in
   wire signed [9:0] m1_43;
   assign m1_43 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_44 = W*in
   wire signed [9:0] m1_44;
   assign m1_44 =10'b0;

   // m1_45 = W*in
   wire signed [9:0] m1_45;
   assign m1_45 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_46 = W*in
   wire signed [9:0] m1_46;
   assign m1_46 =10'b0;

   // m1_47 = W*in
   wire signed [9:0] m1_47;
   assign m1_47 =10'b0;

   // m1_48 = W*in
   wire signed [9:0] m1_48;
   assign m1_48 =10'b0;

   // m1_49 = W*in
   wire signed [9:0] m1_49;
   assign m1_49 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_50 = W*in
   wire signed [9:0] m1_50;
   assign m1_50 =10'b0;

   // m1_51 = W*in
   wire signed [9:0] m1_51;
   assign m1_51 =10'b0;

   // m1_52 = W*in
   wire signed [9:0] m1_52;
   assign m1_52 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_53 = W*in
   wire signed [9:0] m1_53;
   assign m1_53 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_54 = W*in
   wire signed [9:0] m1_54;
   assign m1_54 =10'b0;

   // m1_55 = W*in
   wire signed [9:0] m1_55;
   assign m1_55 ={ {3{in1[5]}} , in1 , {1{1'b0}} };

   // m1_56 = W*in
   wire signed [9:0] m1_56;
   assign m1_56 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_57 = W*in
   wire signed [9:0] m1_57;
   assign m1_57 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_58 = W*in
   wire signed [9:0] m1_58;
   assign m1_58 =10'b0;

   // m1_59 = W*in
   wire signed [9:0] m1_59;
   assign m1_59 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_60 = W*in
   wire signed [9:0] m1_60;
   assign m1_60 =10'b0;

   // m1_61 = W*in
   wire signed [9:0] m1_61;
   assign m1_61 =10'b0;

   // m1_62 = W*in
   wire signed [9:0] m1_62;
   assign m1_62 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_63 = W*in
   wire signed [9:0] m1_63;
   assign m1_63 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_64 = W*in
   wire signed [9:0] m1_64;
   assign m1_64 =10'b0;

   // m1_65 = W*in
   wire signed [9:0] m1_65;
   assign m1_65 =10'b0;

   // m1_66 = W*in
   wire signed [9:0] m1_66;
   assign m1_66 ={ {2{in1[5]}} , in1 , {2{1'b0}} };

   // m1_67 = W*in
   wire signed [9:0] m1_67;
   assign m1_67 =10'b0;

   // m1_68 = W*in
   wire signed [9:0] m1_68;
   assign m1_68 =10'b0;

   // m1_69 = W*in
   wire signed [9:0] m1_69;
   assign m1_69 =10'b0;

   // m1_70 = W*in
   wire signed [9:0] m1_70;
   assign m1_70 =10'b0;

   // m1_71 = W*in
   wire signed [9:0] m1_71;
   assign m1_71 =10'b0;

   // m1_72 = W*in
   wire signed [9:0] m1_72;
   assign m1_72 =10'b0;

   // m1_73 = W*in
   wire signed [9:0] m1_73;
   assign m1_73 =10'b0;

   // m1_74 = W*in
   wire signed [9:0] m1_74;
   assign m1_74 =10'b0;

   // m1_75 = W*in
   wire signed [9:0] m1_75;
   assign m1_75 =10'b0;

   // m1_76 = W*in
   wire signed [9:0] m1_76;
   assign m1_76 =10'b0;

   // m1_77 = W*in
   wire signed [9:0] m1_77;
   assign m1_77 =10'b0;

   // m1_78 = W*in
   wire signed [9:0] m1_78;
   assign m1_78 =10'b0;

   // m1_79 = W*in
   wire signed [9:0] m1_79;
   assign m1_79 ={ {3{neg1[5]}} , neg1 , {1{1'b0}} };

   // m1_80 = W*in
   wire signed [9:0] m1_80;
   assign m1_80 =10'b0;

   // m1_81 = W*in
   wire signed [9:0] m1_81;
   assign m1_81 =10'b0;

   // m2_1 = W*in
   wire signed [9:0] m2_1;
   assign m2_1 =10'b0;

   // m2_2 = W*in
   wire signed [9:0] m2_2;
   assign m2_2 =10'b0;

   // m2_3 = W*in
   wire signed [9:0] m2_3;
   assign m2_3 =10'b0;

   // m2_4 = W*in
   wire signed [9:0] m2_4;
   assign m2_4 =10'b0;

   // m2_5 = W*in
   wire signed [9:0] m2_5;
   assign m2_5 =10'b0;

   // m2_6 = W*in
   wire signed [9:0] m2_6;
   assign m2_6 =10'b0;

   // m2_7 = W*in
   wire signed [9:0] m2_7;
   assign m2_7 =10'b0;

   // m2_8 = W*in
   wire signed [9:0] m2_8;
   assign m2_8 =10'b0;

   // m2_9 = W*in
   wire signed [9:0] m2_9;
   assign m2_9 =10'b0;

   // m2_10 = W*in
   wire signed [9:0] m2_10;
   assign m2_10 =10'b0;

   // m2_11 = W*in
   wire signed [9:0] m2_11;
   assign m2_11 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_12 = W*in
   wire signed [9:0] m2_12;
   assign m2_12 =10'b0;

   // m2_13 = W*in
   wire signed [9:0] m2_13;
   assign m2_13 =10'b0;

   // m2_14 = W*in
   wire signed [9:0] m2_14;
   assign m2_14 =10'b0;

   // m2_15 = W*in
   wire signed [9:0] m2_15;
   assign m2_15 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_16 = W*in
   wire signed [9:0] m2_16;
   assign m2_16 =10'b0;

   // m2_17 = W*in
   wire signed [9:0] m2_17;
   assign m2_17 =10'b0;

   // m2_18 = W*in
   wire signed [9:0] m2_18;
   assign m2_18 =10'b0;

   // m2_19 = W*in
   wire signed [9:0] m2_19;
   assign m2_19 =10'b0;

   // m2_20 = W*in
   wire signed [9:0] m2_20;
   assign m2_20 =10'b0;

   // m2_21 = W*in
   wire signed [9:0] m2_21;
   assign m2_21 =10'b0;

   // m2_22 = W*in
   wire signed [9:0] m2_22;
   assign m2_22 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_23 = W*in
   wire signed [9:0] m2_23;
   assign m2_23 =10'b0;

   // m2_24 = W*in
   wire signed [9:0] m2_24;
   assign m2_24 =10'b0;

   // m2_25 = W*in
   wire signed [9:0] m2_25;
   assign m2_25 =10'b0;

   // m2_26 = W*in
   wire signed [9:0] m2_26;
   assign m2_26 =10'b0;

   // m2_27 = W*in
   wire signed [9:0] m2_27;
   assign m2_27 =10'b0;

   // m2_28 = W*in
   wire signed [9:0] m2_28;
   assign m2_28 =10'b0;

   // m2_29 = W*in
   wire signed [9:0] m2_29;
   assign m2_29 =10'b0;

   // m2_30 = W*in
   wire signed [9:0] m2_30;
   assign m2_30 =10'b0;

   // m2_31 = W*in
   wire signed [9:0] m2_31;
   assign m2_31 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_32 = W*in
   wire signed [9:0] m2_32;
   assign m2_32 =10'b0;

   // m2_33 = W*in
   wire signed [9:0] m2_33;
   assign m2_33 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_34 = W*in
   wire signed [9:0] m2_34;
   assign m2_34 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_35 = W*in
   wire signed [9:0] m2_35;
   assign m2_35 =10'b0;

   // m2_36 = W*in
   wire signed [9:0] m2_36;
   assign m2_36 =10'b0;

   // m2_37 = W*in
   wire signed [9:0] m2_37;
   assign m2_37 =10'b0;

   // m2_38 = W*in
   wire signed [9:0] m2_38;
   assign m2_38 =10'b0;

   // m2_39 = W*in
   wire signed [9:0] m2_39;
   assign m2_39 =10'b0;

   // m2_40 = W*in
   wire signed [9:0] m2_40;
   assign m2_40 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_41 = W*in
   wire signed [9:0] m2_41;
   assign m2_41 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_42 = W*in
   wire signed [9:0] m2_42;
   assign m2_42 =10'b0;

   // m2_43 = W*in
   wire signed [9:0] m2_43;
   assign m2_43 =10'b0;

   // m2_44 = W*in
   wire signed [9:0] m2_44;
   assign m2_44 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_45 = W*in
   wire signed [9:0] m2_45;
   assign m2_45 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_46 = W*in
   wire signed [9:0] m2_46;
   assign m2_46 =10'b0;

   // m2_47 = W*in
   wire signed [9:0] m2_47;
   assign m2_47 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_48 = W*in
   wire signed [9:0] m2_48;
   assign m2_48 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_49 = W*in
   wire signed [9:0] m2_49;
   assign m2_49 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_50 = W*in
   wire signed [9:0] m2_50;
   assign m2_50 =10'b0;

   // m2_51 = W*in
   wire signed [9:0] m2_51;
   assign m2_51 =10'b0;

   // m2_52 = W*in
   wire signed [9:0] m2_52;
   assign m2_52 =10'b0;

   // m2_53 = W*in
   wire signed [9:0] m2_53;
   assign m2_53 =10'b0;

   // m2_54 = W*in
   wire signed [9:0] m2_54;
   assign m2_54 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_55 = W*in
   wire signed [9:0] m2_55;
   assign m2_55 ={ {2{in2[5]}} , in2 , {2{1'b0}} };

   // m2_56 = W*in
   wire signed [9:0] m2_56;
   assign m2_56 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_57 = W*in
   wire signed [9:0] m2_57;
   assign m2_57 =10'b0;

   // m2_58 = W*in
   wire signed [9:0] m2_58;
   assign m2_58 =10'b0;

   // m2_59 = W*in
   wire signed [9:0] m2_59;
   assign m2_59 =10'b0;

   // m2_60 = W*in
   wire signed [9:0] m2_60;
   assign m2_60 =10'b0;

   // m2_61 = W*in
   wire signed [9:0] m2_61;
   assign m2_61 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_62 = W*in
   wire signed [9:0] m2_62;
   assign m2_62 =10'b0;

   // m2_63 = W*in
   wire signed [9:0] m2_63;
   assign m2_63 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_64 = W*in
   wire signed [9:0] m2_64;
   assign m2_64 =10'b0;

   // m2_65 = W*in
   wire signed [9:0] m2_65;
   assign m2_65 =10'b0;

   // m2_66 = W*in
   wire signed [9:0] m2_66;
   assign m2_66 =10'b0;

   // m2_67 = W*in
   wire signed [9:0] m2_67;
   assign m2_67 =10'b0;

   // m2_68 = W*in
   wire signed [9:0] m2_68;
   assign m2_68 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_69 = W*in
   wire signed [9:0] m2_69;
   assign m2_69 =10'b0;

   // m2_70 = W*in
   wire signed [9:0] m2_70;
   assign m2_70 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_71 = W*in
   wire signed [9:0] m2_71;
   assign m2_71 =10'b0;

   // m2_72 = W*in
   wire signed [9:0] m2_72;
   assign m2_72 =10'b0;

   // m2_73 = W*in
   wire signed [9:0] m2_73;
   assign m2_73 =10'b0;

   // m2_74 = W*in
   wire signed [9:0] m2_74;
   assign m2_74 =10'b0;

   // m2_75 = W*in
   wire signed [9:0] m2_75;
   assign m2_75 =10'b0;

   // m2_76 = W*in
   wire signed [9:0] m2_76;
   assign m2_76 =10'b0;

   // m2_77 = W*in
   wire signed [9:0] m2_77;
   assign m2_77 =10'b0;

   // m2_78 = W*in
   wire signed [9:0] m2_78;
   assign m2_78 =10'b0;

   // m2_79 = W*in
   wire signed [9:0] m2_79;
   assign m2_79 =10'b0;

   // m2_80 = W*in
   wire signed [9:0] m2_80;
   assign m2_80 =10'b0;

   // m2_81 = W*in
   wire signed [9:0] m2_81;
   assign m2_81 =10'b0;

   // m3_1 = W*in
   wire signed [9:0] m3_1;
   assign m3_1 =10'b0;

   // m3_2 = W*in
   wire signed [9:0] m3_2;
   assign m3_2 =10'b0;

   // m3_3 = W*in
   wire signed [9:0] m3_3;
   assign m3_3 =10'b0;

   // m3_4 = W*in
   wire signed [9:0] m3_4;
   assign m3_4 =10'b0;

   // m3_5 = W*in
   wire signed [9:0] m3_5;
   assign m3_5 =10'b0;

   // m3_6 = W*in
   wire signed [9:0] m3_6;
   assign m3_6 =10'b0;

   // m3_7 = W*in
   wire signed [9:0] m3_7;
   assign m3_7 =10'b0;

   // m3_8 = W*in
   wire signed [9:0] m3_8;
   assign m3_8 =10'b0;

   // m3_9 = W*in
   wire signed [9:0] m3_9;
   assign m3_9 =10'b0;

   // m3_10 = W*in
   wire signed [9:0] m3_10;
   assign m3_10 =10'b0;

   // m3_11 = W*in
   wire signed [9:0] m3_11;
   assign m3_11 =10'b0;

   // m3_12 = W*in
   wire signed [9:0] m3_12;
   assign m3_12 =10'b0;

   // m3_13 = W*in
   wire signed [9:0] m3_13;
   assign m3_13 =10'b0;

   // m3_14 = W*in
   wire signed [9:0] m3_14;
   assign m3_14 =10'b0;

   // m3_15 = W*in
   wire signed [9:0] m3_15;
   assign m3_15 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_16 = W*in
   wire signed [9:0] m3_16;
   assign m3_16 =10'b0;

   // m3_17 = W*in
   wire signed [9:0] m3_17;
   assign m3_17 =10'b0;

   // m3_18 = W*in
   wire signed [9:0] m3_18;
   assign m3_18 =10'b0;

   // m3_19 = W*in
   wire signed [9:0] m3_19;
   assign m3_19 =10'b0;

   // m3_20 = W*in
   wire signed [9:0] m3_20;
   assign m3_20 =10'b0;

   // m3_21 = W*in
   wire signed [9:0] m3_21;
   assign m3_21 =10'b0;

   // m3_22 = W*in
   wire signed [9:0] m3_22;
   assign m3_22 =10'b0;

   // m3_23 = W*in
   wire signed [9:0] m3_23;
   assign m3_23 =10'b0;

   // m3_24 = W*in
   wire signed [9:0] m3_24;
   assign m3_24 =10'b0;

   // m3_25 = W*in
   wire signed [9:0] m3_25;
   assign m3_25 =10'b0;

   // m3_26 = W*in
   wire signed [9:0] m3_26;
   assign m3_26 =10'b0;

   // m3_27 = W*in
   wire signed [9:0] m3_27;
   assign m3_27 =10'b0;

   // m3_28 = W*in
   wire signed [9:0] m3_28;
   assign m3_28 =10'b0;

   // m3_29 = W*in
   wire signed [9:0] m3_29;
   assign m3_29 =10'b0;

   // m3_30 = W*in
   wire signed [9:0] m3_30;
   assign m3_30 =10'b0;

   // m3_31 = W*in
   wire signed [9:0] m3_31;
   assign m3_31 =10'b0;

   // m3_32 = W*in
   wire signed [9:0] m3_32;
   assign m3_32 =10'b0;

   // m3_33 = W*in
   wire signed [9:0] m3_33;
   assign m3_33 =10'b0;

   // m3_34 = W*in
   wire signed [9:0] m3_34;
   assign m3_34 =10'b0;

   // m3_35 = W*in
   wire signed [9:0] m3_35;
   assign m3_35 =10'b0;

   // m3_36 = W*in
   wire signed [9:0] m3_36;
   assign m3_36 =10'b0;

   // m3_37 = W*in
   wire signed [9:0] m3_37;
   assign m3_37 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_38 = W*in
   wire signed [9:0] m3_38;
   assign m3_38 =10'b0;

   // m3_39 = W*in
   wire signed [9:0] m3_39;
   assign m3_39 =10'b0;

   // m3_40 = W*in
   wire signed [9:0] m3_40;
   assign m3_40 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_41 = W*in
   wire signed [9:0] m3_41;
   assign m3_41 =10'b0;

   // m3_42 = W*in
   wire signed [9:0] m3_42;
   assign m3_42 =10'b0;

   // m3_43 = W*in
   wire signed [9:0] m3_43;
   assign m3_43 =10'b0;

   // m3_44 = W*in
   wire signed [9:0] m3_44;
   assign m3_44 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_45 = W*in
   wire signed [9:0] m3_45;
   assign m3_45 =10'b0;

   // m3_46 = W*in
   wire signed [9:0] m3_46;
   assign m3_46 =10'b0;

   // m3_47 = W*in
   wire signed [9:0] m3_47;
   assign m3_47 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_48 = W*in
   wire signed [9:0] m3_48;
   assign m3_48 =10'b0;

   // m3_49 = W*in
   wire signed [9:0] m3_49;
   assign m3_49 =10'b0;

   // m3_50 = W*in
   wire signed [9:0] m3_50;
   assign m3_50 =10'b0;

   // m3_51 = W*in
   wire signed [9:0] m3_51;
   assign m3_51 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_52 = W*in
   wire signed [9:0] m3_52;
   assign m3_52 =10'b0;

   // m3_53 = W*in
   wire signed [9:0] m3_53;
   assign m3_53 =10'b0;

   // m3_54 = W*in
   wire signed [9:0] m3_54;
   assign m3_54 =10'b0;

   // m3_55 = W*in
   wire signed [9:0] m3_55;
   assign m3_55 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_56 = W*in
   wire signed [9:0] m3_56;
   assign m3_56 =10'b0;

   // m3_57 = W*in
   wire signed [9:0] m3_57;
   assign m3_57 =10'b0;

   // m3_58 = W*in
   wire signed [9:0] m3_58;
   assign m3_58 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_59 = W*in
   wire signed [9:0] m3_59;
   assign m3_59 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_60 = W*in
   wire signed [9:0] m3_60;
   assign m3_60 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_61 = W*in
   wire signed [9:0] m3_61;
   assign m3_61 =10'b0;

   // m3_62 = W*in
   wire signed [9:0] m3_62;
   assign m3_62 =10'b0;

   // m3_63 = W*in
   wire signed [9:0] m3_63;
   assign m3_63 =10'b0;

   // m3_64 = W*in
   wire signed [9:0] m3_64;
   assign m3_64 =10'b0;

   // m3_65 = W*in
   wire signed [9:0] m3_65;
   assign m3_65 =10'b0;

   // m3_66 = W*in
   wire signed [9:0] m3_66;
   assign m3_66 =10'b0;

   // m3_67 = W*in
   wire signed [9:0] m3_67;
   assign m3_67 =10'b0;

   // m3_68 = W*in
   wire signed [9:0] m3_68;
   assign m3_68 =10'b0;

   // m3_69 = W*in
   wire signed [9:0] m3_69;
   assign m3_69 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_70 = W*in
   wire signed [9:0] m3_70;
   assign m3_70 =10'b0;

   // m3_71 = W*in
   wire signed [9:0] m3_71;
   assign m3_71 =10'b0;

   // m3_72 = W*in
   wire signed [9:0] m3_72;
   assign m3_72 =10'b0;

   // m3_73 = W*in
   wire signed [9:0] m3_73;
   assign m3_73 =10'b0;

   // m3_74 = W*in
   wire signed [9:0] m3_74;
   assign m3_74 =10'b0;

   // m3_75 = W*in
   wire signed [9:0] m3_75;
   assign m3_75 =10'b0;

   // m3_76 = W*in
   wire signed [9:0] m3_76;
   assign m3_76 =10'b0;

   // m3_77 = W*in
   wire signed [9:0] m3_77;
   assign m3_77 =10'b0;

   // m3_78 = W*in
   wire signed [9:0] m3_78;
   assign m3_78 =10'b0;

   // m3_79 = W*in
   wire signed [9:0] m3_79;
   assign m3_79 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_80 = W*in
   wire signed [9:0] m3_80;
   assign m3_80 =10'b0;

   // m3_81 = W*in
   wire signed [9:0] m3_81;
   assign m3_81 =10'b0;

   // m4_1 = W*in
   wire signed [9:0] m4_1;
   assign m4_1 =10'b0;

   // m4_2 = W*in
   wire signed [9:0] m4_2;
   assign m4_2 =10'b0;

   // m4_3 = W*in
   wire signed [9:0] m4_3;
   assign m4_3 =10'b0;

   // m4_4 = W*in
   wire signed [9:0] m4_4;
   assign m4_4 =10'b0;

   // m4_5 = W*in
   wire signed [9:0] m4_5;
   assign m4_5 =10'b0;

   // m4_6 = W*in
   wire signed [9:0] m4_6;
   assign m4_6 =10'b0;

   // m4_7 = W*in
   wire signed [9:0] m4_7;
   assign m4_7 =10'b0;

   // m4_8 = W*in
   wire signed [9:0] m4_8;
   assign m4_8 =10'b0;

   // m4_9 = W*in
   wire signed [9:0] m4_9;
   assign m4_9 =10'b0;

   // m4_10 = W*in
   wire signed [9:0] m4_10;
   assign m4_10 =10'b0;

   // m4_11 = W*in
   wire signed [9:0] m4_11;
   assign m4_11 =10'b0;

   // m4_12 = W*in
   wire signed [9:0] m4_12;
   assign m4_12 =10'b0;

   // m4_13 = W*in
   wire signed [9:0] m4_13;
   assign m4_13 =10'b0;

   // m4_14 = W*in
   wire signed [9:0] m4_14;
   assign m4_14 =10'b0;

   // m4_15 = W*in
   wire signed [9:0] m4_15;
   assign m4_15 =10'b0;

   // m4_16 = W*in
   wire signed [9:0] m4_16;
   assign m4_16 =10'b0;

   // m4_17 = W*in
   wire signed [9:0] m4_17;
   assign m4_17 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_18 = W*in
   wire signed [9:0] m4_18;
   assign m4_18 =10'b0;

   // m4_19 = W*in
   wire signed [9:0] m4_19;
   assign m4_19 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_20 = W*in
   wire signed [9:0] m4_20;
   assign m4_20 =10'b0;

   // m4_21 = W*in
   wire signed [9:0] m4_21;
   assign m4_21 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_22 = W*in
   wire signed [9:0] m4_22;
   assign m4_22 =10'b0;

   // m4_23 = W*in
   wire signed [9:0] m4_23;
   assign m4_23 =10'b0;

   // m4_24 = W*in
   wire signed [9:0] m4_24;
   assign m4_24 =10'b0;

   // m4_25 = W*in
   wire signed [9:0] m4_25;
   assign m4_25 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_26 = W*in
   wire signed [9:0] m4_26;
   assign m4_26 =10'b0;

   // m4_27 = W*in
   wire signed [9:0] m4_27;
   assign m4_27 =10'b0;

   // m4_28 = W*in
   wire signed [9:0] m4_28;
   assign m4_28 =10'b0;

   // m4_29 = W*in
   wire signed [9:0] m4_29;
   assign m4_29 =10'b0;

   // m4_30 = W*in
   wire signed [9:0] m4_30;
   assign m4_30 =10'b0;

   // m4_31 = W*in
   wire signed [9:0] m4_31;
   assign m4_31 =10'b0;

   // m4_32 = W*in
   wire signed [9:0] m4_32;
   assign m4_32 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_33 = W*in
   wire signed [9:0] m4_33;
   assign m4_33 =10'b0;

   // m4_34 = W*in
   wire signed [9:0] m4_34;
   assign m4_34 =10'b0;

   // m4_35 = W*in
   wire signed [9:0] m4_35;
   assign m4_35 =10'b0;

   // m4_36 = W*in
   wire signed [9:0] m4_36;
   assign m4_36 =10'b0;

   // m4_37 = W*in
   wire signed [9:0] m4_37;
   assign m4_37 =10'b0;

   // m4_38 = W*in
   wire signed [9:0] m4_38;
   assign m4_38 =10'b0;

   // m4_39 = W*in
   wire signed [9:0] m4_39;
   assign m4_39 =10'b0;

   // m4_40 = W*in
   wire signed [9:0] m4_40;
   assign m4_40 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_41 = W*in
   wire signed [9:0] m4_41;
   assign m4_41 =10'b0;

   // m4_42 = W*in
   wire signed [9:0] m4_42;
   assign m4_42 =10'b0;

   // m4_43 = W*in
   wire signed [9:0] m4_43;
   assign m4_43 =10'b0;

   // m4_44 = W*in
   wire signed [9:0] m4_44;
   assign m4_44 =10'b0;

   // m4_45 = W*in
   wire signed [9:0] m4_45;
   assign m4_45 =10'b0;

   // m4_46 = W*in
   wire signed [9:0] m4_46;
   assign m4_46 =10'b0;

   // m4_47 = W*in
   wire signed [9:0] m4_47;
   assign m4_47 =10'b0;

   // m4_48 = W*in
   wire signed [9:0] m4_48;
   assign m4_48 =10'b0;

   // m4_49 = W*in
   wire signed [9:0] m4_49;
   assign m4_49 =10'b0;

   // m4_50 = W*in
   wire signed [9:0] m4_50;
   assign m4_50 =10'b0;

   // m4_51 = W*in
   wire signed [9:0] m4_51;
   assign m4_51 =10'b0;

   // m4_52 = W*in
   wire signed [9:0] m4_52;
   assign m4_52 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_53 = W*in
   wire signed [9:0] m4_53;
   assign m4_53 =10'b0;

   // m4_54 = W*in
   wire signed [9:0] m4_54;
   assign m4_54 =10'b0;

   // m4_55 = W*in
   wire signed [9:0] m4_55;
   assign m4_55 =10'b0;

   // m4_56 = W*in
   wire signed [9:0] m4_56;
   assign m4_56 =10'b0;

   // m4_57 = W*in
   wire signed [9:0] m4_57;
   assign m4_57 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_58 = W*in
   wire signed [9:0] m4_58;
   assign m4_58 =10'b0;

   // m4_59 = W*in
   wire signed [9:0] m4_59;
   assign m4_59 =10'b0;

   // m4_60 = W*in
   wire signed [9:0] m4_60;
   assign m4_60 =10'b0;

   // m4_61 = W*in
   wire signed [9:0] m4_61;
   assign m4_61 =10'b0;

   // m4_62 = W*in
   wire signed [9:0] m4_62;
   assign m4_62 =10'b0;

   // m4_63 = W*in
   wire signed [9:0] m4_63;
   assign m4_63 =10'b0;

   // m4_64 = W*in
   wire signed [9:0] m4_64;
   assign m4_64 =10'b0;

   // m4_65 = W*in
   wire signed [9:0] m4_65;
   assign m4_65 =10'b0;

   // m4_66 = W*in
   wire signed [9:0] m4_66;
   assign m4_66 =10'b0;

   // m4_67 = W*in
   wire signed [9:0] m4_67;
   assign m4_67 =10'b0;

   // m4_68 = W*in
   wire signed [9:0] m4_68;
   assign m4_68 =10'b0;

   // m4_69 = W*in
   wire signed [9:0] m4_69;
   assign m4_69 =10'b0;

   // m4_70 = W*in
   wire signed [9:0] m4_70;
   assign m4_70 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_71 = W*in
   wire signed [9:0] m4_71;
   assign m4_71 =10'b0;

   // m4_72 = W*in
   wire signed [9:0] m4_72;
   assign m4_72 =10'b0;

   // m4_73 = W*in
   wire signed [9:0] m4_73;
   assign m4_73 =10'b0;

   // m4_74 = W*in
   wire signed [9:0] m4_74;
   assign m4_74 =10'b0;

   // m4_75 = W*in
   wire signed [9:0] m4_75;
   assign m4_75 =10'b0;

   // m4_76 = W*in
   wire signed [9:0] m4_76;
   assign m4_76 =10'b0;

   // m4_77 = W*in
   wire signed [9:0] m4_77;
   assign m4_77 =10'b0;

   // m4_78 = W*in
   wire signed [9:0] m4_78;
   assign m4_78 =10'b0;

   // m4_79 = W*in
   wire signed [9:0] m4_79;
   assign m4_79 =10'b0;

   // m4_80 = W*in
   wire signed [9:0] m4_80;
   assign m4_80 =10'b0;

   // m4_81 = W*in
   wire signed [9:0] m4_81;
   assign m4_81 =10'b0;

   // m5_1 = W*in
   wire signed [9:0] m5_1;
   assign m5_1 ={ {2{neg5[5]}} , neg5 , {2{1'b0}} };

   // m5_2 = W*in
   wire signed [9:0] m5_2;
   assign m5_2 =10'b0;

   // m5_3 = W*in
   wire signed [9:0] m5_3;
   assign m5_3 =10'b0;

   // m5_4 = W*in
   wire signed [9:0] m5_4;
   assign m5_4 =10'b0;

   // m5_5 = W*in
   wire signed [9:0] m5_5;
   assign m5_5 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_6 = W*in
   wire signed [9:0] m5_6;
   assign m5_6 =10'b0;

   // m5_7 = W*in
   wire signed [9:0] m5_7;
   assign m5_7 =10'b0;

   // m5_8 = W*in
   wire signed [9:0] m5_8;
   assign m5_8 =10'b0;

   // m5_9 = W*in
   wire signed [9:0] m5_9;
   assign m5_9 =10'b0;

   // m5_10 = W*in
   wire signed [9:0] m5_10;
   assign m5_10 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_11 = W*in
   wire signed [9:0] m5_11;
   assign m5_11 =10'b0;

   // m5_12 = W*in
   wire signed [9:0] m5_12;
   assign m5_12 ={ {2{in5[5]}} , in5 , {2{1'b0}} };

   // m5_13 = W*in
   wire signed [9:0] m5_13;
   assign m5_13 =10'b0;

   // m5_14 = W*in
   wire signed [9:0] m5_14;
   assign m5_14 =10'b0;

   // m5_15 = W*in
   wire signed [9:0] m5_15;
   assign m5_15 ={ {2{in5[5]}} , in5 , {2{1'b0}} };

   // m5_16 = W*in
   wire signed [9:0] m5_16;
   assign m5_16 =10'b0;

   // m5_17 = W*in
   wire signed [9:0] m5_17;
   assign m5_17 =10'b0;

   // m5_18 = W*in
   wire signed [9:0] m5_18;
   assign m5_18 ={ {2{neg5[5]}} , neg5 , {2{1'b0}} };

   // m5_19 = W*in
   wire signed [9:0] m5_19;
   assign m5_19 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_20 = W*in
   wire signed [9:0] m5_20;
   assign m5_20 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_21 = W*in
   wire signed [9:0] m5_21;
   assign m5_21 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_22 = W*in
   wire signed [9:0] m5_22;
   assign m5_22 =10'b0;

   // m5_23 = W*in
   wire signed [9:0] m5_23;
   assign m5_23 =10'b0;

   // m5_24 = W*in
   wire signed [9:0] m5_24;
   assign m5_24 =10'b0;

   // m5_25 = W*in
   wire signed [9:0] m5_25;
   assign m5_25 =10'b0;

   // m5_26 = W*in
   wire signed [9:0] m5_26;
   assign m5_26 =10'b0;

   // m5_27 = W*in
   wire signed [9:0] m5_27;
   assign m5_27 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_28 = W*in
   wire signed [9:0] m5_28;
   assign m5_28 =10'b0;

   // m5_29 = W*in
   wire signed [9:0] m5_29;
   assign m5_29 =10'b0;

   // m5_30 = W*in
   wire signed [9:0] m5_30;
   assign m5_30 =10'b0;

   // m5_31 = W*in
   wire signed [9:0] m5_31;
   assign m5_31 =10'b0;

   // m5_32 = W*in
   wire signed [9:0] m5_32;
   assign m5_32 =10'b0;

   // m5_33 = W*in
   wire signed [9:0] m5_33;
   assign m5_33 =10'b0;

   // m5_34 = W*in
   wire signed [9:0] m5_34;
   assign m5_34 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_35 = W*in
   wire signed [9:0] m5_35;
   assign m5_35 =10'b0;

   // m5_36 = W*in
   wire signed [9:0] m5_36;
   assign m5_36 =10'b0;

   // m5_37 = W*in
   wire signed [9:0] m5_37;
   assign m5_37 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_38 = W*in
   wire signed [9:0] m5_38;
   assign m5_38 =10'b0;

   // m5_39 = W*in
   wire signed [9:0] m5_39;
   assign m5_39 =10'b0;

   // m5_40 = W*in
   wire signed [9:0] m5_40;
   assign m5_40 =10'b0;

   // m5_41 = W*in
   wire signed [9:0] m5_41;
   assign m5_41 =10'b0;

   // m5_42 = W*in
   wire signed [9:0] m5_42;
   assign m5_42 =10'b0;

   // m5_43 = W*in
   wire signed [9:0] m5_43;
   assign m5_43 =10'b0;

   // m5_44 = W*in
   wire signed [9:0] m5_44;
   assign m5_44 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_45 = W*in
   wire signed [9:0] m5_45;
   assign m5_45 =10'b0;

   // m5_46 = W*in
   wire signed [9:0] m5_46;
   assign m5_46 =10'b0;

   // m5_47 = W*in
   wire signed [9:0] m5_47;
   assign m5_47 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_48 = W*in
   wire signed [9:0] m5_48;
   assign m5_48 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_49 = W*in
   wire signed [9:0] m5_49;
   assign m5_49 ={ {2{in5[5]}} , in5 , {2{1'b0}} };

   // m5_50 = W*in
   wire signed [9:0] m5_50;
   assign m5_50 =10'b0;

   // m5_51 = W*in
   wire signed [9:0] m5_51;
   assign m5_51 =10'b0;

   // m5_52 = W*in
   wire signed [9:0] m5_52;
   assign m5_52 =10'b0;

   // m5_53 = W*in
   wire signed [9:0] m5_53;
   assign m5_53 =10'b0;

   // m5_54 = W*in
   wire signed [9:0] m5_54;
   assign m5_54 =10'b0;

   // m5_55 = W*in
   wire signed [9:0] m5_55;
   assign m5_55 =10'b0;

   // m5_56 = W*in
   wire signed [9:0] m5_56;
   assign m5_56 =10'b0;

   // m5_57 = W*in
   wire signed [9:0] m5_57;
   assign m5_57 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_58 = W*in
   wire signed [9:0] m5_58;
   assign m5_58 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_59 = W*in
   wire signed [9:0] m5_59;
   assign m5_59 =10'b0;

   // m5_60 = W*in
   wire signed [9:0] m5_60;
   assign m5_60 =10'b0;

   // m5_61 = W*in
   wire signed [9:0] m5_61;
   assign m5_61 =10'b0;

   // m5_62 = W*in
   wire signed [9:0] m5_62;
   assign m5_62 =10'b0;

   // m5_63 = W*in
   wire signed [9:0] m5_63;
   assign m5_63 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_64 = W*in
   wire signed [9:0] m5_64;
   assign m5_64 =10'b0;

   // m5_65 = W*in
   wire signed [9:0] m5_65;
   assign m5_65 =10'b0;

   // m5_66 = W*in
   wire signed [9:0] m5_66;
   assign m5_66 =10'b0;

   // m5_67 = W*in
   wire signed [9:0] m5_67;
   assign m5_67 =10'b0;

   // m5_68 = W*in
   wire signed [9:0] m5_68;
   assign m5_68 =10'b0;

   // m5_69 = W*in
   wire signed [9:0] m5_69;
   assign m5_69 ={ {3{in5[5]}} , in5 , {1{1'b0}} };

   // m5_70 = W*in
   wire signed [9:0] m5_70;
   assign m5_70 =10'b0;

   // m5_71 = W*in
   wire signed [9:0] m5_71;
   assign m5_71 =10'b0;

   // m5_72 = W*in
   wire signed [9:0] m5_72;
   assign m5_72 =10'b0;

   // m5_73 = W*in
   wire signed [9:0] m5_73;
   assign m5_73 =10'b0;

   // m5_74 = W*in
   wire signed [9:0] m5_74;
   assign m5_74 =10'b0;

   // m5_75 = W*in
   wire signed [9:0] m5_75;
   assign m5_75 =10'b0;

   // m5_76 = W*in
   wire signed [9:0] m5_76;
   assign m5_76 =10'b0;

   // m5_77 = W*in
   wire signed [9:0] m5_77;
   assign m5_77 =10'b0;

   // m5_78 = W*in
   wire signed [9:0] m5_78;
   assign m5_78 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_79 = W*in
   wire signed [9:0] m5_79;
   assign m5_79 =10'b0;

   // m5_80 = W*in
   wire signed [9:0] m5_80;
   assign m5_80 =10'b0;

   // m5_81 = W*in
   wire signed [9:0] m5_81;
   assign m5_81 =10'b0;

   // m6_1 = W*in
   wire signed [9:0] m6_1;
   assign m6_1 =10'b0;

   // m6_2 = W*in
   wire signed [9:0] m6_2;
   assign m6_2 =10'b0;

   // m6_3 = W*in
   wire signed [9:0] m6_3;
   assign m6_3 =10'b0;

   // m6_4 = W*in
   wire signed [9:0] m6_4;
   assign m6_4 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_5 = W*in
   wire signed [9:0] m6_5;
   assign m6_5 =10'b0;

   // m6_6 = W*in
   wire signed [9:0] m6_6;
   assign m6_6 ={ {2{in6[5]}} , in6 , {2{1'b0}} };

   // m6_7 = W*in
   wire signed [9:0] m6_7;
   assign m6_7 =10'b0;

   // m6_8 = W*in
   wire signed [9:0] m6_8;
   assign m6_8 =10'b0;

   // m6_9 = W*in
   wire signed [9:0] m6_9;
   assign m6_9 =10'b0;

   // m6_10 = W*in
   wire signed [9:0] m6_10;
   assign m6_10 =10'b0;

   // m6_11 = W*in
   wire signed [9:0] m6_11;
   assign m6_11 =10'b0;

   // m6_12 = W*in
   wire signed [9:0] m6_12;
   assign m6_12 =10'b0;

   // m6_13 = W*in
   wire signed [9:0] m6_13;
   assign m6_13 =10'b0;

   // m6_14 = W*in
   wire signed [9:0] m6_14;
   assign m6_14 =10'b0;

   // m6_15 = W*in
   wire signed [9:0] m6_15;
   assign m6_15 =10'b0;

   // m6_16 = W*in
   wire signed [9:0] m6_16;
   assign m6_16 =10'b0;

   // m6_17 = W*in
   wire signed [9:0] m6_17;
   assign m6_17 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_18 = W*in
   wire signed [9:0] m6_18;
   assign m6_18 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_19 = W*in
   wire signed [9:0] m6_19;
   assign m6_19 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_20 = W*in
   wire signed [9:0] m6_20;
   assign m6_20 =10'b0;

   // m6_21 = W*in
   wire signed [9:0] m6_21;
   assign m6_21 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_22 = W*in
   wire signed [9:0] m6_22;
   assign m6_22 =10'b0;

   // m6_23 = W*in
   wire signed [9:0] m6_23;
   assign m6_23 =10'b0;

   // m6_24 = W*in
   wire signed [9:0] m6_24;
   assign m6_24 =10'b0;

   // m6_25 = W*in
   wire signed [9:0] m6_25;
   assign m6_25 =10'b0;

   // m6_26 = W*in
   wire signed [9:0] m6_26;
   assign m6_26 =10'b0;

   // m6_27 = W*in
   wire signed [9:0] m6_27;
   assign m6_27 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_28 = W*in
   wire signed [9:0] m6_28;
   assign m6_28 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_29 = W*in
   wire signed [9:0] m6_29;
   assign m6_29 =10'b0;

   // m6_30 = W*in
   wire signed [9:0] m6_30;
   assign m6_30 =10'b0;

   // m6_31 = W*in
   wire signed [9:0] m6_31;
   assign m6_31 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_32 = W*in
   wire signed [9:0] m6_32;
   assign m6_32 =10'b0;

   // m6_33 = W*in
   wire signed [9:0] m6_33;
   assign m6_33 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_34 = W*in
   wire signed [9:0] m6_34;
   assign m6_34 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_35 = W*in
   wire signed [9:0] m6_35;
   assign m6_35 =10'b0;

   // m6_36 = W*in
   wire signed [9:0] m6_36;
   assign m6_36 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_37 = W*in
   wire signed [9:0] m6_37;
   assign m6_37 =10'b0;

   // m6_38 = W*in
   wire signed [9:0] m6_38;
   assign m6_38 =10'b0;

   // m6_39 = W*in
   wire signed [9:0] m6_39;
   assign m6_39 =10'b0;

   // m6_40 = W*in
   wire signed [9:0] m6_40;
   assign m6_40 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_41 = W*in
   wire signed [9:0] m6_41;
   assign m6_41 =10'b0;

   // m6_42 = W*in
   wire signed [9:0] m6_42;
   assign m6_42 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_43 = W*in
   wire signed [9:0] m6_43;
   assign m6_43 =10'b0;

   // m6_44 = W*in
   wire signed [9:0] m6_44;
   assign m6_44 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_45 = W*in
   wire signed [9:0] m6_45;
   assign m6_45 =10'b0;

   // m6_46 = W*in
   wire signed [9:0] m6_46;
   assign m6_46 =10'b0;

   // m6_47 = W*in
   wire signed [9:0] m6_47;
   assign m6_47 =10'b0;

   // m6_48 = W*in
   wire signed [9:0] m6_48;
   assign m6_48 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_49 = W*in
   wire signed [9:0] m6_49;
   assign m6_49 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_50 = W*in
   wire signed [9:0] m6_50;
   assign m6_50 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_51 = W*in
   wire signed [9:0] m6_51;
   assign m6_51 =10'b0;

   // m6_52 = W*in
   wire signed [9:0] m6_52;
   assign m6_52 =10'b0;

   // m6_53 = W*in
   wire signed [9:0] m6_53;
   assign m6_53 ={ {2{in6[5]}} , in6 , {2{1'b0}} };

   // m6_54 = W*in
   wire signed [9:0] m6_54;
   assign m6_54 =10'b0;

   // m6_55 = W*in
   wire signed [9:0] m6_55;
   assign m6_55 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_56 = W*in
   wire signed [9:0] m6_56;
   assign m6_56 =10'b0;

   // m6_57 = W*in
   wire signed [9:0] m6_57;
   assign m6_57 =10'b0;

   // m6_58 = W*in
   wire signed [9:0] m6_58;
   assign m6_58 =10'b0;

   // m6_59 = W*in
   wire signed [9:0] m6_59;
   assign m6_59 =10'b0;

   // m6_60 = W*in
   wire signed [9:0] m6_60;
   assign m6_60 ={ {3{in6[5]}} , in6 , {1{1'b0}} };

   // m6_61 = W*in
   wire signed [9:0] m6_61;
   assign m6_61 ={ {2{in6[5]}} , in6 , {2{1'b0}} };

   // m6_62 = W*in
   wire signed [9:0] m6_62;
   assign m6_62 =10'b0;

   // m6_63 = W*in
   wire signed [9:0] m6_63;
   assign m6_63 =10'b0;

   // m6_64 = W*in
   wire signed [9:0] m6_64;
   assign m6_64 ={ {3{neg6[5]}} , neg6 , {1{1'b0}} };

   // m6_65 = W*in
   wire signed [9:0] m6_65;
   assign m6_65 =10'b0;

   // m6_66 = W*in
   wire signed [9:0] m6_66;
   assign m6_66 =10'b0;

   // m6_67 = W*in
   wire signed [9:0] m6_67;
   assign m6_67 =10'b0;

   // m6_68 = W*in
   wire signed [9:0] m6_68;
   assign m6_68 ={ {2{in6[5]}} , in6 , {2{1'b0}} };

   // m6_69 = W*in
   wire signed [9:0] m6_69;
   assign m6_69 =10'b0;

   // m6_70 = W*in
   wire signed [9:0] m6_70;
   assign m6_70 =10'b0;

   // m6_71 = W*in
   wire signed [9:0] m6_71;
   assign m6_71 =10'b0;

   // m6_72 = W*in
   wire signed [9:0] m6_72;
   assign m6_72 =10'b0;

   // m6_73 = W*in
   wire signed [9:0] m6_73;
   assign m6_73 =10'b0;

   // m6_74 = W*in
   wire signed [9:0] m6_74;
   assign m6_74 =10'b0;

   // m6_75 = W*in
   wire signed [9:0] m6_75;
   assign m6_75 =10'b0;

   // m6_76 = W*in
   wire signed [9:0] m6_76;
   assign m6_76 ={ {2{in6[5]}} , in6 , {2{1'b0}} };

   // m6_77 = W*in
   wire signed [9:0] m6_77;
   assign m6_77 =10'b0;

   // m6_78 = W*in
   wire signed [9:0] m6_78;
   assign m6_78 =10'b0;

   // m6_79 = W*in
   wire signed [9:0] m6_79;
   assign m6_79 =10'b0;

   // m6_80 = W*in
   wire signed [9:0] m6_80;
   assign m6_80 =10'b0;

   // m6_81 = W*in
   wire signed [9:0] m6_81;
   assign m6_81 =10'b0;

   // m7_1 = W*in
   wire signed [9:0] m7_1;
   assign m7_1 =10'b0;

   // m7_2 = W*in
   wire signed [9:0] m7_2;
   assign m7_2 =10'b0;

   // m7_3 = W*in
   wire signed [9:0] m7_3;
   assign m7_3 =10'b0;

   // m7_4 = W*in
   wire signed [9:0] m7_4;
   assign m7_4 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_5 = W*in
   wire signed [9:0] m7_5;
   assign m7_5 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_6 = W*in
   wire signed [9:0] m7_6;
   assign m7_6 ={ {2{neg7[5]}} , neg7 , {2{1'b0}} };

   // m7_7 = W*in
   wire signed [9:0] m7_7;
   assign m7_7 =10'b0;

   // m7_8 = W*in
   wire signed [9:0] m7_8;
   assign m7_8 =10'b0;

   // m7_9 = W*in
   wire signed [9:0] m7_9;
   assign m7_9 =10'b0;

   // m7_10 = W*in
   wire signed [9:0] m7_10;
   assign m7_10 =10'b0;

   // m7_11 = W*in
   wire signed [9:0] m7_11;
   assign m7_11 =10'b0;

   // m7_12 = W*in
   wire signed [9:0] m7_12;
   assign m7_12 =10'b0;

   // m7_13 = W*in
   wire signed [9:0] m7_13;
   assign m7_13 =10'b0;

   // m7_14 = W*in
   wire signed [9:0] m7_14;
   assign m7_14 =10'b0;

   // m7_15 = W*in
   wire signed [9:0] m7_15;
   assign m7_15 ={ {2{in7[5]}} , in7 , {2{1'b0}} };

   // m7_16 = W*in
   wire signed [9:0] m7_16;
   assign m7_16 =10'b0;

   // m7_17 = W*in
   wire signed [9:0] m7_17;
   assign m7_17 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_18 = W*in
   wire signed [9:0] m7_18;
   assign m7_18 =10'b0;

   // m7_19 = W*in
   wire signed [9:0] m7_19;
   assign m7_19 =10'b0;

   // m7_20 = W*in
   wire signed [9:0] m7_20;
   assign m7_20 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_21 = W*in
   wire signed [9:0] m7_21;
   assign m7_21 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_22 = W*in
   wire signed [9:0] m7_22;
   assign m7_22 =10'b0;

   // m7_23 = W*in
   wire signed [9:0] m7_23;
   assign m7_23 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_24 = W*in
   wire signed [9:0] m7_24;
   assign m7_24 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_25 = W*in
   wire signed [9:0] m7_25;
   assign m7_25 =10'b0;

   // m7_26 = W*in
   wire signed [9:0] m7_26;
   assign m7_26 =10'b0;

   // m7_27 = W*in
   wire signed [9:0] m7_27;
   assign m7_27 =10'b0;

   // m7_28 = W*in
   wire signed [9:0] m7_28;
   assign m7_28 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_29 = W*in
   wire signed [9:0] m7_29;
   assign m7_29 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_30 = W*in
   wire signed [9:0] m7_30;
   assign m7_30 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_31 = W*in
   wire signed [9:0] m7_31;
   assign m7_31 =10'b0;

   // m7_32 = W*in
   wire signed [9:0] m7_32;
   assign m7_32 =10'b0;

   // m7_33 = W*in
   wire signed [9:0] m7_33;
   assign m7_33 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_34 = W*in
   wire signed [9:0] m7_34;
   assign m7_34 =10'b0;

   // m7_35 = W*in
   wire signed [9:0] m7_35;
   assign m7_35 =10'b0;

   // m7_36 = W*in
   wire signed [9:0] m7_36;
   assign m7_36 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_37 = W*in
   wire signed [9:0] m7_37;
   assign m7_37 =10'b0;

   // m7_38 = W*in
   wire signed [9:0] m7_38;
   assign m7_38 =10'b0;

   // m7_39 = W*in
   wire signed [9:0] m7_39;
   assign m7_39 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_40 = W*in
   wire signed [9:0] m7_40;
   assign m7_40 =10'b0;

   // m7_41 = W*in
   wire signed [9:0] m7_41;
   assign m7_41 =10'b0;

   // m7_42 = W*in
   wire signed [9:0] m7_42;
   assign m7_42 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_43 = W*in
   wire signed [9:0] m7_43;
   assign m7_43 ={ {2{in7[5]}} , in7 , {2{1'b0}} };

   // m7_44 = W*in
   wire signed [9:0] m7_44;
   assign m7_44 ={ {2{in7[5]}} , in7 , {2{1'b0}} };

   // m7_45 = W*in
   wire signed [9:0] m7_45;
   assign m7_45 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_46 = W*in
   wire signed [9:0] m7_46;
   assign m7_46 =10'b0;

   // m7_47 = W*in
   wire signed [9:0] m7_47;
   assign m7_47 =10'b0;

   // m7_48 = W*in
   wire signed [9:0] m7_48;
   assign m7_48 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_49 = W*in
   wire signed [9:0] m7_49;
   assign m7_49 =10'b0;

   // m7_50 = W*in
   wire signed [9:0] m7_50;
   assign m7_50 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_51 = W*in
   wire signed [9:0] m7_51;
   assign m7_51 =10'b0;

   // m7_52 = W*in
   wire signed [9:0] m7_52;
   assign m7_52 =10'b0;

   // m7_53 = W*in
   wire signed [9:0] m7_53;
   assign m7_53 =10'b0;

   // m7_54 = W*in
   wire signed [9:0] m7_54;
   assign m7_54 =10'b0;

   // m7_55 = W*in
   wire signed [9:0] m7_55;
   assign m7_55 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_56 = W*in
   wire signed [9:0] m7_56;
   assign m7_56 ={ {3{neg7[5]}} , neg7 , {1{1'b0}} };

   // m7_57 = W*in
   wire signed [9:0] m7_57;
   assign m7_57 =10'b0;

   // m7_58 = W*in
   wire signed [9:0] m7_58;
   assign m7_58 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_59 = W*in
   wire signed [9:0] m7_59;
   assign m7_59 =10'b0;

   // m7_60 = W*in
   wire signed [9:0] m7_60;
   assign m7_60 =10'b0;

   // m7_61 = W*in
   wire signed [9:0] m7_61;
   assign m7_61 =10'b0;

   // m7_62 = W*in
   wire signed [9:0] m7_62;
   assign m7_62 ={ {2{in7[5]}} , in7 , {2{1'b0}} };

   // m7_63 = W*in
   wire signed [9:0] m7_63;
   assign m7_63 =10'b0;

   // m7_64 = W*in
   wire signed [9:0] m7_64;
   assign m7_64 =10'b0;

   // m7_65 = W*in
   wire signed [9:0] m7_65;
   assign m7_65 =10'b0;

   // m7_66 = W*in
   wire signed [9:0] m7_66;
   assign m7_66 ={ {2{in7[5]}} , in7 , {2{1'b0}} };

   // m7_67 = W*in
   wire signed [9:0] m7_67;
   assign m7_67 =10'b0;

   // m7_68 = W*in
   wire signed [9:0] m7_68;
   assign m7_68 ={ {2{neg7[5]}} , neg7 , {2{1'b0}} };

   // m7_69 = W*in
   wire signed [9:0] m7_69;
   assign m7_69 =10'b0;

   // m7_70 = W*in
   wire signed [9:0] m7_70;
   assign m7_70 =10'b0;

   // m7_71 = W*in
   wire signed [9:0] m7_71;
   assign m7_71 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_72 = W*in
   wire signed [9:0] m7_72;
   assign m7_72 =10'b0;

   // m7_73 = W*in
   wire signed [9:0] m7_73;
   assign m7_73 =10'b0;

   // m7_74 = W*in
   wire signed [9:0] m7_74;
   assign m7_74 =10'b0;

   // m7_75 = W*in
   wire signed [9:0] m7_75;
   assign m7_75 =10'b0;

   // m7_76 = W*in
   wire signed [9:0] m7_76;
   assign m7_76 =10'b0;

   // m7_77 = W*in
   wire signed [9:0] m7_77;
   assign m7_77 =10'b0;

   // m7_78 = W*in
   wire signed [9:0] m7_78;
   assign m7_78 =10'b0;

   // m7_79 = W*in
   wire signed [9:0] m7_79;
   assign m7_79 =10'b0;

   // m7_80 = W*in
   wire signed [9:0] m7_80;
   assign m7_80 ={ {2{in7[5]}} , in7 , {2{1'b0}} };

   // m7_81 = W*in
   wire signed [9:0] m7_81;
   assign m7_81 =10'b0;

   // m8_1 = W*in
   wire signed [9:0] m8_1;
   assign m8_1 =10'b0;

   // m8_2 = W*in
   wire signed [9:0] m8_2;
   assign m8_2 =10'b0;

   // m8_3 = W*in
   wire signed [9:0] m8_3;
   assign m8_3 =10'b0;

   // m8_4 = W*in
   wire signed [9:0] m8_4;
   assign m8_4 =10'b0;

   // m8_5 = W*in
   wire signed [9:0] m8_5;
   assign m8_5 =10'b0;

   // m8_6 = W*in
   wire signed [9:0] m8_6;
   assign m8_6 =10'b0;

   // m8_7 = W*in
   wire signed [9:0] m8_7;
   assign m8_7 =10'b0;

   // m8_8 = W*in
   wire signed [9:0] m8_8;
   assign m8_8 =10'b0;

   // m8_9 = W*in
   wire signed [9:0] m8_9;
   assign m8_9 =10'b0;

   // m8_10 = W*in
   wire signed [9:0] m8_10;
   assign m8_10 =10'b0;

   // m8_11 = W*in
   wire signed [9:0] m8_11;
   assign m8_11 =10'b0;

   // m8_12 = W*in
   wire signed [9:0] m8_12;
   assign m8_12 =10'b0;

   // m8_13 = W*in
   wire signed [9:0] m8_13;
   assign m8_13 =10'b0;

   // m8_14 = W*in
   wire signed [9:0] m8_14;
   assign m8_14 =10'b0;

   // m8_15 = W*in
   wire signed [9:0] m8_15;
   assign m8_15 ={ {3{in8[5]}} , in8 , {1{1'b0}} };

   // m8_16 = W*in
   wire signed [9:0] m8_16;
   assign m8_16 =10'b0;

   // m8_17 = W*in
   wire signed [9:0] m8_17;
   assign m8_17 =10'b0;

   // m8_18 = W*in
   wire signed [9:0] m8_18;
   assign m8_18 =10'b0;

   // m8_19 = W*in
   wire signed [9:0] m8_19;
   assign m8_19 =10'b0;

   // m8_20 = W*in
   wire signed [9:0] m8_20;
   assign m8_20 ={ {3{in8[5]}} , in8 , {1{1'b0}} };

   // m8_21 = W*in
   wire signed [9:0] m8_21;
   assign m8_21 =10'b0;

   // m8_22 = W*in
   wire signed [9:0] m8_22;
   assign m8_22 ={ {3{in8[5]}} , in8 , {1{1'b0}} };

   // m8_23 = W*in
   wire signed [9:0] m8_23;
   assign m8_23 =10'b0;

   // m8_24 = W*in
   wire signed [9:0] m8_24;
   assign m8_24 ={ {3{in8[5]}} , in8 , {1{1'b0}} };

   // m8_25 = W*in
   wire signed [9:0] m8_25;
   assign m8_25 =10'b0;

   // m8_26 = W*in
   wire signed [9:0] m8_26;
   assign m8_26 =10'b0;

   // m8_27 = W*in
   wire signed [9:0] m8_27;
   assign m8_27 =10'b0;

   // m8_28 = W*in
   wire signed [9:0] m8_28;
   assign m8_28 =10'b0;

   // m8_29 = W*in
   wire signed [9:0] m8_29;
   assign m8_29 ={ {3{in8[5]}} , in8 , {1{1'b0}} };

   // m8_30 = W*in
   wire signed [9:0] m8_30;
   assign m8_30 =10'b0;

   // m8_31 = W*in
   wire signed [9:0] m8_31;
   assign m8_31 =10'b0;

   // m8_32 = W*in
   wire signed [9:0] m8_32;
   assign m8_32 =10'b0;

   // m8_33 = W*in
   wire signed [9:0] m8_33;
   assign m8_33 ={ {3{neg8[5]}} , neg8 , {1{1'b0}} };

   // m8_34 = W*in
   wire signed [9:0] m8_34;
   assign m8_34 =10'b0;

   // m8_35 = W*in
   wire signed [9:0] m8_35;
   assign m8_35 =10'b0;

   // m8_36 = W*in
   wire signed [9:0] m8_36;
   assign m8_36 =10'b0;

   // m8_37 = W*in
   wire signed [9:0] m8_37;
   assign m8_37 =10'b0;

   // m8_38 = W*in
   wire signed [9:0] m8_38;
   assign m8_38 =10'b0;

   // m8_39 = W*in
   wire signed [9:0] m8_39;
   assign m8_39 =10'b0;

   // m8_40 = W*in
   wire signed [9:0] m8_40;
   assign m8_40 ={ {3{in8[5]}} , in8 , {1{1'b0}} };

   // m8_41 = W*in
   wire signed [9:0] m8_41;
   assign m8_41 =10'b0;

   // m8_42 = W*in
   wire signed [9:0] m8_42;
   assign m8_42 =10'b0;

   // m8_43 = W*in
   wire signed [9:0] m8_43;
   assign m8_43 =10'b0;

   // m8_44 = W*in
   wire signed [9:0] m8_44;
   assign m8_44 ={ {2{in8[5]}} , in8 , {2{1'b0}} };

   // m8_45 = W*in
   wire signed [9:0] m8_45;
   assign m8_45 =10'b0;

   // m8_46 = W*in
   wire signed [9:0] m8_46;
   assign m8_46 =10'b0;

   // m8_47 = W*in
   wire signed [9:0] m8_47;
   assign m8_47 =10'b0;

   // m8_48 = W*in
   wire signed [9:0] m8_48;
   assign m8_48 =10'b0;

   // m8_49 = W*in
   wire signed [9:0] m8_49;
   assign m8_49 =10'b0;

   // m8_50 = W*in
   wire signed [9:0] m8_50;
   assign m8_50 =10'b0;

   // m8_51 = W*in
   wire signed [9:0] m8_51;
   assign m8_51 =10'b0;

   // m8_52 = W*in
   wire signed [9:0] m8_52;
   assign m8_52 =10'b0;

   // m8_53 = W*in
   wire signed [9:0] m8_53;
   assign m8_53 =10'b0;

   // m8_54 = W*in
   wire signed [9:0] m8_54;
   assign m8_54 =10'b0;

   // m8_55 = W*in
   wire signed [9:0] m8_55;
   assign m8_55 =10'b0;

   // m8_56 = W*in
   wire signed [9:0] m8_56;
   assign m8_56 =10'b0;

   // m8_57 = W*in
   wire signed [9:0] m8_57;
   assign m8_57 =10'b0;

   // m8_58 = W*in
   wire signed [9:0] m8_58;
   assign m8_58 =10'b0;

   // m8_59 = W*in
   wire signed [9:0] m8_59;
   assign m8_59 =10'b0;

   // m8_60 = W*in
   wire signed [9:0] m8_60;
   assign m8_60 =10'b0;

   // m8_61 = W*in
   wire signed [9:0] m8_61;
   assign m8_61 =10'b0;

   // m8_62 = W*in
   wire signed [9:0] m8_62;
   assign m8_62 =10'b0;

   // m8_63 = W*in
   wire signed [9:0] m8_63;
   assign m8_63 =10'b0;

   // m8_64 = W*in
   wire signed [9:0] m8_64;
   assign m8_64 =10'b0;

   // m8_65 = W*in
   wire signed [9:0] m8_65;
   assign m8_65 =10'b0;

   // m8_66 = W*in
   wire signed [9:0] m8_66;
   assign m8_66 =10'b0;

   // m8_67 = W*in
   wire signed [9:0] m8_67;
   assign m8_67 =10'b0;

   // m8_68 = W*in
   wire signed [9:0] m8_68;
   assign m8_68 =10'b0;

   // m8_69 = W*in
   wire signed [9:0] m8_69;
   assign m8_69 =10'b0;

   // m8_70 = W*in
   wire signed [9:0] m8_70;
   assign m8_70 =10'b0;

   // m8_71 = W*in
   wire signed [9:0] m8_71;
   assign m8_71 =10'b0;

   // m8_72 = W*in
   wire signed [9:0] m8_72;
   assign m8_72 =10'b0;

   // m8_73 = W*in
   wire signed [9:0] m8_73;
   assign m8_73 =10'b0;

   // m8_74 = W*in
   wire signed [9:0] m8_74;
   assign m8_74 =10'b0;

   // m8_75 = W*in
   wire signed [9:0] m8_75;
   assign m8_75 =10'b0;

   // m8_76 = W*in
   wire signed [9:0] m8_76;
   assign m8_76 =10'b0;

   // m8_77 = W*in
   wire signed [9:0] m8_77;
   assign m8_77 =10'b0;

   // m8_78 = W*in
   wire signed [9:0] m8_78;
   assign m8_78 =10'b0;

   // m8_79 = W*in
   wire signed [9:0] m8_79;
   assign m8_79 =10'b0;

   // m8_80 = W*in
   wire signed [9:0] m8_80;
   assign m8_80 =10'b0;

   // m8_81 = W*in
   wire signed [9:0] m8_81;
   assign m8_81 =10'b0;

   // m9_1 = W*in
   wire signed [9:0] m9_1;
   assign m9_1 =10'b0;

   // m9_2 = W*in
   wire signed [9:0] m9_2;
   assign m9_2 =10'b0;

   // m9_3 = W*in
   wire signed [9:0] m9_3;
   assign m9_3 =10'b0;

   // m9_4 = W*in
   wire signed [9:0] m9_4;
   assign m9_4 =10'b0;

   // m9_5 = W*in
   wire signed [9:0] m9_5;
   assign m9_5 =10'b0;

   // m9_6 = W*in
   wire signed [9:0] m9_6;
   assign m9_6 =10'b0;

   // m9_7 = W*in
   wire signed [9:0] m9_7;
   assign m9_7 =10'b0;

   // m9_8 = W*in
   wire signed [9:0] m9_8;
   assign m9_8 =10'b0;

   // m9_9 = W*in
   wire signed [9:0] m9_9;
   assign m9_9 =10'b0;

   // m9_10 = W*in
   wire signed [9:0] m9_10;
   assign m9_10 =10'b0;

   // m9_11 = W*in
   wire signed [9:0] m9_11;
   assign m9_11 =10'b0;

   // m9_12 = W*in
   wire signed [9:0] m9_12;
   assign m9_12 =10'b0;

   // m9_13 = W*in
   wire signed [9:0] m9_13;
   assign m9_13 =10'b0;

   // m9_14 = W*in
   wire signed [9:0] m9_14;
   assign m9_14 =10'b0;

   // m9_15 = W*in
   wire signed [9:0] m9_15;
   assign m9_15 =10'b0;

   // m9_16 = W*in
   wire signed [9:0] m9_16;
   assign m9_16 =10'b0;

   // m9_17 = W*in
   wire signed [9:0] m9_17;
   assign m9_17 =10'b0;

   // m9_18 = W*in
   wire signed [9:0] m9_18;
   assign m9_18 =10'b0;

   // m9_19 = W*in
   wire signed [9:0] m9_19;
   assign m9_19 =10'b0;

   // m9_20 = W*in
   wire signed [9:0] m9_20;
   assign m9_20 =10'b0;

   // m9_21 = W*in
   wire signed [9:0] m9_21;
   assign m9_21 =10'b0;

   // m9_22 = W*in
   wire signed [9:0] m9_22;
   assign m9_22 =10'b0;

   // m9_23 = W*in
   wire signed [9:0] m9_23;
   assign m9_23 =10'b0;

   // m9_24 = W*in
   wire signed [9:0] m9_24;
   assign m9_24 =10'b0;

   // m9_25 = W*in
   wire signed [9:0] m9_25;
   assign m9_25 ={ {3{in9[5]}} , in9 , {1{1'b0}} };

   // m9_26 = W*in
   wire signed [9:0] m9_26;
   assign m9_26 =10'b0;

   // m9_27 = W*in
   wire signed [9:0] m9_27;
   assign m9_27 =10'b0;

   // m9_28 = W*in
   wire signed [9:0] m9_28;
   assign m9_28 =10'b0;

   // m9_29 = W*in
   wire signed [9:0] m9_29;
   assign m9_29 =10'b0;

   // m9_30 = W*in
   wire signed [9:0] m9_30;
   assign m9_30 =10'b0;

   // m9_31 = W*in
   wire signed [9:0] m9_31;
   assign m9_31 =10'b0;

   // m9_32 = W*in
   wire signed [9:0] m9_32;
   assign m9_32 =10'b0;

   // m9_33 = W*in
   wire signed [9:0] m9_33;
   assign m9_33 =10'b0;

   // m9_34 = W*in
   wire signed [9:0] m9_34;
   assign m9_34 =10'b0;

   // m9_35 = W*in
   wire signed [9:0] m9_35;
   assign m9_35 =10'b0;

   // m9_36 = W*in
   wire signed [9:0] m9_36;
   assign m9_36 =10'b0;

   // m9_37 = W*in
   wire signed [9:0] m9_37;
   assign m9_37 =10'b0;

   // m9_38 = W*in
   wire signed [9:0] m9_38;
   assign m9_38 =10'b0;

   // m9_39 = W*in
   wire signed [9:0] m9_39;
   assign m9_39 =10'b0;

   // m9_40 = W*in
   wire signed [9:0] m9_40;
   assign m9_40 =10'b0;

   // m9_41 = W*in
   wire signed [9:0] m9_41;
   assign m9_41 =10'b0;

   // m9_42 = W*in
   wire signed [9:0] m9_42;
   assign m9_42 =10'b0;

   // m9_43 = W*in
   wire signed [9:0] m9_43;
   assign m9_43 =10'b0;

   // m9_44 = W*in
   wire signed [9:0] m9_44;
   assign m9_44 =10'b0;

   // m9_45 = W*in
   wire signed [9:0] m9_45;
   assign m9_45 =10'b0;

   // m9_46 = W*in
   wire signed [9:0] m9_46;
   assign m9_46 =10'b0;

   // m9_47 = W*in
   wire signed [9:0] m9_47;
   assign m9_47 =10'b0;

   // m9_48 = W*in
   wire signed [9:0] m9_48;
   assign m9_48 =10'b0;

   // m9_49 = W*in
   wire signed [9:0] m9_49;
   assign m9_49 =10'b0;

   // m9_50 = W*in
   wire signed [9:0] m9_50;
   assign m9_50 =10'b0;

   // m9_51 = W*in
   wire signed [9:0] m9_51;
   assign m9_51 =10'b0;

   // m9_52 = W*in
   wire signed [9:0] m9_52;
   assign m9_52 =10'b0;

   // m9_53 = W*in
   wire signed [9:0] m9_53;
   assign m9_53 =10'b0;

   // m9_54 = W*in
   wire signed [9:0] m9_54;
   assign m9_54 =10'b0;

   // m9_55 = W*in
   wire signed [9:0] m9_55;
   assign m9_55 =10'b0;

   // m9_56 = W*in
   wire signed [9:0] m9_56;
   assign m9_56 =10'b0;

   // m9_57 = W*in
   wire signed [9:0] m9_57;
   assign m9_57 =10'b0;

   // m9_58 = W*in
   wire signed [9:0] m9_58;
   assign m9_58 =10'b0;

   // m9_59 = W*in
   wire signed [9:0] m9_59;
   assign m9_59 =10'b0;

   // m9_60 = W*in
   wire signed [9:0] m9_60;
   assign m9_60 =10'b0;

   // m9_61 = W*in
   wire signed [9:0] m9_61;
   assign m9_61 =10'b0;

   // m9_62 = W*in
   wire signed [9:0] m9_62;
   assign m9_62 =10'b0;

   // m9_63 = W*in
   wire signed [9:0] m9_63;
   assign m9_63 =10'b0;

   // m9_64 = W*in
   wire signed [9:0] m9_64;
   assign m9_64 =10'b0;

   // m9_65 = W*in
   wire signed [9:0] m9_65;
   assign m9_65 =10'b0;

   // m9_66 = W*in
   wire signed [9:0] m9_66;
   assign m9_66 =10'b0;

   // m9_67 = W*in
   wire signed [9:0] m9_67;
   assign m9_67 =10'b0;

   // m9_68 = W*in
   wire signed [9:0] m9_68;
   assign m9_68 =10'b0;

   // m9_69 = W*in
   wire signed [9:0] m9_69;
   assign m9_69 =10'b0;

   // m9_70 = W*in
   wire signed [9:0] m9_70;
   assign m9_70 =10'b0;

   // m9_71 = W*in
   wire signed [9:0] m9_71;
   assign m9_71 =10'b0;

   // m9_72 = W*in
   wire signed [9:0] m9_72;
   assign m9_72 =10'b0;

   // m9_73 = W*in
   wire signed [9:0] m9_73;
   assign m9_73 =10'b0;

   // m9_74 = W*in
   wire signed [9:0] m9_74;
   assign m9_74 =10'b0;

   // m9_75 = W*in
   wire signed [9:0] m9_75;
   assign m9_75 =10'b0;

   // m9_76 = W*in
   wire signed [9:0] m9_76;
   assign m9_76 =10'b0;

   // m9_77 = W*in
   wire signed [9:0] m9_77;
   assign m9_77 =10'b0;

   // m9_78 = W*in
   wire signed [9:0] m9_78;
   assign m9_78 =10'b0;

   // m9_79 = W*in
   wire signed [9:0] m9_79;
   assign m9_79 =10'b0;

   // m9_80 = W*in
   wire signed [9:0] m9_80;
   assign m9_80 =10'b0;

   // m9_81 = W*in
   wire signed [9:0] m9_81;
   assign m9_81 =10'b0;

   // m10_1 = W*in
   wire signed [9:0] m10_1;
   assign m10_1 =10'b0;

   // m10_2 = W*in
   wire signed [9:0] m10_2;
   assign m10_2 =10'b0;

   // m10_3 = W*in
   wire signed [9:0] m10_3;
   assign m10_3 =10'b0;

   // m10_4 = W*in
   wire signed [9:0] m10_4;
   assign m10_4 =10'b0;

   // m10_5 = W*in
   wire signed [9:0] m10_5;
   assign m10_5 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_6 = W*in
   wire signed [9:0] m10_6;
   assign m10_6 =10'b0;

   // m10_7 = W*in
   wire signed [9:0] m10_7;
   assign m10_7 =10'b0;

   // m10_8 = W*in
   wire signed [9:0] m10_8;
   assign m10_8 =10'b0;

   // m10_9 = W*in
   wire signed [9:0] m10_9;
   assign m10_9 =10'b0;

   // m10_10 = W*in
   wire signed [9:0] m10_10;
   assign m10_10 =10'b0;

   // m10_11 = W*in
   wire signed [9:0] m10_11;
   assign m10_11 =10'b0;

   // m10_12 = W*in
   wire signed [9:0] m10_12;
   assign m10_12 =10'b0;

   // m10_13 = W*in
   wire signed [9:0] m10_13;
   assign m10_13 =10'b0;

   // m10_14 = W*in
   wire signed [9:0] m10_14;
   assign m10_14 =10'b0;

   // m10_15 = W*in
   wire signed [9:0] m10_15;
   assign m10_15 =10'b0;

   // m10_16 = W*in
   wire signed [9:0] m10_16;
   assign m10_16 =10'b0;

   // m10_17 = W*in
   wire signed [9:0] m10_17;
   assign m10_17 =10'b0;

   // m10_18 = W*in
   wire signed [9:0] m10_18;
   assign m10_18 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_19 = W*in
   wire signed [9:0] m10_19;
   assign m10_19 =10'b0;

   // m10_20 = W*in
   wire signed [9:0] m10_20;
   assign m10_20 =10'b0;

   // m10_21 = W*in
   wire signed [9:0] m10_21;
   assign m10_21 =10'b0;

   // m10_22 = W*in
   wire signed [9:0] m10_22;
   assign m10_22 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_23 = W*in
   wire signed [9:0] m10_23;
   assign m10_23 =10'b0;

   // m10_24 = W*in
   wire signed [9:0] m10_24;
   assign m10_24 =10'b0;

   // m10_25 = W*in
   wire signed [9:0] m10_25;
   assign m10_25 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_26 = W*in
   wire signed [9:0] m10_26;
   assign m10_26 =10'b0;

   // m10_27 = W*in
   wire signed [9:0] m10_27;
   assign m10_27 ={ {3{neg10[5]}} , neg10 , {1{1'b0}} };

   // m10_28 = W*in
   wire signed [9:0] m10_28;
   assign m10_28 =10'b0;

   // m10_29 = W*in
   wire signed [9:0] m10_29;
   assign m10_29 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_30 = W*in
   wire signed [9:0] m10_30;
   assign m10_30 ={ {3{neg10[5]}} , neg10 , {1{1'b0}} };

   // m10_31 = W*in
   wire signed [9:0] m10_31;
   assign m10_31 =10'b0;

   // m10_32 = W*in
   wire signed [9:0] m10_32;
   assign m10_32 =10'b0;

   // m10_33 = W*in
   wire signed [9:0] m10_33;
   assign m10_33 =10'b0;

   // m10_34 = W*in
   wire signed [9:0] m10_34;
   assign m10_34 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_35 = W*in
   wire signed [9:0] m10_35;
   assign m10_35 ={ {3{neg10[5]}} , neg10 , {1{1'b0}} };

   // m10_36 = W*in
   wire signed [9:0] m10_36;
   assign m10_36 =10'b0;

   // m10_37 = W*in
   wire signed [9:0] m10_37;
   assign m10_37 =10'b0;

   // m10_38 = W*in
   wire signed [9:0] m10_38;
   assign m10_38 =10'b0;

   // m10_39 = W*in
   wire signed [9:0] m10_39;
   assign m10_39 =10'b0;

   // m10_40 = W*in
   wire signed [9:0] m10_40;
   assign m10_40 =10'b0;

   // m10_41 = W*in
   wire signed [9:0] m10_41;
   assign m10_41 =10'b0;

   // m10_42 = W*in
   wire signed [9:0] m10_42;
   assign m10_42 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_43 = W*in
   wire signed [9:0] m10_43;
   assign m10_43 =10'b0;

   // m10_44 = W*in
   wire signed [9:0] m10_44;
   assign m10_44 =10'b0;

   // m10_45 = W*in
   wire signed [9:0] m10_45;
   assign m10_45 =10'b0;

   // m10_46 = W*in
   wire signed [9:0] m10_46;
   assign m10_46 ={ {3{neg10[5]}} , neg10 , {1{1'b0}} };

   // m10_47 = W*in
   wire signed [9:0] m10_47;
   assign m10_47 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_48 = W*in
   wire signed [9:0] m10_48;
   assign m10_48 =10'b0;

   // m10_49 = W*in
   wire signed [9:0] m10_49;
   assign m10_49 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_50 = W*in
   wire signed [9:0] m10_50;
   assign m10_50 =10'b0;

   // m10_51 = W*in
   wire signed [9:0] m10_51;
   assign m10_51 =10'b0;

   // m10_52 = W*in
   wire signed [9:0] m10_52;
   assign m10_52 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_53 = W*in
   wire signed [9:0] m10_53;
   assign m10_53 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_54 = W*in
   wire signed [9:0] m10_54;
   assign m10_54 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_55 = W*in
   wire signed [9:0] m10_55;
   assign m10_55 =10'b0;

   // m10_56 = W*in
   wire signed [9:0] m10_56;
   assign m10_56 =10'b0;

   // m10_57 = W*in
   wire signed [9:0] m10_57;
   assign m10_57 =10'b0;

   // m10_58 = W*in
   wire signed [9:0] m10_58;
   assign m10_58 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_59 = W*in
   wire signed [9:0] m10_59;
   assign m10_59 =10'b0;

   // m10_60 = W*in
   wire signed [9:0] m10_60;
   assign m10_60 =10'b0;

   // m10_61 = W*in
   wire signed [9:0] m10_61;
   assign m10_61 =10'b0;

   // m10_62 = W*in
   wire signed [9:0] m10_62;
   assign m10_62 ={ {3{neg10[5]}} , neg10 , {1{1'b0}} };

   // m10_63 = W*in
   wire signed [9:0] m10_63;
   assign m10_63 =10'b0;

   // m10_64 = W*in
   wire signed [9:0] m10_64;
   assign m10_64 =10'b0;

   // m10_65 = W*in
   wire signed [9:0] m10_65;
   assign m10_65 =10'b0;

   // m10_66 = W*in
   wire signed [9:0] m10_66;
   assign m10_66 =10'b0;

   // m10_67 = W*in
   wire signed [9:0] m10_67;
   assign m10_67 =10'b0;

   // m10_68 = W*in
   wire signed [9:0] m10_68;
   assign m10_68 =10'b0;

   // m10_69 = W*in
   wire signed [9:0] m10_69;
   assign m10_69 =10'b0;

   // m10_70 = W*in
   wire signed [9:0] m10_70;
   assign m10_70 =10'b0;

   // m10_71 = W*in
   wire signed [9:0] m10_71;
   assign m10_71 =10'b0;

   // m10_72 = W*in
   wire signed [9:0] m10_72;
   assign m10_72 =10'b0;

   // m10_73 = W*in
   wire signed [9:0] m10_73;
   assign m10_73 =10'b0;

   // m10_74 = W*in
   wire signed [9:0] m10_74;
   assign m10_74 =10'b0;

   // m10_75 = W*in
   wire signed [9:0] m10_75;
   assign m10_75 =10'b0;

   // m10_76 = W*in
   wire signed [9:0] m10_76;
   assign m10_76 =10'b0;

   // m10_77 = W*in
   wire signed [9:0] m10_77;
   assign m10_77 ={ {2{in10[5]}} , in10 , {2{1'b0}} };

   // m10_78 = W*in
   wire signed [9:0] m10_78;
   assign m10_78 =10'b0;

   // m10_79 = W*in
   wire signed [9:0] m10_79;
   assign m10_79 ={ {3{neg10[5]}} , neg10 , {1{1'b0}} };

   // m10_80 = W*in
   wire signed [9:0] m10_80;
   assign m10_80 =10'b0;

   // m10_81 = W*in
   wire signed [9:0] m10_81;
   assign m10_81 =10'b0;

   // m11_1 = W*in
   wire signed [9:0] m11_1;
   assign m11_1 =10'b0;

   // m11_2 = W*in
   wire signed [9:0] m11_2;
   assign m11_2 =10'b0;

   // m11_3 = W*in
   wire signed [9:0] m11_3;
   assign m11_3 =10'b0;

   // m11_4 = W*in
   wire signed [9:0] m11_4;
   assign m11_4 =10'b0;

   // m11_5 = W*in
   wire signed [9:0] m11_5;
   assign m11_5 =10'b0;

   // m11_6 = W*in
   wire signed [9:0] m11_6;
   assign m11_6 =10'b0;

   // m11_7 = W*in
   wire signed [9:0] m11_7;
   assign m11_7 =10'b0;

   // m11_8 = W*in
   wire signed [9:0] m11_8;
   assign m11_8 =10'b0;

   // m11_9 = W*in
   wire signed [9:0] m11_9;
   assign m11_9 =10'b0;

   // m11_10 = W*in
   wire signed [9:0] m11_10;
   assign m11_10 =10'b0;

   // m11_11 = W*in
   wire signed [9:0] m11_11;
   assign m11_11 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_12 = W*in
   wire signed [9:0] m11_12;
   assign m11_12 =10'b0;

   // m11_13 = W*in
   wire signed [9:0] m11_13;
   assign m11_13 =10'b0;

   // m11_14 = W*in
   wire signed [9:0] m11_14;
   assign m11_14 =10'b0;

   // m11_15 = W*in
   wire signed [9:0] m11_15;
   assign m11_15 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_16 = W*in
   wire signed [9:0] m11_16;
   assign m11_16 =10'b0;

   // m11_17 = W*in
   wire signed [9:0] m11_17;
   assign m11_17 ={ {2{in11[5]}} , in11 , {2{1'b0}} };

   // m11_18 = W*in
   wire signed [9:0] m11_18;
   assign m11_18 =10'b0;

   // m11_19 = W*in
   wire signed [9:0] m11_19;
   assign m11_19 =10'b0;

   // m11_20 = W*in
   wire signed [9:0] m11_20;
   assign m11_20 =10'b0;

   // m11_21 = W*in
   wire signed [9:0] m11_21;
   assign m11_21 =10'b0;

   // m11_22 = W*in
   wire signed [9:0] m11_22;
   assign m11_22 =10'b0;

   // m11_23 = W*in
   wire signed [9:0] m11_23;
   assign m11_23 =10'b0;

   // m11_24 = W*in
   wire signed [9:0] m11_24;
   assign m11_24 =10'b0;

   // m11_25 = W*in
   wire signed [9:0] m11_25;
   assign m11_25 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_26 = W*in
   wire signed [9:0] m11_26;
   assign m11_26 =10'b0;

   // m11_27 = W*in
   wire signed [9:0] m11_27;
   assign m11_27 =10'b0;

   // m11_28 = W*in
   wire signed [9:0] m11_28;
   assign m11_28 =10'b0;

   // m11_29 = W*in
   wire signed [9:0] m11_29;
   assign m11_29 =10'b0;

   // m11_30 = W*in
   wire signed [9:0] m11_30;
   assign m11_30 =10'b0;

   // m11_31 = W*in
   wire signed [9:0] m11_31;
   assign m11_31 =10'b0;

   // m11_32 = W*in
   wire signed [9:0] m11_32;
   assign m11_32 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_33 = W*in
   wire signed [9:0] m11_33;
   assign m11_33 =10'b0;

   // m11_34 = W*in
   wire signed [9:0] m11_34;
   assign m11_34 =10'b0;

   // m11_35 = W*in
   wire signed [9:0] m11_35;
   assign m11_35 =10'b0;

   // m11_36 = W*in
   wire signed [9:0] m11_36;
   assign m11_36 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_37 = W*in
   wire signed [9:0] m11_37;
   assign m11_37 =10'b0;

   // m11_38 = W*in
   wire signed [9:0] m11_38;
   assign m11_38 =10'b0;

   // m11_39 = W*in
   wire signed [9:0] m11_39;
   assign m11_39 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_40 = W*in
   wire signed [9:0] m11_40;
   assign m11_40 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_41 = W*in
   wire signed [9:0] m11_41;
   assign m11_41 =10'b0;

   // m11_42 = W*in
   wire signed [9:0] m11_42;
   assign m11_42 =10'b0;

   // m11_43 = W*in
   wire signed [9:0] m11_43;
   assign m11_43 =10'b0;

   // m11_44 = W*in
   wire signed [9:0] m11_44;
   assign m11_44 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_45 = W*in
   wire signed [9:0] m11_45;
   assign m11_45 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_46 = W*in
   wire signed [9:0] m11_46;
   assign m11_46 =10'b0;

   // m11_47 = W*in
   wire signed [9:0] m11_47;
   assign m11_47 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_48 = W*in
   wire signed [9:0] m11_48;
   assign m11_48 =10'b0;

   // m11_49 = W*in
   wire signed [9:0] m11_49;
   assign m11_49 =10'b0;

   // m11_50 = W*in
   wire signed [9:0] m11_50;
   assign m11_50 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_51 = W*in
   wire signed [9:0] m11_51;
   assign m11_51 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_52 = W*in
   wire signed [9:0] m11_52;
   assign m11_52 =10'b0;

   // m11_53 = W*in
   wire signed [9:0] m11_53;
   assign m11_53 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_54 = W*in
   wire signed [9:0] m11_54;
   assign m11_54 ={ {2{in11[5]}} , in11 , {2{1'b0}} };

   // m11_55 = W*in
   wire signed [9:0] m11_55;
   assign m11_55 =10'b0;

   // m11_56 = W*in
   wire signed [9:0] m11_56;
   assign m11_56 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_57 = W*in
   wire signed [9:0] m11_57;
   assign m11_57 ={ {2{in11[5]}} , in11 , {2{1'b0}} };

   // m11_58 = W*in
   wire signed [9:0] m11_58;
   assign m11_58 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_59 = W*in
   wire signed [9:0] m11_59;
   assign m11_59 =10'b0;

   // m11_60 = W*in
   wire signed [9:0] m11_60;
   assign m11_60 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_61 = W*in
   wire signed [9:0] m11_61;
   assign m11_61 =10'b0;

   // m11_62 = W*in
   wire signed [9:0] m11_62;
   assign m11_62 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_63 = W*in
   wire signed [9:0] m11_63;
   assign m11_63 =10'b0;

   // m11_64 = W*in
   wire signed [9:0] m11_64;
   assign m11_64 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_65 = W*in
   wire signed [9:0] m11_65;
   assign m11_65 =10'b0;

   // m11_66 = W*in
   wire signed [9:0] m11_66;
   assign m11_66 =10'b0;

   // m11_67 = W*in
   wire signed [9:0] m11_67;
   assign m11_67 =10'b0;

   // m11_68 = W*in
   wire signed [9:0] m11_68;
   assign m11_68 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_69 = W*in
   wire signed [9:0] m11_69;
   assign m11_69 ={ {3{in11[5]}} , in11 , {1{1'b0}} };

   // m11_70 = W*in
   wire signed [9:0] m11_70;
   assign m11_70 =10'b0;

   // m11_71 = W*in
   wire signed [9:0] m11_71;
   assign m11_71 =10'b0;

   // m11_72 = W*in
   wire signed [9:0] m11_72;
   assign m11_72 =10'b0;

   // m11_73 = W*in
   wire signed [9:0] m11_73;
   assign m11_73 =10'b0;

   // m11_74 = W*in
   wire signed [9:0] m11_74;
   assign m11_74 =10'b0;

   // m11_75 = W*in
   wire signed [9:0] m11_75;
   assign m11_75 =10'b0;

   // m11_76 = W*in
   wire signed [9:0] m11_76;
   assign m11_76 =10'b0;

   // m11_77 = W*in
   wire signed [9:0] m11_77;
   assign m11_77 =10'b0;

   // m11_78 = W*in
   wire signed [9:0] m11_78;
   assign m11_78 ={ {3{neg11[5]}} , neg11 , {1{1'b0}} };

   // m11_79 = W*in
   wire signed [9:0] m11_79;
   assign m11_79 =10'b0;

   // m11_80 = W*in
   wire signed [9:0] m11_80;
   assign m11_80 =10'b0;

   // m11_81 = W*in
   wire signed [9:0] m11_81;
   assign m11_81 =10'b0;

   // m12_1 = W*in
   wire signed [9:0] m12_1;
   assign m12_1 =10'b0;

   // m12_2 = W*in
   wire signed [9:0] m12_2;
   assign m12_2 =10'b0;

   // m12_3 = W*in
   wire signed [9:0] m12_3;
   assign m12_3 =10'b0;

   // m12_4 = W*in
   wire signed [9:0] m12_4;
   assign m12_4 =10'b0;

   // m12_5 = W*in
   wire signed [9:0] m12_5;
   assign m12_5 =10'b0;

   // m12_6 = W*in
   wire signed [9:0] m12_6;
   assign m12_6 =10'b0;

   // m12_7 = W*in
   wire signed [9:0] m12_7;
   assign m12_7 =10'b0;

   // m12_8 = W*in
   wire signed [9:0] m12_8;
   assign m12_8 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_9 = W*in
   wire signed [9:0] m12_9;
   assign m12_9 =10'b0;

   // m12_10 = W*in
   wire signed [9:0] m12_10;
   assign m12_10 =10'b0;

   // m12_11 = W*in
   wire signed [9:0] m12_11;
   assign m12_11 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_12 = W*in
   wire signed [9:0] m12_12;
   assign m12_12 =10'b0;

   // m12_13 = W*in
   wire signed [9:0] m12_13;
   assign m12_13 =10'b0;

   // m12_14 = W*in
   wire signed [9:0] m12_14;
   assign m12_14 =10'b0;

   // m12_15 = W*in
   wire signed [9:0] m12_15;
   assign m12_15 =10'b0;

   // m12_16 = W*in
   wire signed [9:0] m12_16;
   assign m12_16 =10'b0;

   // m12_17 = W*in
   wire signed [9:0] m12_17;
   assign m12_17 =10'b0;

   // m12_18 = W*in
   wire signed [9:0] m12_18;
   assign m12_18 =10'b0;

   // m12_19 = W*in
   wire signed [9:0] m12_19;
   assign m12_19 =10'b0;

   // m12_20 = W*in
   wire signed [9:0] m12_20;
   assign m12_20 =10'b0;

   // m12_21 = W*in
   wire signed [9:0] m12_21;
   assign m12_21 =10'b0;

   // m12_22 = W*in
   wire signed [9:0] m12_22;
   assign m12_22 =10'b0;

   // m12_23 = W*in
   wire signed [9:0] m12_23;
   assign m12_23 ={ {3{neg12[5]}} , neg12 , {1{1'b0}} };

   // m12_24 = W*in
   wire signed [9:0] m12_24;
   assign m12_24 =10'b0;

   // m12_25 = W*in
   wire signed [9:0] m12_25;
   assign m12_25 =10'b0;

   // m12_26 = W*in
   wire signed [9:0] m12_26;
   assign m12_26 =10'b0;

   // m12_27 = W*in
   wire signed [9:0] m12_27;
   assign m12_27 =10'b0;

   // m12_28 = W*in
   wire signed [9:0] m12_28;
   assign m12_28 =10'b0;

   // m12_29 = W*in
   wire signed [9:0] m12_29;
   assign m12_29 =10'b0;

   // m12_30 = W*in
   wire signed [9:0] m12_30;
   assign m12_30 =10'b0;

   // m12_31 = W*in
   wire signed [9:0] m12_31;
   assign m12_31 =10'b0;

   // m12_32 = W*in
   wire signed [9:0] m12_32;
   assign m12_32 =10'b0;

   // m12_33 = W*in
   wire signed [9:0] m12_33;
   assign m12_33 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_34 = W*in
   wire signed [9:0] m12_34;
   assign m12_34 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_35 = W*in
   wire signed [9:0] m12_35;
   assign m12_35 ={ {3{neg12[5]}} , neg12 , {1{1'b0}} };

   // m12_36 = W*in
   wire signed [9:0] m12_36;
   assign m12_36 =10'b0;

   // m12_37 = W*in
   wire signed [9:0] m12_37;
   assign m12_37 ={ {2{in12[5]}} , in12 , {2{1'b0}} };

   // m12_38 = W*in
   wire signed [9:0] m12_38;
   assign m12_38 =10'b0;

   // m12_39 = W*in
   wire signed [9:0] m12_39;
   assign m12_39 =10'b0;

   // m12_40 = W*in
   wire signed [9:0] m12_40;
   assign m12_40 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_41 = W*in
   wire signed [9:0] m12_41;
   assign m12_41 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_42 = W*in
   wire signed [9:0] m12_42;
   assign m12_42 =10'b0;

   // m12_43 = W*in
   wire signed [9:0] m12_43;
   assign m12_43 =10'b0;

   // m12_44 = W*in
   wire signed [9:0] m12_44;
   assign m12_44 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_45 = W*in
   wire signed [9:0] m12_45;
   assign m12_45 =10'b0;

   // m12_46 = W*in
   wire signed [9:0] m12_46;
   assign m12_46 ={ {3{neg12[5]}} , neg12 , {1{1'b0}} };

   // m12_47 = W*in
   wire signed [9:0] m12_47;
   assign m12_47 =10'b0;

   // m12_48 = W*in
   wire signed [9:0] m12_48;
   assign m12_48 =10'b0;

   // m12_49 = W*in
   wire signed [9:0] m12_49;
   assign m12_49 =10'b0;

   // m12_50 = W*in
   wire signed [9:0] m12_50;
   assign m12_50 =10'b0;

   // m12_51 = W*in
   wire signed [9:0] m12_51;
   assign m12_51 ={ {2{in12[5]}} , in12 , {2{1'b0}} };

   // m12_52 = W*in
   wire signed [9:0] m12_52;
   assign m12_52 =10'b0;

   // m12_53 = W*in
   wire signed [9:0] m12_53;
   assign m12_53 =10'b0;

   // m12_54 = W*in
   wire signed [9:0] m12_54;
   assign m12_54 =10'b0;

   // m12_55 = W*in
   wire signed [9:0] m12_55;
   assign m12_55 =10'b0;

   // m12_56 = W*in
   wire signed [9:0] m12_56;
   assign m12_56 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_57 = W*in
   wire signed [9:0] m12_57;
   assign m12_57 =10'b0;

   // m12_58 = W*in
   wire signed [9:0] m12_58;
   assign m12_58 ={ {2{in12[5]}} , in12 , {2{1'b0}} };

   // m12_59 = W*in
   wire signed [9:0] m12_59;
   assign m12_59 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_60 = W*in
   wire signed [9:0] m12_60;
   assign m12_60 ={ {2{in12[5]}} , in12 , {2{1'b0}} };

   // m12_61 = W*in
   wire signed [9:0] m12_61;
   assign m12_61 =10'b0;

   // m12_62 = W*in
   wire signed [9:0] m12_62;
   assign m12_62 =10'b0;

   // m12_63 = W*in
   wire signed [9:0] m12_63;
   assign m12_63 =10'b0;

   // m12_64 = W*in
   wire signed [9:0] m12_64;
   assign m12_64 =10'b0;

   // m12_65 = W*in
   wire signed [9:0] m12_65;
   assign m12_65 =10'b0;

   // m12_66 = W*in
   wire signed [9:0] m12_66;
   assign m12_66 =10'b0;

   // m12_67 = W*in
   wire signed [9:0] m12_67;
   assign m12_67 =10'b0;

   // m12_68 = W*in
   wire signed [9:0] m12_68;
   assign m12_68 =10'b0;

   // m12_69 = W*in
   wire signed [9:0] m12_69;
   assign m12_69 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_70 = W*in
   wire signed [9:0] m12_70;
   assign m12_70 =10'b0;

   // m12_71 = W*in
   wire signed [9:0] m12_71;
   assign m12_71 ={ {3{neg12[5]}} , neg12 , {1{1'b0}} };

   // m12_72 = W*in
   wire signed [9:0] m12_72;
   assign m12_72 =10'b0;

   // m12_73 = W*in
   wire signed [9:0] m12_73;
   assign m12_73 =10'b0;

   // m12_74 = W*in
   wire signed [9:0] m12_74;
   assign m12_74 =10'b0;

   // m12_75 = W*in
   wire signed [9:0] m12_75;
   assign m12_75 =10'b0;

   // m12_76 = W*in
   wire signed [9:0] m12_76;
   assign m12_76 =10'b0;

   // m12_77 = W*in
   wire signed [9:0] m12_77;
   assign m12_77 =10'b0;

   // m12_78 = W*in
   wire signed [9:0] m12_78;
   assign m12_78 =10'b0;

   // m12_79 = W*in
   wire signed [9:0] m12_79;
   assign m12_79 =10'b0;

   // m12_80 = W*in
   wire signed [9:0] m12_80;
   assign m12_80 =10'b0;

   // m12_81 = W*in
   wire signed [9:0] m12_81;
   assign m12_81 =10'b0;

   // m13_1 = W*in
   wire signed [9:0] m13_1;
   assign m13_1 =10'b0;

   // m13_2 = W*in
   wire signed [9:0] m13_2;
   assign m13_2 =10'b0;

   // m13_3 = W*in
   wire signed [9:0] m13_3;
   assign m13_3 ={ {2{in13[5]}} , in13 , {2{1'b0}} };

   // m13_4 = W*in
   wire signed [9:0] m13_4;
   assign m13_4 =10'b0;

   // m13_5 = W*in
   wire signed [9:0] m13_5;
   assign m13_5 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_6 = W*in
   wire signed [9:0] m13_6;
   assign m13_6 =10'b0;

   // m13_7 = W*in
   wire signed [9:0] m13_7;
   assign m13_7 =10'b0;

   // m13_8 = W*in
   wire signed [9:0] m13_8;
   assign m13_8 =10'b0;

   // m13_9 = W*in
   wire signed [9:0] m13_9;
   assign m13_9 =10'b0;

   // m13_10 = W*in
   wire signed [9:0] m13_10;
   assign m13_10 =10'b0;

   // m13_11 = W*in
   wire signed [9:0] m13_11;
   assign m13_11 =10'b0;

   // m13_12 = W*in
   wire signed [9:0] m13_12;
   assign m13_12 =10'b0;

   // m13_13 = W*in
   wire signed [9:0] m13_13;
   assign m13_13 =10'b0;

   // m13_14 = W*in
   wire signed [9:0] m13_14;
   assign m13_14 =10'b0;

   // m13_15 = W*in
   wire signed [9:0] m13_15;
   assign m13_15 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_16 = W*in
   wire signed [9:0] m13_16;
   assign m13_16 =10'b0;

   // m13_17 = W*in
   wire signed [9:0] m13_17;
   assign m13_17 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_18 = W*in
   wire signed [9:0] m13_18;
   assign m13_18 =10'b0;

   // m13_19 = W*in
   wire signed [9:0] m13_19;
   assign m13_19 =10'b0;

   // m13_20 = W*in
   wire signed [9:0] m13_20;
   assign m13_20 =10'b0;

   // m13_21 = W*in
   wire signed [9:0] m13_21;
   assign m13_21 =10'b0;

   // m13_22 = W*in
   wire signed [9:0] m13_22;
   assign m13_22 =10'b0;

   // m13_23 = W*in
   wire signed [9:0] m13_23;
   assign m13_23 =10'b0;

   // m13_24 = W*in
   wire signed [9:0] m13_24;
   assign m13_24 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_25 = W*in
   wire signed [9:0] m13_25;
   assign m13_25 =10'b0;

   // m13_26 = W*in
   wire signed [9:0] m13_26;
   assign m13_26 =10'b0;

   // m13_27 = W*in
   wire signed [9:0] m13_27;
   assign m13_27 =10'b0;

   // m13_28 = W*in
   wire signed [9:0] m13_28;
   assign m13_28 =10'b0;

   // m13_29 = W*in
   wire signed [9:0] m13_29;
   assign m13_29 =10'b0;

   // m13_30 = W*in
   wire signed [9:0] m13_30;
   assign m13_30 =10'b0;

   // m13_31 = W*in
   wire signed [9:0] m13_31;
   assign m13_31 =10'b0;

   // m13_32 = W*in
   wire signed [9:0] m13_32;
   assign m13_32 =10'b0;

   // m13_33 = W*in
   wire signed [9:0] m13_33;
   assign m13_33 =10'b0;

   // m13_34 = W*in
   wire signed [9:0] m13_34;
   assign m13_34 =10'b0;

   // m13_35 = W*in
   wire signed [9:0] m13_35;
   assign m13_35 =10'b0;

   // m13_36 = W*in
   wire signed [9:0] m13_36;
   assign m13_36 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_37 = W*in
   wire signed [9:0] m13_37;
   assign m13_37 =10'b0;

   // m13_38 = W*in
   wire signed [9:0] m13_38;
   assign m13_38 =10'b0;

   // m13_39 = W*in
   wire signed [9:0] m13_39;
   assign m13_39 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_40 = W*in
   wire signed [9:0] m13_40;
   assign m13_40 =10'b0;

   // m13_41 = W*in
   wire signed [9:0] m13_41;
   assign m13_41 =10'b0;

   // m13_42 = W*in
   wire signed [9:0] m13_42;
   assign m13_42 =10'b0;

   // m13_43 = W*in
   wire signed [9:0] m13_43;
   assign m13_43 =10'b0;

   // m13_44 = W*in
   wire signed [9:0] m13_44;
   assign m13_44 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_45 = W*in
   wire signed [9:0] m13_45;
   assign m13_45 =10'b0;

   // m13_46 = W*in
   wire signed [9:0] m13_46;
   assign m13_46 =10'b0;

   // m13_47 = W*in
   wire signed [9:0] m13_47;
   assign m13_47 =10'b0;

   // m13_48 = W*in
   wire signed [9:0] m13_48;
   assign m13_48 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_49 = W*in
   wire signed [9:0] m13_49;
   assign m13_49 =10'b0;

   // m13_50 = W*in
   wire signed [9:0] m13_50;
   assign m13_50 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_51 = W*in
   wire signed [9:0] m13_51;
   assign m13_51 =10'b0;

   // m13_52 = W*in
   wire signed [9:0] m13_52;
   assign m13_52 =10'b0;

   // m13_53 = W*in
   wire signed [9:0] m13_53;
   assign m13_53 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_54 = W*in
   wire signed [9:0] m13_54;
   assign m13_54 =10'b0;

   // m13_55 = W*in
   wire signed [9:0] m13_55;
   assign m13_55 =10'b0;

   // m13_56 = W*in
   wire signed [9:0] m13_56;
   assign m13_56 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_57 = W*in
   wire signed [9:0] m13_57;
   assign m13_57 =10'b0;

   // m13_58 = W*in
   wire signed [9:0] m13_58;
   assign m13_58 =10'b0;

   // m13_59 = W*in
   wire signed [9:0] m13_59;
   assign m13_59 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_60 = W*in
   wire signed [9:0] m13_60;
   assign m13_60 =10'b0;

   // m13_61 = W*in
   wire signed [9:0] m13_61;
   assign m13_61 =10'b0;

   // m13_62 = W*in
   wire signed [9:0] m13_62;
   assign m13_62 =10'b0;

   // m13_63 = W*in
   wire signed [9:0] m13_63;
   assign m13_63 =10'b0;

   // m13_64 = W*in
   wire signed [9:0] m13_64;
   assign m13_64 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_65 = W*in
   wire signed [9:0] m13_65;
   assign m13_65 =10'b0;

   // m13_66 = W*in
   wire signed [9:0] m13_66;
   assign m13_66 =10'b0;

   // m13_67 = W*in
   wire signed [9:0] m13_67;
   assign m13_67 =10'b0;

   // m13_68 = W*in
   wire signed [9:0] m13_68;
   assign m13_68 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_69 = W*in
   wire signed [9:0] m13_69;
   assign m13_69 =10'b0;

   // m13_70 = W*in
   wire signed [9:0] m13_70;
   assign m13_70 =10'b0;

   // m13_71 = W*in
   wire signed [9:0] m13_71;
   assign m13_71 =10'b0;

   // m13_72 = W*in
   wire signed [9:0] m13_72;
   assign m13_72 =10'b0;

   // m13_73 = W*in
   wire signed [9:0] m13_73;
   assign m13_73 =10'b0;

   // m13_74 = W*in
   wire signed [9:0] m13_74;
   assign m13_74 =10'b0;

   // m13_75 = W*in
   wire signed [9:0] m13_75;
   assign m13_75 =10'b0;

   // m13_76 = W*in
   wire signed [9:0] m13_76;
   assign m13_76 =10'b0;

   // m13_77 = W*in
   wire signed [9:0] m13_77;
   assign m13_77 =10'b0;

   // m13_78 = W*in
   wire signed [9:0] m13_78;
   assign m13_78 ={ {3{in13[5]}} , in13 , {1{1'b0}} };

   // m13_79 = W*in
   wire signed [9:0] m13_79;
   assign m13_79 =10'b0;

   // m13_80 = W*in
   wire signed [9:0] m13_80;
   assign m13_80 =10'b0;

   // m13_81 = W*in
   wire signed [9:0] m13_81;
   assign m13_81 =10'b0;

   // m14_1 = W*in
   wire signed [9:0] m14_1;
   assign m14_1 =10'b0;

   // m14_2 = W*in
   wire signed [9:0] m14_2;
   assign m14_2 ={ {2{in14[5]}} , in14 , {2{1'b0}} };

   // m14_3 = W*in
   wire signed [9:0] m14_3;
   assign m14_3 =10'b0;

   // m14_4 = W*in
   wire signed [9:0] m14_4;
   assign m14_4 =10'b0;

   // m14_5 = W*in
   wire signed [9:0] m14_5;
   assign m14_5 =10'b0;

   // m14_6 = W*in
   wire signed [9:0] m14_6;
   assign m14_6 =10'b0;

   // m14_7 = W*in
   wire signed [9:0] m14_7;
   assign m14_7 =10'b0;

   // m14_8 = W*in
   wire signed [9:0] m14_8;
   assign m14_8 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_9 = W*in
   wire signed [9:0] m14_9;
   assign m14_9 =10'b0;

   // m14_10 = W*in
   wire signed [9:0] m14_10;
   assign m14_10 =10'b0;

   // m14_11 = W*in
   wire signed [9:0] m14_11;
   assign m14_11 =10'b0;

   // m14_12 = W*in
   wire signed [9:0] m14_12;
   assign m14_12 =10'b0;

   // m14_13 = W*in
   wire signed [9:0] m14_13;
   assign m14_13 =10'b0;

   // m14_14 = W*in
   wire signed [9:0] m14_14;
   assign m14_14 =10'b0;

   // m14_15 = W*in
   wire signed [9:0] m14_15;
   assign m14_15 =10'b0;

   // m14_16 = W*in
   wire signed [9:0] m14_16;
   assign m14_16 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_17 = W*in
   wire signed [9:0] m14_17;
   assign m14_17 =10'b0;

   // m14_18 = W*in
   wire signed [9:0] m14_18;
   assign m14_18 =10'b0;

   // m14_19 = W*in
   wire signed [9:0] m14_19;
   assign m14_19 =10'b0;

   // m14_20 = W*in
   wire signed [9:0] m14_20;
   assign m14_20 =10'b0;

   // m14_21 = W*in
   wire signed [9:0] m14_21;
   assign m14_21 =10'b0;

   // m14_22 = W*in
   wire signed [9:0] m14_22;
   assign m14_22 =10'b0;

   // m14_23 = W*in
   wire signed [9:0] m14_23;
   assign m14_23 =10'b0;

   // m14_24 = W*in
   wire signed [9:0] m14_24;
   assign m14_24 =10'b0;

   // m14_25 = W*in
   wire signed [9:0] m14_25;
   assign m14_25 =10'b0;

   // m14_26 = W*in
   wire signed [9:0] m14_26;
   assign m14_26 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_27 = W*in
   wire signed [9:0] m14_27;
   assign m14_27 =10'b0;

   // m14_28 = W*in
   wire signed [9:0] m14_28;
   assign m14_28 =10'b0;

   // m14_29 = W*in
   wire signed [9:0] m14_29;
   assign m14_29 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_30 = W*in
   wire signed [9:0] m14_30;
   assign m14_30 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_31 = W*in
   wire signed [9:0] m14_31;
   assign m14_31 =10'b0;

   // m14_32 = W*in
   wire signed [9:0] m14_32;
   assign m14_32 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_33 = W*in
   wire signed [9:0] m14_33;
   assign m14_33 =10'b0;

   // m14_34 = W*in
   wire signed [9:0] m14_34;
   assign m14_34 =10'b0;

   // m14_35 = W*in
   wire signed [9:0] m14_35;
   assign m14_35 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_36 = W*in
   wire signed [9:0] m14_36;
   assign m14_36 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_37 = W*in
   wire signed [9:0] m14_37;
   assign m14_37 =10'b0;

   // m14_38 = W*in
   wire signed [9:0] m14_38;
   assign m14_38 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_39 = W*in
   wire signed [9:0] m14_39;
   assign m14_39 =10'b0;

   // m14_40 = W*in
   wire signed [9:0] m14_40;
   assign m14_40 =10'b0;

   // m14_41 = W*in
   wire signed [9:0] m14_41;
   assign m14_41 =10'b0;

   // m14_42 = W*in
   wire signed [9:0] m14_42;
   assign m14_42 =10'b0;

   // m14_43 = W*in
   wire signed [9:0] m14_43;
   assign m14_43 =10'b0;

   // m14_44 = W*in
   wire signed [9:0] m14_44;
   assign m14_44 =10'b0;

   // m14_45 = W*in
   wire signed [9:0] m14_45;
   assign m14_45 =10'b0;

   // m14_46 = W*in
   wire signed [9:0] m14_46;
   assign m14_46 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_47 = W*in
   wire signed [9:0] m14_47;
   assign m14_47 =10'b0;

   // m14_48 = W*in
   wire signed [9:0] m14_48;
   assign m14_48 =10'b0;

   // m14_49 = W*in
   wire signed [9:0] m14_49;
   assign m14_49 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_50 = W*in
   wire signed [9:0] m14_50;
   assign m14_50 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_51 = W*in
   wire signed [9:0] m14_51;
   assign m14_51 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_52 = W*in
   wire signed [9:0] m14_52;
   assign m14_52 =10'b0;

   // m14_53 = W*in
   wire signed [9:0] m14_53;
   assign m14_53 =10'b0;

   // m14_54 = W*in
   wire signed [9:0] m14_54;
   assign m14_54 =10'b0;

   // m14_55 = W*in
   wire signed [9:0] m14_55;
   assign m14_55 =10'b0;

   // m14_56 = W*in
   wire signed [9:0] m14_56;
   assign m14_56 =10'b0;

   // m14_57 = W*in
   wire signed [9:0] m14_57;
   assign m14_57 =10'b0;

   // m14_58 = W*in
   wire signed [9:0] m14_58;
   assign m14_58 =10'b0;

   // m14_59 = W*in
   wire signed [9:0] m14_59;
   assign m14_59 =10'b0;

   // m14_60 = W*in
   wire signed [9:0] m14_60;
   assign m14_60 =10'b0;

   // m14_61 = W*in
   wire signed [9:0] m14_61;
   assign m14_61 =10'b0;

   // m14_62 = W*in
   wire signed [9:0] m14_62;
   assign m14_62 =10'b0;

   // m14_63 = W*in
   wire signed [9:0] m14_63;
   assign m14_63 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_64 = W*in
   wire signed [9:0] m14_64;
   assign m14_64 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_65 = W*in
   wire signed [9:0] m14_65;
   assign m14_65 =10'b0;

   // m14_66 = W*in
   wire signed [9:0] m14_66;
   assign m14_66 =10'b0;

   // m14_67 = W*in
   wire signed [9:0] m14_67;
   assign m14_67 =10'b0;

   // m14_68 = W*in
   wire signed [9:0] m14_68;
   assign m14_68 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_69 = W*in
   wire signed [9:0] m14_69;
   assign m14_69 =10'b0;

   // m14_70 = W*in
   wire signed [9:0] m14_70;
   assign m14_70 =10'b0;

   // m14_71 = W*in
   wire signed [9:0] m14_71;
   assign m14_71 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_72 = W*in
   wire signed [9:0] m14_72;
   assign m14_72 =10'b0;

   // m14_73 = W*in
   wire signed [9:0] m14_73;
   assign m14_73 ={ {2{in14[5]}} , in14 , {2{1'b0}} };

   // m14_74 = W*in
   wire signed [9:0] m14_74;
   assign m14_74 =10'b0;

   // m14_75 = W*in
   wire signed [9:0] m14_75;
   assign m14_75 =10'b0;

   // m14_76 = W*in
   wire signed [9:0] m14_76;
   assign m14_76 =10'b0;

   // m14_77 = W*in
   wire signed [9:0] m14_77;
   assign m14_77 =10'b0;

   // m14_78 = W*in
   wire signed [9:0] m14_78;
   assign m14_78 =10'b0;

   // m14_79 = W*in
   wire signed [9:0] m14_79;
   assign m14_79 =10'b0;

   // m14_80 = W*in
   wire signed [9:0] m14_80;
   assign m14_80 =10'b0;

   // m14_81 = W*in
   wire signed [9:0] m14_81;
   assign m14_81 =10'b0;

   // m15_1 = W*in
   wire signed [9:0] m15_1;
   assign m15_1 =10'b0;

   // m15_2 = W*in
   wire signed [9:0] m15_2;
   assign m15_2 =10'b0;

   // m15_3 = W*in
   wire signed [9:0] m15_3;
   assign m15_3 =10'b0;

   // m15_4 = W*in
   wire signed [9:0] m15_4;
   assign m15_4 =10'b0;

   // m15_5 = W*in
   wire signed [9:0] m15_5;
   assign m15_5 =10'b0;

   // m15_6 = W*in
   wire signed [9:0] m15_6;
   assign m15_6 =10'b0;

   // m15_7 = W*in
   wire signed [9:0] m15_7;
   assign m15_7 =10'b0;

   // m15_8 = W*in
   wire signed [9:0] m15_8;
   assign m15_8 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_9 = W*in
   wire signed [9:0] m15_9;
   assign m15_9 =10'b0;

   // m15_10 = W*in
   wire signed [9:0] m15_10;
   assign m15_10 =10'b0;

   // m15_11 = W*in
   wire signed [9:0] m15_11;
   assign m15_11 =10'b0;

   // m15_12 = W*in
   wire signed [9:0] m15_12;
   assign m15_12 =10'b0;

   // m15_13 = W*in
   wire signed [9:0] m15_13;
   assign m15_13 =10'b0;

   // m15_14 = W*in
   wire signed [9:0] m15_14;
   assign m15_14 =10'b0;

   // m15_15 = W*in
   wire signed [9:0] m15_15;
   assign m15_15 =10'b0;

   // m15_16 = W*in
   wire signed [9:0] m15_16;
   assign m15_16 =10'b0;

   // m15_17 = W*in
   wire signed [9:0] m15_17;
   assign m15_17 =10'b0;

   // m15_18 = W*in
   wire signed [9:0] m15_18;
   assign m15_18 =10'b0;

   // m15_19 = W*in
   wire signed [9:0] m15_19;
   assign m15_19 =10'b0;

   // m15_20 = W*in
   wire signed [9:0] m15_20;
   assign m15_20 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_21 = W*in
   wire signed [9:0] m15_21;
   assign m15_21 =10'b0;

   // m15_22 = W*in
   wire signed [9:0] m15_22;
   assign m15_22 =10'b0;

   // m15_23 = W*in
   wire signed [9:0] m15_23;
   assign m15_23 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_24 = W*in
   wire signed [9:0] m15_24;
   assign m15_24 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_25 = W*in
   wire signed [9:0] m15_25;
   assign m15_25 =10'b0;

   // m15_26 = W*in
   wire signed [9:0] m15_26;
   assign m15_26 =10'b0;

   // m15_27 = W*in
   wire signed [9:0] m15_27;
   assign m15_27 =10'b0;

   // m15_28 = W*in
   wire signed [9:0] m15_28;
   assign m15_28 =10'b0;

   // m15_29 = W*in
   wire signed [9:0] m15_29;
   assign m15_29 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_30 = W*in
   wire signed [9:0] m15_30;
   assign m15_30 =10'b0;

   // m15_31 = W*in
   wire signed [9:0] m15_31;
   assign m15_31 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_32 = W*in
   wire signed [9:0] m15_32;
   assign m15_32 =10'b0;

   // m15_33 = W*in
   wire signed [9:0] m15_33;
   assign m15_33 =10'b0;

   // m15_34 = W*in
   wire signed [9:0] m15_34;
   assign m15_34 =10'b0;

   // m15_35 = W*in
   wire signed [9:0] m15_35;
   assign m15_35 =10'b0;

   // m15_36 = W*in
   wire signed [9:0] m15_36;
   assign m15_36 =10'b0;

   // m15_37 = W*in
   wire signed [9:0] m15_37;
   assign m15_37 =10'b0;

   // m15_38 = W*in
   wire signed [9:0] m15_38;
   assign m15_38 =10'b0;

   // m15_39 = W*in
   wire signed [9:0] m15_39;
   assign m15_39 =10'b0;

   // m15_40 = W*in
   wire signed [9:0] m15_40;
   assign m15_40 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_41 = W*in
   wire signed [9:0] m15_41;
   assign m15_41 =10'b0;

   // m15_42 = W*in
   wire signed [9:0] m15_42;
   assign m15_42 =10'b0;

   // m15_43 = W*in
   wire signed [9:0] m15_43;
   assign m15_43 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_44 = W*in
   wire signed [9:0] m15_44;
   assign m15_44 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_45 = W*in
   wire signed [9:0] m15_45;
   assign m15_45 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_46 = W*in
   wire signed [9:0] m15_46;
   assign m15_46 =10'b0;

   // m15_47 = W*in
   wire signed [9:0] m15_47;
   assign m15_47 =10'b0;

   // m15_48 = W*in
   wire signed [9:0] m15_48;
   assign m15_48 ={ {2{in15[5]}} , in15 , {2{1'b0}} };

   // m15_49 = W*in
   wire signed [9:0] m15_49;
   assign m15_49 =10'b0;

   // m15_50 = W*in
   wire signed [9:0] m15_50;
   assign m15_50 =10'b0;

   // m15_51 = W*in
   wire signed [9:0] m15_51;
   assign m15_51 =10'b0;

   // m15_52 = W*in
   wire signed [9:0] m15_52;
   assign m15_52 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_53 = W*in
   wire signed [9:0] m15_53;
   assign m15_53 =10'b0;

   // m15_54 = W*in
   wire signed [9:0] m15_54;
   assign m15_54 =10'b0;

   // m15_55 = W*in
   wire signed [9:0] m15_55;
   assign m15_55 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_56 = W*in
   wire signed [9:0] m15_56;
   assign m15_56 =10'b0;

   // m15_57 = W*in
   wire signed [9:0] m15_57;
   assign m15_57 =10'b0;

   // m15_58 = W*in
   wire signed [9:0] m15_58;
   assign m15_58 =10'b0;

   // m15_59 = W*in
   wire signed [9:0] m15_59;
   assign m15_59 =10'b0;

   // m15_60 = W*in
   wire signed [9:0] m15_60;
   assign m15_60 =10'b0;

   // m15_61 = W*in
   wire signed [9:0] m15_61;
   assign m15_61 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_62 = W*in
   wire signed [9:0] m15_62;
   assign m15_62 =10'b0;

   // m15_63 = W*in
   wire signed [9:0] m15_63;
   assign m15_63 =10'b0;

   // m15_64 = W*in
   wire signed [9:0] m15_64;
   assign m15_64 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_65 = W*in
   wire signed [9:0] m15_65;
   assign m15_65 =10'b0;

   // m15_66 = W*in
   wire signed [9:0] m15_66;
   assign m15_66 =10'b0;

   // m15_67 = W*in
   wire signed [9:0] m15_67;
   assign m15_67 ={ {2{in15[5]}} , in15 , {2{1'b0}} };

   // m15_68 = W*in
   wire signed [9:0] m15_68;
   assign m15_68 =10'b0;

   // m15_69 = W*in
   wire signed [9:0] m15_69;
   assign m15_69 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_70 = W*in
   wire signed [9:0] m15_70;
   assign m15_70 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_71 = W*in
   wire signed [9:0] m15_71;
   assign m15_71 =10'b0;

   // m15_72 = W*in
   wire signed [9:0] m15_72;
   assign m15_72 =10'b0;

   // m15_73 = W*in
   wire signed [9:0] m15_73;
   assign m15_73 =10'b0;

   // m15_74 = W*in
   wire signed [9:0] m15_74;
   assign m15_74 =10'b0;

   // m15_75 = W*in
   wire signed [9:0] m15_75;
   assign m15_75 ={ {2{in15[5]}} , in15 , {2{1'b0}} };

   // m15_76 = W*in
   wire signed [9:0] m15_76;
   assign m15_76 =10'b0;

   // m15_77 = W*in
   wire signed [9:0] m15_77;
   assign m15_77 =10'b0;

   // m15_78 = W*in
   wire signed [9:0] m15_78;
   assign m15_78 =10'b0;

   // m15_79 = W*in
   wire signed [9:0] m15_79;
   assign m15_79 =10'b0;

   // m15_80 = W*in
   wire signed [9:0] m15_80;
   assign m15_80 =10'b0;

   // m15_81 = W*in
   wire signed [9:0] m15_81;
   assign m15_81 =10'b0;

   // m16_1 = W*in
   wire signed [9:0] m16_1;
   assign m16_1 =10'b0;

   // m16_2 = W*in
   wire signed [9:0] m16_2;
   assign m16_2 =10'b0;

   // m16_3 = W*in
   wire signed [9:0] m16_3;
   assign m16_3 =10'b0;

   // m16_4 = W*in
   wire signed [9:0] m16_4;
   assign m16_4 =10'b0;

   // m16_5 = W*in
   wire signed [9:0] m16_5;
   assign m16_5 =10'b0;

   // m16_6 = W*in
   wire signed [9:0] m16_6;
   assign m16_6 =10'b0;

   // m16_7 = W*in
   wire signed [9:0] m16_7;
   assign m16_7 =10'b0;

   // m16_8 = W*in
   wire signed [9:0] m16_8;
   assign m16_8 =10'b0;

   // m16_9 = W*in
   wire signed [9:0] m16_9;
   assign m16_9 ={ {2{in16[5]}} , in16 , {2{1'b0}} };

   // m16_10 = W*in
   wire signed [9:0] m16_10;
   assign m16_10 =10'b0;

   // m16_11 = W*in
   wire signed [9:0] m16_11;
   assign m16_11 =10'b0;

   // m16_12 = W*in
   wire signed [9:0] m16_12;
   assign m16_12 =10'b0;

   // m16_13 = W*in
   wire signed [9:0] m16_13;
   assign m16_13 =10'b0;

   // m16_14 = W*in
   wire signed [9:0] m16_14;
   assign m16_14 =10'b0;

   // m16_15 = W*in
   wire signed [9:0] m16_15;
   assign m16_15 ={ {2{in16[5]}} , in16 , {2{1'b0}} };

   // m16_16 = W*in
   wire signed [9:0] m16_16;
   assign m16_16 =10'b0;

   // m16_17 = W*in
   wire signed [9:0] m16_17;
   assign m16_17 =10'b0;

   // m16_18 = W*in
   wire signed [9:0] m16_18;
   assign m16_18 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_19 = W*in
   wire signed [9:0] m16_19;
   assign m16_19 =10'b0;

   // m16_20 = W*in
   wire signed [9:0] m16_20;
   assign m16_20 ={ {3{neg16[5]}} , neg16 , {1{1'b0}} };

   // m16_21 = W*in
   wire signed [9:0] m16_21;
   assign m16_21 =10'b0;

   // m16_22 = W*in
   wire signed [9:0] m16_22;
   assign m16_22 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_23 = W*in
   wire signed [9:0] m16_23;
   assign m16_23 =10'b0;

   // m16_24 = W*in
   wire signed [9:0] m16_24;
   assign m16_24 ={ {3{neg16[5]}} , neg16 , {1{1'b0}} };

   // m16_25 = W*in
   wire signed [9:0] m16_25;
   assign m16_25 =10'b0;

   // m16_26 = W*in
   wire signed [9:0] m16_26;
   assign m16_26 =10'b0;

   // m16_27 = W*in
   wire signed [9:0] m16_27;
   assign m16_27 =10'b0;

   // m16_28 = W*in
   wire signed [9:0] m16_28;
   assign m16_28 ={ {3{neg16[5]}} , neg16 , {1{1'b0}} };

   // m16_29 = W*in
   wire signed [9:0] m16_29;
   assign m16_29 ={ {3{neg16[5]}} , neg16 , {1{1'b0}} };

   // m16_30 = W*in
   wire signed [9:0] m16_30;
   assign m16_30 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_31 = W*in
   wire signed [9:0] m16_31;
   assign m16_31 =10'b0;

   // m16_32 = W*in
   wire signed [9:0] m16_32;
   assign m16_32 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_33 = W*in
   wire signed [9:0] m16_33;
   assign m16_33 =10'b0;

   // m16_34 = W*in
   wire signed [9:0] m16_34;
   assign m16_34 ={ {3{neg16[5]}} , neg16 , {1{1'b0}} };

   // m16_35 = W*in
   wire signed [9:0] m16_35;
   assign m16_35 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_36 = W*in
   wire signed [9:0] m16_36;
   assign m16_36 =10'b0;

   // m16_37 = W*in
   wire signed [9:0] m16_37;
   assign m16_37 ={ {3{neg16[5]}} , neg16 , {1{1'b0}} };

   // m16_38 = W*in
   wire signed [9:0] m16_38;
   assign m16_38 =10'b0;

   // m16_39 = W*in
   wire signed [9:0] m16_39;
   assign m16_39 =10'b0;

   // m16_40 = W*in
   wire signed [9:0] m16_40;
   assign m16_40 =10'b0;

   // m16_41 = W*in
   wire signed [9:0] m16_41;
   assign m16_41 =10'b0;

   // m16_42 = W*in
   wire signed [9:0] m16_42;
   assign m16_42 ={ {2{in16[5]}} , in16 , {2{1'b0}} };

   // m16_43 = W*in
   wire signed [9:0] m16_43;
   assign m16_43 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_44 = W*in
   wire signed [9:0] m16_44;
   assign m16_44 =10'b0;

   // m16_45 = W*in
   wire signed [9:0] m16_45;
   assign m16_45 ={ {2{neg16[5]}} , neg16 , {2{1'b0}} };

   // m16_46 = W*in
   wire signed [9:0] m16_46;
   assign m16_46 =10'b0;

   // m16_47 = W*in
   wire signed [9:0] m16_47;
   assign m16_47 =10'b0;

   // m16_48 = W*in
   wire signed [9:0] m16_48;
   assign m16_48 =10'b0;

   // m16_49 = W*in
   wire signed [9:0] m16_49;
   assign m16_49 =10'b0;

   // m16_50 = W*in
   wire signed [9:0] m16_50;
   assign m16_50 =10'b0;

   // m16_51 = W*in
   wire signed [9:0] m16_51;
   assign m16_51 =10'b0;

   // m16_52 = W*in
   wire signed [9:0] m16_52;
   assign m16_52 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_53 = W*in
   wire signed [9:0] m16_53;
   assign m16_53 =10'b0;

   // m16_54 = W*in
   wire signed [9:0] m16_54;
   assign m16_54 =10'b0;

   // m16_55 = W*in
   wire signed [9:0] m16_55;
   assign m16_55 =10'b0;

   // m16_56 = W*in
   wire signed [9:0] m16_56;
   assign m16_56 =10'b0;

   // m16_57 = W*in
   wire signed [9:0] m16_57;
   assign m16_57 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_58 = W*in
   wire signed [9:0] m16_58;
   assign m16_58 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_59 = W*in
   wire signed [9:0] m16_59;
   assign m16_59 =10'b0;

   // m16_60 = W*in
   wire signed [9:0] m16_60;
   assign m16_60 =10'b0;

   // m16_61 = W*in
   wire signed [9:0] m16_61;
   assign m16_61 =10'b0;

   // m16_62 = W*in
   wire signed [9:0] m16_62;
   assign m16_62 ={ {2{in16[5]}} , in16 , {2{1'b0}} };

   // m16_63 = W*in
   wire signed [9:0] m16_63;
   assign m16_63 =10'b0;

   // m16_64 = W*in
   wire signed [9:0] m16_64;
   assign m16_64 =10'b0;

   // m16_65 = W*in
   wire signed [9:0] m16_65;
   assign m16_65 =10'b0;

   // m16_66 = W*in
   wire signed [9:0] m16_66;
   assign m16_66 ={ {2{in16[5]}} , in16 , {2{1'b0}} };

   // m16_67 = W*in
   wire signed [9:0] m16_67;
   assign m16_67 =10'b0;

   // m16_68 = W*in
   wire signed [9:0] m16_68;
   assign m16_68 =10'b0;

   // m16_69 = W*in
   wire signed [9:0] m16_69;
   assign m16_69 =10'b0;

   // m16_70 = W*in
   wire signed [9:0] m16_70;
   assign m16_70 =10'b0;

   // m16_71 = W*in
   wire signed [9:0] m16_71;
   assign m16_71 =10'b0;

   // m16_72 = W*in
   wire signed [9:0] m16_72;
   assign m16_72 =10'b0;

   // m16_73 = W*in
   wire signed [9:0] m16_73;
   assign m16_73 =10'b0;

   // m16_74 = W*in
   wire signed [9:0] m16_74;
   assign m16_74 =10'b0;

   // m16_75 = W*in
   wire signed [9:0] m16_75;
   assign m16_75 =10'b0;

   // m16_76 = W*in
   wire signed [9:0] m16_76;
   assign m16_76 =10'b0;

   // m16_77 = W*in
   wire signed [9:0] m16_77;
   assign m16_77 =10'b0;

   // m16_78 = W*in
   wire signed [9:0] m16_78;
   assign m16_78 =10'b0;

   // m16_79 = W*in
   wire signed [9:0] m16_79;
   assign m16_79 =10'b0;

   // m16_80 = W*in
   wire signed [9:0] m16_80;
   assign m16_80 =10'b0;

   // m16_81 = W*in
   wire signed [9:0] m16_81;
   assign m16_81 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m17_1 = W*in
   wire signed [9:0] m17_1;
   assign m17_1 =10'b0;

   // m17_2 = W*in
   wire signed [9:0] m17_2;
   assign m17_2 =10'b0;

   // m17_3 = W*in
   wire signed [9:0] m17_3;
   assign m17_3 =10'b0;

   // m17_4 = W*in
   wire signed [9:0] m17_4;
   assign m17_4 ={ {3{neg17[5]}} , neg17 , {1{1'b0}} };

   // m17_5 = W*in
   wire signed [9:0] m17_5;
   assign m17_5 =10'b0;

   // m17_6 = W*in
   wire signed [9:0] m17_6;
   assign m17_6 =10'b0;

   // m17_7 = W*in
   wire signed [9:0] m17_7;
   assign m17_7 =10'b0;

   // m17_8 = W*in
   wire signed [9:0] m17_8;
   assign m17_8 =10'b0;

   // m17_9 = W*in
   wire signed [9:0] m17_9;
   assign m17_9 =10'b0;

   // m17_10 = W*in
   wire signed [9:0] m17_10;
   assign m17_10 =10'b0;

   // m17_11 = W*in
   wire signed [9:0] m17_11;
   assign m17_11 ={ {3{neg17[5]}} , neg17 , {1{1'b0}} };

   // m17_12 = W*in
   wire signed [9:0] m17_12;
   assign m17_12 =10'b0;

   // m17_13 = W*in
   wire signed [9:0] m17_13;
   assign m17_13 =10'b0;

   // m17_14 = W*in
   wire signed [9:0] m17_14;
   assign m17_14 =10'b0;

   // m17_15 = W*in
   wire signed [9:0] m17_15;
   assign m17_15 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_16 = W*in
   wire signed [9:0] m17_16;
   assign m17_16 =10'b0;

   // m17_17 = W*in
   wire signed [9:0] m17_17;
   assign m17_17 =10'b0;

   // m17_18 = W*in
   wire signed [9:0] m17_18;
   assign m17_18 =10'b0;

   // m17_19 = W*in
   wire signed [9:0] m17_19;
   assign m17_19 =10'b0;

   // m17_20 = W*in
   wire signed [9:0] m17_20;
   assign m17_20 =10'b0;

   // m17_21 = W*in
   wire signed [9:0] m17_21;
   assign m17_21 =10'b0;

   // m17_22 = W*in
   wire signed [9:0] m17_22;
   assign m17_22 =10'b0;

   // m17_23 = W*in
   wire signed [9:0] m17_23;
   assign m17_23 =10'b0;

   // m17_24 = W*in
   wire signed [9:0] m17_24;
   assign m17_24 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_25 = W*in
   wire signed [9:0] m17_25;
   assign m17_25 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_26 = W*in
   wire signed [9:0] m17_26;
   assign m17_26 =10'b0;

   // m17_27 = W*in
   wire signed [9:0] m17_27;
   assign m17_27 =10'b0;

   // m17_28 = W*in
   wire signed [9:0] m17_28;
   assign m17_28 =10'b0;

   // m17_29 = W*in
   wire signed [9:0] m17_29;
   assign m17_29 =10'b0;

   // m17_30 = W*in
   wire signed [9:0] m17_30;
   assign m17_30 =10'b0;

   // m17_31 = W*in
   wire signed [9:0] m17_31;
   assign m17_31 =10'b0;

   // m17_32 = W*in
   wire signed [9:0] m17_32;
   assign m17_32 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_33 = W*in
   wire signed [9:0] m17_33;
   assign m17_33 =10'b0;

   // m17_34 = W*in
   wire signed [9:0] m17_34;
   assign m17_34 =10'b0;

   // m17_35 = W*in
   wire signed [9:0] m17_35;
   assign m17_35 =10'b0;

   // m17_36 = W*in
   wire signed [9:0] m17_36;
   assign m17_36 ={ {3{neg17[5]}} , neg17 , {1{1'b0}} };

   // m17_37 = W*in
   wire signed [9:0] m17_37;
   assign m17_37 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_38 = W*in
   wire signed [9:0] m17_38;
   assign m17_38 ={ {3{neg17[5]}} , neg17 , {1{1'b0}} };

   // m17_39 = W*in
   wire signed [9:0] m17_39;
   assign m17_39 =10'b0;

   // m17_40 = W*in
   wire signed [9:0] m17_40;
   assign m17_40 ={ {2{in17[5]}} , in17 , {2{1'b0}} };

   // m17_41 = W*in
   wire signed [9:0] m17_41;
   assign m17_41 =10'b0;

   // m17_42 = W*in
   wire signed [9:0] m17_42;
   assign m17_42 =10'b0;

   // m17_43 = W*in
   wire signed [9:0] m17_43;
   assign m17_43 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_44 = W*in
   wire signed [9:0] m17_44;
   assign m17_44 =10'b0;

   // m17_45 = W*in
   wire signed [9:0] m17_45;
   assign m17_45 =10'b0;

   // m17_46 = W*in
   wire signed [9:0] m17_46;
   assign m17_46 =10'b0;

   // m17_47 = W*in
   wire signed [9:0] m17_47;
   assign m17_47 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_48 = W*in
   wire signed [9:0] m17_48;
   assign m17_48 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_49 = W*in
   wire signed [9:0] m17_49;
   assign m17_49 =10'b0;

   // m17_50 = W*in
   wire signed [9:0] m17_50;
   assign m17_50 ={ {3{neg17[5]}} , neg17 , {1{1'b0}} };

   // m17_51 = W*in
   wire signed [9:0] m17_51;
   assign m17_51 =10'b0;

   // m17_52 = W*in
   wire signed [9:0] m17_52;
   assign m17_52 =10'b0;

   // m17_53 = W*in
   wire signed [9:0] m17_53;
   assign m17_53 =10'b0;

   // m17_54 = W*in
   wire signed [9:0] m17_54;
   assign m17_54 =10'b0;

   // m17_55 = W*in
   wire signed [9:0] m17_55;
   assign m17_55 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_56 = W*in
   wire signed [9:0] m17_56;
   assign m17_56 =10'b0;

   // m17_57 = W*in
   wire signed [9:0] m17_57;
   assign m17_57 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_58 = W*in
   wire signed [9:0] m17_58;
   assign m17_58 =10'b0;

   // m17_59 = W*in
   wire signed [9:0] m17_59;
   assign m17_59 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_60 = W*in
   wire signed [9:0] m17_60;
   assign m17_60 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_61 = W*in
   wire signed [9:0] m17_61;
   assign m17_61 =10'b0;

   // m17_62 = W*in
   wire signed [9:0] m17_62;
   assign m17_62 =10'b0;

   // m17_63 = W*in
   wire signed [9:0] m17_63;
   assign m17_63 =10'b0;

   // m17_64 = W*in
   wire signed [9:0] m17_64;
   assign m17_64 =10'b0;

   // m17_65 = W*in
   wire signed [9:0] m17_65;
   assign m17_65 =10'b0;

   // m17_66 = W*in
   wire signed [9:0] m17_66;
   assign m17_66 =10'b0;

   // m17_67 = W*in
   wire signed [9:0] m17_67;
   assign m17_67 =10'b0;

   // m17_68 = W*in
   wire signed [9:0] m17_68;
   assign m17_68 ={ {3{neg17[5]}} , neg17 , {1{1'b0}} };

   // m17_69 = W*in
   wire signed [9:0] m17_69;
   assign m17_69 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_70 = W*in
   wire signed [9:0] m17_70;
   assign m17_70 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_71 = W*in
   wire signed [9:0] m17_71;
   assign m17_71 =10'b0;

   // m17_72 = W*in
   wire signed [9:0] m17_72;
   assign m17_72 =10'b0;

   // m17_73 = W*in
   wire signed [9:0] m17_73;
   assign m17_73 =10'b0;

   // m17_74 = W*in
   wire signed [9:0] m17_74;
   assign m17_74 ={ {2{in17[5]}} , in17 , {2{1'b0}} };

   // m17_75 = W*in
   wire signed [9:0] m17_75;
   assign m17_75 =10'b0;

   // m17_76 = W*in
   wire signed [9:0] m17_76;
   assign m17_76 =10'b0;

   // m17_77 = W*in
   wire signed [9:0] m17_77;
   assign m17_77 =10'b0;

   // m17_78 = W*in
   wire signed [9:0] m17_78;
   assign m17_78 =10'b0;

   // m17_79 = W*in
   wire signed [9:0] m17_79;
   assign m17_79 ={ {3{in17[5]}} , in17 , {1{1'b0}} };

   // m17_80 = W*in
   wire signed [9:0] m17_80;
   assign m17_80 =10'b0;

   // m17_81 = W*in
   wire signed [9:0] m17_81;
   assign m17_81 =10'b0;

   // m18_1 = W*in
   wire signed [9:0] m18_1;
   assign m18_1 =10'b0;

   // m18_2 = W*in
   wire signed [9:0] m18_2;
   assign m18_2 ={ {2{in18[5]}} , in18 , {2{1'b0}} };

   // m18_3 = W*in
   wire signed [9:0] m18_3;
   assign m18_3 =10'b0;

   // m18_4 = W*in
   wire signed [9:0] m18_4;
   assign m18_4 =10'b0;

   // m18_5 = W*in
   wire signed [9:0] m18_5;
   assign m18_5 ={ {2{in18[5]}} , in18 , {2{1'b0}} };

   // m18_6 = W*in
   wire signed [9:0] m18_6;
   assign m18_6 =10'b0;

   // m18_7 = W*in
   wire signed [9:0] m18_7;
   assign m18_7 =10'b0;

   // m18_8 = W*in
   wire signed [9:0] m18_8;
   assign m18_8 ={ {2{in18[5]}} , in18 , {2{1'b0}} };

   // m18_9 = W*in
   wire signed [9:0] m18_9;
   assign m18_9 =10'b0;

   // m18_10 = W*in
   wire signed [9:0] m18_10;
   assign m18_10 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_11 = W*in
   wire signed [9:0] m18_11;
   assign m18_11 =10'b0;

   // m18_12 = W*in
   wire signed [9:0] m18_12;
   assign m18_12 =10'b0;

   // m18_13 = W*in
   wire signed [9:0] m18_13;
   assign m18_13 =10'b0;

   // m18_14 = W*in
   wire signed [9:0] m18_14;
   assign m18_14 =10'b0;

   // m18_15 = W*in
   wire signed [9:0] m18_15;
   assign m18_15 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_16 = W*in
   wire signed [9:0] m18_16;
   assign m18_16 =10'b0;

   // m18_17 = W*in
   wire signed [9:0] m18_17;
   assign m18_17 =10'b0;

   // m18_18 = W*in
   wire signed [9:0] m18_18;
   assign m18_18 =10'b0;

   // m18_19 = W*in
   wire signed [9:0] m18_19;
   assign m18_19 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_20 = W*in
   wire signed [9:0] m18_20;
   assign m18_20 =10'b0;

   // m18_21 = W*in
   wire signed [9:0] m18_21;
   assign m18_21 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_22 = W*in
   wire signed [9:0] m18_22;
   assign m18_22 =10'b0;

   // m18_23 = W*in
   wire signed [9:0] m18_23;
   assign m18_23 =10'b0;

   // m18_24 = W*in
   wire signed [9:0] m18_24;
   assign m18_24 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_25 = W*in
   wire signed [9:0] m18_25;
   assign m18_25 =10'b0;

   // m18_26 = W*in
   wire signed [9:0] m18_26;
   assign m18_26 =10'b0;

   // m18_27 = W*in
   wire signed [9:0] m18_27;
   assign m18_27 =10'b0;

   // m18_28 = W*in
   wire signed [9:0] m18_28;
   assign m18_28 =10'b0;

   // m18_29 = W*in
   wire signed [9:0] m18_29;
   assign m18_29 =10'b0;

   // m18_30 = W*in
   wire signed [9:0] m18_30;
   assign m18_30 =10'b0;

   // m18_31 = W*in
   wire signed [9:0] m18_31;
   assign m18_31 =10'b0;

   // m18_32 = W*in
   wire signed [9:0] m18_32;
   assign m18_32 =10'b0;

   // m18_33 = W*in
   wire signed [9:0] m18_33;
   assign m18_33 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_34 = W*in
   wire signed [9:0] m18_34;
   assign m18_34 =10'b0;

   // m18_35 = W*in
   wire signed [9:0] m18_35;
   assign m18_35 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_36 = W*in
   wire signed [9:0] m18_36;
   assign m18_36 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_37 = W*in
   wire signed [9:0] m18_37;
   assign m18_37 =10'b0;

   // m18_38 = W*in
   wire signed [9:0] m18_38;
   assign m18_38 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_39 = W*in
   wire signed [9:0] m18_39;
   assign m18_39 =10'b0;

   // m18_40 = W*in
   wire signed [9:0] m18_40;
   assign m18_40 =10'b0;

   // m18_41 = W*in
   wire signed [9:0] m18_41;
   assign m18_41 =10'b0;

   // m18_42 = W*in
   wire signed [9:0] m18_42;
   assign m18_42 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_43 = W*in
   wire signed [9:0] m18_43;
   assign m18_43 =10'b0;

   // m18_44 = W*in
   wire signed [9:0] m18_44;
   assign m18_44 =10'b0;

   // m18_45 = W*in
   wire signed [9:0] m18_45;
   assign m18_45 =10'b0;

   // m18_46 = W*in
   wire signed [9:0] m18_46;
   assign m18_46 =10'b0;

   // m18_47 = W*in
   wire signed [9:0] m18_47;
   assign m18_47 =10'b0;

   // m18_48 = W*in
   wire signed [9:0] m18_48;
   assign m18_48 =10'b0;

   // m18_49 = W*in
   wire signed [9:0] m18_49;
   assign m18_49 ={ {2{in18[5]}} , in18 , {2{1'b0}} };

   // m18_50 = W*in
   wire signed [9:0] m18_50;
   assign m18_50 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_51 = W*in
   wire signed [9:0] m18_51;
   assign m18_51 =10'b0;

   // m18_52 = W*in
   wire signed [9:0] m18_52;
   assign m18_52 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_53 = W*in
   wire signed [9:0] m18_53;
   assign m18_53 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_54 = W*in
   wire signed [9:0] m18_54;
   assign m18_54 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_55 = W*in
   wire signed [9:0] m18_55;
   assign m18_55 =10'b0;

   // m18_56 = W*in
   wire signed [9:0] m18_56;
   assign m18_56 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_57 = W*in
   wire signed [9:0] m18_57;
   assign m18_57 =10'b0;

   // m18_58 = W*in
   wire signed [9:0] m18_58;
   assign m18_58 =10'b0;

   // m18_59 = W*in
   wire signed [9:0] m18_59;
   assign m18_59 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_60 = W*in
   wire signed [9:0] m18_60;
   assign m18_60 =10'b0;

   // m18_61 = W*in
   wire signed [9:0] m18_61;
   assign m18_61 =10'b0;

   // m18_62 = W*in
   wire signed [9:0] m18_62;
   assign m18_62 =10'b0;

   // m18_63 = W*in
   wire signed [9:0] m18_63;
   assign m18_63 =10'b0;

   // m18_64 = W*in
   wire signed [9:0] m18_64;
   assign m18_64 =10'b0;

   // m18_65 = W*in
   wire signed [9:0] m18_65;
   assign m18_65 =10'b0;

   // m18_66 = W*in
   wire signed [9:0] m18_66;
   assign m18_66 =10'b0;

   // m18_67 = W*in
   wire signed [9:0] m18_67;
   assign m18_67 =10'b0;

   // m18_68 = W*in
   wire signed [9:0] m18_68;
   assign m18_68 =10'b0;

   // m18_69 = W*in
   wire signed [9:0] m18_69;
   assign m18_69 =10'b0;

   // m18_70 = W*in
   wire signed [9:0] m18_70;
   assign m18_70 =10'b0;

   // m18_71 = W*in
   wire signed [9:0] m18_71;
   assign m18_71 ={ {3{in18[5]}} , in18 , {1{1'b0}} };

   // m18_72 = W*in
   wire signed [9:0] m18_72;
   assign m18_72 =10'b0;

   // m18_73 = W*in
   wire signed [9:0] m18_73;
   assign m18_73 ={ {2{in18[5]}} , in18 , {2{1'b0}} };

   // m18_74 = W*in
   wire signed [9:0] m18_74;
   assign m18_74 =10'b0;

   // m18_75 = W*in
   wire signed [9:0] m18_75;
   assign m18_75 =10'b0;

   // m18_76 = W*in
   wire signed [9:0] m18_76;
   assign m18_76 =10'b0;

   // m18_77 = W*in
   wire signed [9:0] m18_77;
   assign m18_77 =10'b0;

   // m18_78 = W*in
   wire signed [9:0] m18_78;
   assign m18_78 ={ {3{neg18[5]}} , neg18 , {1{1'b0}} };

   // m18_79 = W*in
   wire signed [9:0] m18_79;
   assign m18_79 =10'b0;

   // m18_80 = W*in
   wire signed [9:0] m18_80;
   assign m18_80 =10'b0;

   // m18_81 = W*in
   wire signed [9:0] m18_81;
   assign m18_81 =10'b0;

   // m19_1 = W*in
   wire signed [9:0] m19_1;
   assign m19_1 =10'b0;

   // m19_2 = W*in
   wire signed [9:0] m19_2;
   assign m19_2 =10'b0;

   // m19_3 = W*in
   wire signed [9:0] m19_3;
   assign m19_3 =10'b0;

   // m19_4 = W*in
   wire signed [9:0] m19_4;
   assign m19_4 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_5 = W*in
   wire signed [9:0] m19_5;
   assign m19_5 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_6 = W*in
   wire signed [9:0] m19_6;
   assign m19_6 =10'b0;

   // m19_7 = W*in
   wire signed [9:0] m19_7;
   assign m19_7 ={ {2{in19[5]}} , in19 , {2{1'b0}} };

   // m19_8 = W*in
   wire signed [9:0] m19_8;
   assign m19_8 =10'b0;

   // m19_9 = W*in
   wire signed [9:0] m19_9;
   assign m19_9 =10'b0;

   // m19_10 = W*in
   wire signed [9:0] m19_10;
   assign m19_10 =10'b0;

   // m19_11 = W*in
   wire signed [9:0] m19_11;
   assign m19_11 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_12 = W*in
   wire signed [9:0] m19_12;
   assign m19_12 =10'b0;

   // m19_13 = W*in
   wire signed [9:0] m19_13;
   assign m19_13 =10'b0;

   // m19_14 = W*in
   wire signed [9:0] m19_14;
   assign m19_14 =10'b0;

   // m19_15 = W*in
   wire signed [9:0] m19_15;
   assign m19_15 ={ {2{in19[5]}} , in19 , {2{1'b0}} };

   // m19_16 = W*in
   wire signed [9:0] m19_16;
   assign m19_16 =10'b0;

   // m19_17 = W*in
   wire signed [9:0] m19_17;
   assign m19_17 =10'b0;

   // m19_18 = W*in
   wire signed [9:0] m19_18;
   assign m19_18 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_19 = W*in
   wire signed [9:0] m19_19;
   assign m19_19 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_20 = W*in
   wire signed [9:0] m19_20;
   assign m19_20 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_21 = W*in
   wire signed [9:0] m19_21;
   assign m19_21 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_22 = W*in
   wire signed [9:0] m19_22;
   assign m19_22 =10'b0;

   // m19_23 = W*in
   wire signed [9:0] m19_23;
   assign m19_23 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_24 = W*in
   wire signed [9:0] m19_24;
   assign m19_24 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_25 = W*in
   wire signed [9:0] m19_25;
   assign m19_25 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_26 = W*in
   wire signed [9:0] m19_26;
   assign m19_26 =10'b0;

   // m19_27 = W*in
   wire signed [9:0] m19_27;
   assign m19_27 =10'b0;

   // m19_28 = W*in
   wire signed [9:0] m19_28;
   assign m19_28 =10'b0;

   // m19_29 = W*in
   wire signed [9:0] m19_29;
   assign m19_29 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_30 = W*in
   wire signed [9:0] m19_30;
   assign m19_30 =10'b0;

   // m19_31 = W*in
   wire signed [9:0] m19_31;
   assign m19_31 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_32 = W*in
   wire signed [9:0] m19_32;
   assign m19_32 =10'b0;

   // m19_33 = W*in
   wire signed [9:0] m19_33;
   assign m19_33 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_34 = W*in
   wire signed [9:0] m19_34;
   assign m19_34 =10'b0;

   // m19_35 = W*in
   wire signed [9:0] m19_35;
   assign m19_35 =10'b0;

   // m19_36 = W*in
   wire signed [9:0] m19_36;
   assign m19_36 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_37 = W*in
   wire signed [9:0] m19_37;
   assign m19_37 =10'b0;

   // m19_38 = W*in
   wire signed [9:0] m19_38;
   assign m19_38 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_39 = W*in
   wire signed [9:0] m19_39;
   assign m19_39 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_40 = W*in
   wire signed [9:0] m19_40;
   assign m19_40 =10'b0;

   // m19_41 = W*in
   wire signed [9:0] m19_41;
   assign m19_41 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_42 = W*in
   wire signed [9:0] m19_42;
   assign m19_42 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_43 = W*in
   wire signed [9:0] m19_43;
   assign m19_43 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_44 = W*in
   wire signed [9:0] m19_44;
   assign m19_44 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_45 = W*in
   wire signed [9:0] m19_45;
   assign m19_45 =10'b0;

   // m19_46 = W*in
   wire signed [9:0] m19_46;
   assign m19_46 =10'b0;

   // m19_47 = W*in
   wire signed [9:0] m19_47;
   assign m19_47 ={ {2{in19[5]}} , in19 , {2{1'b0}} };

   // m19_48 = W*in
   wire signed [9:0] m19_48;
   assign m19_48 =10'b0;

   // m19_49 = W*in
   wire signed [9:0] m19_49;
   assign m19_49 =10'b0;

   // m19_50 = W*in
   wire signed [9:0] m19_50;
   assign m19_50 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_51 = W*in
   wire signed [9:0] m19_51;
   assign m19_51 ={ {2{in19[5]}} , in19 , {2{1'b0}} };

   // m19_52 = W*in
   wire signed [9:0] m19_52;
   assign m19_52 =10'b0;

   // m19_53 = W*in
   wire signed [9:0] m19_53;
   assign m19_53 =10'b0;

   // m19_54 = W*in
   wire signed [9:0] m19_54;
   assign m19_54 =10'b0;

   // m19_55 = W*in
   wire signed [9:0] m19_55;
   assign m19_55 =10'b0;

   // m19_56 = W*in
   wire signed [9:0] m19_56;
   assign m19_56 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_57 = W*in
   wire signed [9:0] m19_57;
   assign m19_57 =10'b0;

   // m19_58 = W*in
   wire signed [9:0] m19_58;
   assign m19_58 ={ {2{in19[5]}} , in19 , {2{1'b0}} };

   // m19_59 = W*in
   wire signed [9:0] m19_59;
   assign m19_59 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_60 = W*in
   wire signed [9:0] m19_60;
   assign m19_60 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_61 = W*in
   wire signed [9:0] m19_61;
   assign m19_61 =10'b0;

   // m19_62 = W*in
   wire signed [9:0] m19_62;
   assign m19_62 =10'b0;

   // m19_63 = W*in
   wire signed [9:0] m19_63;
   assign m19_63 =10'b0;

   // m19_64 = W*in
   wire signed [9:0] m19_64;
   assign m19_64 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_65 = W*in
   wire signed [9:0] m19_65;
   assign m19_65 =10'b0;

   // m19_66 = W*in
   wire signed [9:0] m19_66;
   assign m19_66 =10'b0;

   // m19_67 = W*in
   wire signed [9:0] m19_67;
   assign m19_67 =10'b0;

   // m19_68 = W*in
   wire signed [9:0] m19_68;
   assign m19_68 =10'b0;

   // m19_69 = W*in
   wire signed [9:0] m19_69;
   assign m19_69 ={ {2{in19[5]}} , in19 , {2{1'b0}} };

   // m19_70 = W*in
   wire signed [9:0] m19_70;
   assign m19_70 =10'b0;

   // m19_71 = W*in
   wire signed [9:0] m19_71;
   assign m19_71 =10'b0;

   // m19_72 = W*in
   wire signed [9:0] m19_72;
   assign m19_72 =10'b0;

   // m19_73 = W*in
   wire signed [9:0] m19_73;
   assign m19_73 =10'b0;

   // m19_74 = W*in
   wire signed [9:0] m19_74;
   assign m19_74 =10'b0;

   // m19_75 = W*in
   wire signed [9:0] m19_75;
   assign m19_75 =10'b0;

   // m19_76 = W*in
   wire signed [9:0] m19_76;
   assign m19_76 =10'b0;

   // m19_77 = W*in
   wire signed [9:0] m19_77;
   assign m19_77 =10'b0;

   // m19_78 = W*in
   wire signed [9:0] m19_78;
   assign m19_78 =10'b0;

   // m19_79 = W*in
   wire signed [9:0] m19_79;
   assign m19_79 ={ {3{in19[5]}} , in19 , {1{1'b0}} };

   // m19_80 = W*in
   wire signed [9:0] m19_80;
   assign m19_80 =10'b0;

   // m19_81 = W*in
   wire signed [9:0] m19_81;
   assign m19_81 =10'b0;

   // m20_1 = W*in
   wire signed [9:0] m20_1;
   assign m20_1 =10'b0;

   // m20_2 = W*in
   wire signed [9:0] m20_2;
   assign m20_2 =10'b0;

   // m20_3 = W*in
   wire signed [9:0] m20_3;
   assign m20_3 =10'b0;

   // m20_4 = W*in
   wire signed [9:0] m20_4;
   assign m20_4 =10'b0;

   // m20_5 = W*in
   wire signed [9:0] m20_5;
   assign m20_5 =10'b0;

   // m20_6 = W*in
   wire signed [9:0] m20_6;
   assign m20_6 =10'b0;

   // m20_7 = W*in
   wire signed [9:0] m20_7;
   assign m20_7 =10'b0;

   // m20_8 = W*in
   wire signed [9:0] m20_8;
   assign m20_8 =10'b0;

   // m20_9 = W*in
   wire signed [9:0] m20_9;
   assign m20_9 =10'b0;

   // m20_10 = W*in
   wire signed [9:0] m20_10;
   assign m20_10 =10'b0;

   // m20_11 = W*in
   wire signed [9:0] m20_11;
   assign m20_11 =10'b0;

   // m20_12 = W*in
   wire signed [9:0] m20_12;
   assign m20_12 =10'b0;

   // m20_13 = W*in
   wire signed [9:0] m20_13;
   assign m20_13 ={ {2{in20[5]}} , in20 , {2{1'b0}} };

   // m20_14 = W*in
   wire signed [9:0] m20_14;
   assign m20_14 =10'b0;

   // m20_15 = W*in
   wire signed [9:0] m20_15;
   assign m20_15 =10'b0;

   // m20_16 = W*in
   wire signed [9:0] m20_16;
   assign m20_16 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_17 = W*in
   wire signed [9:0] m20_17;
   assign m20_17 =10'b0;

   // m20_18 = W*in
   wire signed [9:0] m20_18;
   assign m20_18 =10'b0;

   // m20_19 = W*in
   wire signed [9:0] m20_19;
   assign m20_19 ={ {2{neg20[5]}} , neg20 , {2{1'b0}} };

   // m20_20 = W*in
   wire signed [9:0] m20_20;
   assign m20_20 =10'b0;

   // m20_21 = W*in
   wire signed [9:0] m20_21;
   assign m20_21 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_22 = W*in
   wire signed [9:0] m20_22;
   assign m20_22 =10'b0;

   // m20_23 = W*in
   wire signed [9:0] m20_23;
   assign m20_23 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_24 = W*in
   wire signed [9:0] m20_24;
   assign m20_24 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_25 = W*in
   wire signed [9:0] m20_25;
   assign m20_25 =10'b0;

   // m20_26 = W*in
   wire signed [9:0] m20_26;
   assign m20_26 =10'b0;

   // m20_27 = W*in
   wire signed [9:0] m20_27;
   assign m20_27 ={ {2{in20[5]}} , in20 , {2{1'b0}} };

   // m20_28 = W*in
   wire signed [9:0] m20_28;
   assign m20_28 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_29 = W*in
   wire signed [9:0] m20_29;
   assign m20_29 =10'b0;

   // m20_30 = W*in
   wire signed [9:0] m20_30;
   assign m20_30 ={ {2{in20[5]}} , in20 , {2{1'b0}} };

   // m20_31 = W*in
   wire signed [9:0] m20_31;
   assign m20_31 =10'b0;

   // m20_32 = W*in
   wire signed [9:0] m20_32;
   assign m20_32 ={ {2{in20[5]}} , in20 , {2{1'b0}} };

   // m20_33 = W*in
   wire signed [9:0] m20_33;
   assign m20_33 =10'b0;

   // m20_34 = W*in
   wire signed [9:0] m20_34;
   assign m20_34 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_35 = W*in
   wire signed [9:0] m20_35;
   assign m20_35 ={ {2{in20[5]}} , in20 , {2{1'b0}} };

   // m20_36 = W*in
   wire signed [9:0] m20_36;
   assign m20_36 =10'b0;

   // m20_37 = W*in
   wire signed [9:0] m20_37;
   assign m20_37 =10'b0;

   // m20_38 = W*in
   wire signed [9:0] m20_38;
   assign m20_38 =10'b0;

   // m20_39 = W*in
   wire signed [9:0] m20_39;
   assign m20_39 =10'b0;

   // m20_40 = W*in
   wire signed [9:0] m20_40;
   assign m20_40 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_41 = W*in
   wire signed [9:0] m20_41;
   assign m20_41 =10'b0;

   // m20_42 = W*in
   wire signed [9:0] m20_42;
   assign m20_42 =10'b0;

   // m20_43 = W*in
   wire signed [9:0] m20_43;
   assign m20_43 =10'b0;

   // m20_44 = W*in
   wire signed [9:0] m20_44;
   assign m20_44 =10'b0;

   // m20_45 = W*in
   wire signed [9:0] m20_45;
   assign m20_45 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_46 = W*in
   wire signed [9:0] m20_46;
   assign m20_46 ={ {2{in20[5]}} , in20 , {2{1'b0}} };

   // m20_47 = W*in
   wire signed [9:0] m20_47;
   assign m20_47 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_48 = W*in
   wire signed [9:0] m20_48;
   assign m20_48 =10'b0;

   // m20_49 = W*in
   wire signed [9:0] m20_49;
   assign m20_49 =10'b0;

   // m20_50 = W*in
   wire signed [9:0] m20_50;
   assign m20_50 =10'b0;

   // m20_51 = W*in
   wire signed [9:0] m20_51;
   assign m20_51 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_52 = W*in
   wire signed [9:0] m20_52;
   assign m20_52 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_53 = W*in
   wire signed [9:0] m20_53;
   assign m20_53 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_54 = W*in
   wire signed [9:0] m20_54;
   assign m20_54 =10'b0;

   // m20_55 = W*in
   wire signed [9:0] m20_55;
   assign m20_55 =10'b0;

   // m20_56 = W*in
   wire signed [9:0] m20_56;
   assign m20_56 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_57 = W*in
   wire signed [9:0] m20_57;
   assign m20_57 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_58 = W*in
   wire signed [9:0] m20_58;
   assign m20_58 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_59 = W*in
   wire signed [9:0] m20_59;
   assign m20_59 ={ {3{neg20[5]}} , neg20 , {1{1'b0}} };

   // m20_60 = W*in
   wire signed [9:0] m20_60;
   assign m20_60 =10'b0;

   // m20_61 = W*in
   wire signed [9:0] m20_61;
   assign m20_61 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_62 = W*in
   wire signed [9:0] m20_62;
   assign m20_62 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_63 = W*in
   wire signed [9:0] m20_63;
   assign m20_63 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_64 = W*in
   wire signed [9:0] m20_64;
   assign m20_64 =10'b0;

   // m20_65 = W*in
   wire signed [9:0] m20_65;
   assign m20_65 =10'b0;

   // m20_66 = W*in
   wire signed [9:0] m20_66;
   assign m20_66 =10'b0;

   // m20_67 = W*in
   wire signed [9:0] m20_67;
   assign m20_67 =10'b0;

   // m20_68 = W*in
   wire signed [9:0] m20_68;
   assign m20_68 =10'b0;

   // m20_69 = W*in
   wire signed [9:0] m20_69;
   assign m20_69 =10'b0;

   // m20_70 = W*in
   wire signed [9:0] m20_70;
   assign m20_70 =10'b0;

   // m20_71 = W*in
   wire signed [9:0] m20_71;
   assign m20_71 =10'b0;

   // m20_72 = W*in
   wire signed [9:0] m20_72;
   assign m20_72 =10'b0;

   // m20_73 = W*in
   wire signed [9:0] m20_73;
   assign m20_73 =10'b0;

   // m20_74 = W*in
   wire signed [9:0] m20_74;
   assign m20_74 =10'b0;

   // m20_75 = W*in
   wire signed [9:0] m20_75;
   assign m20_75 =10'b0;

   // m20_76 = W*in
   wire signed [9:0] m20_76;
   assign m20_76 =10'b0;

   // m20_77 = W*in
   wire signed [9:0] m20_77;
   assign m20_77 =10'b0;

   // m20_78 = W*in
   wire signed [9:0] m20_78;
   assign m20_78 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_79 = W*in
   wire signed [9:0] m20_79;
   assign m20_79 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_80 = W*in
   wire signed [9:0] m20_80;
   assign m20_80 =10'b0;

   // m20_81 = W*in
   wire signed [9:0] m20_81;
   assign m20_81 =10'b0;

   // m21_1 = W*in
   wire signed [9:0] m21_1;
   assign m21_1 =10'b0;

   // m21_2 = W*in
   wire signed [9:0] m21_2;
   assign m21_2 =10'b0;

   // m21_3 = W*in
   wire signed [9:0] m21_3;
   assign m21_3 =10'b0;

   // m21_4 = W*in
   wire signed [9:0] m21_4;
   assign m21_4 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_5 = W*in
   wire signed [9:0] m21_5;
   assign m21_5 =10'b0;

   // m21_6 = W*in
   wire signed [9:0] m21_6;
   assign m21_6 =10'b0;

   // m21_7 = W*in
   wire signed [9:0] m21_7;
   assign m21_7 =10'b0;

   // m21_8 = W*in
   wire signed [9:0] m21_8;
   assign m21_8 =10'b0;

   // m21_9 = W*in
   wire signed [9:0] m21_9;
   assign m21_9 =10'b0;

   // m21_10 = W*in
   wire signed [9:0] m21_10;
   assign m21_10 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_11 = W*in
   wire signed [9:0] m21_11;
   assign m21_11 =10'b0;

   // m21_12 = W*in
   wire signed [9:0] m21_12;
   assign m21_12 =10'b0;

   // m21_13 = W*in
   wire signed [9:0] m21_13;
   assign m21_13 =10'b0;

   // m21_14 = W*in
   wire signed [9:0] m21_14;
   assign m21_14 =10'b0;

   // m21_15 = W*in
   wire signed [9:0] m21_15;
   assign m21_15 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_16 = W*in
   wire signed [9:0] m21_16;
   assign m21_16 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_17 = W*in
   wire signed [9:0] m21_17;
   assign m21_17 ={ {4{in21[5]}} , in21[5:0] };

   // m21_18 = W*in
   wire signed [9:0] m21_18;
   assign m21_18 =10'b0;

   // m21_19 = W*in
   wire signed [9:0] m21_19;
   assign m21_19 =10'b0;

   // m21_20 = W*in
   wire signed [9:0] m21_20;
   assign m21_20 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_21 = W*in
   wire signed [9:0] m21_21;
   assign m21_21 =10'b0;

   // m21_22 = W*in
   wire signed [9:0] m21_22;
   assign m21_22 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_23 = W*in
   wire signed [9:0] m21_23;
   assign m21_23 =10'b0;

   // m21_24 = W*in
   wire signed [9:0] m21_24;
   assign m21_24 =10'b0;

   // m21_25 = W*in
   wire signed [9:0] m21_25;
   assign m21_25 =10'b0;

   // m21_26 = W*in
   wire signed [9:0] m21_26;
   assign m21_26 =10'b0;

   // m21_27 = W*in
   wire signed [9:0] m21_27;
   assign m21_27 =10'b0;

   // m21_28 = W*in
   wire signed [9:0] m21_28;
   assign m21_28 =10'b0;

   // m21_29 = W*in
   wire signed [9:0] m21_29;
   assign m21_29 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_30 = W*in
   wire signed [9:0] m21_30;
   assign m21_30 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_31 = W*in
   wire signed [9:0] m21_31;
   assign m21_31 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_32 = W*in
   wire signed [9:0] m21_32;
   assign m21_32 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_33 = W*in
   wire signed [9:0] m21_33;
   assign m21_33 =10'b0;

   // m21_34 = W*in
   wire signed [9:0] m21_34;
   assign m21_34 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_35 = W*in
   wire signed [9:0] m21_35;
   assign m21_35 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_36 = W*in
   wire signed [9:0] m21_36;
   assign m21_36 ={ {2{in21[5]}} , in21 , {2{1'b0}} };

   // m21_37 = W*in
   wire signed [9:0] m21_37;
   assign m21_37 =10'b0;

   // m21_38 = W*in
   wire signed [9:0] m21_38;
   assign m21_38 ={ {2{in21[5]}} , in21 , {2{1'b0}} };

   // m21_39 = W*in
   wire signed [9:0] m21_39;
   assign m21_39 =10'b0;

   // m21_40 = W*in
   wire signed [9:0] m21_40;
   assign m21_40 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_41 = W*in
   wire signed [9:0] m21_41;
   assign m21_41 =10'b0;

   // m21_42 = W*in
   wire signed [9:0] m21_42;
   assign m21_42 =10'b0;

   // m21_43 = W*in
   wire signed [9:0] m21_43;
   assign m21_43 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_44 = W*in
   wire signed [9:0] m21_44;
   assign m21_44 =10'b0;

   // m21_45 = W*in
   wire signed [9:0] m21_45;
   assign m21_45 =10'b0;

   // m21_46 = W*in
   wire signed [9:0] m21_46;
   assign m21_46 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_47 = W*in
   wire signed [9:0] m21_47;
   assign m21_47 =10'b0;

   // m21_48 = W*in
   wire signed [9:0] m21_48;
   assign m21_48 =10'b0;

   // m21_49 = W*in
   wire signed [9:0] m21_49;
   assign m21_49 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_50 = W*in
   wire signed [9:0] m21_50;
   assign m21_50 =10'b0;

   // m21_51 = W*in
   wire signed [9:0] m21_51;
   assign m21_51 =10'b0;

   // m21_52 = W*in
   wire signed [9:0] m21_52;
   assign m21_52 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_53 = W*in
   wire signed [9:0] m21_53;
   assign m21_53 =10'b0;

   // m21_54 = W*in
   wire signed [9:0] m21_54;
   assign m21_54 =10'b0;

   // m21_55 = W*in
   wire signed [9:0] m21_55;
   assign m21_55 =10'b0;

   // m21_56 = W*in
   wire signed [9:0] m21_56;
   assign m21_56 =10'b0;

   // m21_57 = W*in
   wire signed [9:0] m21_57;
   assign m21_57 =10'b0;

   // m21_58 = W*in
   wire signed [9:0] m21_58;
   assign m21_58 =10'b0;

   // m21_59 = W*in
   wire signed [9:0] m21_59;
   assign m21_59 =10'b0;

   // m21_60 = W*in
   wire signed [9:0] m21_60;
   assign m21_60 =10'b0;

   // m21_61 = W*in
   wire signed [9:0] m21_61;
   assign m21_61 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_62 = W*in
   wire signed [9:0] m21_62;
   assign m21_62 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_63 = W*in
   wire signed [9:0] m21_63;
   assign m21_63 =10'b0;

   // m21_64 = W*in
   wire signed [9:0] m21_64;
   assign m21_64 =10'b0;

   // m21_65 = W*in
   wire signed [9:0] m21_65;
   assign m21_65 =10'b0;

   // m21_66 = W*in
   wire signed [9:0] m21_66;
   assign m21_66 =10'b0;

   // m21_67 = W*in
   wire signed [9:0] m21_67;
   assign m21_67 =10'b0;

   // m21_68 = W*in
   wire signed [9:0] m21_68;
   assign m21_68 ={ {3{in21[5]}} , in21 , {1{1'b0}} };

   // m21_69 = W*in
   wire signed [9:0] m21_69;
   assign m21_69 =10'b0;

   // m21_70 = W*in
   wire signed [9:0] m21_70;
   assign m21_70 =10'b0;

   // m21_71 = W*in
   wire signed [9:0] m21_71;
   assign m21_71 =10'b0;

   // m21_72 = W*in
   wire signed [9:0] m21_72;
   assign m21_72 =10'b0;

   // m21_73 = W*in
   wire signed [9:0] m21_73;
   assign m21_73 =10'b0;

   // m21_74 = W*in
   wire signed [9:0] m21_74;
   assign m21_74 =10'b0;

   // m21_75 = W*in
   wire signed [9:0] m21_75;
   assign m21_75 =10'b0;

   // m21_76 = W*in
   wire signed [9:0] m21_76;
   assign m21_76 =10'b0;

   // m21_77 = W*in
   wire signed [9:0] m21_77;
   assign m21_77 ={ {2{in21[5]}} , in21 , {2{1'b0}} };

   // m21_78 = W*in
   wire signed [9:0] m21_78;
   assign m21_78 =10'b0;

   // m21_79 = W*in
   wire signed [9:0] m21_79;
   assign m21_79 ={ {3{neg21[5]}} , neg21 , {1{1'b0}} };

   // m21_80 = W*in
   wire signed [9:0] m21_80;
   assign m21_80 =10'b0;

   // m21_81 = W*in
   wire signed [9:0] m21_81;
   assign m21_81 =10'b0;

   // m22_1 = W*in
   wire signed [9:0] m22_1;
   assign m22_1 =10'b0;

   // m22_2 = W*in
   wire signed [9:0] m22_2;
   assign m22_2 =10'b0;

   // m22_3 = W*in
   wire signed [9:0] m22_3;
   assign m22_3 =10'b0;

   // m22_4 = W*in
   wire signed [9:0] m22_4;
   assign m22_4 =10'b0;

   // m22_5 = W*in
   wire signed [9:0] m22_5;
   assign m22_5 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_6 = W*in
   wire signed [9:0] m22_6;
   assign m22_6 =10'b0;

   // m22_7 = W*in
   wire signed [9:0] m22_7;
   assign m22_7 =10'b0;

   // m22_8 = W*in
   wire signed [9:0] m22_8;
   assign m22_8 =10'b0;

   // m22_9 = W*in
   wire signed [9:0] m22_9;
   assign m22_9 =10'b0;

   // m22_10 = W*in
   wire signed [9:0] m22_10;
   assign m22_10 =10'b0;

   // m22_11 = W*in
   wire signed [9:0] m22_11;
   assign m22_11 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_12 = W*in
   wire signed [9:0] m22_12;
   assign m22_12 =10'b0;

   // m22_13 = W*in
   wire signed [9:0] m22_13;
   assign m22_13 =10'b0;

   // m22_14 = W*in
   wire signed [9:0] m22_14;
   assign m22_14 =10'b0;

   // m22_15 = W*in
   wire signed [9:0] m22_15;
   assign m22_15 =10'b0;

   // m22_16 = W*in
   wire signed [9:0] m22_16;
   assign m22_16 =10'b0;

   // m22_17 = W*in
   wire signed [9:0] m22_17;
   assign m22_17 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_18 = W*in
   wire signed [9:0] m22_18;
   assign m22_18 =10'b0;

   // m22_19 = W*in
   wire signed [9:0] m22_19;
   assign m22_19 =10'b0;

   // m22_20 = W*in
   wire signed [9:0] m22_20;
   assign m22_20 =10'b0;

   // m22_21 = W*in
   wire signed [9:0] m22_21;
   assign m22_21 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_22 = W*in
   wire signed [9:0] m22_22;
   assign m22_22 =10'b0;

   // m22_23 = W*in
   wire signed [9:0] m22_23;
   assign m22_23 =10'b0;

   // m22_24 = W*in
   wire signed [9:0] m22_24;
   assign m22_24 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_25 = W*in
   wire signed [9:0] m22_25;
   assign m22_25 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_26 = W*in
   wire signed [9:0] m22_26;
   assign m22_26 =10'b0;

   // m22_27 = W*in
   wire signed [9:0] m22_27;
   assign m22_27 =10'b0;

   // m22_28 = W*in
   wire signed [9:0] m22_28;
   assign m22_28 ={ {2{in22[5]}} , in22 , {2{1'b0}} };

   // m22_29 = W*in
   wire signed [9:0] m22_29;
   assign m22_29 =10'b0;

   // m22_30 = W*in
   wire signed [9:0] m22_30;
   assign m22_30 =10'b0;

   // m22_31 = W*in
   wire signed [9:0] m22_31;
   assign m22_31 =10'b0;

   // m22_32 = W*in
   wire signed [9:0] m22_32;
   assign m22_32 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_33 = W*in
   wire signed [9:0] m22_33;
   assign m22_33 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_34 = W*in
   wire signed [9:0] m22_34;
   assign m22_34 =10'b0;

   // m22_35 = W*in
   wire signed [9:0] m22_35;
   assign m22_35 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_36 = W*in
   wire signed [9:0] m22_36;
   assign m22_36 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_37 = W*in
   wire signed [9:0] m22_37;
   assign m22_37 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_38 = W*in
   wire signed [9:0] m22_38;
   assign m22_38 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_39 = W*in
   wire signed [9:0] m22_39;
   assign m22_39 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_40 = W*in
   wire signed [9:0] m22_40;
   assign m22_40 =10'b0;

   // m22_41 = W*in
   wire signed [9:0] m22_41;
   assign m22_41 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_42 = W*in
   wire signed [9:0] m22_42;
   assign m22_42 =10'b0;

   // m22_43 = W*in
   wire signed [9:0] m22_43;
   assign m22_43 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_44 = W*in
   wire signed [9:0] m22_44;
   assign m22_44 =10'b0;

   // m22_45 = W*in
   wire signed [9:0] m22_45;
   assign m22_45 =10'b0;

   // m22_46 = W*in
   wire signed [9:0] m22_46;
   assign m22_46 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_47 = W*in
   wire signed [9:0] m22_47;
   assign m22_47 =10'b0;

   // m22_48 = W*in
   wire signed [9:0] m22_48;
   assign m22_48 =10'b0;

   // m22_49 = W*in
   wire signed [9:0] m22_49;
   assign m22_49 =10'b0;

   // m22_50 = W*in
   wire signed [9:0] m22_50;
   assign m22_50 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_51 = W*in
   wire signed [9:0] m22_51;
   assign m22_51 =10'b0;

   // m22_52 = W*in
   wire signed [9:0] m22_52;
   assign m22_52 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_53 = W*in
   wire signed [9:0] m22_53;
   assign m22_53 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_54 = W*in
   wire signed [9:0] m22_54;
   assign m22_54 =10'b0;

   // m22_55 = W*in
   wire signed [9:0] m22_55;
   assign m22_55 =10'b0;

   // m22_56 = W*in
   wire signed [9:0] m22_56;
   assign m22_56 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_57 = W*in
   wire signed [9:0] m22_57;
   assign m22_57 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_58 = W*in
   wire signed [9:0] m22_58;
   assign m22_58 =10'b0;

   // m22_59 = W*in
   wire signed [9:0] m22_59;
   assign m22_59 =10'b0;

   // m22_60 = W*in
   wire signed [9:0] m22_60;
   assign m22_60 =10'b0;

   // m22_61 = W*in
   wire signed [9:0] m22_61;
   assign m22_61 =10'b0;

   // m22_62 = W*in
   wire signed [9:0] m22_62;
   assign m22_62 =10'b0;

   // m22_63 = W*in
   wire signed [9:0] m22_63;
   assign m22_63 =10'b0;

   // m22_64 = W*in
   wire signed [9:0] m22_64;
   assign m22_64 =10'b0;

   // m22_65 = W*in
   wire signed [9:0] m22_65;
   assign m22_65 ={ {2{in22[5]}} , in22 , {2{1'b0}} };

   // m22_66 = W*in
   wire signed [9:0] m22_66;
   assign m22_66 =10'b0;

   // m22_67 = W*in
   wire signed [9:0] m22_67;
   assign m22_67 =10'b0;

   // m22_68 = W*in
   wire signed [9:0] m22_68;
   assign m22_68 =10'b0;

   // m22_69 = W*in
   wire signed [9:0] m22_69;
   assign m22_69 ={ {3{neg22[5]}} , neg22 , {1{1'b0}} };

   // m22_70 = W*in
   wire signed [9:0] m22_70;
   assign m22_70 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_71 = W*in
   wire signed [9:0] m22_71;
   assign m22_71 =10'b0;

   // m22_72 = W*in
   wire signed [9:0] m22_72;
   assign m22_72 ={ {2{in22[5]}} , in22 , {2{1'b0}} };

   // m22_73 = W*in
   wire signed [9:0] m22_73;
   assign m22_73 =10'b0;

   // m22_74 = W*in
   wire signed [9:0] m22_74;
   assign m22_74 =10'b0;

   // m22_75 = W*in
   wire signed [9:0] m22_75;
   assign m22_75 =10'b0;

   // m22_76 = W*in
   wire signed [9:0] m22_76;
   assign m22_76 =10'b0;

   // m22_77 = W*in
   wire signed [9:0] m22_77;
   assign m22_77 =10'b0;

   // m22_78 = W*in
   wire signed [9:0] m22_78;
   assign m22_78 ={ {3{in22[5]}} , in22 , {1{1'b0}} };

   // m22_79 = W*in
   wire signed [9:0] m22_79;
   assign m22_79 =10'b0;

   // m22_80 = W*in
   wire signed [9:0] m22_80;
   assign m22_80 =10'b0;

   // m22_81 = W*in
   wire signed [9:0] m22_81;
   assign m22_81 =10'b0;

   // m23_1 = W*in
   wire signed [9:0] m23_1;
   assign m23_1 =10'b0;

   // m23_2 = W*in
   wire signed [9:0] m23_2;
   assign m23_2 =10'b0;

   // m23_3 = W*in
   wire signed [9:0] m23_3;
   assign m23_3 =10'b0;

   // m23_4 = W*in
   wire signed [9:0] m23_4;
   assign m23_4 =10'b0;

   // m23_5 = W*in
   wire signed [9:0] m23_5;
   assign m23_5 =10'b0;

   // m23_6 = W*in
   wire signed [9:0] m23_6;
   assign m23_6 =10'b0;

   // m23_7 = W*in
   wire signed [9:0] m23_7;
   assign m23_7 =10'b0;

   // m23_8 = W*in
   wire signed [9:0] m23_8;
   assign m23_8 =10'b0;

   // m23_9 = W*in
   wire signed [9:0] m23_9;
   assign m23_9 =10'b0;

   // m23_10 = W*in
   wire signed [9:0] m23_10;
   assign m23_10 =10'b0;

   // m23_11 = W*in
   wire signed [9:0] m23_11;
   assign m23_11 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_12 = W*in
   wire signed [9:0] m23_12;
   assign m23_12 =10'b0;

   // m23_13 = W*in
   wire signed [9:0] m23_13;
   assign m23_13 =10'b0;

   // m23_14 = W*in
   wire signed [9:0] m23_14;
   assign m23_14 =10'b0;

   // m23_15 = W*in
   wire signed [9:0] m23_15;
   assign m23_15 =10'b0;

   // m23_16 = W*in
   wire signed [9:0] m23_16;
   assign m23_16 =10'b0;

   // m23_17 = W*in
   wire signed [9:0] m23_17;
   assign m23_17 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_18 = W*in
   wire signed [9:0] m23_18;
   assign m23_18 =10'b0;

   // m23_19 = W*in
   wire signed [9:0] m23_19;
   assign m23_19 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_20 = W*in
   wire signed [9:0] m23_20;
   assign m23_20 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_21 = W*in
   wire signed [9:0] m23_21;
   assign m23_21 =10'b0;

   // m23_22 = W*in
   wire signed [9:0] m23_22;
   assign m23_22 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_23 = W*in
   wire signed [9:0] m23_23;
   assign m23_23 =10'b0;

   // m23_24 = W*in
   wire signed [9:0] m23_24;
   assign m23_24 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_25 = W*in
   wire signed [9:0] m23_25;
   assign m23_25 =10'b0;

   // m23_26 = W*in
   wire signed [9:0] m23_26;
   assign m23_26 =10'b0;

   // m23_27 = W*in
   wire signed [9:0] m23_27;
   assign m23_27 =10'b0;

   // m23_28 = W*in
   wire signed [9:0] m23_28;
   assign m23_28 =10'b0;

   // m23_29 = W*in
   wire signed [9:0] m23_29;
   assign m23_29 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_30 = W*in
   wire signed [9:0] m23_30;
   assign m23_30 =10'b0;

   // m23_31 = W*in
   wire signed [9:0] m23_31;
   assign m23_31 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_32 = W*in
   wire signed [9:0] m23_32;
   assign m23_32 =10'b0;

   // m23_33 = W*in
   wire signed [9:0] m23_33;
   assign m23_33 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_34 = W*in
   wire signed [9:0] m23_34;
   assign m23_34 =10'b0;

   // m23_35 = W*in
   wire signed [9:0] m23_35;
   assign m23_35 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_36 = W*in
   wire signed [9:0] m23_36;
   assign m23_36 =10'b0;

   // m23_37 = W*in
   wire signed [9:0] m23_37;
   assign m23_37 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_38 = W*in
   wire signed [9:0] m23_38;
   assign m23_38 =10'b0;

   // m23_39 = W*in
   wire signed [9:0] m23_39;
   assign m23_39 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_40 = W*in
   wire signed [9:0] m23_40;
   assign m23_40 =10'b0;

   // m23_41 = W*in
   wire signed [9:0] m23_41;
   assign m23_41 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_42 = W*in
   wire signed [9:0] m23_42;
   assign m23_42 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_43 = W*in
   wire signed [9:0] m23_43;
   assign m23_43 =10'b0;

   // m23_44 = W*in
   wire signed [9:0] m23_44;
   assign m23_44 =10'b0;

   // m23_45 = W*in
   wire signed [9:0] m23_45;
   assign m23_45 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_46 = W*in
   wire signed [9:0] m23_46;
   assign m23_46 =10'b0;

   // m23_47 = W*in
   wire signed [9:0] m23_47;
   assign m23_47 =10'b0;

   // m23_48 = W*in
   wire signed [9:0] m23_48;
   assign m23_48 =10'b0;

   // m23_49 = W*in
   wire signed [9:0] m23_49;
   assign m23_49 =10'b0;

   // m23_50 = W*in
   wire signed [9:0] m23_50;
   assign m23_50 =10'b0;

   // m23_51 = W*in
   wire signed [9:0] m23_51;
   assign m23_51 =10'b0;

   // m23_52 = W*in
   wire signed [9:0] m23_52;
   assign m23_52 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_53 = W*in
   wire signed [9:0] m23_53;
   assign m23_53 =10'b0;

   // m23_54 = W*in
   wire signed [9:0] m23_54;
   assign m23_54 =10'b0;

   // m23_55 = W*in
   wire signed [9:0] m23_55;
   assign m23_55 =10'b0;

   // m23_56 = W*in
   wire signed [9:0] m23_56;
   assign m23_56 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_57 = W*in
   wire signed [9:0] m23_57;
   assign m23_57 =10'b0;

   // m23_58 = W*in
   wire signed [9:0] m23_58;
   assign m23_58 =10'b0;

   // m23_59 = W*in
   wire signed [9:0] m23_59;
   assign m23_59 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_60 = W*in
   wire signed [9:0] m23_60;
   assign m23_60 =10'b0;

   // m23_61 = W*in
   wire signed [9:0] m23_61;
   assign m23_61 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_62 = W*in
   wire signed [9:0] m23_62;
   assign m23_62 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_63 = W*in
   wire signed [9:0] m23_63;
   assign m23_63 =10'b0;

   // m23_64 = W*in
   wire signed [9:0] m23_64;
   assign m23_64 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_65 = W*in
   wire signed [9:0] m23_65;
   assign m23_65 ={ {2{in23[5]}} , in23 , {2{1'b0}} };

   // m23_66 = W*in
   wire signed [9:0] m23_66;
   assign m23_66 =10'b0;

   // m23_67 = W*in
   wire signed [9:0] m23_67;
   assign m23_67 =10'b0;

   // m23_68 = W*in
   wire signed [9:0] m23_68;
   assign m23_68 ={ {3{neg23[5]}} , neg23 , {1{1'b0}} };

   // m23_69 = W*in
   wire signed [9:0] m23_69;
   assign m23_69 =10'b0;

   // m23_70 = W*in
   wire signed [9:0] m23_70;
   assign m23_70 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_71 = W*in
   wire signed [9:0] m23_71;
   assign m23_71 =10'b0;

   // m23_72 = W*in
   wire signed [9:0] m23_72;
   assign m23_72 ={ {2{in23[5]}} , in23 , {2{1'b0}} };

   // m23_73 = W*in
   wire signed [9:0] m23_73;
   assign m23_73 =10'b0;

   // m23_74 = W*in
   wire signed [9:0] m23_74;
   assign m23_74 =10'b0;

   // m23_75 = W*in
   wire signed [9:0] m23_75;
   assign m23_75 =10'b0;

   // m23_76 = W*in
   wire signed [9:0] m23_76;
   assign m23_76 =10'b0;

   // m23_77 = W*in
   wire signed [9:0] m23_77;
   assign m23_77 =10'b0;

   // m23_78 = W*in
   wire signed [9:0] m23_78;
   assign m23_78 ={ {2{in23[5]}} , in23 , {2{1'b0}} };

   // m23_79 = W*in
   wire signed [9:0] m23_79;
   assign m23_79 ={ {3{in23[5]}} , in23 , {1{1'b0}} };

   // m23_80 = W*in
   wire signed [9:0] m23_80;
   assign m23_80 =10'b0;

   // m23_81 = W*in
   wire signed [9:0] m23_81;
   assign m23_81 =10'b0;

   // m24_1 = W*in
   wire signed [9:0] m24_1;
   assign m24_1 =10'b0;

   // m24_2 = W*in
   wire signed [9:0] m24_2;
   assign m24_2 =10'b0;

   // m24_3 = W*in
   wire signed [9:0] m24_3;
   assign m24_3 =10'b0;

   // m24_4 = W*in
   wire signed [9:0] m24_4;
   assign m24_4 =10'b0;

   // m24_5 = W*in
   wire signed [9:0] m24_5;
   assign m24_5 =10'b0;

   // m24_6 = W*in
   wire signed [9:0] m24_6;
   assign m24_6 =10'b0;

   // m24_7 = W*in
   wire signed [9:0] m24_7;
   assign m24_7 =10'b0;

   // m24_8 = W*in
   wire signed [9:0] m24_8;
   assign m24_8 =10'b0;

   // m24_9 = W*in
   wire signed [9:0] m24_9;
   assign m24_9 =10'b0;

   // m24_10 = W*in
   wire signed [9:0] m24_10;
   assign m24_10 =10'b0;

   // m24_11 = W*in
   wire signed [9:0] m24_11;
   assign m24_11 ={ {3{neg24[5]}} , neg24 , {1{1'b0}} };

   // m24_12 = W*in
   wire signed [9:0] m24_12;
   assign m24_12 =10'b0;

   // m24_13 = W*in
   wire signed [9:0] m24_13;
   assign m24_13 =10'b0;

   // m24_14 = W*in
   wire signed [9:0] m24_14;
   assign m24_14 ={ {2{in24[5]}} , in24 , {2{1'b0}} };

   // m24_15 = W*in
   wire signed [9:0] m24_15;
   assign m24_15 =10'b0;

   // m24_16 = W*in
   wire signed [9:0] m24_16;
   assign m24_16 =10'b0;

   // m24_17 = W*in
   wire signed [9:0] m24_17;
   assign m24_17 =10'b0;

   // m24_18 = W*in
   wire signed [9:0] m24_18;
   assign m24_18 =10'b0;

   // m24_19 = W*in
   wire signed [9:0] m24_19;
   assign m24_19 =10'b0;

   // m24_20 = W*in
   wire signed [9:0] m24_20;
   assign m24_20 =10'b0;

   // m24_21 = W*in
   wire signed [9:0] m24_21;
   assign m24_21 =10'b0;

   // m24_22 = W*in
   wire signed [9:0] m24_22;
   assign m24_22 =10'b0;

   // m24_23 = W*in
   wire signed [9:0] m24_23;
   assign m24_23 =10'b0;

   // m24_24 = W*in
   wire signed [9:0] m24_24;
   assign m24_24 =10'b0;

   // m24_25 = W*in
   wire signed [9:0] m24_25;
   assign m24_25 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_26 = W*in
   wire signed [9:0] m24_26;
   assign m24_26 =10'b0;

   // m24_27 = W*in
   wire signed [9:0] m24_27;
   assign m24_27 =10'b0;

   // m24_28 = W*in
   wire signed [9:0] m24_28;
   assign m24_28 =10'b0;

   // m24_29 = W*in
   wire signed [9:0] m24_29;
   assign m24_29 =10'b0;

   // m24_30 = W*in
   wire signed [9:0] m24_30;
   assign m24_30 =10'b0;

   // m24_31 = W*in
   wire signed [9:0] m24_31;
   assign m24_31 =10'b0;

   // m24_32 = W*in
   wire signed [9:0] m24_32;
   assign m24_32 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_33 = W*in
   wire signed [9:0] m24_33;
   assign m24_33 =10'b0;

   // m24_34 = W*in
   wire signed [9:0] m24_34;
   assign m24_34 =10'b0;

   // m24_35 = W*in
   wire signed [9:0] m24_35;
   assign m24_35 =10'b0;

   // m24_36 = W*in
   wire signed [9:0] m24_36;
   assign m24_36 ={ {3{neg24[5]}} , neg24 , {1{1'b0}} };

   // m24_37 = W*in
   wire signed [9:0] m24_37;
   assign m24_37 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_38 = W*in
   wire signed [9:0] m24_38;
   assign m24_38 ={ {3{neg24[5]}} , neg24 , {1{1'b0}} };

   // m24_39 = W*in
   wire signed [9:0] m24_39;
   assign m24_39 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_40 = W*in
   wire signed [9:0] m24_40;
   assign m24_40 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_41 = W*in
   wire signed [9:0] m24_41;
   assign m24_41 =10'b0;

   // m24_42 = W*in
   wire signed [9:0] m24_42;
   assign m24_42 =10'b0;

   // m24_43 = W*in
   wire signed [9:0] m24_43;
   assign m24_43 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_44 = W*in
   wire signed [9:0] m24_44;
   assign m24_44 =10'b0;

   // m24_45 = W*in
   wire signed [9:0] m24_45;
   assign m24_45 =10'b0;

   // m24_46 = W*in
   wire signed [9:0] m24_46;
   assign m24_46 =10'b0;

   // m24_47 = W*in
   wire signed [9:0] m24_47;
   assign m24_47 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_48 = W*in
   wire signed [9:0] m24_48;
   assign m24_48 =10'b0;

   // m24_49 = W*in
   wire signed [9:0] m24_49;
   assign m24_49 ={ {3{neg24[5]}} , neg24 , {1{1'b0}} };

   // m24_50 = W*in
   wire signed [9:0] m24_50;
   assign m24_50 ={ {3{neg24[5]}} , neg24 , {1{1'b0}} };

   // m24_51 = W*in
   wire signed [9:0] m24_51;
   assign m24_51 =10'b0;

   // m24_52 = W*in
   wire signed [9:0] m24_52;
   assign m24_52 =10'b0;

   // m24_53 = W*in
   wire signed [9:0] m24_53;
   assign m24_53 =10'b0;

   // m24_54 = W*in
   wire signed [9:0] m24_54;
   assign m24_54 =10'b0;

   // m24_55 = W*in
   wire signed [9:0] m24_55;
   assign m24_55 =10'b0;

   // m24_56 = W*in
   wire signed [9:0] m24_56;
   assign m24_56 =10'b0;

   // m24_57 = W*in
   wire signed [9:0] m24_57;
   assign m24_57 =10'b0;

   // m24_58 = W*in
   wire signed [9:0] m24_58;
   assign m24_58 =10'b0;

   // m24_59 = W*in
   wire signed [9:0] m24_59;
   assign m24_59 =10'b0;

   // m24_60 = W*in
   wire signed [9:0] m24_60;
   assign m24_60 =10'b0;

   // m24_61 = W*in
   wire signed [9:0] m24_61;
   assign m24_61 =10'b0;

   // m24_62 = W*in
   wire signed [9:0] m24_62;
   assign m24_62 =10'b0;

   // m24_63 = W*in
   wire signed [9:0] m24_63;
   assign m24_63 =10'b0;

   // m24_64 = W*in
   wire signed [9:0] m24_64;
   assign m24_64 =10'b0;

   // m24_65 = W*in
   wire signed [9:0] m24_65;
   assign m24_65 ={ {2{in24[5]}} , in24 , {2{1'b0}} };

   // m24_66 = W*in
   wire signed [9:0] m24_66;
   assign m24_66 =10'b0;

   // m24_67 = W*in
   wire signed [9:0] m24_67;
   assign m24_67 =10'b0;

   // m24_68 = W*in
   wire signed [9:0] m24_68;
   assign m24_68 ={ {3{neg24[5]}} , neg24 , {1{1'b0}} };

   // m24_69 = W*in
   wire signed [9:0] m24_69;
   assign m24_69 =10'b0;

   // m24_70 = W*in
   wire signed [9:0] m24_70;
   assign m24_70 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_71 = W*in
   wire signed [9:0] m24_71;
   assign m24_71 =10'b0;

   // m24_72 = W*in
   wire signed [9:0] m24_72;
   assign m24_72 =10'b0;

   // m24_73 = W*in
   wire signed [9:0] m24_73;
   assign m24_73 =10'b0;

   // m24_74 = W*in
   wire signed [9:0] m24_74;
   assign m24_74 =10'b0;

   // m24_75 = W*in
   wire signed [9:0] m24_75;
   assign m24_75 =10'b0;

   // m24_76 = W*in
   wire signed [9:0] m24_76;
   assign m24_76 =10'b0;

   // m24_77 = W*in
   wire signed [9:0] m24_77;
   assign m24_77 =10'b0;

   // m24_78 = W*in
   wire signed [9:0] m24_78;
   assign m24_78 ={ {3{in24[5]}} , in24 , {1{1'b0}} };

   // m24_79 = W*in
   wire signed [9:0] m24_79;
   assign m24_79 =10'b0;

   // m24_80 = W*in
   wire signed [9:0] m24_80;
   assign m24_80 =10'b0;

   // m24_81 = W*in
   wire signed [9:0] m24_81;
   assign m24_81 =10'b0;

   // m25_1 = W*in
   wire signed [9:0] m25_1;
   assign m25_1 =10'b0;

   // m25_2 = W*in
   wire signed [9:0] m25_2;
   assign m25_2 =10'b0;

   // m25_3 = W*in
   wire signed [9:0] m25_3;
   assign m25_3 =10'b0;

   // m25_4 = W*in
   wire signed [9:0] m25_4;
   assign m25_4 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_5 = W*in
   wire signed [9:0] m25_5;
   assign m25_5 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_6 = W*in
   wire signed [9:0] m25_6;
   assign m25_6 =10'b0;

   // m25_7 = W*in
   wire signed [9:0] m25_7;
   assign m25_7 =10'b0;

   // m25_8 = W*in
   wire signed [9:0] m25_8;
   assign m25_8 =10'b0;

   // m25_9 = W*in
   wire signed [9:0] m25_9;
   assign m25_9 =10'b0;

   // m25_10 = W*in
   wire signed [9:0] m25_10;
   assign m25_10 =10'b0;

   // m25_11 = W*in
   wire signed [9:0] m25_11;
   assign m25_11 =10'b0;

   // m25_12 = W*in
   wire signed [9:0] m25_12;
   assign m25_12 =10'b0;

   // m25_13 = W*in
   wire signed [9:0] m25_13;
   assign m25_13 =10'b0;

   // m25_14 = W*in
   wire signed [9:0] m25_14;
   assign m25_14 =10'b0;

   // m25_15 = W*in
   wire signed [9:0] m25_15;
   assign m25_15 ={ {3{in25[5]}} , in25 , {1{1'b0}} };

   // m25_16 = W*in
   wire signed [9:0] m25_16;
   assign m25_16 =10'b0;

   // m25_17 = W*in
   wire signed [9:0] m25_17;
   assign m25_17 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_18 = W*in
   wire signed [9:0] m25_18;
   assign m25_18 =10'b0;

   // m25_19 = W*in
   wire signed [9:0] m25_19;
   assign m25_19 =10'b0;

   // m25_20 = W*in
   wire signed [9:0] m25_20;
   assign m25_20 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_21 = W*in
   wire signed [9:0] m25_21;
   assign m25_21 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_22 = W*in
   wire signed [9:0] m25_22;
   assign m25_22 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_23 = W*in
   wire signed [9:0] m25_23;
   assign m25_23 ={ {3{in25[5]}} , in25 , {1{1'b0}} };

   // m25_24 = W*in
   wire signed [9:0] m25_24;
   assign m25_24 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_25 = W*in
   wire signed [9:0] m25_25;
   assign m25_25 ={ {3{in25[5]}} , in25 , {1{1'b0}} };

   // m25_26 = W*in
   wire signed [9:0] m25_26;
   assign m25_26 =10'b0;

   // m25_27 = W*in
   wire signed [9:0] m25_27;
   assign m25_27 =10'b0;

   // m25_28 = W*in
   wire signed [9:0] m25_28;
   assign m25_28 =10'b0;

   // m25_29 = W*in
   wire signed [9:0] m25_29;
   assign m25_29 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_30 = W*in
   wire signed [9:0] m25_30;
   assign m25_30 ={ {3{in25[5]}} , in25 , {1{1'b0}} };

   // m25_31 = W*in
   wire signed [9:0] m25_31;
   assign m25_31 =10'b0;

   // m25_32 = W*in
   wire signed [9:0] m25_32;
   assign m25_32 =10'b0;

   // m25_33 = W*in
   wire signed [9:0] m25_33;
   assign m25_33 =10'b0;

   // m25_34 = W*in
   wire signed [9:0] m25_34;
   assign m25_34 =10'b0;

   // m25_35 = W*in
   wire signed [9:0] m25_35;
   assign m25_35 =10'b0;

   // m25_36 = W*in
   wire signed [9:0] m25_36;
   assign m25_36 =10'b0;

   // m25_37 = W*in
   wire signed [9:0] m25_37;
   assign m25_37 =10'b0;

   // m25_38 = W*in
   wire signed [9:0] m25_38;
   assign m25_38 =10'b0;

   // m25_39 = W*in
   wire signed [9:0] m25_39;
   assign m25_39 ={ {3{in25[5]}} , in25 , {1{1'b0}} };

   // m25_40 = W*in
   wire signed [9:0] m25_40;
   assign m25_40 =10'b0;

   // m25_41 = W*in
   wire signed [9:0] m25_41;
   assign m25_41 =10'b0;

   // m25_42 = W*in
   wire signed [9:0] m25_42;
   assign m25_42 =10'b0;

   // m25_43 = W*in
   wire signed [9:0] m25_43;
   assign m25_43 ={ {2{in25[5]}} , in25 , {2{1'b0}} };

   // m25_44 = W*in
   wire signed [9:0] m25_44;
   assign m25_44 ={ {2{in25[5]}} , in25 , {2{1'b0}} };

   // m25_45 = W*in
   wire signed [9:0] m25_45;
   assign m25_45 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_46 = W*in
   wire signed [9:0] m25_46;
   assign m25_46 =10'b0;

   // m25_47 = W*in
   wire signed [9:0] m25_47;
   assign m25_47 =10'b0;

   // m25_48 = W*in
   wire signed [9:0] m25_48;
   assign m25_48 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_49 = W*in
   wire signed [9:0] m25_49;
   assign m25_49 =10'b0;

   // m25_50 = W*in
   wire signed [9:0] m25_50;
   assign m25_50 =10'b0;

   // m25_51 = W*in
   wire signed [9:0] m25_51;
   assign m25_51 =10'b0;

   // m25_52 = W*in
   wire signed [9:0] m25_52;
   assign m25_52 =10'b0;

   // m25_53 = W*in
   wire signed [9:0] m25_53;
   assign m25_53 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_54 = W*in
   wire signed [9:0] m25_54;
   assign m25_54 =10'b0;

   // m25_55 = W*in
   wire signed [9:0] m25_55;
   assign m25_55 ={ {2{in25[5]}} , in25 , {2{1'b0}} };

   // m25_56 = W*in
   wire signed [9:0] m25_56;
   assign m25_56 =10'b0;

   // m25_57 = W*in
   wire signed [9:0] m25_57;
   assign m25_57 =10'b0;

   // m25_58 = W*in
   wire signed [9:0] m25_58;
   assign m25_58 ={ {3{in25[5]}} , in25 , {1{1'b0}} };

   // m25_59 = W*in
   wire signed [9:0] m25_59;
   assign m25_59 =10'b0;

   // m25_60 = W*in
   wire signed [9:0] m25_60;
   assign m25_60 =10'b0;

   // m25_61 = W*in
   wire signed [9:0] m25_61;
   assign m25_61 =10'b0;

   // m25_62 = W*in
   wire signed [9:0] m25_62;
   assign m25_62 ={ {2{in25[5]}} , in25 , {2{1'b0}} };

   // m25_63 = W*in
   wire signed [9:0] m25_63;
   assign m25_63 =10'b0;

   // m25_64 = W*in
   wire signed [9:0] m25_64;
   assign m25_64 =10'b0;

   // m25_65 = W*in
   wire signed [9:0] m25_65;
   assign m25_65 =10'b0;

   // m25_66 = W*in
   wire signed [9:0] m25_66;
   assign m25_66 =10'b0;

   // m25_67 = W*in
   wire signed [9:0] m25_67;
   assign m25_67 =10'b0;

   // m25_68 = W*in
   wire signed [9:0] m25_68;
   assign m25_68 ={ {3{neg25[5]}} , neg25 , {1{1'b0}} };

   // m25_69 = W*in
   wire signed [9:0] m25_69;
   assign m25_69 =10'b0;

   // m25_70 = W*in
   wire signed [9:0] m25_70;
   assign m25_70 =10'b0;

   // m25_71 = W*in
   wire signed [9:0] m25_71;
   assign m25_71 =10'b0;

   // m25_72 = W*in
   wire signed [9:0] m25_72;
   assign m25_72 =10'b0;

   // m25_73 = W*in
   wire signed [9:0] m25_73;
   assign m25_73 =10'b0;

   // m25_74 = W*in
   wire signed [9:0] m25_74;
   assign m25_74 =10'b0;

   // m25_75 = W*in
   wire signed [9:0] m25_75;
   assign m25_75 =10'b0;

   // m25_76 = W*in
   wire signed [9:0] m25_76;
   assign m25_76 =10'b0;

   // m25_77 = W*in
   wire signed [9:0] m25_77;
   assign m25_77 =10'b0;

   // m25_78 = W*in
   wire signed [9:0] m25_78;
   assign m25_78 =10'b0;

   // m25_79 = W*in
   wire signed [9:0] m25_79;
   assign m25_79 =10'b0;

   // m25_80 = W*in
   wire signed [9:0] m25_80;
   assign m25_80 ={ {2{in25[5]}} , in25 , {2{1'b0}} };

   // m25_81 = W*in
   wire signed [9:0] m25_81;
   assign m25_81 ={ {2{in25[5]}} , in25 , {2{1'b0}} };

   // m26_1 = W*in
   wire signed [9:0] m26_1;
   assign m26_1 =10'b0;

   // m26_2 = W*in
   wire signed [9:0] m26_2;
   assign m26_2 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_3 = W*in
   wire signed [9:0] m26_3;
   assign m26_3 =10'b0;

   // m26_4 = W*in
   wire signed [9:0] m26_4;
   assign m26_4 =10'b0;

   // m26_5 = W*in
   wire signed [9:0] m26_5;
   assign m26_5 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_6 = W*in
   wire signed [9:0] m26_6;
   assign m26_6 =10'b0;

   // m26_7 = W*in
   wire signed [9:0] m26_7;
   assign m26_7 =10'b0;

   // m26_8 = W*in
   wire signed [9:0] m26_8;
   assign m26_8 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_9 = W*in
   wire signed [9:0] m26_9;
   assign m26_9 =10'b0;

   // m26_10 = W*in
   wire signed [9:0] m26_10;
   assign m26_10 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_11 = W*in
   wire signed [9:0] m26_11;
   assign m26_11 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_12 = W*in
   wire signed [9:0] m26_12;
   assign m26_12 =10'b0;

   // m26_13 = W*in
   wire signed [9:0] m26_13;
   assign m26_13 =10'b0;

   // m26_14 = W*in
   wire signed [9:0] m26_14;
   assign m26_14 =10'b0;

   // m26_15 = W*in
   wire signed [9:0] m26_15;
   assign m26_15 =10'b0;

   // m26_16 = W*in
   wire signed [9:0] m26_16;
   assign m26_16 =10'b0;

   // m26_17 = W*in
   wire signed [9:0] m26_17;
   assign m26_17 =10'b0;

   // m26_18 = W*in
   wire signed [9:0] m26_18;
   assign m26_18 =10'b0;

   // m26_19 = W*in
   wire signed [9:0] m26_19;
   assign m26_19 =10'b0;

   // m26_20 = W*in
   wire signed [9:0] m26_20;
   assign m26_20 =10'b0;

   // m26_21 = W*in
   wire signed [9:0] m26_21;
   assign m26_21 =10'b0;

   // m26_22 = W*in
   wire signed [9:0] m26_22;
   assign m26_22 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_23 = W*in
   wire signed [9:0] m26_23;
   assign m26_23 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_24 = W*in
   wire signed [9:0] m26_24;
   assign m26_24 =10'b0;

   // m26_25 = W*in
   wire signed [9:0] m26_25;
   assign m26_25 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_26 = W*in
   wire signed [9:0] m26_26;
   assign m26_26 =10'b0;

   // m26_27 = W*in
   wire signed [9:0] m26_27;
   assign m26_27 =10'b0;

   // m26_28 = W*in
   wire signed [9:0] m26_28;
   assign m26_28 =10'b0;

   // m26_29 = W*in
   wire signed [9:0] m26_29;
   assign m26_29 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_30 = W*in
   wire signed [9:0] m26_30;
   assign m26_30 =10'b0;

   // m26_31 = W*in
   wire signed [9:0] m26_31;
   assign m26_31 =10'b0;

   // m26_32 = W*in
   wire signed [9:0] m26_32;
   assign m26_32 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_33 = W*in
   wire signed [9:0] m26_33;
   assign m26_33 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_34 = W*in
   wire signed [9:0] m26_34;
   assign m26_34 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_35 = W*in
   wire signed [9:0] m26_35;
   assign m26_35 =10'b0;

   // m26_36 = W*in
   wire signed [9:0] m26_36;
   assign m26_36 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_37 = W*in
   wire signed [9:0] m26_37;
   assign m26_37 =10'b0;

   // m26_38 = W*in
   wire signed [9:0] m26_38;
   assign m26_38 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_39 = W*in
   wire signed [9:0] m26_39;
   assign m26_39 =10'b0;

   // m26_40 = W*in
   wire signed [9:0] m26_40;
   assign m26_40 =10'b0;

   // m26_41 = W*in
   wire signed [9:0] m26_41;
   assign m26_41 =10'b0;

   // m26_42 = W*in
   wire signed [9:0] m26_42;
   assign m26_42 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_43 = W*in
   wire signed [9:0] m26_43;
   assign m26_43 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_44 = W*in
   wire signed [9:0] m26_44;
   assign m26_44 =10'b0;

   // m26_45 = W*in
   wire signed [9:0] m26_45;
   assign m26_45 =10'b0;

   // m26_46 = W*in
   wire signed [9:0] m26_46;
   assign m26_46 =10'b0;

   // m26_47 = W*in
   wire signed [9:0] m26_47;
   assign m26_47 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_48 = W*in
   wire signed [9:0] m26_48;
   assign m26_48 =10'b0;

   // m26_49 = W*in
   wire signed [9:0] m26_49;
   assign m26_49 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_50 = W*in
   wire signed [9:0] m26_50;
   assign m26_50 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_51 = W*in
   wire signed [9:0] m26_51;
   assign m26_51 =10'b0;

   // m26_52 = W*in
   wire signed [9:0] m26_52;
   assign m26_52 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_53 = W*in
   wire signed [9:0] m26_53;
   assign m26_53 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_54 = W*in
   wire signed [9:0] m26_54;
   assign m26_54 =10'b0;

   // m26_55 = W*in
   wire signed [9:0] m26_55;
   assign m26_55 =10'b0;

   // m26_56 = W*in
   wire signed [9:0] m26_56;
   assign m26_56 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_57 = W*in
   wire signed [9:0] m26_57;
   assign m26_57 =10'b0;

   // m26_58 = W*in
   wire signed [9:0] m26_58;
   assign m26_58 =10'b0;

   // m26_59 = W*in
   wire signed [9:0] m26_59;
   assign m26_59 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_60 = W*in
   wire signed [9:0] m26_60;
   assign m26_60 =10'b0;

   // m26_61 = W*in
   wire signed [9:0] m26_61;
   assign m26_61 =10'b0;

   // m26_62 = W*in
   wire signed [9:0] m26_62;
   assign m26_62 =10'b0;

   // m26_63 = W*in
   wire signed [9:0] m26_63;
   assign m26_63 =10'b0;

   // m26_64 = W*in
   wire signed [9:0] m26_64;
   assign m26_64 =10'b0;

   // m26_65 = W*in
   wire signed [9:0] m26_65;
   assign m26_65 =10'b0;

   // m26_66 = W*in
   wire signed [9:0] m26_66;
   assign m26_66 =10'b0;

   // m26_67 = W*in
   wire signed [9:0] m26_67;
   assign m26_67 =10'b0;

   // m26_68 = W*in
   wire signed [9:0] m26_68;
   assign m26_68 ={ {3{in26[5]}} , in26 , {1{1'b0}} };

   // m26_69 = W*in
   wire signed [9:0] m26_69;
   assign m26_69 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_70 = W*in
   wire signed [9:0] m26_70;
   assign m26_70 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_71 = W*in
   wire signed [9:0] m26_71;
   assign m26_71 =10'b0;

   // m26_72 = W*in
   wire signed [9:0] m26_72;
   assign m26_72 =10'b0;

   // m26_73 = W*in
   wire signed [9:0] m26_73;
   assign m26_73 ={ {2{in26[5]}} , in26 , {2{1'b0}} };

   // m26_74 = W*in
   wire signed [9:0] m26_74;
   assign m26_74 =10'b0;

   // m26_75 = W*in
   wire signed [9:0] m26_75;
   assign m26_75 =10'b0;

   // m26_76 = W*in
   wire signed [9:0] m26_76;
   assign m26_76 =10'b0;

   // m26_77 = W*in
   wire signed [9:0] m26_77;
   assign m26_77 =10'b0;

   // m26_78 = W*in
   wire signed [9:0] m26_78;
   assign m26_78 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_79 = W*in
   wire signed [9:0] m26_79;
   assign m26_79 ={ {3{neg26[5]}} , neg26 , {1{1'b0}} };

   // m26_80 = W*in
   wire signed [9:0] m26_80;
   assign m26_80 =10'b0;

   // m26_81 = W*in
   wire signed [9:0] m26_81;
   assign m26_81 =10'b0;

   // m27_1 = W*in
   wire signed [9:0] m27_1;
   assign m27_1 =10'b0;

   // m27_2 = W*in
   wire signed [9:0] m27_2;
   assign m27_2 =10'b0;

   // m27_3 = W*in
   wire signed [9:0] m27_3;
   assign m27_3 =10'b0;

   // m27_4 = W*in
   wire signed [9:0] m27_4;
   assign m27_4 =10'b0;

   // m27_5 = W*in
   wire signed [9:0] m27_5;
   assign m27_5 =10'b0;

   // m27_6 = W*in
   wire signed [9:0] m27_6;
   assign m27_6 =10'b0;

   // m27_7 = W*in
   wire signed [9:0] m27_7;
   assign m27_7 =10'b0;

   // m27_8 = W*in
   wire signed [9:0] m27_8;
   assign m27_8 ={ {2{in27[5]}} , in27 , {2{1'b0}} };

   // m27_9 = W*in
   wire signed [9:0] m27_9;
   assign m27_9 =10'b0;

   // m27_10 = W*in
   wire signed [9:0] m27_10;
   assign m27_10 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_11 = W*in
   wire signed [9:0] m27_11;
   assign m27_11 =10'b0;

   // m27_12 = W*in
   wire signed [9:0] m27_12;
   assign m27_12 =10'b0;

   // m27_13 = W*in
   wire signed [9:0] m27_13;
   assign m27_13 =10'b0;

   // m27_14 = W*in
   wire signed [9:0] m27_14;
   assign m27_14 =10'b0;

   // m27_15 = W*in
   wire signed [9:0] m27_15;
   assign m27_15 =10'b0;

   // m27_16 = W*in
   wire signed [9:0] m27_16;
   assign m27_16 =10'b0;

   // m27_17 = W*in
   wire signed [9:0] m27_17;
   assign m27_17 ={ {2{neg27[5]}} , neg27 , {2{1'b0}} };

   // m27_18 = W*in
   wire signed [9:0] m27_18;
   assign m27_18 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_19 = W*in
   wire signed [9:0] m27_19;
   assign m27_19 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_20 = W*in
   wire signed [9:0] m27_20;
   assign m27_20 =10'b0;

   // m27_21 = W*in
   wire signed [9:0] m27_21;
   assign m27_21 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_22 = W*in
   wire signed [9:0] m27_22;
   assign m27_22 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_23 = W*in
   wire signed [9:0] m27_23;
   assign m27_23 =10'b0;

   // m27_24 = W*in
   wire signed [9:0] m27_24;
   assign m27_24 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_25 = W*in
   wire signed [9:0] m27_25;
   assign m27_25 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_26 = W*in
   wire signed [9:0] m27_26;
   assign m27_26 =10'b0;

   // m27_27 = W*in
   wire signed [9:0] m27_27;
   assign m27_27 =10'b0;

   // m27_28 = W*in
   wire signed [9:0] m27_28;
   assign m27_28 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_29 = W*in
   wire signed [9:0] m27_29;
   assign m27_29 =10'b0;

   // m27_30 = W*in
   wire signed [9:0] m27_30;
   assign m27_30 ={ {2{in27[5]}} , in27 , {2{1'b0}} };

   // m27_31 = W*in
   wire signed [9:0] m27_31;
   assign m27_31 =10'b0;

   // m27_32 = W*in
   wire signed [9:0] m27_32;
   assign m27_32 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_33 = W*in
   wire signed [9:0] m27_33;
   assign m27_33 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_34 = W*in
   wire signed [9:0] m27_34;
   assign m27_34 =10'b0;

   // m27_35 = W*in
   wire signed [9:0] m27_35;
   assign m27_35 =10'b0;

   // m27_36 = W*in
   wire signed [9:0] m27_36;
   assign m27_36 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_37 = W*in
   wire signed [9:0] m27_37;
   assign m27_37 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_38 = W*in
   wire signed [9:0] m27_38;
   assign m27_38 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_39 = W*in
   wire signed [9:0] m27_39;
   assign m27_39 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_40 = W*in
   wire signed [9:0] m27_40;
   assign m27_40 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_41 = W*in
   wire signed [9:0] m27_41;
   assign m27_41 =10'b0;

   // m27_42 = W*in
   wire signed [9:0] m27_42;
   assign m27_42 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_43 = W*in
   wire signed [9:0] m27_43;
   assign m27_43 ={ {2{in27[5]}} , in27 , {2{1'b0}} };

   // m27_44 = W*in
   wire signed [9:0] m27_44;
   assign m27_44 ={ {2{in27[5]}} , in27 , {2{1'b0}} };

   // m27_45 = W*in
   wire signed [9:0] m27_45;
   assign m27_45 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_46 = W*in
   wire signed [9:0] m27_46;
   assign m27_46 =10'b0;

   // m27_47 = W*in
   wire signed [9:0] m27_47;
   assign m27_47 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_48 = W*in
   wire signed [9:0] m27_48;
   assign m27_48 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_49 = W*in
   wire signed [9:0] m27_49;
   assign m27_49 =10'b0;

   // m27_50 = W*in
   wire signed [9:0] m27_50;
   assign m27_50 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_51 = W*in
   wire signed [9:0] m27_51;
   assign m27_51 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_52 = W*in
   wire signed [9:0] m27_52;
   assign m27_52 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_53 = W*in
   wire signed [9:0] m27_53;
   assign m27_53 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_54 = W*in
   wire signed [9:0] m27_54;
   assign m27_54 =10'b0;

   // m27_55 = W*in
   wire signed [9:0] m27_55;
   assign m27_55 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_56 = W*in
   wire signed [9:0] m27_56;
   assign m27_56 =10'b0;

   // m27_57 = W*in
   wire signed [9:0] m27_57;
   assign m27_57 =10'b0;

   // m27_58 = W*in
   wire signed [9:0] m27_58;
   assign m27_58 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_59 = W*in
   wire signed [9:0] m27_59;
   assign m27_59 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_60 = W*in
   wire signed [9:0] m27_60;
   assign m27_60 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_61 = W*in
   wire signed [9:0] m27_61;
   assign m27_61 =10'b0;

   // m27_62 = W*in
   wire signed [9:0] m27_62;
   assign m27_62 =10'b0;

   // m27_63 = W*in
   wire signed [9:0] m27_63;
   assign m27_63 =10'b0;

   // m27_64 = W*in
   wire signed [9:0] m27_64;
   assign m27_64 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_65 = W*in
   wire signed [9:0] m27_65;
   assign m27_65 =10'b0;

   // m27_66 = W*in
   wire signed [9:0] m27_66;
   assign m27_66 =10'b0;

   // m27_67 = W*in
   wire signed [9:0] m27_67;
   assign m27_67 =10'b0;

   // m27_68 = W*in
   wire signed [9:0] m27_68;
   assign m27_68 ={ {3{neg27[5]}} , neg27 , {1{1'b0}} };

   // m27_69 = W*in
   wire signed [9:0] m27_69;
   assign m27_69 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_70 = W*in
   wire signed [9:0] m27_70;
   assign m27_70 =10'b0;

   // m27_71 = W*in
   wire signed [9:0] m27_71;
   assign m27_71 =10'b0;

   // m27_72 = W*in
   wire signed [9:0] m27_72;
   assign m27_72 =10'b0;

   // m27_73 = W*in
   wire signed [9:0] m27_73;
   assign m27_73 =10'b0;

   // m27_74 = W*in
   wire signed [9:0] m27_74;
   assign m27_74 =10'b0;

   // m27_75 = W*in
   wire signed [9:0] m27_75;
   assign m27_75 =10'b0;

   // m27_76 = W*in
   wire signed [9:0] m27_76;
   assign m27_76 =10'b0;

   // m27_77 = W*in
   wire signed [9:0] m27_77;
   assign m27_77 =10'b0;

   // m27_78 = W*in
   wire signed [9:0] m27_78;
   assign m27_78 ={ {3{in27[5]}} , in27 , {1{1'b0}} };

   // m27_79 = W*in
   wire signed [9:0] m27_79;
   assign m27_79 ={ {2{in27[5]}} , in27 , {2{1'b0}} };

   // m27_80 = W*in
   wire signed [9:0] m27_80;
   assign m27_80 =10'b0;

   // m27_81 = W*in
   wire signed [9:0] m27_81;
   assign m27_81 =10'b0;

   // m28_1 = W*in
   wire signed [9:0] m28_1;
   assign m28_1 =10'b0;

   // m28_2 = W*in
   wire signed [9:0] m28_2;
   assign m28_2 =10'b0;

   // m28_3 = W*in
   wire signed [9:0] m28_3;
   assign m28_3 =10'b0;

   // m28_4 = W*in
   wire signed [9:0] m28_4;
   assign m28_4 =10'b0;

   // m28_5 = W*in
   wire signed [9:0] m28_5;
   assign m28_5 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_6 = W*in
   wire signed [9:0] m28_6;
   assign m28_6 =10'b0;

   // m28_7 = W*in
   wire signed [9:0] m28_7;
   assign m28_7 =10'b0;

   // m28_8 = W*in
   wire signed [9:0] m28_8;
   assign m28_8 =10'b0;

   // m28_9 = W*in
   wire signed [9:0] m28_9;
   assign m28_9 =10'b0;

   // m28_10 = W*in
   wire signed [9:0] m28_10;
   assign m28_10 =10'b0;

   // m28_11 = W*in
   wire signed [9:0] m28_11;
   assign m28_11 =10'b0;

   // m28_12 = W*in
   wire signed [9:0] m28_12;
   assign m28_12 =10'b0;

   // m28_13 = W*in
   wire signed [9:0] m28_13;
   assign m28_13 =10'b0;

   // m28_14 = W*in
   wire signed [9:0] m28_14;
   assign m28_14 =10'b0;

   // m28_15 = W*in
   wire signed [9:0] m28_15;
   assign m28_15 ={ {3{in28[5]}} , in28 , {1{1'b0}} };

   // m28_16 = W*in
   wire signed [9:0] m28_16;
   assign m28_16 =10'b0;

   // m28_17 = W*in
   wire signed [9:0] m28_17;
   assign m28_17 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_18 = W*in
   wire signed [9:0] m28_18;
   assign m28_18 =10'b0;

   // m28_19 = W*in
   wire signed [9:0] m28_19;
   assign m28_19 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_20 = W*in
   wire signed [9:0] m28_20;
   assign m28_20 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_21 = W*in
   wire signed [9:0] m28_21;
   assign m28_21 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_22 = W*in
   wire signed [9:0] m28_22;
   assign m28_22 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_23 = W*in
   wire signed [9:0] m28_23;
   assign m28_23 =10'b0;

   // m28_24 = W*in
   wire signed [9:0] m28_24;
   assign m28_24 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_25 = W*in
   wire signed [9:0] m28_25;
   assign m28_25 ={ {3{in28[5]}} , in28 , {1{1'b0}} };

   // m28_26 = W*in
   wire signed [9:0] m28_26;
   assign m28_26 =10'b0;

   // m28_27 = W*in
   wire signed [9:0] m28_27;
   assign m28_27 =10'b0;

   // m28_28 = W*in
   wire signed [9:0] m28_28;
   assign m28_28 =10'b0;

   // m28_29 = W*in
   wire signed [9:0] m28_29;
   assign m28_29 =10'b0;

   // m28_30 = W*in
   wire signed [9:0] m28_30;
   assign m28_30 ={ {2{in28[5]}} , in28 , {2{1'b0}} };

   // m28_31 = W*in
   wire signed [9:0] m28_31;
   assign m28_31 =10'b0;

   // m28_32 = W*in
   wire signed [9:0] m28_32;
   assign m28_32 =10'b0;

   // m28_33 = W*in
   wire signed [9:0] m28_33;
   assign m28_33 ={ {3{in28[5]}} , in28 , {1{1'b0}} };

   // m28_34 = W*in
   wire signed [9:0] m28_34;
   assign m28_34 =10'b0;

   // m28_35 = W*in
   wire signed [9:0] m28_35;
   assign m28_35 =10'b0;

   // m28_36 = W*in
   wire signed [9:0] m28_36;
   assign m28_36 =10'b0;

   // m28_37 = W*in
   wire signed [9:0] m28_37;
   assign m28_37 =10'b0;

   // m28_38 = W*in
   wire signed [9:0] m28_38;
   assign m28_38 =10'b0;

   // m28_39 = W*in
   wire signed [9:0] m28_39;
   assign m28_39 =10'b0;

   // m28_40 = W*in
   wire signed [9:0] m28_40;
   assign m28_40 =10'b0;

   // m28_41 = W*in
   wire signed [9:0] m28_41;
   assign m28_41 =10'b0;

   // m28_42 = W*in
   wire signed [9:0] m28_42;
   assign m28_42 =10'b0;

   // m28_43 = W*in
   wire signed [9:0] m28_43;
   assign m28_43 ={ {2{in28[5]}} , in28 , {2{1'b0}} };

   // m28_44 = W*in
   wire signed [9:0] m28_44;
   assign m28_44 ={ {3{in28[5]}} , in28 , {1{1'b0}} };

   // m28_45 = W*in
   wire signed [9:0] m28_45;
   assign m28_45 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_46 = W*in
   wire signed [9:0] m28_46;
   assign m28_46 =10'b0;

   // m28_47 = W*in
   wire signed [9:0] m28_47;
   assign m28_47 =10'b0;

   // m28_48 = W*in
   wire signed [9:0] m28_48;
   assign m28_48 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_49 = W*in
   wire signed [9:0] m28_49;
   assign m28_49 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_50 = W*in
   wire signed [9:0] m28_50;
   assign m28_50 =10'b0;

   // m28_51 = W*in
   wire signed [9:0] m28_51;
   assign m28_51 =10'b0;

   // m28_52 = W*in
   wire signed [9:0] m28_52;
   assign m28_52 =10'b0;

   // m28_53 = W*in
   wire signed [9:0] m28_53;
   assign m28_53 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_54 = W*in
   wire signed [9:0] m28_54;
   assign m28_54 =10'b0;

   // m28_55 = W*in
   wire signed [9:0] m28_55;
   assign m28_55 ={ {3{in28[5]}} , in28 , {1{1'b0}} };

   // m28_56 = W*in
   wire signed [9:0] m28_56;
   assign m28_56 =10'b0;

   // m28_57 = W*in
   wire signed [9:0] m28_57;
   assign m28_57 =10'b0;

   // m28_58 = W*in
   wire signed [9:0] m28_58;
   assign m28_58 =10'b0;

   // m28_59 = W*in
   wire signed [9:0] m28_59;
   assign m28_59 =10'b0;

   // m28_60 = W*in
   wire signed [9:0] m28_60;
   assign m28_60 =10'b0;

   // m28_61 = W*in
   wire signed [9:0] m28_61;
   assign m28_61 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_62 = W*in
   wire signed [9:0] m28_62;
   assign m28_62 ={ {2{in28[5]}} , in28 , {2{1'b0}} };

   // m28_63 = W*in
   wire signed [9:0] m28_63;
   assign m28_63 =10'b0;

   // m28_64 = W*in
   wire signed [9:0] m28_64;
   assign m28_64 =10'b0;

   // m28_65 = W*in
   wire signed [9:0] m28_65;
   assign m28_65 =10'b0;

   // m28_66 = W*in
   wire signed [9:0] m28_66;
   assign m28_66 =10'b0;

   // m28_67 = W*in
   wire signed [9:0] m28_67;
   assign m28_67 =10'b0;

   // m28_68 = W*in
   wire signed [9:0] m28_68;
   assign m28_68 ={ {3{neg28[5]}} , neg28 , {1{1'b0}} };

   // m28_69 = W*in
   wire signed [9:0] m28_69;
   assign m28_69 =10'b0;

   // m28_70 = W*in
   wire signed [9:0] m28_70;
   assign m28_70 =10'b0;

   // m28_71 = W*in
   wire signed [9:0] m28_71;
   assign m28_71 =10'b0;

   // m28_72 = W*in
   wire signed [9:0] m28_72;
   assign m28_72 =10'b0;

   // m28_73 = W*in
   wire signed [9:0] m28_73;
   assign m28_73 =10'b0;

   // m28_74 = W*in
   wire signed [9:0] m28_74;
   assign m28_74 =10'b0;

   // m28_75 = W*in
   wire signed [9:0] m28_75;
   assign m28_75 =10'b0;

   // m28_76 = W*in
   wire signed [9:0] m28_76;
   assign m28_76 =10'b0;

   // m28_77 = W*in
   wire signed [9:0] m28_77;
   assign m28_77 =10'b0;

   // m28_78 = W*in
   wire signed [9:0] m28_78;
   assign m28_78 =10'b0;

   // m28_79 = W*in
   wire signed [9:0] m28_79;
   assign m28_79 ={ {3{in28[5]}} , in28 , {1{1'b0}} };

   // m28_80 = W*in
   wire signed [9:0] m28_80;
   assign m28_80 =10'b0;

   // m28_81 = W*in
   wire signed [9:0] m28_81;
   assign m28_81 ={ {2{in28[5]}} , in28 , {2{1'b0}} };

   // m29_1 = W*in
   wire signed [9:0] m29_1;
   assign m29_1 =10'b0;

   // m29_2 = W*in
   wire signed [9:0] m29_2;
   assign m29_2 =10'b0;

   // m29_3 = W*in
   wire signed [9:0] m29_3;
   assign m29_3 =10'b0;

   // m29_4 = W*in
   wire signed [9:0] m29_4;
   assign m29_4 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_5 = W*in
   wire signed [9:0] m29_5;
   assign m29_5 =10'b0;

   // m29_6 = W*in
   wire signed [9:0] m29_6;
   assign m29_6 =10'b0;

   // m29_7 = W*in
   wire signed [9:0] m29_7;
   assign m29_7 =10'b0;

   // m29_8 = W*in
   wire signed [9:0] m29_8;
   assign m29_8 =10'b0;

   // m29_9 = W*in
   wire signed [9:0] m29_9;
   assign m29_9 =10'b0;

   // m29_10 = W*in
   wire signed [9:0] m29_10;
   assign m29_10 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_11 = W*in
   wire signed [9:0] m29_11;
   assign m29_11 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_12 = W*in
   wire signed [9:0] m29_12;
   assign m29_12 =10'b0;

   // m29_13 = W*in
   wire signed [9:0] m29_13;
   assign m29_13 =10'b0;

   // m29_14 = W*in
   wire signed [9:0] m29_14;
   assign m29_14 =10'b0;

   // m29_15 = W*in
   wire signed [9:0] m29_15;
   assign m29_15 =10'b0;

   // m29_16 = W*in
   wire signed [9:0] m29_16;
   assign m29_16 =10'b0;

   // m29_17 = W*in
   wire signed [9:0] m29_17;
   assign m29_17 =10'b0;

   // m29_18 = W*in
   wire signed [9:0] m29_18;
   assign m29_18 =10'b0;

   // m29_19 = W*in
   wire signed [9:0] m29_19;
   assign m29_19 =10'b0;

   // m29_20 = W*in
   wire signed [9:0] m29_20;
   assign m29_20 ={ {2{in29[5]}} , in29 , {2{1'b0}} };

   // m29_21 = W*in
   wire signed [9:0] m29_21;
   assign m29_21 =10'b0;

   // m29_22 = W*in
   wire signed [9:0] m29_22;
   assign m29_22 ={ {2{in29[5]}} , in29 , {2{1'b0}} };

   // m29_23 = W*in
   wire signed [9:0] m29_23;
   assign m29_23 =10'b0;

   // m29_24 = W*in
   wire signed [9:0] m29_24;
   assign m29_24 =10'b0;

   // m29_25 = W*in
   wire signed [9:0] m29_25;
   assign m29_25 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_26 = W*in
   wire signed [9:0] m29_26;
   assign m29_26 =10'b0;

   // m29_27 = W*in
   wire signed [9:0] m29_27;
   assign m29_27 =10'b0;

   // m29_28 = W*in
   wire signed [9:0] m29_28;
   assign m29_28 =10'b0;

   // m29_29 = W*in
   wire signed [9:0] m29_29;
   assign m29_29 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_30 = W*in
   wire signed [9:0] m29_30;
   assign m29_30 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_31 = W*in
   wire signed [9:0] m29_31;
   assign m29_31 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_32 = W*in
   wire signed [9:0] m29_32;
   assign m29_32 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_33 = W*in
   wire signed [9:0] m29_33;
   assign m29_33 =10'b0;

   // m29_34 = W*in
   wire signed [9:0] m29_34;
   assign m29_34 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_35 = W*in
   wire signed [9:0] m29_35;
   assign m29_35 =10'b0;

   // m29_36 = W*in
   wire signed [9:0] m29_36;
   assign m29_36 =10'b0;

   // m29_37 = W*in
   wire signed [9:0] m29_37;
   assign m29_37 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_38 = W*in
   wire signed [9:0] m29_38;
   assign m29_38 =10'b0;

   // m29_39 = W*in
   wire signed [9:0] m29_39;
   assign m29_39 =10'b0;

   // m29_40 = W*in
   wire signed [9:0] m29_40;
   assign m29_40 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_41 = W*in
   wire signed [9:0] m29_41;
   assign m29_41 ={ {2{in29[5]}} , in29 , {2{1'b0}} };

   // m29_42 = W*in
   wire signed [9:0] m29_42;
   assign m29_42 =10'b0;

   // m29_43 = W*in
   wire signed [9:0] m29_43;
   assign m29_43 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_44 = W*in
   wire signed [9:0] m29_44;
   assign m29_44 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_45 = W*in
   wire signed [9:0] m29_45;
   assign m29_45 =10'b0;

   // m29_46 = W*in
   wire signed [9:0] m29_46;
   assign m29_46 =10'b0;

   // m29_47 = W*in
   wire signed [9:0] m29_47;
   assign m29_47 =10'b0;

   // m29_48 = W*in
   wire signed [9:0] m29_48;
   assign m29_48 =10'b0;

   // m29_49 = W*in
   wire signed [9:0] m29_49;
   assign m29_49 =10'b0;

   // m29_50 = W*in
   wire signed [9:0] m29_50;
   assign m29_50 =10'b0;

   // m29_51 = W*in
   wire signed [9:0] m29_51;
   assign m29_51 =10'b0;

   // m29_52 = W*in
   wire signed [9:0] m29_52;
   assign m29_52 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_53 = W*in
   wire signed [9:0] m29_53;
   assign m29_53 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_54 = W*in
   wire signed [9:0] m29_54;
   assign m29_54 =10'b0;

   // m29_55 = W*in
   wire signed [9:0] m29_55;
   assign m29_55 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_56 = W*in
   wire signed [9:0] m29_56;
   assign m29_56 =10'b0;

   // m29_57 = W*in
   wire signed [9:0] m29_57;
   assign m29_57 =10'b0;

   // m29_58 = W*in
   wire signed [9:0] m29_58;
   assign m29_58 =10'b0;

   // m29_59 = W*in
   wire signed [9:0] m29_59;
   assign m29_59 ={ {3{in29[5]}} , in29 , {1{1'b0}} };

   // m29_60 = W*in
   wire signed [9:0] m29_60;
   assign m29_60 =10'b0;

   // m29_61 = W*in
   wire signed [9:0] m29_61;
   assign m29_61 ={ {2{in29[5]}} , in29 , {2{1'b0}} };

   // m29_62 = W*in
   wire signed [9:0] m29_62;
   assign m29_62 ={ {3{neg29[5]}} , neg29 , {1{1'b0}} };

   // m29_63 = W*in
   wire signed [9:0] m29_63;
   assign m29_63 =10'b0;

   // m29_64 = W*in
   wire signed [9:0] m29_64;
   assign m29_64 =10'b0;

   // m29_65 = W*in
   wire signed [9:0] m29_65;
   assign m29_65 =10'b0;

   // m29_66 = W*in
   wire signed [9:0] m29_66;
   assign m29_66 =10'b0;

   // m29_67 = W*in
   wire signed [9:0] m29_67;
   assign m29_67 =10'b0;

   // m29_68 = W*in
   wire signed [9:0] m29_68;
   assign m29_68 =10'b0;

   // m29_69 = W*in
   wire signed [9:0] m29_69;
   assign m29_69 =10'b0;

   // m29_70 = W*in
   wire signed [9:0] m29_70;
   assign m29_70 =10'b0;

   // m29_71 = W*in
   wire signed [9:0] m29_71;
   assign m29_71 =10'b0;

   // m29_72 = W*in
   wire signed [9:0] m29_72;
   assign m29_72 =10'b0;

   // m29_73 = W*in
   wire signed [9:0] m29_73;
   assign m29_73 =10'b0;

   // m29_74 = W*in
   wire signed [9:0] m29_74;
   assign m29_74 =10'b0;

   // m29_75 = W*in
   wire signed [9:0] m29_75;
   assign m29_75 =10'b0;

   // m29_76 = W*in
   wire signed [9:0] m29_76;
   assign m29_76 =10'b0;

   // m29_77 = W*in
   wire signed [9:0] m29_77;
   assign m29_77 ={ {2{in29[5]}} , in29 , {2{1'b0}} };

   // m29_78 = W*in
   wire signed [9:0] m29_78;
   assign m29_78 =10'b0;

   // m29_79 = W*in
   wire signed [9:0] m29_79;
   assign m29_79 =10'b0;

   // m29_80 = W*in
   wire signed [9:0] m29_80;
   assign m29_80 =10'b0;

   // m29_81 = W*in
   wire signed [9:0] m29_81;
   assign m29_81 =10'b0;

   // m30_1 = W*in
   wire signed [9:0] m30_1;
   assign m30_1 =10'b0;

   // m30_2 = W*in
   wire signed [9:0] m30_2;
   assign m30_2 =10'b0;

   // m30_3 = W*in
   wire signed [9:0] m30_3;
   assign m30_3 =10'b0;

   // m30_4 = W*in
   wire signed [9:0] m30_4;
   assign m30_4 =10'b0;

   // m30_5 = W*in
   wire signed [9:0] m30_5;
   assign m30_5 =10'b0;

   // m30_6 = W*in
   wire signed [9:0] m30_6;
   assign m30_6 =10'b0;

   // m30_7 = W*in
   wire signed [9:0] m30_7;
   assign m30_7 =10'b0;

   // m30_8 = W*in
   wire signed [9:0] m30_8;
   assign m30_8 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_9 = W*in
   wire signed [9:0] m30_9;
   assign m30_9 =10'b0;

   // m30_10 = W*in
   wire signed [9:0] m30_10;
   assign m30_10 =10'b0;

   // m30_11 = W*in
   wire signed [9:0] m30_11;
   assign m30_11 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_12 = W*in
   wire signed [9:0] m30_12;
   assign m30_12 =10'b0;

   // m30_13 = W*in
   wire signed [9:0] m30_13;
   assign m30_13 =10'b0;

   // m30_14 = W*in
   wire signed [9:0] m30_14;
   assign m30_14 =10'b0;

   // m30_15 = W*in
   wire signed [9:0] m30_15;
   assign m30_15 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_16 = W*in
   wire signed [9:0] m30_16;
   assign m30_16 ={ {2{in30[5]}} , in30 , {2{1'b0}} };

   // m30_17 = W*in
   wire signed [9:0] m30_17;
   assign m30_17 =10'b0;

   // m30_18 = W*in
   wire signed [9:0] m30_18;
   assign m30_18 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_19 = W*in
   wire signed [9:0] m30_19;
   assign m30_19 =10'b0;

   // m30_20 = W*in
   wire signed [9:0] m30_20;
   assign m30_20 =10'b0;

   // m30_21 = W*in
   wire signed [9:0] m30_21;
   assign m30_21 =10'b0;

   // m30_22 = W*in
   wire signed [9:0] m30_22;
   assign m30_22 =10'b0;

   // m30_23 = W*in
   wire signed [9:0] m30_23;
   assign m30_23 =10'b0;

   // m30_24 = W*in
   wire signed [9:0] m30_24;
   assign m30_24 =10'b0;

   // m30_25 = W*in
   wire signed [9:0] m30_25;
   assign m30_25 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_26 = W*in
   wire signed [9:0] m30_26;
   assign m30_26 =10'b0;

   // m30_27 = W*in
   wire signed [9:0] m30_27;
   assign m30_27 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_28 = W*in
   wire signed [9:0] m30_28;
   assign m30_28 =10'b0;

   // m30_29 = W*in
   wire signed [9:0] m30_29;
   assign m30_29 =10'b0;

   // m30_30 = W*in
   wire signed [9:0] m30_30;
   assign m30_30 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_31 = W*in
   wire signed [9:0] m30_31;
   assign m30_31 =10'b0;

   // m30_32 = W*in
   wire signed [9:0] m30_32;
   assign m30_32 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_33 = W*in
   wire signed [9:0] m30_33;
   assign m30_33 =10'b0;

   // m30_34 = W*in
   wire signed [9:0] m30_34;
   assign m30_34 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_35 = W*in
   wire signed [9:0] m30_35;
   assign m30_35 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_36 = W*in
   wire signed [9:0] m30_36;
   assign m30_36 =10'b0;

   // m30_37 = W*in
   wire signed [9:0] m30_37;
   assign m30_37 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_38 = W*in
   wire signed [9:0] m30_38;
   assign m30_38 =10'b0;

   // m30_39 = W*in
   wire signed [9:0] m30_39;
   assign m30_39 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_40 = W*in
   wire signed [9:0] m30_40;
   assign m30_40 =10'b0;

   // m30_41 = W*in
   wire signed [9:0] m30_41;
   assign m30_41 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_42 = W*in
   wire signed [9:0] m30_42;
   assign m30_42 =10'b0;

   // m30_43 = W*in
   wire signed [9:0] m30_43;
   assign m30_43 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_44 = W*in
   wire signed [9:0] m30_44;
   assign m30_44 =10'b0;

   // m30_45 = W*in
   wire signed [9:0] m30_45;
   assign m30_45 =10'b0;

   // m30_46 = W*in
   wire signed [9:0] m30_46;
   assign m30_46 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_47 = W*in
   wire signed [9:0] m30_47;
   assign m30_47 =10'b0;

   // m30_48 = W*in
   wire signed [9:0] m30_48;
   assign m30_48 =10'b0;

   // m30_49 = W*in
   wire signed [9:0] m30_49;
   assign m30_49 =10'b0;

   // m30_50 = W*in
   wire signed [9:0] m30_50;
   assign m30_50 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_51 = W*in
   wire signed [9:0] m30_51;
   assign m30_51 =10'b0;

   // m30_52 = W*in
   wire signed [9:0] m30_52;
   assign m30_52 =10'b0;

   // m30_53 = W*in
   wire signed [9:0] m30_53;
   assign m30_53 =10'b0;

   // m30_54 = W*in
   wire signed [9:0] m30_54;
   assign m30_54 =10'b0;

   // m30_55 = W*in
   wire signed [9:0] m30_55;
   assign m30_55 =10'b0;

   // m30_56 = W*in
   wire signed [9:0] m30_56;
   assign m30_56 =10'b0;

   // m30_57 = W*in
   wire signed [9:0] m30_57;
   assign m30_57 =10'b0;

   // m30_58 = W*in
   wire signed [9:0] m30_58;
   assign m30_58 ={ {3{neg30[5]}} , neg30 , {1{1'b0}} };

   // m30_59 = W*in
   wire signed [9:0] m30_59;
   assign m30_59 =10'b0;

   // m30_60 = W*in
   wire signed [9:0] m30_60;
   assign m30_60 =10'b0;

   // m30_61 = W*in
   wire signed [9:0] m30_61;
   assign m30_61 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_62 = W*in
   wire signed [9:0] m30_62;
   assign m30_62 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_63 = W*in
   wire signed [9:0] m30_63;
   assign m30_63 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_64 = W*in
   wire signed [9:0] m30_64;
   assign m30_64 =10'b0;

   // m30_65 = W*in
   wire signed [9:0] m30_65;
   assign m30_65 =10'b0;

   // m30_66 = W*in
   wire signed [9:0] m30_66;
   assign m30_66 =10'b0;

   // m30_67 = W*in
   wire signed [9:0] m30_67;
   assign m30_67 =10'b0;

   // m30_68 = W*in
   wire signed [9:0] m30_68;
   assign m30_68 =10'b0;

   // m30_69 = W*in
   wire signed [9:0] m30_69;
   assign m30_69 =10'b0;

   // m30_70 = W*in
   wire signed [9:0] m30_70;
   assign m30_70 =10'b0;

   // m30_71 = W*in
   wire signed [9:0] m30_71;
   assign m30_71 =10'b0;

   // m30_72 = W*in
   wire signed [9:0] m30_72;
   assign m30_72 =10'b0;

   // m30_73 = W*in
   wire signed [9:0] m30_73;
   assign m30_73 =10'b0;

   // m30_74 = W*in
   wire signed [9:0] m30_74;
   assign m30_74 =10'b0;

   // m30_75 = W*in
   wire signed [9:0] m30_75;
   assign m30_75 =10'b0;

   // m30_76 = W*in
   wire signed [9:0] m30_76;
   assign m30_76 =10'b0;

   // m30_77 = W*in
   wire signed [9:0] m30_77;
   assign m30_77 =10'b0;

   // m30_78 = W*in
   wire signed [9:0] m30_78;
   assign m30_78 =10'b0;

   // m30_79 = W*in
   wire signed [9:0] m30_79;
   assign m30_79 ={ {3{in30[5]}} , in30 , {1{1'b0}} };

   // m30_80 = W*in
   wire signed [9:0] m30_80;
   assign m30_80 =10'b0;

   // m30_81 = W*in
   wire signed [9:0] m30_81;
   assign m30_81 =10'b0;

   // m31_1 = W*in
   wire signed [9:0] m31_1;
   assign m31_1 =10'b0;

   // m31_2 = W*in
   wire signed [9:0] m31_2;
   assign m31_2 =10'b0;

   // m31_3 = W*in
   wire signed [9:0] m31_3;
   assign m31_3 =10'b0;

   // m31_4 = W*in
   wire signed [9:0] m31_4;
   assign m31_4 =10'b0;

   // m31_5 = W*in
   wire signed [9:0] m31_5;
   assign m31_5 =10'b0;

   // m31_6 = W*in
   wire signed [9:0] m31_6;
   assign m31_6 =10'b0;

   // m31_7 = W*in
   wire signed [9:0] m31_7;
   assign m31_7 =10'b0;

   // m31_8 = W*in
   wire signed [9:0] m31_8;
   assign m31_8 =10'b0;

   // m31_9 = W*in
   wire signed [9:0] m31_9;
   assign m31_9 =10'b0;

   // m31_10 = W*in
   wire signed [9:0] m31_10;
   assign m31_10 =10'b0;

   // m31_11 = W*in
   wire signed [9:0] m31_11;
   assign m31_11 =10'b0;

   // m31_12 = W*in
   wire signed [9:0] m31_12;
   assign m31_12 =10'b0;

   // m31_13 = W*in
   wire signed [9:0] m31_13;
   assign m31_13 =10'b0;

   // m31_14 = W*in
   wire signed [9:0] m31_14;
   assign m31_14 =10'b0;

   // m31_15 = W*in
   wire signed [9:0] m31_15;
   assign m31_15 =10'b0;

   // m31_16 = W*in
   wire signed [9:0] m31_16;
   assign m31_16 =10'b0;

   // m31_17 = W*in
   wire signed [9:0] m31_17;
   assign m31_17 =10'b0;

   // m31_18 = W*in
   wire signed [9:0] m31_18;
   assign m31_18 =10'b0;

   // m31_19 = W*in
   wire signed [9:0] m31_19;
   assign m31_19 =10'b0;

   // m31_20 = W*in
   wire signed [9:0] m31_20;
   assign m31_20 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_21 = W*in
   wire signed [9:0] m31_21;
   assign m31_21 =10'b0;

   // m31_22 = W*in
   wire signed [9:0] m31_22;
   assign m31_22 =10'b0;

   // m31_23 = W*in
   wire signed [9:0] m31_23;
   assign m31_23 ={ {3{neg31[5]}} , neg31 , {1{1'b0}} };

   // m31_24 = W*in
   wire signed [9:0] m31_24;
   assign m31_24 =10'b0;

   // m31_25 = W*in
   wire signed [9:0] m31_25;
   assign m31_25 ={ {3{neg31[5]}} , neg31 , {1{1'b0}} };

   // m31_26 = W*in
   wire signed [9:0] m31_26;
   assign m31_26 =10'b0;

   // m31_27 = W*in
   wire signed [9:0] m31_27;
   assign m31_27 =10'b0;

   // m31_28 = W*in
   wire signed [9:0] m31_28;
   assign m31_28 =10'b0;

   // m31_29 = W*in
   wire signed [9:0] m31_29;
   assign m31_29 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_30 = W*in
   wire signed [9:0] m31_30;
   assign m31_30 =10'b0;

   // m31_31 = W*in
   wire signed [9:0] m31_31;
   assign m31_31 =10'b0;

   // m31_32 = W*in
   wire signed [9:0] m31_32;
   assign m31_32 =10'b0;

   // m31_33 = W*in
   wire signed [9:0] m31_33;
   assign m31_33 =10'b0;

   // m31_34 = W*in
   wire signed [9:0] m31_34;
   assign m31_34 ={ {3{neg31[5]}} , neg31 , {1{1'b0}} };

   // m31_35 = W*in
   wire signed [9:0] m31_35;
   assign m31_35 =10'b0;

   // m31_36 = W*in
   wire signed [9:0] m31_36;
   assign m31_36 =10'b0;

   // m31_37 = W*in
   wire signed [9:0] m31_37;
   assign m31_37 =10'b0;

   // m31_38 = W*in
   wire signed [9:0] m31_38;
   assign m31_38 =10'b0;

   // m31_39 = W*in
   wire signed [9:0] m31_39;
   assign m31_39 =10'b0;

   // m31_40 = W*in
   wire signed [9:0] m31_40;
   assign m31_40 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_41 = W*in
   wire signed [9:0] m31_41;
   assign m31_41 =10'b0;

   // m31_42 = W*in
   wire signed [9:0] m31_42;
   assign m31_42 ={ {3{neg31[5]}} , neg31 , {1{1'b0}} };

   // m31_43 = W*in
   wire signed [9:0] m31_43;
   assign m31_43 ={ {3{neg31[5]}} , neg31 , {1{1'b0}} };

   // m31_44 = W*in
   wire signed [9:0] m31_44;
   assign m31_44 ={ {2{in31[5]}} , in31 , {2{1'b0}} };

   // m31_45 = W*in
   wire signed [9:0] m31_45;
   assign m31_45 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_46 = W*in
   wire signed [9:0] m31_46;
   assign m31_46 =10'b0;

   // m31_47 = W*in
   wire signed [9:0] m31_47;
   assign m31_47 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_48 = W*in
   wire signed [9:0] m31_48;
   assign m31_48 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_49 = W*in
   wire signed [9:0] m31_49;
   assign m31_49 =10'b0;

   // m31_50 = W*in
   wire signed [9:0] m31_50;
   assign m31_50 =10'b0;

   // m31_51 = W*in
   wire signed [9:0] m31_51;
   assign m31_51 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_52 = W*in
   wire signed [9:0] m31_52;
   assign m31_52 =10'b0;

   // m31_53 = W*in
   wire signed [9:0] m31_53;
   assign m31_53 =10'b0;

   // m31_54 = W*in
   wire signed [9:0] m31_54;
   assign m31_54 =10'b0;

   // m31_55 = W*in
   wire signed [9:0] m31_55;
   assign m31_55 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_56 = W*in
   wire signed [9:0] m31_56;
   assign m31_56 =10'b0;

   // m31_57 = W*in
   wire signed [9:0] m31_57;
   assign m31_57 =10'b0;

   // m31_58 = W*in
   wire signed [9:0] m31_58;
   assign m31_58 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_59 = W*in
   wire signed [9:0] m31_59;
   assign m31_59 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_60 = W*in
   wire signed [9:0] m31_60;
   assign m31_60 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_61 = W*in
   wire signed [9:0] m31_61;
   assign m31_61 =10'b0;

   // m31_62 = W*in
   wire signed [9:0] m31_62;
   assign m31_62 =10'b0;

   // m31_63 = W*in
   wire signed [9:0] m31_63;
   assign m31_63 =10'b0;

   // m31_64 = W*in
   wire signed [9:0] m31_64;
   assign m31_64 =10'b0;

   // m31_65 = W*in
   wire signed [9:0] m31_65;
   assign m31_65 =10'b0;

   // m31_66 = W*in
   wire signed [9:0] m31_66;
   assign m31_66 =10'b0;

   // m31_67 = W*in
   wire signed [9:0] m31_67;
   assign m31_67 =10'b0;

   // m31_68 = W*in
   wire signed [9:0] m31_68;
   assign m31_68 =10'b0;

   // m31_69 = W*in
   wire signed [9:0] m31_69;
   assign m31_69 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_70 = W*in
   wire signed [9:0] m31_70;
   assign m31_70 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_71 = W*in
   wire signed [9:0] m31_71;
   assign m31_71 =10'b0;

   // m31_72 = W*in
   wire signed [9:0] m31_72;
   assign m31_72 =10'b0;

   // m31_73 = W*in
   wire signed [9:0] m31_73;
   assign m31_73 =10'b0;

   // m31_74 = W*in
   wire signed [9:0] m31_74;
   assign m31_74 =10'b0;

   // m31_75 = W*in
   wire signed [9:0] m31_75;
   assign m31_75 =10'b0;

   // m31_76 = W*in
   wire signed [9:0] m31_76;
   assign m31_76 =10'b0;

   // m31_77 = W*in
   wire signed [9:0] m31_77;
   assign m31_77 =10'b0;

   // m31_78 = W*in
   wire signed [9:0] m31_78;
   assign m31_78 =10'b0;

   // m31_79 = W*in
   wire signed [9:0] m31_79;
   assign m31_79 ={ {3{in31[5]}} , in31 , {1{1'b0}} };

   // m31_80 = W*in
   wire signed [9:0] m31_80;
   assign m31_80 =10'b0;

   // m31_81 = W*in
   wire signed [9:0] m31_81;
   assign m31_81 =10'b0;

   // m32_1 = W*in
   wire signed [9:0] m32_1;
   assign m32_1 =10'b0;

   // m32_2 = W*in
   wire signed [9:0] m32_2;
   assign m32_2 =10'b0;

   // m32_3 = W*in
   wire signed [9:0] m32_3;
   assign m32_3 =10'b0;

   // m32_4 = W*in
   wire signed [9:0] m32_4;
   assign m32_4 =10'b0;

   // m32_5 = W*in
   wire signed [9:0] m32_5;
   assign m32_5 =10'b0;

   // m32_6 = W*in
   wire signed [9:0] m32_6;
   assign m32_6 =10'b0;

   // m32_7 = W*in
   wire signed [9:0] m32_7;
   assign m32_7 =10'b0;

   // m32_8 = W*in
   wire signed [9:0] m32_8;
   assign m32_8 =10'b0;

   // m32_9 = W*in
   wire signed [9:0] m32_9;
   assign m32_9 =10'b0;

   // m32_10 = W*in
   wire signed [9:0] m32_10;
   assign m32_10 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_11 = W*in
   wire signed [9:0] m32_11;
   assign m32_11 ={ {3{neg32[5]}} , neg32 , {1{1'b0}} };

   // m32_12 = W*in
   wire signed [9:0] m32_12;
   assign m32_12 =10'b0;

   // m32_13 = W*in
   wire signed [9:0] m32_13;
   assign m32_13 =10'b0;

   // m32_14 = W*in
   wire signed [9:0] m32_14;
   assign m32_14 =10'b0;

   // m32_15 = W*in
   wire signed [9:0] m32_15;
   assign m32_15 =10'b0;

   // m32_16 = W*in
   wire signed [9:0] m32_16;
   assign m32_16 =10'b0;

   // m32_17 = W*in
   wire signed [9:0] m32_17;
   assign m32_17 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_18 = W*in
   wire signed [9:0] m32_18;
   assign m32_18 =10'b0;

   // m32_19 = W*in
   wire signed [9:0] m32_19;
   assign m32_19 =10'b0;

   // m32_20 = W*in
   wire signed [9:0] m32_20;
   assign m32_20 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_21 = W*in
   wire signed [9:0] m32_21;
   assign m32_21 =10'b0;

   // m32_22 = W*in
   wire signed [9:0] m32_22;
   assign m32_22 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_23 = W*in
   wire signed [9:0] m32_23;
   assign m32_23 =10'b0;

   // m32_24 = W*in
   wire signed [9:0] m32_24;
   assign m32_24 =10'b0;

   // m32_25 = W*in
   wire signed [9:0] m32_25;
   assign m32_25 =10'b0;

   // m32_26 = W*in
   wire signed [9:0] m32_26;
   assign m32_26 =10'b0;

   // m32_27 = W*in
   wire signed [9:0] m32_27;
   assign m32_27 =10'b0;

   // m32_28 = W*in
   wire signed [9:0] m32_28;
   assign m32_28 =10'b0;

   // m32_29 = W*in
   wire signed [9:0] m32_29;
   assign m32_29 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_30 = W*in
   wire signed [9:0] m32_30;
   assign m32_30 ={ {3{neg32[5]}} , neg32 , {1{1'b0}} };

   // m32_31 = W*in
   wire signed [9:0] m32_31;
   assign m32_31 =10'b0;

   // m32_32 = W*in
   wire signed [9:0] m32_32;
   assign m32_32 =10'b0;

   // m32_33 = W*in
   wire signed [9:0] m32_33;
   assign m32_33 =10'b0;

   // m32_34 = W*in
   wire signed [9:0] m32_34;
   assign m32_34 =10'b0;

   // m32_35 = W*in
   wire signed [9:0] m32_35;
   assign m32_35 =10'b0;

   // m32_36 = W*in
   wire signed [9:0] m32_36;
   assign m32_36 =10'b0;

   // m32_37 = W*in
   wire signed [9:0] m32_37;
   assign m32_37 =10'b0;

   // m32_38 = W*in
   wire signed [9:0] m32_38;
   assign m32_38 =10'b0;

   // m32_39 = W*in
   wire signed [9:0] m32_39;
   assign m32_39 =10'b0;

   // m32_40 = W*in
   wire signed [9:0] m32_40;
   assign m32_40 =10'b0;

   // m32_41 = W*in
   wire signed [9:0] m32_41;
   assign m32_41 ={ {3{neg32[5]}} , neg32 , {1{1'b0}} };

   // m32_42 = W*in
   wire signed [9:0] m32_42;
   assign m32_42 =10'b0;

   // m32_43 = W*in
   wire signed [9:0] m32_43;
   assign m32_43 =10'b0;

   // m32_44 = W*in
   wire signed [9:0] m32_44;
   assign m32_44 =10'b0;

   // m32_45 = W*in
   wire signed [9:0] m32_45;
   assign m32_45 =10'b0;

   // m32_46 = W*in
   wire signed [9:0] m32_46;
   assign m32_46 =10'b0;

   // m32_47 = W*in
   wire signed [9:0] m32_47;
   assign m32_47 =10'b0;

   // m32_48 = W*in
   wire signed [9:0] m32_48;
   assign m32_48 ={ {2{in32[5]}} , in32 , {2{1'b0}} };

   // m32_49 = W*in
   wire signed [9:0] m32_49;
   assign m32_49 ={ {2{in32[5]}} , in32 , {2{1'b0}} };

   // m32_50 = W*in
   wire signed [9:0] m32_50;
   assign m32_50 ={ {3{neg32[5]}} , neg32 , {1{1'b0}} };

   // m32_51 = W*in
   wire signed [9:0] m32_51;
   assign m32_51 =10'b0;

   // m32_52 = W*in
   wire signed [9:0] m32_52;
   assign m32_52 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_53 = W*in
   wire signed [9:0] m32_53;
   assign m32_53 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_54 = W*in
   wire signed [9:0] m32_54;
   assign m32_54 =10'b0;

   // m32_55 = W*in
   wire signed [9:0] m32_55;
   assign m32_55 =10'b0;

   // m32_56 = W*in
   wire signed [9:0] m32_56;
   assign m32_56 =10'b0;

   // m32_57 = W*in
   wire signed [9:0] m32_57;
   assign m32_57 =10'b0;

   // m32_58 = W*in
   wire signed [9:0] m32_58;
   assign m32_58 =10'b0;

   // m32_59 = W*in
   wire signed [9:0] m32_59;
   assign m32_59 =10'b0;

   // m32_60 = W*in
   wire signed [9:0] m32_60;
   assign m32_60 =10'b0;

   // m32_61 = W*in
   wire signed [9:0] m32_61;
   assign m32_61 =10'b0;

   // m32_62 = W*in
   wire signed [9:0] m32_62;
   assign m32_62 =10'b0;

   // m32_63 = W*in
   wire signed [9:0] m32_63;
   assign m32_63 ={ {3{neg32[5]}} , neg32 , {1{1'b0}} };

   // m32_64 = W*in
   wire signed [9:0] m32_64;
   assign m32_64 =10'b0;

   // m32_65 = W*in
   wire signed [9:0] m32_65;
   assign m32_65 =10'b0;

   // m32_66 = W*in
   wire signed [9:0] m32_66;
   assign m32_66 =10'b0;

   // m32_67 = W*in
   wire signed [9:0] m32_67;
   assign m32_67 =10'b0;

   // m32_68 = W*in
   wire signed [9:0] m32_68;
   assign m32_68 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_69 = W*in
   wire signed [9:0] m32_69;
   assign m32_69 =10'b0;

   // m32_70 = W*in
   wire signed [9:0] m32_70;
   assign m32_70 ={ {3{in32[5]}} , in32 , {1{1'b0}} };

   // m32_71 = W*in
   wire signed [9:0] m32_71;
   assign m32_71 =10'b0;

   // m32_72 = W*in
   wire signed [9:0] m32_72;
   assign m32_72 =10'b0;

   // m32_73 = W*in
   wire signed [9:0] m32_73;
   assign m32_73 =10'b0;

   // m32_74 = W*in
   wire signed [9:0] m32_74;
   assign m32_74 =10'b0;

   // m32_75 = W*in
   wire signed [9:0] m32_75;
   assign m32_75 =10'b0;

   // m32_76 = W*in
   wire signed [9:0] m32_76;
   assign m32_76 =10'b0;

   // m32_77 = W*in
   wire signed [9:0] m32_77;
   assign m32_77 =10'b0;

   // m32_78 = W*in
   wire signed [9:0] m32_78;
   assign m32_78 =10'b0;

   // m32_79 = W*in
   wire signed [9:0] m32_79;
   assign m32_79 =10'b0;

   // m32_80 = W*in
   wire signed [9:0] m32_80;
   assign m32_80 =10'b0;

   // m32_81 = W*in
   wire signed [9:0] m32_81;
   assign m32_81 =10'b0;

   // m33_1 = W*in
   wire signed [9:0] m33_1;
   assign m33_1 =10'b0;

   // m33_2 = W*in
   wire signed [9:0] m33_2;
   assign m33_2 =10'b0;

   // m33_3 = W*in
   wire signed [9:0] m33_3;
   assign m33_3 =10'b0;

   // m33_4 = W*in
   wire signed [9:0] m33_4;
   assign m33_4 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_5 = W*in
   wire signed [9:0] m33_5;
   assign m33_5 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_6 = W*in
   wire signed [9:0] m33_6;
   assign m33_6 =10'b0;

   // m33_7 = W*in
   wire signed [9:0] m33_7;
   assign m33_7 =10'b0;

   // m33_8 = W*in
   wire signed [9:0] m33_8;
   assign m33_8 =10'b0;

   // m33_9 = W*in
   wire signed [9:0] m33_9;
   assign m33_9 =10'b0;

   // m33_10 = W*in
   wire signed [9:0] m33_10;
   assign m33_10 =10'b0;

   // m33_11 = W*in
   wire signed [9:0] m33_11;
   assign m33_11 =10'b0;

   // m33_12 = W*in
   wire signed [9:0] m33_12;
   assign m33_12 =10'b0;

   // m33_13 = W*in
   wire signed [9:0] m33_13;
   assign m33_13 =10'b0;

   // m33_14 = W*in
   wire signed [9:0] m33_14;
   assign m33_14 =10'b0;

   // m33_15 = W*in
   wire signed [9:0] m33_15;
   assign m33_15 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_16 = W*in
   wire signed [9:0] m33_16;
   assign m33_16 =10'b0;

   // m33_17 = W*in
   wire signed [9:0] m33_17;
   assign m33_17 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_18 = W*in
   wire signed [9:0] m33_18;
   assign m33_18 =10'b0;

   // m33_19 = W*in
   wire signed [9:0] m33_19;
   assign m33_19 =10'b0;

   // m33_20 = W*in
   wire signed [9:0] m33_20;
   assign m33_20 =10'b0;

   // m33_21 = W*in
   wire signed [9:0] m33_21;
   assign m33_21 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_22 = W*in
   wire signed [9:0] m33_22;
   assign m33_22 =10'b0;

   // m33_23 = W*in
   wire signed [9:0] m33_23;
   assign m33_23 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_24 = W*in
   wire signed [9:0] m33_24;
   assign m33_24 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_25 = W*in
   wire signed [9:0] m33_25;
   assign m33_25 =10'b0;

   // m33_26 = W*in
   wire signed [9:0] m33_26;
   assign m33_26 =10'b0;

   // m33_27 = W*in
   wire signed [9:0] m33_27;
   assign m33_27 =10'b0;

   // m33_28 = W*in
   wire signed [9:0] m33_28;
   assign m33_28 =10'b0;

   // m33_29 = W*in
   wire signed [9:0] m33_29;
   assign m33_29 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_30 = W*in
   wire signed [9:0] m33_30;
   assign m33_30 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_31 = W*in
   wire signed [9:0] m33_31;
   assign m33_31 =10'b0;

   // m33_32 = W*in
   wire signed [9:0] m33_32;
   assign m33_32 =10'b0;

   // m33_33 = W*in
   wire signed [9:0] m33_33;
   assign m33_33 =10'b0;

   // m33_34 = W*in
   wire signed [9:0] m33_34;
   assign m33_34 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_35 = W*in
   wire signed [9:0] m33_35;
   assign m33_35 =10'b0;

   // m33_36 = W*in
   wire signed [9:0] m33_36;
   assign m33_36 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_37 = W*in
   wire signed [9:0] m33_37;
   assign m33_37 =10'b0;

   // m33_38 = W*in
   wire signed [9:0] m33_38;
   assign m33_38 =10'b0;

   // m33_39 = W*in
   wire signed [9:0] m33_39;
   assign m33_39 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_40 = W*in
   wire signed [9:0] m33_40;
   assign m33_40 =10'b0;

   // m33_41 = W*in
   wire signed [9:0] m33_41;
   assign m33_41 =10'b0;

   // m33_42 = W*in
   wire signed [9:0] m33_42;
   assign m33_42 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_43 = W*in
   wire signed [9:0] m33_43;
   assign m33_43 ={ {2{in33[5]}} , in33 , {2{1'b0}} };

   // m33_44 = W*in
   wire signed [9:0] m33_44;
   assign m33_44 ={ {2{in33[5]}} , in33 , {2{1'b0}} };

   // m33_45 = W*in
   wire signed [9:0] m33_45;
   assign m33_45 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_46 = W*in
   wire signed [9:0] m33_46;
   assign m33_46 =10'b0;

   // m33_47 = W*in
   wire signed [9:0] m33_47;
   assign m33_47 =10'b0;

   // m33_48 = W*in
   wire signed [9:0] m33_48;
   assign m33_48 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_49 = W*in
   wire signed [9:0] m33_49;
   assign m33_49 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_50 = W*in
   wire signed [9:0] m33_50;
   assign m33_50 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_51 = W*in
   wire signed [9:0] m33_51;
   assign m33_51 =10'b0;

   // m33_52 = W*in
   wire signed [9:0] m33_52;
   assign m33_52 =10'b0;

   // m33_53 = W*in
   wire signed [9:0] m33_53;
   assign m33_53 =10'b0;

   // m33_54 = W*in
   wire signed [9:0] m33_54;
   assign m33_54 =10'b0;

   // m33_55 = W*in
   wire signed [9:0] m33_55;
   assign m33_55 =10'b0;

   // m33_56 = W*in
   wire signed [9:0] m33_56;
   assign m33_56 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_57 = W*in
   wire signed [9:0] m33_57;
   assign m33_57 =10'b0;

   // m33_58 = W*in
   wire signed [9:0] m33_58;
   assign m33_58 ={ {3{in33[5]}} , in33 , {1{1'b0}} };

   // m33_59 = W*in
   wire signed [9:0] m33_59;
   assign m33_59 =10'b0;

   // m33_60 = W*in
   wire signed [9:0] m33_60;
   assign m33_60 =10'b0;

   // m33_61 = W*in
   wire signed [9:0] m33_61;
   assign m33_61 =10'b0;

   // m33_62 = W*in
   wire signed [9:0] m33_62;
   assign m33_62 ={ {2{in33[5]}} , in33 , {2{1'b0}} };

   // m33_63 = W*in
   wire signed [9:0] m33_63;
   assign m33_63 =10'b0;

   // m33_64 = W*in
   wire signed [9:0] m33_64;
   assign m33_64 =10'b0;

   // m33_65 = W*in
   wire signed [9:0] m33_65;
   assign m33_65 =10'b0;

   // m33_66 = W*in
   wire signed [9:0] m33_66;
   assign m33_66 =10'b0;

   // m33_67 = W*in
   wire signed [9:0] m33_67;
   assign m33_67 =10'b0;

   // m33_68 = W*in
   wire signed [9:0] m33_68;
   assign m33_68 ={ {3{neg33[5]}} , neg33 , {1{1'b0}} };

   // m33_69 = W*in
   wire signed [9:0] m33_69;
   assign m33_69 =10'b0;

   // m33_70 = W*in
   wire signed [9:0] m33_70;
   assign m33_70 =10'b0;

   // m33_71 = W*in
   wire signed [9:0] m33_71;
   assign m33_71 =10'b0;

   // m33_72 = W*in
   wire signed [9:0] m33_72;
   assign m33_72 =10'b0;

   // m33_73 = W*in
   wire signed [9:0] m33_73;
   assign m33_73 =10'b0;

   // m33_74 = W*in
   wire signed [9:0] m33_74;
   assign m33_74 =10'b0;

   // m33_75 = W*in
   wire signed [9:0] m33_75;
   assign m33_75 =10'b0;

   // m33_76 = W*in
   wire signed [9:0] m33_76;
   assign m33_76 =10'b0;

   // m33_77 = W*in
   wire signed [9:0] m33_77;
   assign m33_77 =10'b0;

   // m33_78 = W*in
   wire signed [9:0] m33_78;
   assign m33_78 =10'b0;

   // m33_79 = W*in
   wire signed [9:0] m33_79;
   assign m33_79 =10'b0;

   // m33_80 = W*in
   wire signed [9:0] m33_80;
   assign m33_80 =10'b0;

   // m33_81 = W*in
   wire signed [9:0] m33_81;
   assign m33_81 =10'b0;

   // m34_1 = W*in
   wire signed [9:0] m34_1;
   assign m34_1 =10'b0;

   // m34_2 = W*in
   wire signed [9:0] m34_2;
   assign m34_2 =10'b0;

   // m34_3 = W*in
   wire signed [9:0] m34_3;
   assign m34_3 =10'b0;

   // m34_4 = W*in
   wire signed [9:0] m34_4;
   assign m34_4 =10'b0;

   // m34_5 = W*in
   wire signed [9:0] m34_5;
   assign m34_5 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_6 = W*in
   wire signed [9:0] m34_6;
   assign m34_6 =10'b0;

   // m34_7 = W*in
   wire signed [9:0] m34_7;
   assign m34_7 =10'b0;

   // m34_8 = W*in
   wire signed [9:0] m34_8;
   assign m34_8 =10'b0;

   // m34_9 = W*in
   wire signed [9:0] m34_9;
   assign m34_9 =10'b0;

   // m34_10 = W*in
   wire signed [9:0] m34_10;
   assign m34_10 =10'b0;

   // m34_11 = W*in
   wire signed [9:0] m34_11;
   assign m34_11 ={ {3{neg34[5]}} , neg34 , {1{1'b0}} };

   // m34_12 = W*in
   wire signed [9:0] m34_12;
   assign m34_12 =10'b0;

   // m34_13 = W*in
   wire signed [9:0] m34_13;
   assign m34_13 =10'b0;

   // m34_14 = W*in
   wire signed [9:0] m34_14;
   assign m34_14 =10'b0;

   // m34_15 = W*in
   wire signed [9:0] m34_15;
   assign m34_15 ={ {3{neg34[5]}} , neg34 , {1{1'b0}} };

   // m34_16 = W*in
   wire signed [9:0] m34_16;
   assign m34_16 =10'b0;

   // m34_17 = W*in
   wire signed [9:0] m34_17;
   assign m34_17 =10'b0;

   // m34_18 = W*in
   wire signed [9:0] m34_18;
   assign m34_18 =10'b0;

   // m34_19 = W*in
   wire signed [9:0] m34_19;
   assign m34_19 =10'b0;

   // m34_20 = W*in
   wire signed [9:0] m34_20;
   assign m34_20 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_21 = W*in
   wire signed [9:0] m34_21;
   assign m34_21 =10'b0;

   // m34_22 = W*in
   wire signed [9:0] m34_22;
   assign m34_22 =10'b0;

   // m34_23 = W*in
   wire signed [9:0] m34_23;
   assign m34_23 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_24 = W*in
   wire signed [9:0] m34_24;
   assign m34_24 ={ {2{in34[5]}} , in34 , {2{1'b0}} };

   // m34_25 = W*in
   wire signed [9:0] m34_25;
   assign m34_25 =10'b0;

   // m34_26 = W*in
   wire signed [9:0] m34_26;
   assign m34_26 =10'b0;

   // m34_27 = W*in
   wire signed [9:0] m34_27;
   assign m34_27 =10'b0;

   // m34_28 = W*in
   wire signed [9:0] m34_28;
   assign m34_28 ={ {2{in34[5]}} , in34 , {2{1'b0}} };

   // m34_29 = W*in
   wire signed [9:0] m34_29;
   assign m34_29 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_30 = W*in
   wire signed [9:0] m34_30;
   assign m34_30 =10'b0;

   // m34_31 = W*in
   wire signed [9:0] m34_31;
   assign m34_31 =10'b0;

   // m34_32 = W*in
   wire signed [9:0] m34_32;
   assign m34_32 =10'b0;

   // m34_33 = W*in
   wire signed [9:0] m34_33;
   assign m34_33 =10'b0;

   // m34_34 = W*in
   wire signed [9:0] m34_34;
   assign m34_34 =10'b0;

   // m34_35 = W*in
   wire signed [9:0] m34_35;
   assign m34_35 =10'b0;

   // m34_36 = W*in
   wire signed [9:0] m34_36;
   assign m34_36 =10'b0;

   // m34_37 = W*in
   wire signed [9:0] m34_37;
   assign m34_37 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_38 = W*in
   wire signed [9:0] m34_38;
   assign m34_38 =10'b0;

   // m34_39 = W*in
   wire signed [9:0] m34_39;
   assign m34_39 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_40 = W*in
   wire signed [9:0] m34_40;
   assign m34_40 =10'b0;

   // m34_41 = W*in
   wire signed [9:0] m34_41;
   assign m34_41 ={ {3{neg34[5]}} , neg34 , {1{1'b0}} };

   // m34_42 = W*in
   wire signed [9:0] m34_42;
   assign m34_42 =10'b0;

   // m34_43 = W*in
   wire signed [9:0] m34_43;
   assign m34_43 =10'b0;

   // m34_44 = W*in
   wire signed [9:0] m34_44;
   assign m34_44 =10'b0;

   // m34_45 = W*in
   wire signed [9:0] m34_45;
   assign m34_45 ={ {2{in34[5]}} , in34 , {2{1'b0}} };

   // m34_46 = W*in
   wire signed [9:0] m34_46;
   assign m34_46 =10'b0;

   // m34_47 = W*in
   wire signed [9:0] m34_47;
   assign m34_47 =10'b0;

   // m34_48 = W*in
   wire signed [9:0] m34_48;
   assign m34_48 =10'b0;

   // m34_49 = W*in
   wire signed [9:0] m34_49;
   assign m34_49 =10'b0;

   // m34_50 = W*in
   wire signed [9:0] m34_50;
   assign m34_50 =10'b0;

   // m34_51 = W*in
   wire signed [9:0] m34_51;
   assign m34_51 =10'b0;

   // m34_52 = W*in
   wire signed [9:0] m34_52;
   assign m34_52 =10'b0;

   // m34_53 = W*in
   wire signed [9:0] m34_53;
   assign m34_53 =10'b0;

   // m34_54 = W*in
   wire signed [9:0] m34_54;
   assign m34_54 =10'b0;

   // m34_55 = W*in
   wire signed [9:0] m34_55;
   assign m34_55 =10'b0;

   // m34_56 = W*in
   wire signed [9:0] m34_56;
   assign m34_56 =10'b0;

   // m34_57 = W*in
   wire signed [9:0] m34_57;
   assign m34_57 =10'b0;

   // m34_58 = W*in
   wire signed [9:0] m34_58;
   assign m34_58 ={ {3{neg34[5]}} , neg34 , {1{1'b0}} };

   // m34_59 = W*in
   wire signed [9:0] m34_59;
   assign m34_59 =10'b0;

   // m34_60 = W*in
   wire signed [9:0] m34_60;
   assign m34_60 =10'b0;

   // m34_61 = W*in
   wire signed [9:0] m34_61;
   assign m34_61 =10'b0;

   // m34_62 = W*in
   wire signed [9:0] m34_62;
   assign m34_62 ={ {3{neg34[5]}} , neg34 , {1{1'b0}} };

   // m34_63 = W*in
   wire signed [9:0] m34_63;
   assign m34_63 =10'b0;

   // m34_64 = W*in
   wire signed [9:0] m34_64;
   assign m34_64 ={ {2{in34[5]}} , in34 , {2{1'b0}} };

   // m34_65 = W*in
   wire signed [9:0] m34_65;
   assign m34_65 =10'b0;

   // m34_66 = W*in
   wire signed [9:0] m34_66;
   assign m34_66 =10'b0;

   // m34_67 = W*in
   wire signed [9:0] m34_67;
   assign m34_67 =10'b0;

   // m34_68 = W*in
   wire signed [9:0] m34_68;
   assign m34_68 =10'b0;

   // m34_69 = W*in
   wire signed [9:0] m34_69;
   assign m34_69 =10'b0;

   // m34_70 = W*in
   wire signed [9:0] m34_70;
   assign m34_70 =10'b0;

   // m34_71 = W*in
   wire signed [9:0] m34_71;
   assign m34_71 =10'b0;

   // m34_72 = W*in
   wire signed [9:0] m34_72;
   assign m34_72 =10'b0;

   // m34_73 = W*in
   wire signed [9:0] m34_73;
   assign m34_73 =10'b0;

   // m34_74 = W*in
   wire signed [9:0] m34_74;
   assign m34_74 =10'b0;

   // m34_75 = W*in
   wire signed [9:0] m34_75;
   assign m34_75 =10'b0;

   // m34_76 = W*in
   wire signed [9:0] m34_76;
   assign m34_76 =10'b0;

   // m34_77 = W*in
   wire signed [9:0] m34_77;
   assign m34_77 =10'b0;

   // m34_78 = W*in
   wire signed [9:0] m34_78;
   assign m34_78 ={ {2{in34[5]}} , in34 , {2{1'b0}} };

   // m34_79 = W*in
   wire signed [9:0] m34_79;
   assign m34_79 ={ {3{in34[5]}} , in34 , {1{1'b0}} };

   // m34_80 = W*in
   wire signed [9:0] m34_80;
   assign m34_80 =10'b0;

   // m34_81 = W*in
   wire signed [9:0] m34_81;
   assign m34_81 =10'b0;

   // m35_1 = W*in
   wire signed [9:0] m35_1;
   assign m35_1 =10'b0;

   // m35_2 = W*in
   wire signed [9:0] m35_2;
   assign m35_2 =10'b0;

   // m35_3 = W*in
   wire signed [9:0] m35_3;
   assign m35_3 =10'b0;

   // m35_4 = W*in
   wire signed [9:0] m35_4;
   assign m35_4 =10'b0;

   // m35_5 = W*in
   wire signed [9:0] m35_5;
   assign m35_5 ={ {3{neg35[5]}} , neg35 , {1{1'b0}} };

   // m35_6 = W*in
   wire signed [9:0] m35_6;
   assign m35_6 =10'b0;

   // m35_7 = W*in
   wire signed [9:0] m35_7;
   assign m35_7 =10'b0;

   // m35_8 = W*in
   wire signed [9:0] m35_8;
   assign m35_8 =10'b0;

   // m35_9 = W*in
   wire signed [9:0] m35_9;
   assign m35_9 =10'b0;

   // m35_10 = W*in
   wire signed [9:0] m35_10;
   assign m35_10 =10'b0;

   // m35_11 = W*in
   wire signed [9:0] m35_11;
   assign m35_11 =10'b0;

   // m35_12 = W*in
   wire signed [9:0] m35_12;
   assign m35_12 =10'b0;

   // m35_13 = W*in
   wire signed [9:0] m35_13;
   assign m35_13 =10'b0;

   // m35_14 = W*in
   wire signed [9:0] m35_14;
   assign m35_14 =10'b0;

   // m35_15 = W*in
   wire signed [9:0] m35_15;
   assign m35_15 ={ {3{in35[5]}} , in35 , {1{1'b0}} };

   // m35_16 = W*in
   wire signed [9:0] m35_16;
   assign m35_16 ={ {3{in35[5]}} , in35 , {1{1'b0}} };

   // m35_17 = W*in
   wire signed [9:0] m35_17;
   assign m35_17 =10'b0;

   // m35_18 = W*in
   wire signed [9:0] m35_18;
   assign m35_18 =10'b0;

   // m35_19 = W*in
   wire signed [9:0] m35_19;
   assign m35_19 ={ {3{neg35[5]}} , neg35 , {1{1'b0}} };

   // m35_20 = W*in
   wire signed [9:0] m35_20;
   assign m35_20 =10'b0;

   // m35_21 = W*in
   wire signed [9:0] m35_21;
   assign m35_21 ={ {3{neg35[5]}} , neg35 , {1{1'b0}} };

   // m35_22 = W*in
   wire signed [9:0] m35_22;
   assign m35_22 =10'b0;

   // m35_23 = W*in
   wire signed [9:0] m35_23;
   assign m35_23 =10'b0;

   // m35_24 = W*in
   wire signed [9:0] m35_24;
   assign m35_24 =10'b0;

   // m35_25 = W*in
   wire signed [9:0] m35_25;
   assign m35_25 =10'b0;

   // m35_26 = W*in
   wire signed [9:0] m35_26;
   assign m35_26 =10'b0;

   // m35_27 = W*in
   wire signed [9:0] m35_27;
   assign m35_27 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_28 = W*in
   wire signed [9:0] m35_28;
   assign m35_28 =10'b0;

   // m35_29 = W*in
   wire signed [9:0] m35_29;
   assign m35_29 =10'b0;

   // m35_30 = W*in
   wire signed [9:0] m35_30;
   assign m35_30 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_31 = W*in
   wire signed [9:0] m35_31;
   assign m35_31 =10'b0;

   // m35_32 = W*in
   wire signed [9:0] m35_32;
   assign m35_32 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_33 = W*in
   wire signed [9:0] m35_33;
   assign m35_33 =10'b0;

   // m35_34 = W*in
   wire signed [9:0] m35_34;
   assign m35_34 =10'b0;

   // m35_35 = W*in
   wire signed [9:0] m35_35;
   assign m35_35 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_36 = W*in
   wire signed [9:0] m35_36;
   assign m35_36 =10'b0;

   // m35_37 = W*in
   wire signed [9:0] m35_37;
   assign m35_37 =10'b0;

   // m35_38 = W*in
   wire signed [9:0] m35_38;
   assign m35_38 =10'b0;

   // m35_39 = W*in
   wire signed [9:0] m35_39;
   assign m35_39 =10'b0;

   // m35_40 = W*in
   wire signed [9:0] m35_40;
   assign m35_40 =10'b0;

   // m35_41 = W*in
   wire signed [9:0] m35_41;
   assign m35_41 =10'b0;

   // m35_42 = W*in
   wire signed [9:0] m35_42;
   assign m35_42 =10'b0;

   // m35_43 = W*in
   wire signed [9:0] m35_43;
   assign m35_43 =10'b0;

   // m35_44 = W*in
   wire signed [9:0] m35_44;
   assign m35_44 =10'b0;

   // m35_45 = W*in
   wire signed [9:0] m35_45;
   assign m35_45 =10'b0;

   // m35_46 = W*in
   wire signed [9:0] m35_46;
   assign m35_46 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_47 = W*in
   wire signed [9:0] m35_47;
   assign m35_47 =10'b0;

   // m35_48 = W*in
   wire signed [9:0] m35_48;
   assign m35_48 =10'b0;

   // m35_49 = W*in
   wire signed [9:0] m35_49;
   assign m35_49 =10'b0;

   // m35_50 = W*in
   wire signed [9:0] m35_50;
   assign m35_50 =10'b0;

   // m35_51 = W*in
   wire signed [9:0] m35_51;
   assign m35_51 =10'b0;

   // m35_52 = W*in
   wire signed [9:0] m35_52;
   assign m35_52 ={ {3{neg35[5]}} , neg35 , {1{1'b0}} };

   // m35_53 = W*in
   wire signed [9:0] m35_53;
   assign m35_53 ={ {3{neg35[5]}} , neg35 , {1{1'b0}} };

   // m35_54 = W*in
   wire signed [9:0] m35_54;
   assign m35_54 =10'b0;

   // m35_55 = W*in
   wire signed [9:0] m35_55;
   assign m35_55 =10'b0;

   // m35_56 = W*in
   wire signed [9:0] m35_56;
   assign m35_56 =10'b0;

   // m35_57 = W*in
   wire signed [9:0] m35_57;
   assign m35_57 =10'b0;

   // m35_58 = W*in
   wire signed [9:0] m35_58;
   assign m35_58 =10'b0;

   // m35_59 = W*in
   wire signed [9:0] m35_59;
   assign m35_59 =10'b0;

   // m35_60 = W*in
   wire signed [9:0] m35_60;
   assign m35_60 =10'b0;

   // m35_61 = W*in
   wire signed [9:0] m35_61;
   assign m35_61 ={ {3{in35[5]}} , in35 , {1{1'b0}} };

   // m35_62 = W*in
   wire signed [9:0] m35_62;
   assign m35_62 ={ {3{in35[5]}} , in35 , {1{1'b0}} };

   // m35_63 = W*in
   wire signed [9:0] m35_63;
   assign m35_63 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_64 = W*in
   wire signed [9:0] m35_64;
   assign m35_64 =10'b0;

   // m35_65 = W*in
   wire signed [9:0] m35_65;
   assign m35_65 =10'b0;

   // m35_66 = W*in
   wire signed [9:0] m35_66;
   assign m35_66 =10'b0;

   // m35_67 = W*in
   wire signed [9:0] m35_67;
   assign m35_67 =10'b0;

   // m35_68 = W*in
   wire signed [9:0] m35_68;
   assign m35_68 =10'b0;

   // m35_69 = W*in
   wire signed [9:0] m35_69;
   assign m35_69 =10'b0;

   // m35_70 = W*in
   wire signed [9:0] m35_70;
   assign m35_70 =10'b0;

   // m35_71 = W*in
   wire signed [9:0] m35_71;
   assign m35_71 =10'b0;

   // m35_72 = W*in
   wire signed [9:0] m35_72;
   assign m35_72 =10'b0;

   // m35_73 = W*in
   wire signed [9:0] m35_73;
   assign m35_73 =10'b0;

   // m35_74 = W*in
   wire signed [9:0] m35_74;
   assign m35_74 =10'b0;

   // m35_75 = W*in
   wire signed [9:0] m35_75;
   assign m35_75 =10'b0;

   // m35_76 = W*in
   wire signed [9:0] m35_76;
   assign m35_76 =10'b0;

   // m35_77 = W*in
   wire signed [9:0] m35_77;
   assign m35_77 ={ {3{neg35[5]}} , neg35 , {1{1'b0}} };

   // m35_78 = W*in
   wire signed [9:0] m35_78;
   assign m35_78 ={ {3{in35[5]}} , in35 , {1{1'b0}} };

   // m35_79 = W*in
   wire signed [9:0] m35_79;
   assign m35_79 ={ {2{in35[5]}} , in35 , {2{1'b0}} };

   // m35_80 = W*in
   wire signed [9:0] m35_80;
   assign m35_80 =10'b0;

   // m35_81 = W*in
   wire signed [9:0] m35_81;
   assign m35_81 =10'b0;

   // m36_1 = W*in
   wire signed [9:0] m36_1;
   assign m36_1 =10'b0;

   // m36_2 = W*in
   wire signed [9:0] m36_2;
   assign m36_2 =10'b0;

   // m36_3 = W*in
   wire signed [9:0] m36_3;
   assign m36_3 =10'b0;

   // m36_4 = W*in
   wire signed [9:0] m36_4;
   assign m36_4 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_5 = W*in
   wire signed [9:0] m36_5;
   assign m36_5 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_6 = W*in
   wire signed [9:0] m36_6;
   assign m36_6 =10'b0;

   // m36_7 = W*in
   wire signed [9:0] m36_7;
   assign m36_7 =10'b0;

   // m36_8 = W*in
   wire signed [9:0] m36_8;
   assign m36_8 =10'b0;

   // m36_9 = W*in
   wire signed [9:0] m36_9;
   assign m36_9 =10'b0;

   // m36_10 = W*in
   wire signed [9:0] m36_10;
   assign m36_10 =10'b0;

   // m36_11 = W*in
   wire signed [9:0] m36_11;
   assign m36_11 =10'b0;

   // m36_12 = W*in
   wire signed [9:0] m36_12;
   assign m36_12 =10'b0;

   // m36_13 = W*in
   wire signed [9:0] m36_13;
   assign m36_13 =10'b0;

   // m36_14 = W*in
   wire signed [9:0] m36_14;
   assign m36_14 =10'b0;

   // m36_15 = W*in
   wire signed [9:0] m36_15;
   assign m36_15 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_16 = W*in
   wire signed [9:0] m36_16;
   assign m36_16 =10'b0;

   // m36_17 = W*in
   wire signed [9:0] m36_17;
   assign m36_17 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_18 = W*in
   wire signed [9:0] m36_18;
   assign m36_18 =10'b0;

   // m36_19 = W*in
   wire signed [9:0] m36_19;
   assign m36_19 =10'b0;

   // m36_20 = W*in
   wire signed [9:0] m36_20;
   assign m36_20 =10'b0;

   // m36_21 = W*in
   wire signed [9:0] m36_21;
   assign m36_21 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_22 = W*in
   wire signed [9:0] m36_22;
   assign m36_22 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_23 = W*in
   wire signed [9:0] m36_23;
   assign m36_23 =10'b0;

   // m36_24 = W*in
   wire signed [9:0] m36_24;
   assign m36_24 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_25 = W*in
   wire signed [9:0] m36_25;
   assign m36_25 =10'b0;

   // m36_26 = W*in
   wire signed [9:0] m36_26;
   assign m36_26 =10'b0;

   // m36_27 = W*in
   wire signed [9:0] m36_27;
   assign m36_27 =10'b0;

   // m36_28 = W*in
   wire signed [9:0] m36_28;
   assign m36_28 =10'b0;

   // m36_29 = W*in
   wire signed [9:0] m36_29;
   assign m36_29 =10'b0;

   // m36_30 = W*in
   wire signed [9:0] m36_30;
   assign m36_30 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_31 = W*in
   wire signed [9:0] m36_31;
   assign m36_31 =10'b0;

   // m36_32 = W*in
   wire signed [9:0] m36_32;
   assign m36_32 =10'b0;

   // m36_33 = W*in
   wire signed [9:0] m36_33;
   assign m36_33 =10'b0;

   // m36_34 = W*in
   wire signed [9:0] m36_34;
   assign m36_34 =10'b0;

   // m36_35 = W*in
   wire signed [9:0] m36_35;
   assign m36_35 =10'b0;

   // m36_36 = W*in
   wire signed [9:0] m36_36;
   assign m36_36 =10'b0;

   // m36_37 = W*in
   wire signed [9:0] m36_37;
   assign m36_37 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_38 = W*in
   wire signed [9:0] m36_38;
   assign m36_38 =10'b0;

   // m36_39 = W*in
   wire signed [9:0] m36_39;
   assign m36_39 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_40 = W*in
   wire signed [9:0] m36_40;
   assign m36_40 =10'b0;

   // m36_41 = W*in
   wire signed [9:0] m36_41;
   assign m36_41 =10'b0;

   // m36_42 = W*in
   wire signed [9:0] m36_42;
   assign m36_42 =10'b0;

   // m36_43 = W*in
   wire signed [9:0] m36_43;
   assign m36_43 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_44 = W*in
   wire signed [9:0] m36_44;
   assign m36_44 ={ {2{in36[5]}} , in36 , {2{1'b0}} };

   // m36_45 = W*in
   wire signed [9:0] m36_45;
   assign m36_45 =10'b0;

   // m36_46 = W*in
   wire signed [9:0] m36_46;
   assign m36_46 =10'b0;

   // m36_47 = W*in
   wire signed [9:0] m36_47;
   assign m36_47 =10'b0;

   // m36_48 = W*in
   wire signed [9:0] m36_48;
   assign m36_48 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_49 = W*in
   wire signed [9:0] m36_49;
   assign m36_49 =10'b0;

   // m36_50 = W*in
   wire signed [9:0] m36_50;
   assign m36_50 =10'b0;

   // m36_51 = W*in
   wire signed [9:0] m36_51;
   assign m36_51 =10'b0;

   // m36_52 = W*in
   wire signed [9:0] m36_52;
   assign m36_52 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_53 = W*in
   wire signed [9:0] m36_53;
   assign m36_53 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_54 = W*in
   wire signed [9:0] m36_54;
   assign m36_54 =10'b0;

   // m36_55 = W*in
   wire signed [9:0] m36_55;
   assign m36_55 =10'b0;

   // m36_56 = W*in
   wire signed [9:0] m36_56;
   assign m36_56 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_57 = W*in
   wire signed [9:0] m36_57;
   assign m36_57 =10'b0;

   // m36_58 = W*in
   wire signed [9:0] m36_58;
   assign m36_58 ={ {2{in36[5]}} , in36 , {2{1'b0}} };

   // m36_59 = W*in
   wire signed [9:0] m36_59;
   assign m36_59 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_60 = W*in
   wire signed [9:0] m36_60;
   assign m36_60 =10'b0;

   // m36_61 = W*in
   wire signed [9:0] m36_61;
   assign m36_61 =10'b0;

   // m36_62 = W*in
   wire signed [9:0] m36_62;
   assign m36_62 ={ {3{in36[5]}} , in36 , {1{1'b0}} };

   // m36_63 = W*in
   wire signed [9:0] m36_63;
   assign m36_63 =10'b0;

   // m36_64 = W*in
   wire signed [9:0] m36_64;
   assign m36_64 =10'b0;

   // m36_65 = W*in
   wire signed [9:0] m36_65;
   assign m36_65 =10'b0;

   // m36_66 = W*in
   wire signed [9:0] m36_66;
   assign m36_66 =10'b0;

   // m36_67 = W*in
   wire signed [9:0] m36_67;
   assign m36_67 =10'b0;

   // m36_68 = W*in
   wire signed [9:0] m36_68;
   assign m36_68 ={ {3{neg36[5]}} , neg36 , {1{1'b0}} };

   // m36_69 = W*in
   wire signed [9:0] m36_69;
   assign m36_69 =10'b0;

   // m36_70 = W*in
   wire signed [9:0] m36_70;
   assign m36_70 =10'b0;

   // m36_71 = W*in
   wire signed [9:0] m36_71;
   assign m36_71 =10'b0;

   // m36_72 = W*in
   wire signed [9:0] m36_72;
   assign m36_72 =10'b0;

   // m36_73 = W*in
   wire signed [9:0] m36_73;
   assign m36_73 =10'b0;

   // m36_74 = W*in
   wire signed [9:0] m36_74;
   assign m36_74 =10'b0;

   // m36_75 = W*in
   wire signed [9:0] m36_75;
   assign m36_75 =10'b0;

   // m36_76 = W*in
   wire signed [9:0] m36_76;
   assign m36_76 =10'b0;

   // m36_77 = W*in
   wire signed [9:0] m36_77;
   assign m36_77 =10'b0;

   // m36_78 = W*in
   wire signed [9:0] m36_78;
   assign m36_78 =10'b0;

   // m36_79 = W*in
   wire signed [9:0] m36_79;
   assign m36_79 =10'b0;

   // m36_80 = W*in
   wire signed [9:0] m36_80;
   assign m36_80 =10'b0;

   // m36_81 = W*in
   wire signed [9:0] m36_81;
   assign m36_81 =10'b0;

   // m37_1 = W*in
   wire signed [9:0] m37_1;
   assign m37_1 =10'b0;

   // m37_2 = W*in
   wire signed [9:0] m37_2;
   assign m37_2 =10'b0;

   // m37_3 = W*in
   wire signed [9:0] m37_3;
   assign m37_3 =10'b0;

   // m37_4 = W*in
   wire signed [9:0] m37_4;
   assign m37_4 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_5 = W*in
   wire signed [9:0] m37_5;
   assign m37_5 =10'b0;

   // m37_6 = W*in
   wire signed [9:0] m37_6;
   assign m37_6 =10'b0;

   // m37_7 = W*in
   wire signed [9:0] m37_7;
   assign m37_7 =10'b0;

   // m37_8 = W*in
   wire signed [9:0] m37_8;
   assign m37_8 =10'b0;

   // m37_9 = W*in
   wire signed [9:0] m37_9;
   assign m37_9 =10'b0;

   // m37_10 = W*in
   wire signed [9:0] m37_10;
   assign m37_10 ={ {2{in37[5]}} , in37 , {2{1'b0}} };

   // m37_11 = W*in
   wire signed [9:0] m37_11;
   assign m37_11 =10'b0;

   // m37_12 = W*in
   wire signed [9:0] m37_12;
   assign m37_12 =10'b0;

   // m37_13 = W*in
   wire signed [9:0] m37_13;
   assign m37_13 =10'b0;

   // m37_14 = W*in
   wire signed [9:0] m37_14;
   assign m37_14 =10'b0;

   // m37_15 = W*in
   wire signed [9:0] m37_15;
   assign m37_15 =10'b0;

   // m37_16 = W*in
   wire signed [9:0] m37_16;
   assign m37_16 =10'b0;

   // m37_17 = W*in
   wire signed [9:0] m37_17;
   assign m37_17 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_18 = W*in
   wire signed [9:0] m37_18;
   assign m37_18 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_19 = W*in
   wire signed [9:0] m37_19;
   assign m37_19 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_20 = W*in
   wire signed [9:0] m37_20;
   assign m37_20 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_21 = W*in
   wire signed [9:0] m37_21;
   assign m37_21 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_22 = W*in
   wire signed [9:0] m37_22;
   assign m37_22 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_23 = W*in
   wire signed [9:0] m37_23;
   assign m37_23 =10'b0;

   // m37_24 = W*in
   wire signed [9:0] m37_24;
   assign m37_24 =10'b0;

   // m37_25 = W*in
   wire signed [9:0] m37_25;
   assign m37_25 =10'b0;

   // m37_26 = W*in
   wire signed [9:0] m37_26;
   assign m37_26 =10'b0;

   // m37_27 = W*in
   wire signed [9:0] m37_27;
   assign m37_27 =10'b0;

   // m37_28 = W*in
   wire signed [9:0] m37_28;
   assign m37_28 =10'b0;

   // m37_29 = W*in
   wire signed [9:0] m37_29;
   assign m37_29 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_30 = W*in
   wire signed [9:0] m37_30;
   assign m37_30 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_31 = W*in
   wire signed [9:0] m37_31;
   assign m37_31 =10'b0;

   // m37_32 = W*in
   wire signed [9:0] m37_32;
   assign m37_32 =10'b0;

   // m37_33 = W*in
   wire signed [9:0] m37_33;
   assign m37_33 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_34 = W*in
   wire signed [9:0] m37_34;
   assign m37_34 =10'b0;

   // m37_35 = W*in
   wire signed [9:0] m37_35;
   assign m37_35 =10'b0;

   // m37_36 = W*in
   wire signed [9:0] m37_36;
   assign m37_36 =10'b0;

   // m37_37 = W*in
   wire signed [9:0] m37_37;
   assign m37_37 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_38 = W*in
   wire signed [9:0] m37_38;
   assign m37_38 =10'b0;

   // m37_39 = W*in
   wire signed [9:0] m37_39;
   assign m37_39 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_40 = W*in
   wire signed [9:0] m37_40;
   assign m37_40 =10'b0;

   // m37_41 = W*in
   wire signed [9:0] m37_41;
   assign m37_41 =10'b0;

   // m37_42 = W*in
   wire signed [9:0] m37_42;
   assign m37_42 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_43 = W*in
   wire signed [9:0] m37_43;
   assign m37_43 =10'b0;

   // m37_44 = W*in
   wire signed [9:0] m37_44;
   assign m37_44 =10'b0;

   // m37_45 = W*in
   wire signed [9:0] m37_45;
   assign m37_45 =10'b0;

   // m37_46 = W*in
   wire signed [9:0] m37_46;
   assign m37_46 =10'b0;

   // m37_47 = W*in
   wire signed [9:0] m37_47;
   assign m37_47 =10'b0;

   // m37_48 = W*in
   wire signed [9:0] m37_48;
   assign m37_48 =10'b0;

   // m37_49 = W*in
   wire signed [9:0] m37_49;
   assign m37_49 =10'b0;

   // m37_50 = W*in
   wire signed [9:0] m37_50;
   assign m37_50 =10'b0;

   // m37_51 = W*in
   wire signed [9:0] m37_51;
   assign m37_51 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_52 = W*in
   wire signed [9:0] m37_52;
   assign m37_52 ={ {2{in37[5]}} , in37 , {2{1'b0}} };

   // m37_53 = W*in
   wire signed [9:0] m37_53;
   assign m37_53 =10'b0;

   // m37_54 = W*in
   wire signed [9:0] m37_54;
   assign m37_54 =10'b0;

   // m37_55 = W*in
   wire signed [9:0] m37_55;
   assign m37_55 =10'b0;

   // m37_56 = W*in
   wire signed [9:0] m37_56;
   assign m37_56 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_57 = W*in
   wire signed [9:0] m37_57;
   assign m37_57 =10'b0;

   // m37_58 = W*in
   wire signed [9:0] m37_58;
   assign m37_58 =10'b0;

   // m37_59 = W*in
   wire signed [9:0] m37_59;
   assign m37_59 =10'b0;

   // m37_60 = W*in
   wire signed [9:0] m37_60;
   assign m37_60 =10'b0;

   // m37_61 = W*in
   wire signed [9:0] m37_61;
   assign m37_61 =10'b0;

   // m37_62 = W*in
   wire signed [9:0] m37_62;
   assign m37_62 =10'b0;

   // m37_63 = W*in
   wire signed [9:0] m37_63;
   assign m37_63 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_64 = W*in
   wire signed [9:0] m37_64;
   assign m37_64 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_65 = W*in
   wire signed [9:0] m37_65;
   assign m37_65 ={ {2{in37[5]}} , in37 , {2{1'b0}} };

   // m37_66 = W*in
   wire signed [9:0] m37_66;
   assign m37_66 =10'b0;

   // m37_67 = W*in
   wire signed [9:0] m37_67;
   assign m37_67 =10'b0;

   // m37_68 = W*in
   wire signed [9:0] m37_68;
   assign m37_68 =10'b0;

   // m37_69 = W*in
   wire signed [9:0] m37_69;
   assign m37_69 =10'b0;

   // m37_70 = W*in
   wire signed [9:0] m37_70;
   assign m37_70 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_71 = W*in
   wire signed [9:0] m37_71;
   assign m37_71 =10'b0;

   // m37_72 = W*in
   wire signed [9:0] m37_72;
   assign m37_72 =10'b0;

   // m37_73 = W*in
   wire signed [9:0] m37_73;
   assign m37_73 =10'b0;

   // m37_74 = W*in
   wire signed [9:0] m37_74;
   assign m37_74 =10'b0;

   // m37_75 = W*in
   wire signed [9:0] m37_75;
   assign m37_75 =10'b0;

   // m37_76 = W*in
   wire signed [9:0] m37_76;
   assign m37_76 =10'b0;

   // m37_77 = W*in
   wire signed [9:0] m37_77;
   assign m37_77 =10'b0;

   // m37_78 = W*in
   wire signed [9:0] m37_78;
   assign m37_78 ={ {3{in37[5]}} , in37 , {1{1'b0}} };

   // m37_79 = W*in
   wire signed [9:0] m37_79;
   assign m37_79 ={ {3{neg37[5]}} , neg37 , {1{1'b0}} };

   // m37_80 = W*in
   wire signed [9:0] m37_80;
   assign m37_80 =10'b0;

   // m37_81 = W*in
   wire signed [9:0] m37_81;
   assign m37_81 =10'b0;

   // m38_1 = W*in
   wire signed [9:0] m38_1;
   assign m38_1 =10'b0;

   // m38_2 = W*in
   wire signed [9:0] m38_2;
   assign m38_2 =10'b0;

   // m38_3 = W*in
   wire signed [9:0] m38_3;
   assign m38_3 =10'b0;

   // m38_4 = W*in
   wire signed [9:0] m38_4;
   assign m38_4 =10'b0;

   // m38_5 = W*in
   wire signed [9:0] m38_5;
   assign m38_5 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_6 = W*in
   wire signed [9:0] m38_6;
   assign m38_6 ={ {2{in38[5]}} , in38 , {2{1'b0}} };

   // m38_7 = W*in
   wire signed [9:0] m38_7;
   assign m38_7 =10'b0;

   // m38_8 = W*in
   wire signed [9:0] m38_8;
   assign m38_8 ={ {2{in38[5]}} , in38 , {2{1'b0}} };

   // m38_9 = W*in
   wire signed [9:0] m38_9;
   assign m38_9 =10'b0;

   // m38_10 = W*in
   wire signed [9:0] m38_10;
   assign m38_10 =10'b0;

   // m38_11 = W*in
   wire signed [9:0] m38_11;
   assign m38_11 =10'b0;

   // m38_12 = W*in
   wire signed [9:0] m38_12;
   assign m38_12 =10'b0;

   // m38_13 = W*in
   wire signed [9:0] m38_13;
   assign m38_13 =10'b0;

   // m38_14 = W*in
   wire signed [9:0] m38_14;
   assign m38_14 =10'b0;

   // m38_15 = W*in
   wire signed [9:0] m38_15;
   assign m38_15 =10'b0;

   // m38_16 = W*in
   wire signed [9:0] m38_16;
   assign m38_16 =10'b0;

   // m38_17 = W*in
   wire signed [9:0] m38_17;
   assign m38_17 ={ {2{in38[5]}} , in38 , {2{1'b0}} };

   // m38_18 = W*in
   wire signed [9:0] m38_18;
   assign m38_18 =10'b0;

   // m38_19 = W*in
   wire signed [9:0] m38_19;
   assign m38_19 =10'b0;

   // m38_20 = W*in
   wire signed [9:0] m38_20;
   assign m38_20 =10'b0;

   // m38_21 = W*in
   wire signed [9:0] m38_21;
   assign m38_21 =10'b0;

   // m38_22 = W*in
   wire signed [9:0] m38_22;
   assign m38_22 =10'b0;

   // m38_23 = W*in
   wire signed [9:0] m38_23;
   assign m38_23 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_24 = W*in
   wire signed [9:0] m38_24;
   assign m38_24 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_25 = W*in
   wire signed [9:0] m38_25;
   assign m38_25 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_26 = W*in
   wire signed [9:0] m38_26;
   assign m38_26 =10'b0;

   // m38_27 = W*in
   wire signed [9:0] m38_27;
   assign m38_27 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_28 = W*in
   wire signed [9:0] m38_28;
   assign m38_28 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_29 = W*in
   wire signed [9:0] m38_29;
   assign m38_29 =10'b0;

   // m38_30 = W*in
   wire signed [9:0] m38_30;
   assign m38_30 =10'b0;

   // m38_31 = W*in
   wire signed [9:0] m38_31;
   assign m38_31 =10'b0;

   // m38_32 = W*in
   wire signed [9:0] m38_32;
   assign m38_32 =10'b0;

   // m38_33 = W*in
   wire signed [9:0] m38_33;
   assign m38_33 ={ {3{in38[5]}} , in38 , {1{1'b0}} };

   // m38_34 = W*in
   wire signed [9:0] m38_34;
   assign m38_34 ={ {2{in38[5]}} , in38 , {2{1'b0}} };

   // m38_35 = W*in
   wire signed [9:0] m38_35;
   assign m38_35 =10'b0;

   // m38_36 = W*in
   wire signed [9:0] m38_36;
   assign m38_36 =10'b0;

   // m38_37 = W*in
   wire signed [9:0] m38_37;
   assign m38_37 =10'b0;

   // m38_38 = W*in
   wire signed [9:0] m38_38;
   assign m38_38 =10'b0;

   // m38_39 = W*in
   wire signed [9:0] m38_39;
   assign m38_39 =10'b0;

   // m38_40 = W*in
   wire signed [9:0] m38_40;
   assign m38_40 =10'b0;

   // m38_41 = W*in
   wire signed [9:0] m38_41;
   assign m38_41 =10'b0;

   // m38_42 = W*in
   wire signed [9:0] m38_42;
   assign m38_42 =10'b0;

   // m38_43 = W*in
   wire signed [9:0] m38_43;
   assign m38_43 =10'b0;

   // m38_44 = W*in
   wire signed [9:0] m38_44;
   assign m38_44 ={ {3{neg38[5]}} , neg38 , {1{1'b0}} };

   // m38_45 = W*in
   wire signed [9:0] m38_45;
   assign m38_45 =10'b0;

   // m38_46 = W*in
   wire signed [9:0] m38_46;
   assign m38_46 =10'b0;

   // m38_47 = W*in
   wire signed [9:0] m38_47;
   assign m38_47 =10'b0;

   // m38_48 = W*in
   wire signed [9:0] m38_48;
   assign m38_48 =10'b0;

   // m38_49 = W*in
   wire signed [9:0] m38_49;
   assign m38_49 =10'b0;

   // m38_50 = W*in
   wire signed [9:0] m38_50;
   assign m38_50 =10'b0;

   // m38_51 = W*in
   wire signed [9:0] m38_51;
   assign m38_51 =10'b0;

   // m38_52 = W*in
   wire signed [9:0] m38_52;
   assign m38_52 =10'b0;

   // m38_53 = W*in
   wire signed [9:0] m38_53;
   assign m38_53 =10'b0;

   // m38_54 = W*in
   wire signed [9:0] m38_54;
   assign m38_54 =10'b0;

   // m38_55 = W*in
   wire signed [9:0] m38_55;
   assign m38_55 =10'b0;

   // m38_56 = W*in
   wire signed [9:0] m38_56;
   assign m38_56 ={ {2{in38[5]}} , in38 , {2{1'b0}} };

   // m38_57 = W*in
   wire signed [9:0] m38_57;
   assign m38_57 =10'b0;

   // m38_58 = W*in
   wire signed [9:0] m38_58;
   assign m38_58 =10'b0;

   // m38_59 = W*in
   wire signed [9:0] m38_59;
   assign m38_59 =10'b0;

   // m38_60 = W*in
   wire signed [9:0] m38_60;
   assign m38_60 =10'b0;

   // m38_61 = W*in
   wire signed [9:0] m38_61;
   assign m38_61 =10'b0;

   // m38_62 = W*in
   wire signed [9:0] m38_62;
   assign m38_62 =10'b0;

   // m38_63 = W*in
   wire signed [9:0] m38_63;
   assign m38_63 ={ {2{in38[5]}} , in38 , {2{1'b0}} };

   // m38_64 = W*in
   wire signed [9:0] m38_64;
   assign m38_64 =10'b0;

   // m38_65 = W*in
   wire signed [9:0] m38_65;
   assign m38_65 =10'b0;

   // m38_66 = W*in
   wire signed [9:0] m38_66;
   assign m38_66 =10'b0;

   // m38_67 = W*in
   wire signed [9:0] m38_67;
   assign m38_67 =10'b0;

   // m38_68 = W*in
   wire signed [9:0] m38_68;
   assign m38_68 =10'b0;

   // m38_69 = W*in
   wire signed [9:0] m38_69;
   assign m38_69 =10'b0;

   // m38_70 = W*in
   wire signed [9:0] m38_70;
   assign m38_70 =10'b0;

   // m38_71 = W*in
   wire signed [9:0] m38_71;
   assign m38_71 =10'b0;

   // m38_72 = W*in
   wire signed [9:0] m38_72;
   assign m38_72 =10'b0;

   // m38_73 = W*in
   wire signed [9:0] m38_73;
   assign m38_73 =10'b0;

   // m38_74 = W*in
   wire signed [9:0] m38_74;
   assign m38_74 =10'b0;

   // m38_75 = W*in
   wire signed [9:0] m38_75;
   assign m38_75 =10'b0;

   // m38_76 = W*in
   wire signed [9:0] m38_76;
   assign m38_76 =10'b0;

   // m38_77 = W*in
   wire signed [9:0] m38_77;
   assign m38_77 =10'b0;

   // m38_78 = W*in
   wire signed [9:0] m38_78;
   assign m38_78 =10'b0;

   // m38_79 = W*in
   wire signed [9:0] m38_79;
   assign m38_79 =10'b0;

   // m38_80 = W*in
   wire signed [9:0] m38_80;
   assign m38_80 =10'b0;

   // m38_81 = W*in
   wire signed [9:0] m38_81;
   assign m38_81 =10'b0;

   // m39_1 = W*in
   wire signed [9:0] m39_1;
   assign m39_1 =10'b0;

   // m39_2 = W*in
   wire signed [9:0] m39_2;
   assign m39_2 =10'b0;

   // m39_3 = W*in
   wire signed [9:0] m39_3;
   assign m39_3 =10'b0;

   // m39_4 = W*in
   wire signed [9:0] m39_4;
   assign m39_4 =10'b0;

   // m39_5 = W*in
   wire signed [9:0] m39_5;
   assign m39_5 =10'b0;

   // m39_6 = W*in
   wire signed [9:0] m39_6;
   assign m39_6 =10'b0;

   // m39_7 = W*in
   wire signed [9:0] m39_7;
   assign m39_7 =10'b0;

   // m39_8 = W*in
   wire signed [9:0] m39_8;
   assign m39_8 =10'b0;

   // m39_9 = W*in
   wire signed [9:0] m39_9;
   assign m39_9 =10'b0;

   // m39_10 = W*in
   wire signed [9:0] m39_10;
   assign m39_10 =10'b0;

   // m39_11 = W*in
   wire signed [9:0] m39_11;
   assign m39_11 =10'b0;

   // m39_12 = W*in
   wire signed [9:0] m39_12;
   assign m39_12 =10'b0;

   // m39_13 = W*in
   wire signed [9:0] m39_13;
   assign m39_13 =10'b0;

   // m39_14 = W*in
   wire signed [9:0] m39_14;
   assign m39_14 =10'b0;

   // m39_15 = W*in
   wire signed [9:0] m39_15;
   assign m39_15 =10'b0;

   // m39_16 = W*in
   wire signed [9:0] m39_16;
   assign m39_16 =10'b0;

   // m39_17 = W*in
   wire signed [9:0] m39_17;
   assign m39_17 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_18 = W*in
   wire signed [9:0] m39_18;
   assign m39_18 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_19 = W*in
   wire signed [9:0] m39_19;
   assign m39_19 =10'b0;

   // m39_20 = W*in
   wire signed [9:0] m39_20;
   assign m39_20 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_21 = W*in
   wire signed [9:0] m39_21;
   assign m39_21 =10'b0;

   // m39_22 = W*in
   wire signed [9:0] m39_22;
   assign m39_22 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_23 = W*in
   wire signed [9:0] m39_23;
   assign m39_23 =10'b0;

   // m39_24 = W*in
   wire signed [9:0] m39_24;
   assign m39_24 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_25 = W*in
   wire signed [9:0] m39_25;
   assign m39_25 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_26 = W*in
   wire signed [9:0] m39_26;
   assign m39_26 =10'b0;

   // m39_27 = W*in
   wire signed [9:0] m39_27;
   assign m39_27 =10'b0;

   // m39_28 = W*in
   wire signed [9:0] m39_28;
   assign m39_28 =10'b0;

   // m39_29 = W*in
   wire signed [9:0] m39_29;
   assign m39_29 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_30 = W*in
   wire signed [9:0] m39_30;
   assign m39_30 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_31 = W*in
   wire signed [9:0] m39_31;
   assign m39_31 =10'b0;

   // m39_32 = W*in
   wire signed [9:0] m39_32;
   assign m39_32 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_33 = W*in
   wire signed [9:0] m39_33;
   assign m39_33 =10'b0;

   // m39_34 = W*in
   wire signed [9:0] m39_34;
   assign m39_34 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_35 = W*in
   wire signed [9:0] m39_35;
   assign m39_35 =10'b0;

   // m39_36 = W*in
   wire signed [9:0] m39_36;
   assign m39_36 =10'b0;

   // m39_37 = W*in
   wire signed [9:0] m39_37;
   assign m39_37 ={ {2{in39[5]}} , in39 , {2{1'b0}} };

   // m39_38 = W*in
   wire signed [9:0] m39_38;
   assign m39_38 =10'b0;

   // m39_39 = W*in
   wire signed [9:0] m39_39;
   assign m39_39 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_40 = W*in
   wire signed [9:0] m39_40;
   assign m39_40 =10'b0;

   // m39_41 = W*in
   wire signed [9:0] m39_41;
   assign m39_41 =10'b0;

   // m39_42 = W*in
   wire signed [9:0] m39_42;
   assign m39_42 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_43 = W*in
   wire signed [9:0] m39_43;
   assign m39_43 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_44 = W*in
   wire signed [9:0] m39_44;
   assign m39_44 =10'b0;

   // m39_45 = W*in
   wire signed [9:0] m39_45;
   assign m39_45 =10'b0;

   // m39_46 = W*in
   wire signed [9:0] m39_46;
   assign m39_46 =10'b0;

   // m39_47 = W*in
   wire signed [9:0] m39_47;
   assign m39_47 =10'b0;

   // m39_48 = W*in
   wire signed [9:0] m39_48;
   assign m39_48 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_49 = W*in
   wire signed [9:0] m39_49;
   assign m39_49 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_50 = W*in
   wire signed [9:0] m39_50;
   assign m39_50 =10'b0;

   // m39_51 = W*in
   wire signed [9:0] m39_51;
   assign m39_51 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_52 = W*in
   wire signed [9:0] m39_52;
   assign m39_52 =10'b0;

   // m39_53 = W*in
   wire signed [9:0] m39_53;
   assign m39_53 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_54 = W*in
   wire signed [9:0] m39_54;
   assign m39_54 =10'b0;

   // m39_55 = W*in
   wire signed [9:0] m39_55;
   assign m39_55 =10'b0;

   // m39_56 = W*in
   wire signed [9:0] m39_56;
   assign m39_56 =10'b0;

   // m39_57 = W*in
   wire signed [9:0] m39_57;
   assign m39_57 =10'b0;

   // m39_58 = W*in
   wire signed [9:0] m39_58;
   assign m39_58 =10'b0;

   // m39_59 = W*in
   wire signed [9:0] m39_59;
   assign m39_59 =10'b0;

   // m39_60 = W*in
   wire signed [9:0] m39_60;
   assign m39_60 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_61 = W*in
   wire signed [9:0] m39_61;
   assign m39_61 =10'b0;

   // m39_62 = W*in
   wire signed [9:0] m39_62;
   assign m39_62 =10'b0;

   // m39_63 = W*in
   wire signed [9:0] m39_63;
   assign m39_63 ={ {3{in39[5]}} , in39 , {1{1'b0}} };

   // m39_64 = W*in
   wire signed [9:0] m39_64;
   assign m39_64 =10'b0;

   // m39_65 = W*in
   wire signed [9:0] m39_65;
   assign m39_65 =10'b0;

   // m39_66 = W*in
   wire signed [9:0] m39_66;
   assign m39_66 =10'b0;

   // m39_67 = W*in
   wire signed [9:0] m39_67;
   assign m39_67 =10'b0;

   // m39_68 = W*in
   wire signed [9:0] m39_68;
   assign m39_68 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_69 = W*in
   wire signed [9:0] m39_69;
   assign m39_69 =10'b0;

   // m39_70 = W*in
   wire signed [9:0] m39_70;
   assign m39_70 =10'b0;

   // m39_71 = W*in
   wire signed [9:0] m39_71;
   assign m39_71 =10'b0;

   // m39_72 = W*in
   wire signed [9:0] m39_72;
   assign m39_72 =10'b0;

   // m39_73 = W*in
   wire signed [9:0] m39_73;
   assign m39_73 =10'b0;

   // m39_74 = W*in
   wire signed [9:0] m39_74;
   assign m39_74 =10'b0;

   // m39_75 = W*in
   wire signed [9:0] m39_75;
   assign m39_75 =10'b0;

   // m39_76 = W*in
   wire signed [9:0] m39_76;
   assign m39_76 =10'b0;

   // m39_77 = W*in
   wire signed [9:0] m39_77;
   assign m39_77 ={ {3{neg39[5]}} , neg39 , {1{1'b0}} };

   // m39_78 = W*in
   wire signed [9:0] m39_78;
   assign m39_78 =10'b0;

   // m39_79 = W*in
   wire signed [9:0] m39_79;
   assign m39_79 =10'b0;

   // m39_80 = W*in
   wire signed [9:0] m39_80;
   assign m39_80 =10'b0;

   // m39_81 = W*in
   wire signed [9:0] m39_81;
   assign m39_81 =10'b0;

   // m40_1 = W*in
   wire signed [9:0] m40_1;
   assign m40_1 =10'b0;

   // m40_2 = W*in
   wire signed [9:0] m40_2;
   assign m40_2 =10'b0;

   // m40_3 = W*in
   wire signed [9:0] m40_3;
   assign m40_3 =10'b0;

   // m40_4 = W*in
   wire signed [9:0] m40_4;
   assign m40_4 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_5 = W*in
   wire signed [9:0] m40_5;
   assign m40_5 =10'b0;

   // m40_6 = W*in
   wire signed [9:0] m40_6;
   assign m40_6 =10'b0;

   // m40_7 = W*in
   wire signed [9:0] m40_7;
   assign m40_7 =10'b0;

   // m40_8 = W*in
   wire signed [9:0] m40_8;
   assign m40_8 =10'b0;

   // m40_9 = W*in
   wire signed [9:0] m40_9;
   assign m40_9 =10'b0;

   // m40_10 = W*in
   wire signed [9:0] m40_10;
   assign m40_10 =10'b0;

   // m40_11 = W*in
   wire signed [9:0] m40_11;
   assign m40_11 =10'b0;

   // m40_12 = W*in
   wire signed [9:0] m40_12;
   assign m40_12 =10'b0;

   // m40_13 = W*in
   wire signed [9:0] m40_13;
   assign m40_13 =10'b0;

   // m40_14 = W*in
   wire signed [9:0] m40_14;
   assign m40_14 =10'b0;

   // m40_15 = W*in
   wire signed [9:0] m40_15;
   assign m40_15 =10'b0;

   // m40_16 = W*in
   wire signed [9:0] m40_16;
   assign m40_16 =10'b0;

   // m40_17 = W*in
   wire signed [9:0] m40_17;
   assign m40_17 =10'b0;

   // m40_18 = W*in
   wire signed [9:0] m40_18;
   assign m40_18 =10'b0;

   // m40_19 = W*in
   wire signed [9:0] m40_19;
   assign m40_19 =10'b0;

   // m40_20 = W*in
   wire signed [9:0] m40_20;
   assign m40_20 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_21 = W*in
   wire signed [9:0] m40_21;
   assign m40_21 =10'b0;

   // m40_22 = W*in
   wire signed [9:0] m40_22;
   assign m40_22 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_23 = W*in
   wire signed [9:0] m40_23;
   assign m40_23 =10'b0;

   // m40_24 = W*in
   wire signed [9:0] m40_24;
   assign m40_24 =10'b0;

   // m40_25 = W*in
   wire signed [9:0] m40_25;
   assign m40_25 =10'b0;

   // m40_26 = W*in
   wire signed [9:0] m40_26;
   assign m40_26 =10'b0;

   // m40_27 = W*in
   wire signed [9:0] m40_27;
   assign m40_27 =10'b0;

   // m40_28 = W*in
   wire signed [9:0] m40_28;
   assign m40_28 =10'b0;

   // m40_29 = W*in
   wire signed [9:0] m40_29;
   assign m40_29 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_30 = W*in
   wire signed [9:0] m40_30;
   assign m40_30 =10'b0;

   // m40_31 = W*in
   wire signed [9:0] m40_31;
   assign m40_31 =10'b0;

   // m40_32 = W*in
   wire signed [9:0] m40_32;
   assign m40_32 =10'b0;

   // m40_33 = W*in
   wire signed [9:0] m40_33;
   assign m40_33 =10'b0;

   // m40_34 = W*in
   wire signed [9:0] m40_34;
   assign m40_34 =10'b0;

   // m40_35 = W*in
   wire signed [9:0] m40_35;
   assign m40_35 =10'b0;

   // m40_36 = W*in
   wire signed [9:0] m40_36;
   assign m40_36 =10'b0;

   // m40_37 = W*in
   wire signed [9:0] m40_37;
   assign m40_37 =10'b0;

   // m40_38 = W*in
   wire signed [9:0] m40_38;
   assign m40_38 =10'b0;

   // m40_39 = W*in
   wire signed [9:0] m40_39;
   assign m40_39 =10'b0;

   // m40_40 = W*in
   wire signed [9:0] m40_40;
   assign m40_40 =10'b0;

   // m40_41 = W*in
   wire signed [9:0] m40_41;
   assign m40_41 =10'b0;

   // m40_42 = W*in
   wire signed [9:0] m40_42;
   assign m40_42 =10'b0;

   // m40_43 = W*in
   wire signed [9:0] m40_43;
   assign m40_43 =10'b0;

   // m40_44 = W*in
   wire signed [9:0] m40_44;
   assign m40_44 =10'b0;

   // m40_45 = W*in
   wire signed [9:0] m40_45;
   assign m40_45 =10'b0;

   // m40_46 = W*in
   wire signed [9:0] m40_46;
   assign m40_46 =10'b0;

   // m40_47 = W*in
   wire signed [9:0] m40_47;
   assign m40_47 =10'b0;

   // m40_48 = W*in
   wire signed [9:0] m40_48;
   assign m40_48 =10'b0;

   // m40_49 = W*in
   wire signed [9:0] m40_49;
   assign m40_49 =10'b0;

   // m40_50 = W*in
   wire signed [9:0] m40_50;
   assign m40_50 =10'b0;

   // m40_51 = W*in
   wire signed [9:0] m40_51;
   assign m40_51 =10'b0;

   // m40_52 = W*in
   wire signed [9:0] m40_52;
   assign m40_52 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_53 = W*in
   wire signed [9:0] m40_53;
   assign m40_53 =10'b0;

   // m40_54 = W*in
   wire signed [9:0] m40_54;
   assign m40_54 =10'b0;

   // m40_55 = W*in
   wire signed [9:0] m40_55;
   assign m40_55 =10'b0;

   // m40_56 = W*in
   wire signed [9:0] m40_56;
   assign m40_56 =10'b0;

   // m40_57 = W*in
   wire signed [9:0] m40_57;
   assign m40_57 =10'b0;

   // m40_58 = W*in
   wire signed [9:0] m40_58;
   assign m40_58 =10'b0;

   // m40_59 = W*in
   wire signed [9:0] m40_59;
   assign m40_59 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_60 = W*in
   wire signed [9:0] m40_60;
   assign m40_60 =10'b0;

   // m40_61 = W*in
   wire signed [9:0] m40_61;
   assign m40_61 =10'b0;

   // m40_62 = W*in
   wire signed [9:0] m40_62;
   assign m40_62 =10'b0;

   // m40_63 = W*in
   wire signed [9:0] m40_63;
   assign m40_63 =10'b0;

   // m40_64 = W*in
   wire signed [9:0] m40_64;
   assign m40_64 =10'b0;

   // m40_65 = W*in
   wire signed [9:0] m40_65;
   assign m40_65 =10'b0;

   // m40_66 = W*in
   wire signed [9:0] m40_66;
   assign m40_66 =10'b0;

   // m40_67 = W*in
   wire signed [9:0] m40_67;
   assign m40_67 =10'b0;

   // m40_68 = W*in
   wire signed [9:0] m40_68;
   assign m40_68 =10'b0;

   // m40_69 = W*in
   wire signed [9:0] m40_69;
   assign m40_69 =10'b0;

   // m40_70 = W*in
   wire signed [9:0] m40_70;
   assign m40_70 =10'b0;

   // m40_71 = W*in
   wire signed [9:0] m40_71;
   assign m40_71 =10'b0;

   // m40_72 = W*in
   wire signed [9:0] m40_72;
   assign m40_72 =10'b0;

   // m40_73 = W*in
   wire signed [9:0] m40_73;
   assign m40_73 =10'b0;

   // m40_74 = W*in
   wire signed [9:0] m40_74;
   assign m40_74 =10'b0;

   // m40_75 = W*in
   wire signed [9:0] m40_75;
   assign m40_75 =10'b0;

   // m40_76 = W*in
   wire signed [9:0] m40_76;
   assign m40_76 =10'b0;

   // m40_77 = W*in
   wire signed [9:0] m40_77;
   assign m40_77 ={ {3{in40[5]}} , in40 , {1{1'b0}} };

   // m40_78 = W*in
   wire signed [9:0] m40_78;
   assign m40_78 =10'b0;

   // m40_79 = W*in
   wire signed [9:0] m40_79;
   assign m40_79 =10'b0;

   // m40_80 = W*in
   wire signed [9:0] m40_80;
   assign m40_80 =10'b0;

   // m40_81 = W*in
   wire signed [9:0] m40_81;
   assign m40_81 =10'b0;

   // m41_1 = W*in
   wire signed [9:0] m41_1;
   assign m41_1 =10'b0;

   // m41_2 = W*in
   wire signed [9:0] m41_2;
   assign m41_2 =10'b0;

   // m41_3 = W*in
   wire signed [9:0] m41_3;
   assign m41_3 ={ {2{in41[5]}} , in41 , {2{1'b0}} };

   // m41_4 = W*in
   wire signed [9:0] m41_4;
   assign m41_4 =10'b0;

   // m41_5 = W*in
   wire signed [9:0] m41_5;
   assign m41_5 =10'b0;

   // m41_6 = W*in
   wire signed [9:0] m41_6;
   assign m41_6 =10'b0;

   // m41_7 = W*in
   wire signed [9:0] m41_7;
   assign m41_7 =10'b0;

   // m41_8 = W*in
   wire signed [9:0] m41_8;
   assign m41_8 =10'b0;

   // m41_9 = W*in
   wire signed [9:0] m41_9;
   assign m41_9 =10'b0;

   // m41_10 = W*in
   wire signed [9:0] m41_10;
   assign m41_10 =10'b0;

   // m41_11 = W*in
   wire signed [9:0] m41_11;
   assign m41_11 =10'b0;

   // m41_12 = W*in
   wire signed [9:0] m41_12;
   assign m41_12 =10'b0;

   // m41_13 = W*in
   wire signed [9:0] m41_13;
   assign m41_13 =10'b0;

   // m41_14 = W*in
   wire signed [9:0] m41_14;
   assign m41_14 =10'b0;

   // m41_15 = W*in
   wire signed [9:0] m41_15;
   assign m41_15 =10'b0;

   // m41_16 = W*in
   wire signed [9:0] m41_16;
   assign m41_16 =10'b0;

   // m41_17 = W*in
   wire signed [9:0] m41_17;
   assign m41_17 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_18 = W*in
   wire signed [9:0] m41_18;
   assign m41_18 =10'b0;

   // m41_19 = W*in
   wire signed [9:0] m41_19;
   assign m41_19 =10'b0;

   // m41_20 = W*in
   wire signed [9:0] m41_20;
   assign m41_20 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_21 = W*in
   wire signed [9:0] m41_21;
   assign m41_21 =10'b0;

   // m41_22 = W*in
   wire signed [9:0] m41_22;
   assign m41_22 =10'b0;

   // m41_23 = W*in
   wire signed [9:0] m41_23;
   assign m41_23 =10'b0;

   // m41_24 = W*in
   wire signed [9:0] m41_24;
   assign m41_24 =10'b0;

   // m41_25 = W*in
   wire signed [9:0] m41_25;
   assign m41_25 =10'b0;

   // m41_26 = W*in
   wire signed [9:0] m41_26;
   assign m41_26 =10'b0;

   // m41_27 = W*in
   wire signed [9:0] m41_27;
   assign m41_27 =10'b0;

   // m41_28 = W*in
   wire signed [9:0] m41_28;
   assign m41_28 =10'b0;

   // m41_29 = W*in
   wire signed [9:0] m41_29;
   assign m41_29 =10'b0;

   // m41_30 = W*in
   wire signed [9:0] m41_30;
   assign m41_30 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_31 = W*in
   wire signed [9:0] m41_31;
   assign m41_31 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_32 = W*in
   wire signed [9:0] m41_32;
   assign m41_32 =10'b0;

   // m41_33 = W*in
   wire signed [9:0] m41_33;
   assign m41_33 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_34 = W*in
   wire signed [9:0] m41_34;
   assign m41_34 =10'b0;

   // m41_35 = W*in
   wire signed [9:0] m41_35;
   assign m41_35 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_36 = W*in
   wire signed [9:0] m41_36;
   assign m41_36 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_37 = W*in
   wire signed [9:0] m41_37;
   assign m41_37 =10'b0;

   // m41_38 = W*in
   wire signed [9:0] m41_38;
   assign m41_38 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_39 = W*in
   wire signed [9:0] m41_39;
   assign m41_39 =10'b0;

   // m41_40 = W*in
   wire signed [9:0] m41_40;
   assign m41_40 =10'b0;

   // m41_41 = W*in
   wire signed [9:0] m41_41;
   assign m41_41 =10'b0;

   // m41_42 = W*in
   wire signed [9:0] m41_42;
   assign m41_42 =10'b0;

   // m41_43 = W*in
   wire signed [9:0] m41_43;
   assign m41_43 =10'b0;

   // m41_44 = W*in
   wire signed [9:0] m41_44;
   assign m41_44 =10'b0;

   // m41_45 = W*in
   wire signed [9:0] m41_45;
   assign m41_45 =10'b0;

   // m41_46 = W*in
   wire signed [9:0] m41_46;
   assign m41_46 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_47 = W*in
   wire signed [9:0] m41_47;
   assign m41_47 =10'b0;

   // m41_48 = W*in
   wire signed [9:0] m41_48;
   assign m41_48 =10'b0;

   // m41_49 = W*in
   wire signed [9:0] m41_49;
   assign m41_49 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_50 = W*in
   wire signed [9:0] m41_50;
   assign m41_50 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_51 = W*in
   wire signed [9:0] m41_51;
   assign m41_51 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_52 = W*in
   wire signed [9:0] m41_52;
   assign m41_52 =10'b0;

   // m41_53 = W*in
   wire signed [9:0] m41_53;
   assign m41_53 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_54 = W*in
   wire signed [9:0] m41_54;
   assign m41_54 =10'b0;

   // m41_55 = W*in
   wire signed [9:0] m41_55;
   assign m41_55 =10'b0;

   // m41_56 = W*in
   wire signed [9:0] m41_56;
   assign m41_56 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_57 = W*in
   wire signed [9:0] m41_57;
   assign m41_57 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_58 = W*in
   wire signed [9:0] m41_58;
   assign m41_58 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_59 = W*in
   wire signed [9:0] m41_59;
   assign m41_59 =10'b0;

   // m41_60 = W*in
   wire signed [9:0] m41_60;
   assign m41_60 =10'b0;

   // m41_61 = W*in
   wire signed [9:0] m41_61;
   assign m41_61 =10'b0;

   // m41_62 = W*in
   wire signed [9:0] m41_62;
   assign m41_62 =10'b0;

   // m41_63 = W*in
   wire signed [9:0] m41_63;
   assign m41_63 =10'b0;

   // m41_64 = W*in
   wire signed [9:0] m41_64;
   assign m41_64 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_65 = W*in
   wire signed [9:0] m41_65;
   assign m41_65 =10'b0;

   // m41_66 = W*in
   wire signed [9:0] m41_66;
   assign m41_66 =10'b0;

   // m41_67 = W*in
   wire signed [9:0] m41_67;
   assign m41_67 =10'b0;

   // m41_68 = W*in
   wire signed [9:0] m41_68;
   assign m41_68 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_69 = W*in
   wire signed [9:0] m41_69;
   assign m41_69 ={ {3{neg41[5]}} , neg41 , {1{1'b0}} };

   // m41_70 = W*in
   wire signed [9:0] m41_70;
   assign m41_70 =10'b0;

   // m41_71 = W*in
   wire signed [9:0] m41_71;
   assign m41_71 =10'b0;

   // m41_72 = W*in
   wire signed [9:0] m41_72;
   assign m41_72 =10'b0;

   // m41_73 = W*in
   wire signed [9:0] m41_73;
   assign m41_73 =10'b0;

   // m41_74 = W*in
   wire signed [9:0] m41_74;
   assign m41_74 =10'b0;

   // m41_75 = W*in
   wire signed [9:0] m41_75;
   assign m41_75 =10'b0;

   // m41_76 = W*in
   wire signed [9:0] m41_76;
   assign m41_76 =10'b0;

   // m41_77 = W*in
   wire signed [9:0] m41_77;
   assign m41_77 =10'b0;

   // m41_78 = W*in
   wire signed [9:0] m41_78;
   assign m41_78 ={ {2{in41[5]}} , in41 , {2{1'b0}} };

   // m41_79 = W*in
   wire signed [9:0] m41_79;
   assign m41_79 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_80 = W*in
   wire signed [9:0] m41_80;
   assign m41_80 =10'b0;

   // m41_81 = W*in
   wire signed [9:0] m41_81;
   assign m41_81 =10'b0;

   // m42_1 = W*in
   wire signed [9:0] m42_1;
   assign m42_1 ={ {2{in42[5]}} , in42 , {2{1'b0}} };

   // m42_2 = W*in
   wire signed [9:0] m42_2;
   assign m42_2 =10'b0;

   // m42_3 = W*in
   wire signed [9:0] m42_3;
   assign m42_3 =10'b0;

   // m42_4 = W*in
   wire signed [9:0] m42_4;
   assign m42_4 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_5 = W*in
   wire signed [9:0] m42_5;
   assign m42_5 =10'b0;

   // m42_6 = W*in
   wire signed [9:0] m42_6;
   assign m42_6 =10'b0;

   // m42_7 = W*in
   wire signed [9:0] m42_7;
   assign m42_7 =10'b0;

   // m42_8 = W*in
   wire signed [9:0] m42_8;
   assign m42_8 =10'b0;

   // m42_9 = W*in
   wire signed [9:0] m42_9;
   assign m42_9 =10'b0;

   // m42_10 = W*in
   wire signed [9:0] m42_10;
   assign m42_10 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_11 = W*in
   wire signed [9:0] m42_11;
   assign m42_11 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_12 = W*in
   wire signed [9:0] m42_12;
   assign m42_12 =10'b0;

   // m42_13 = W*in
   wire signed [9:0] m42_13;
   assign m42_13 =10'b0;

   // m42_14 = W*in
   wire signed [9:0] m42_14;
   assign m42_14 =10'b0;

   // m42_15 = W*in
   wire signed [9:0] m42_15;
   assign m42_15 =10'b0;

   // m42_16 = W*in
   wire signed [9:0] m42_16;
   assign m42_16 =10'b0;

   // m42_17 = W*in
   wire signed [9:0] m42_17;
   assign m42_17 =10'b0;

   // m42_18 = W*in
   wire signed [9:0] m42_18;
   assign m42_18 ={ {2{in42[5]}} , in42 , {2{1'b0}} };

   // m42_19 = W*in
   wire signed [9:0] m42_19;
   assign m42_19 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_20 = W*in
   wire signed [9:0] m42_20;
   assign m42_20 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_21 = W*in
   wire signed [9:0] m42_21;
   assign m42_21 =10'b0;

   // m42_22 = W*in
   wire signed [9:0] m42_22;
   assign m42_22 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_23 = W*in
   wire signed [9:0] m42_23;
   assign m42_23 =10'b0;

   // m42_24 = W*in
   wire signed [9:0] m42_24;
   assign m42_24 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_25 = W*in
   wire signed [9:0] m42_25;
   assign m42_25 =10'b0;

   // m42_26 = W*in
   wire signed [9:0] m42_26;
   assign m42_26 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_27 = W*in
   wire signed [9:0] m42_27;
   assign m42_27 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_28 = W*in
   wire signed [9:0] m42_28;
   assign m42_28 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_29 = W*in
   wire signed [9:0] m42_29;
   assign m42_29 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_30 = W*in
   wire signed [9:0] m42_30;
   assign m42_30 =10'b0;

   // m42_31 = W*in
   wire signed [9:0] m42_31;
   assign m42_31 =10'b0;

   // m42_32 = W*in
   wire signed [9:0] m42_32;
   assign m42_32 =10'b0;

   // m42_33 = W*in
   wire signed [9:0] m42_33;
   assign m42_33 =10'b0;

   // m42_34 = W*in
   wire signed [9:0] m42_34;
   assign m42_34 =10'b0;

   // m42_35 = W*in
   wire signed [9:0] m42_35;
   assign m42_35 =10'b0;

   // m42_36 = W*in
   wire signed [9:0] m42_36;
   assign m42_36 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_37 = W*in
   wire signed [9:0] m42_37;
   assign m42_37 =10'b0;

   // m42_38 = W*in
   wire signed [9:0] m42_38;
   assign m42_38 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_39 = W*in
   wire signed [9:0] m42_39;
   assign m42_39 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_40 = W*in
   wire signed [9:0] m42_40;
   assign m42_40 =10'b0;

   // m42_41 = W*in
   wire signed [9:0] m42_41;
   assign m42_41 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_42 = W*in
   wire signed [9:0] m42_42;
   assign m42_42 ={ {2{in42[5]}} , in42 , {2{1'b0}} };

   // m42_43 = W*in
   wire signed [9:0] m42_43;
   assign m42_43 =10'b0;

   // m42_44 = W*in
   wire signed [9:0] m42_44;
   assign m42_44 =10'b0;

   // m42_45 = W*in
   wire signed [9:0] m42_45;
   assign m42_45 =10'b0;

   // m42_46 = W*in
   wire signed [9:0] m42_46;
   assign m42_46 =10'b0;

   // m42_47 = W*in
   wire signed [9:0] m42_47;
   assign m42_47 =10'b0;

   // m42_48 = W*in
   wire signed [9:0] m42_48;
   assign m42_48 =10'b0;

   // m42_49 = W*in
   wire signed [9:0] m42_49;
   assign m42_49 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_50 = W*in
   wire signed [9:0] m42_50;
   assign m42_50 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_51 = W*in
   wire signed [9:0] m42_51;
   assign m42_51 =10'b0;

   // m42_52 = W*in
   wire signed [9:0] m42_52;
   assign m42_52 =10'b0;

   // m42_53 = W*in
   wire signed [9:0] m42_53;
   assign m42_53 =10'b0;

   // m42_54 = W*in
   wire signed [9:0] m42_54;
   assign m42_54 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_55 = W*in
   wire signed [9:0] m42_55;
   assign m42_55 =10'b0;

   // m42_56 = W*in
   wire signed [9:0] m42_56;
   assign m42_56 =10'b0;

   // m42_57 = W*in
   wire signed [9:0] m42_57;
   assign m42_57 =10'b0;

   // m42_58 = W*in
   wire signed [9:0] m42_58;
   assign m42_58 =10'b0;

   // m42_59 = W*in
   wire signed [9:0] m42_59;
   assign m42_59 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_60 = W*in
   wire signed [9:0] m42_60;
   assign m42_60 =10'b0;

   // m42_61 = W*in
   wire signed [9:0] m42_61;
   assign m42_61 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_62 = W*in
   wire signed [9:0] m42_62;
   assign m42_62 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_63 = W*in
   wire signed [9:0] m42_63;
   assign m42_63 =10'b0;

   // m42_64 = W*in
   wire signed [9:0] m42_64;
   assign m42_64 =10'b0;

   // m42_65 = W*in
   wire signed [9:0] m42_65;
   assign m42_65 =10'b0;

   // m42_66 = W*in
   wire signed [9:0] m42_66;
   assign m42_66 =10'b0;

   // m42_67 = W*in
   wire signed [9:0] m42_67;
   assign m42_67 =10'b0;

   // m42_68 = W*in
   wire signed [9:0] m42_68;
   assign m42_68 ={ {3{in42[5]}} , in42 , {1{1'b0}} };

   // m42_69 = W*in
   wire signed [9:0] m42_69;
   assign m42_69 =10'b0;

   // m42_70 = W*in
   wire signed [9:0] m42_70;
   assign m42_70 =10'b0;

   // m42_71 = W*in
   wire signed [9:0] m42_71;
   assign m42_71 =10'b0;

   // m42_72 = W*in
   wire signed [9:0] m42_72;
   assign m42_72 =10'b0;

   // m42_73 = W*in
   wire signed [9:0] m42_73;
   assign m42_73 =10'b0;

   // m42_74 = W*in
   wire signed [9:0] m42_74;
   assign m42_74 =10'b0;

   // m42_75 = W*in
   wire signed [9:0] m42_75;
   assign m42_75 =10'b0;

   // m42_76 = W*in
   wire signed [9:0] m42_76;
   assign m42_76 =10'b0;

   // m42_77 = W*in
   wire signed [9:0] m42_77;
   assign m42_77 =10'b0;

   // m42_78 = W*in
   wire signed [9:0] m42_78;
   assign m42_78 =10'b0;

   // m42_79 = W*in
   wire signed [9:0] m42_79;
   assign m42_79 =10'b0;

   // m42_80 = W*in
   wire signed [9:0] m42_80;
   assign m42_80 =10'b0;

   // m42_81 = W*in
   wire signed [9:0] m42_81;
   assign m42_81 =10'b0;

   // m43_1 = W*in
   wire signed [9:0] m43_1;
   assign m43_1 =10'b0;

   // m43_2 = W*in
   wire signed [9:0] m43_2;
   assign m43_2 =10'b0;

   // m43_3 = W*in
   wire signed [9:0] m43_3;
   assign m43_3 =10'b0;

   // m43_4 = W*in
   wire signed [9:0] m43_4;
   assign m43_4 =10'b0;

   // m43_5 = W*in
   wire signed [9:0] m43_5;
   assign m43_5 =10'b0;

   // m43_6 = W*in
   wire signed [9:0] m43_6;
   assign m43_6 =10'b0;

   // m43_7 = W*in
   wire signed [9:0] m43_7;
   assign m43_7 =10'b0;

   // m43_8 = W*in
   wire signed [9:0] m43_8;
   assign m43_8 ={ {2{in43[5]}} , in43 , {2{1'b0}} };

   // m43_9 = W*in
   wire signed [9:0] m43_9;
   assign m43_9 =10'b0;

   // m43_10 = W*in
   wire signed [9:0] m43_10;
   assign m43_10 =10'b0;

   // m43_11 = W*in
   wire signed [9:0] m43_11;
   assign m43_11 =10'b0;

   // m43_12 = W*in
   wire signed [9:0] m43_12;
   assign m43_12 =10'b0;

   // m43_13 = W*in
   wire signed [9:0] m43_13;
   assign m43_13 =10'b0;

   // m43_14 = W*in
   wire signed [9:0] m43_14;
   assign m43_14 =10'b0;

   // m43_15 = W*in
   wire signed [9:0] m43_15;
   assign m43_15 =10'b0;

   // m43_16 = W*in
   wire signed [9:0] m43_16;
   assign m43_16 =10'b0;

   // m43_17 = W*in
   wire signed [9:0] m43_17;
   assign m43_17 =10'b0;

   // m43_18 = W*in
   wire signed [9:0] m43_18;
   assign m43_18 =10'b0;

   // m43_19 = W*in
   wire signed [9:0] m43_19;
   assign m43_19 =10'b0;

   // m43_20 = W*in
   wire signed [9:0] m43_20;
   assign m43_20 =10'b0;

   // m43_21 = W*in
   wire signed [9:0] m43_21;
   assign m43_21 =10'b0;

   // m43_22 = W*in
   wire signed [9:0] m43_22;
   assign m43_22 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_23 = W*in
   wire signed [9:0] m43_23;
   assign m43_23 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_24 = W*in
   wire signed [9:0] m43_24;
   assign m43_24 =10'b0;

   // m43_25 = W*in
   wire signed [9:0] m43_25;
   assign m43_25 ={ {2{in43[5]}} , in43 , {2{1'b0}} };

   // m43_26 = W*in
   wire signed [9:0] m43_26;
   assign m43_26 =10'b0;

   // m43_27 = W*in
   wire signed [9:0] m43_27;
   assign m43_27 =10'b0;

   // m43_28 = W*in
   wire signed [9:0] m43_28;
   assign m43_28 =10'b0;

   // m43_29 = W*in
   wire signed [9:0] m43_29;
   assign m43_29 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_30 = W*in
   wire signed [9:0] m43_30;
   assign m43_30 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_31 = W*in
   wire signed [9:0] m43_31;
   assign m43_31 =10'b0;

   // m43_32 = W*in
   wire signed [9:0] m43_32;
   assign m43_32 =10'b0;

   // m43_33 = W*in
   wire signed [9:0] m43_33;
   assign m43_33 ={ {2{in43[5]}} , in43 , {2{1'b0}} };

   // m43_34 = W*in
   wire signed [9:0] m43_34;
   assign m43_34 =10'b0;

   // m43_35 = W*in
   wire signed [9:0] m43_35;
   assign m43_35 =10'b0;

   // m43_36 = W*in
   wire signed [9:0] m43_36;
   assign m43_36 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_37 = W*in
   wire signed [9:0] m43_37;
   assign m43_37 =10'b0;

   // m43_38 = W*in
   wire signed [9:0] m43_38;
   assign m43_38 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_39 = W*in
   wire signed [9:0] m43_39;
   assign m43_39 =10'b0;

   // m43_40 = W*in
   wire signed [9:0] m43_40;
   assign m43_40 =10'b0;

   // m43_41 = W*in
   wire signed [9:0] m43_41;
   assign m43_41 =10'b0;

   // m43_42 = W*in
   wire signed [9:0] m43_42;
   assign m43_42 =10'b0;

   // m43_43 = W*in
   wire signed [9:0] m43_43;
   assign m43_43 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_44 = W*in
   wire signed [9:0] m43_44;
   assign m43_44 =10'b0;

   // m43_45 = W*in
   wire signed [9:0] m43_45;
   assign m43_45 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_46 = W*in
   wire signed [9:0] m43_46;
   assign m43_46 =10'b0;

   // m43_47 = W*in
   wire signed [9:0] m43_47;
   assign m43_47 =10'b0;

   // m43_48 = W*in
   wire signed [9:0] m43_48;
   assign m43_48 =10'b0;

   // m43_49 = W*in
   wire signed [9:0] m43_49;
   assign m43_49 =10'b0;

   // m43_50 = W*in
   wire signed [9:0] m43_50;
   assign m43_50 =10'b0;

   // m43_51 = W*in
   wire signed [9:0] m43_51;
   assign m43_51 =10'b0;

   // m43_52 = W*in
   wire signed [9:0] m43_52;
   assign m43_52 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_53 = W*in
   wire signed [9:0] m43_53;
   assign m43_53 =10'b0;

   // m43_54 = W*in
   wire signed [9:0] m43_54;
   assign m43_54 =10'b0;

   // m43_55 = W*in
   wire signed [9:0] m43_55;
   assign m43_55 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_56 = W*in
   wire signed [9:0] m43_56;
   assign m43_56 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_57 = W*in
   wire signed [9:0] m43_57;
   assign m43_57 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_58 = W*in
   wire signed [9:0] m43_58;
   assign m43_58 =10'b0;

   // m43_59 = W*in
   wire signed [9:0] m43_59;
   assign m43_59 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_60 = W*in
   wire signed [9:0] m43_60;
   assign m43_60 =10'b0;

   // m43_61 = W*in
   wire signed [9:0] m43_61;
   assign m43_61 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_62 = W*in
   wire signed [9:0] m43_62;
   assign m43_62 ={ {3{in43[5]}} , in43 , {1{1'b0}} };

   // m43_63 = W*in
   wire signed [9:0] m43_63;
   assign m43_63 =10'b0;

   // m43_64 = W*in
   wire signed [9:0] m43_64;
   assign m43_64 =10'b0;

   // m43_65 = W*in
   wire signed [9:0] m43_65;
   assign m43_65 =10'b0;

   // m43_66 = W*in
   wire signed [9:0] m43_66;
   assign m43_66 =10'b0;

   // m43_67 = W*in
   wire signed [9:0] m43_67;
   assign m43_67 =10'b0;

   // m43_68 = W*in
   wire signed [9:0] m43_68;
   assign m43_68 =10'b0;

   // m43_69 = W*in
   wire signed [9:0] m43_69;
   assign m43_69 =10'b0;

   // m43_70 = W*in
   wire signed [9:0] m43_70;
   assign m43_70 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_71 = W*in
   wire signed [9:0] m43_71;
   assign m43_71 =10'b0;

   // m43_72 = W*in
   wire signed [9:0] m43_72;
   assign m43_72 =10'b0;

   // m43_73 = W*in
   wire signed [9:0] m43_73;
   assign m43_73 =10'b0;

   // m43_74 = W*in
   wire signed [9:0] m43_74;
   assign m43_74 =10'b0;

   // m43_75 = W*in
   wire signed [9:0] m43_75;
   assign m43_75 =10'b0;

   // m43_76 = W*in
   wire signed [9:0] m43_76;
   assign m43_76 =10'b0;

   // m43_77 = W*in
   wire signed [9:0] m43_77;
   assign m43_77 =10'b0;

   // m43_78 = W*in
   wire signed [9:0] m43_78;
   assign m43_78 ={ {3{neg43[5]}} , neg43 , {1{1'b0}} };

   // m43_79 = W*in
   wire signed [9:0] m43_79;
   assign m43_79 =10'b0;

   // m43_80 = W*in
   wire signed [9:0] m43_80;
   assign m43_80 =10'b0;

   // m43_81 = W*in
   wire signed [9:0] m43_81;
   assign m43_81 =10'b0;

   // m44_1 = W*in
   wire signed [9:0] m44_1;
   assign m44_1 =10'b0;

   // m44_2 = W*in
   wire signed [9:0] m44_2;
   assign m44_2 =10'b0;

   // m44_3 = W*in
   wire signed [9:0] m44_3;
   assign m44_3 =10'b0;

   // m44_4 = W*in
   wire signed [9:0] m44_4;
   assign m44_4 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_5 = W*in
   wire signed [9:0] m44_5;
   assign m44_5 =10'b0;

   // m44_6 = W*in
   wire signed [9:0] m44_6;
   assign m44_6 =10'b0;

   // m44_7 = W*in
   wire signed [9:0] m44_7;
   assign m44_7 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_8 = W*in
   wire signed [9:0] m44_8;
   assign m44_8 =10'b0;

   // m44_9 = W*in
   wire signed [9:0] m44_9;
   assign m44_9 =10'b0;

   // m44_10 = W*in
   wire signed [9:0] m44_10;
   assign m44_10 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_11 = W*in
   wire signed [9:0] m44_11;
   assign m44_11 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_12 = W*in
   wire signed [9:0] m44_12;
   assign m44_12 =10'b0;

   // m44_13 = W*in
   wire signed [9:0] m44_13;
   assign m44_13 =10'b0;

   // m44_14 = W*in
   wire signed [9:0] m44_14;
   assign m44_14 =10'b0;

   // m44_15 = W*in
   wire signed [9:0] m44_15;
   assign m44_15 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_16 = W*in
   wire signed [9:0] m44_16;
   assign m44_16 =10'b0;

   // m44_17 = W*in
   wire signed [9:0] m44_17;
   assign m44_17 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_18 = W*in
   wire signed [9:0] m44_18;
   assign m44_18 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_19 = W*in
   wire signed [9:0] m44_19;
   assign m44_19 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_20 = W*in
   wire signed [9:0] m44_20;
   assign m44_20 =10'b0;

   // m44_21 = W*in
   wire signed [9:0] m44_21;
   assign m44_21 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_22 = W*in
   wire signed [9:0] m44_22;
   assign m44_22 =10'b0;

   // m44_23 = W*in
   wire signed [9:0] m44_23;
   assign m44_23 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_24 = W*in
   wire signed [9:0] m44_24;
   assign m44_24 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_25 = W*in
   wire signed [9:0] m44_25;
   assign m44_25 =10'b0;

   // m44_26 = W*in
   wire signed [9:0] m44_26;
   assign m44_26 =10'b0;

   // m44_27 = W*in
   wire signed [9:0] m44_27;
   assign m44_27 =10'b0;

   // m44_28 = W*in
   wire signed [9:0] m44_28;
   assign m44_28 =10'b0;

   // m44_29 = W*in
   wire signed [9:0] m44_29;
   assign m44_29 =10'b0;

   // m44_30 = W*in
   wire signed [9:0] m44_30;
   assign m44_30 =10'b0;

   // m44_31 = W*in
   wire signed [9:0] m44_31;
   assign m44_31 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_32 = W*in
   wire signed [9:0] m44_32;
   assign m44_32 =10'b0;

   // m44_33 = W*in
   wire signed [9:0] m44_33;
   assign m44_33 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_34 = W*in
   wire signed [9:0] m44_34;
   assign m44_34 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_35 = W*in
   wire signed [9:0] m44_35;
   assign m44_35 =10'b0;

   // m44_36 = W*in
   wire signed [9:0] m44_36;
   assign m44_36 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_37 = W*in
   wire signed [9:0] m44_37;
   assign m44_37 =10'b0;

   // m44_38 = W*in
   wire signed [9:0] m44_38;
   assign m44_38 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_39 = W*in
   wire signed [9:0] m44_39;
   assign m44_39 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_40 = W*in
   wire signed [9:0] m44_40;
   assign m44_40 =10'b0;

   // m44_41 = W*in
   wire signed [9:0] m44_41;
   assign m44_41 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_42 = W*in
   wire signed [9:0] m44_42;
   assign m44_42 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_43 = W*in
   wire signed [9:0] m44_43;
   assign m44_43 =10'b0;

   // m44_44 = W*in
   wire signed [9:0] m44_44;
   assign m44_44 =10'b0;

   // m44_45 = W*in
   wire signed [9:0] m44_45;
   assign m44_45 =10'b0;

   // m44_46 = W*in
   wire signed [9:0] m44_46;
   assign m44_46 =10'b0;

   // m44_47 = W*in
   wire signed [9:0] m44_47;
   assign m44_47 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_48 = W*in
   wire signed [9:0] m44_48;
   assign m44_48 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_49 = W*in
   wire signed [9:0] m44_49;
   assign m44_49 =10'b0;

   // m44_50 = W*in
   wire signed [9:0] m44_50;
   assign m44_50 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_51 = W*in
   wire signed [9:0] m44_51;
   assign m44_51 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_52 = W*in
   wire signed [9:0] m44_52;
   assign m44_52 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_53 = W*in
   wire signed [9:0] m44_53;
   assign m44_53 =10'b0;

   // m44_54 = W*in
   wire signed [9:0] m44_54;
   assign m44_54 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_55 = W*in
   wire signed [9:0] m44_55;
   assign m44_55 =10'b0;

   // m44_56 = W*in
   wire signed [9:0] m44_56;
   assign m44_56 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_57 = W*in
   wire signed [9:0] m44_57;
   assign m44_57 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_58 = W*in
   wire signed [9:0] m44_58;
   assign m44_58 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_59 = W*in
   wire signed [9:0] m44_59;
   assign m44_59 ={ {3{in44[5]}} , in44 , {1{1'b0}} };

   // m44_60 = W*in
   wire signed [9:0] m44_60;
   assign m44_60 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_61 = W*in
   wire signed [9:0] m44_61;
   assign m44_61 =10'b0;

   // m44_62 = W*in
   wire signed [9:0] m44_62;
   assign m44_62 =10'b0;

   // m44_63 = W*in
   wire signed [9:0] m44_63;
   assign m44_63 =10'b0;

   // m44_64 = W*in
   wire signed [9:0] m44_64;
   assign m44_64 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_65 = W*in
   wire signed [9:0] m44_65;
   assign m44_65 =10'b0;

   // m44_66 = W*in
   wire signed [9:0] m44_66;
   assign m44_66 =10'b0;

   // m44_67 = W*in
   wire signed [9:0] m44_67;
   assign m44_67 =10'b0;

   // m44_68 = W*in
   wire signed [9:0] m44_68;
   assign m44_68 =10'b0;

   // m44_69 = W*in
   wire signed [9:0] m44_69;
   assign m44_69 ={ {2{in44[5]}} , in44 , {2{1'b0}} };

   // m44_70 = W*in
   wire signed [9:0] m44_70;
   assign m44_70 =10'b0;

   // m44_71 = W*in
   wire signed [9:0] m44_71;
   assign m44_71 =10'b0;

   // m44_72 = W*in
   wire signed [9:0] m44_72;
   assign m44_72 =10'b0;

   // m44_73 = W*in
   wire signed [9:0] m44_73;
   assign m44_73 =10'b0;

   // m44_74 = W*in
   wire signed [9:0] m44_74;
   assign m44_74 =10'b0;

   // m44_75 = W*in
   wire signed [9:0] m44_75;
   assign m44_75 =10'b0;

   // m44_76 = W*in
   wire signed [9:0] m44_76;
   assign m44_76 =10'b0;

   // m44_77 = W*in
   wire signed [9:0] m44_77;
   assign m44_77 =10'b0;

   // m44_78 = W*in
   wire signed [9:0] m44_78;
   assign m44_78 ={ {3{neg44[5]}} , neg44 , {1{1'b0}} };

   // m44_79 = W*in
   wire signed [9:0] m44_79;
   assign m44_79 =10'b0;

   // m44_80 = W*in
   wire signed [9:0] m44_80;
   assign m44_80 =10'b0;

   // m44_81 = W*in
   wire signed [9:0] m44_81;
   assign m44_81 =10'b0;

   // m45_1 = W*in
   wire signed [9:0] m45_1;
   assign m45_1 =10'b0;

   // m45_2 = W*in
   wire signed [9:0] m45_2;
   assign m45_2 =10'b0;

   // m45_3 = W*in
   wire signed [9:0] m45_3;
   assign m45_3 =10'b0;

   // m45_4 = W*in
   wire signed [9:0] m45_4;
   assign m45_4 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_5 = W*in
   wire signed [9:0] m45_5;
   assign m45_5 =10'b0;

   // m45_6 = W*in
   wire signed [9:0] m45_6;
   assign m45_6 =10'b0;

   // m45_7 = W*in
   wire signed [9:0] m45_7;
   assign m45_7 =10'b0;

   // m45_8 = W*in
   wire signed [9:0] m45_8;
   assign m45_8 =10'b0;

   // m45_9 = W*in
   wire signed [9:0] m45_9;
   assign m45_9 =10'b0;

   // m45_10 = W*in
   wire signed [9:0] m45_10;
   assign m45_10 =10'b0;

   // m45_11 = W*in
   wire signed [9:0] m45_11;
   assign m45_11 =10'b0;

   // m45_12 = W*in
   wire signed [9:0] m45_12;
   assign m45_12 =10'b0;

   // m45_13 = W*in
   wire signed [9:0] m45_13;
   assign m45_13 =10'b0;

   // m45_14 = W*in
   wire signed [9:0] m45_14;
   assign m45_14 =10'b0;

   // m45_15 = W*in
   wire signed [9:0] m45_15;
   assign m45_15 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_16 = W*in
   wire signed [9:0] m45_16;
   assign m45_16 =10'b0;

   // m45_17 = W*in
   wire signed [9:0] m45_17;
   assign m45_17 =10'b0;

   // m45_18 = W*in
   wire signed [9:0] m45_18;
   assign m45_18 =10'b0;

   // m45_19 = W*in
   wire signed [9:0] m45_19;
   assign m45_19 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_20 = W*in
   wire signed [9:0] m45_20;
   assign m45_20 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_21 = W*in
   wire signed [9:0] m45_21;
   assign m45_21 =10'b0;

   // m45_22 = W*in
   wire signed [9:0] m45_22;
   assign m45_22 =10'b0;

   // m45_23 = W*in
   wire signed [9:0] m45_23;
   assign m45_23 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_24 = W*in
   wire signed [9:0] m45_24;
   assign m45_24 =10'b0;

   // m45_25 = W*in
   wire signed [9:0] m45_25;
   assign m45_25 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_26 = W*in
   wire signed [9:0] m45_26;
   assign m45_26 =10'b0;

   // m45_27 = W*in
   wire signed [9:0] m45_27;
   assign m45_27 =10'b0;

   // m45_28 = W*in
   wire signed [9:0] m45_28;
   assign m45_28 =10'b0;

   // m45_29 = W*in
   wire signed [9:0] m45_29;
   assign m45_29 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_30 = W*in
   wire signed [9:0] m45_30;
   assign m45_30 =10'b0;

   // m45_31 = W*in
   wire signed [9:0] m45_31;
   assign m45_31 =10'b0;

   // m45_32 = W*in
   wire signed [9:0] m45_32;
   assign m45_32 =10'b0;

   // m45_33 = W*in
   wire signed [9:0] m45_33;
   assign m45_33 =10'b0;

   // m45_34 = W*in
   wire signed [9:0] m45_34;
   assign m45_34 =10'b0;

   // m45_35 = W*in
   wire signed [9:0] m45_35;
   assign m45_35 =10'b0;

   // m45_36 = W*in
   wire signed [9:0] m45_36;
   assign m45_36 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_37 = W*in
   wire signed [9:0] m45_37;
   assign m45_37 =10'b0;

   // m45_38 = W*in
   wire signed [9:0] m45_38;
   assign m45_38 =10'b0;

   // m45_39 = W*in
   wire signed [9:0] m45_39;
   assign m45_39 =10'b0;

   // m45_40 = W*in
   wire signed [9:0] m45_40;
   assign m45_40 =10'b0;

   // m45_41 = W*in
   wire signed [9:0] m45_41;
   assign m45_41 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_42 = W*in
   wire signed [9:0] m45_42;
   assign m45_42 ={ {2{in45[5]}} , in45 , {2{1'b0}} };

   // m45_43 = W*in
   wire signed [9:0] m45_43;
   assign m45_43 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_44 = W*in
   wire signed [9:0] m45_44;
   assign m45_44 =10'b0;

   // m45_45 = W*in
   wire signed [9:0] m45_45;
   assign m45_45 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_46 = W*in
   wire signed [9:0] m45_46;
   assign m45_46 =10'b0;

   // m45_47 = W*in
   wire signed [9:0] m45_47;
   assign m45_47 =10'b0;

   // m45_48 = W*in
   wire signed [9:0] m45_48;
   assign m45_48 =10'b0;

   // m45_49 = W*in
   wire signed [9:0] m45_49;
   assign m45_49 ={ {2{in45[5]}} , in45 , {2{1'b0}} };

   // m45_50 = W*in
   wire signed [9:0] m45_50;
   assign m45_50 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_51 = W*in
   wire signed [9:0] m45_51;
   assign m45_51 =10'b0;

   // m45_52 = W*in
   wire signed [9:0] m45_52;
   assign m45_52 =10'b0;

   // m45_53 = W*in
   wire signed [9:0] m45_53;
   assign m45_53 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_54 = W*in
   wire signed [9:0] m45_54;
   assign m45_54 =10'b0;

   // m45_55 = W*in
   wire signed [9:0] m45_55;
   assign m45_55 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_56 = W*in
   wire signed [9:0] m45_56;
   assign m45_56 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_57 = W*in
   wire signed [9:0] m45_57;
   assign m45_57 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_58 = W*in
   wire signed [9:0] m45_58;
   assign m45_58 =10'b0;

   // m45_59 = W*in
   wire signed [9:0] m45_59;
   assign m45_59 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_60 = W*in
   wire signed [9:0] m45_60;
   assign m45_60 =10'b0;

   // m45_61 = W*in
   wire signed [9:0] m45_61;
   assign m45_61 =10'b0;

   // m45_62 = W*in
   wire signed [9:0] m45_62;
   assign m45_62 ={ {2{in45[5]}} , in45 , {2{1'b0}} };

   // m45_63 = W*in
   wire signed [9:0] m45_63;
   assign m45_63 =10'b0;

   // m45_64 = W*in
   wire signed [9:0] m45_64;
   assign m45_64 =10'b0;

   // m45_65 = W*in
   wire signed [9:0] m45_65;
   assign m45_65 =10'b0;

   // m45_66 = W*in
   wire signed [9:0] m45_66;
   assign m45_66 ={ {2{in45[5]}} , in45 , {2{1'b0}} };

   // m45_67 = W*in
   wire signed [9:0] m45_67;
   assign m45_67 =10'b0;

   // m45_68 = W*in
   wire signed [9:0] m45_68;
   assign m45_68 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_69 = W*in
   wire signed [9:0] m45_69;
   assign m45_69 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_70 = W*in
   wire signed [9:0] m45_70;
   assign m45_70 =10'b0;

   // m45_71 = W*in
   wire signed [9:0] m45_71;
   assign m45_71 =10'b0;

   // m45_72 = W*in
   wire signed [9:0] m45_72;
   assign m45_72 =10'b0;

   // m45_73 = W*in
   wire signed [9:0] m45_73;
   assign m45_73 =10'b0;

   // m45_74 = W*in
   wire signed [9:0] m45_74;
   assign m45_74 =10'b0;

   // m45_75 = W*in
   wire signed [9:0] m45_75;
   assign m45_75 =10'b0;

   // m45_76 = W*in
   wire signed [9:0] m45_76;
   assign m45_76 =10'b0;

   // m45_77 = W*in
   wire signed [9:0] m45_77;
   assign m45_77 =10'b0;

   // m45_78 = W*in
   wire signed [9:0] m45_78;
   assign m45_78 =10'b0;

   // m45_79 = W*in
   wire signed [9:0] m45_79;
   assign m45_79 ={ {3{neg45[5]}} , neg45 , {1{1'b0}} };

   // m45_80 = W*in
   wire signed [9:0] m45_80;
   assign m45_80 =10'b0;

   // m45_81 = W*in
   wire signed [9:0] m45_81;
   assign m45_81 =10'b0;

   // m46_1 = W*in
   wire signed [9:0] m46_1;
   assign m46_1 =10'b0;

   // m46_2 = W*in
   wire signed [9:0] m46_2;
   assign m46_2 =10'b0;

   // m46_3 = W*in
   wire signed [9:0] m46_3;
   assign m46_3 =10'b0;

   // m46_4 = W*in
   wire signed [9:0] m46_4;
   assign m46_4 =10'b0;

   // m46_5 = W*in
   wire signed [9:0] m46_5;
   assign m46_5 =10'b0;

   // m46_6 = W*in
   wire signed [9:0] m46_6;
   assign m46_6 =10'b0;

   // m46_7 = W*in
   wire signed [9:0] m46_7;
   assign m46_7 =10'b0;

   // m46_8 = W*in
   wire signed [9:0] m46_8;
   assign m46_8 =10'b0;

   // m46_9 = W*in
   wire signed [9:0] m46_9;
   assign m46_9 =10'b0;

   // m46_10 = W*in
   wire signed [9:0] m46_10;
   assign m46_10 =10'b0;

   // m46_11 = W*in
   wire signed [9:0] m46_11;
   assign m46_11 =10'b0;

   // m46_12 = W*in
   wire signed [9:0] m46_12;
   assign m46_12 =10'b0;

   // m46_13 = W*in
   wire signed [9:0] m46_13;
   assign m46_13 =10'b0;

   // m46_14 = W*in
   wire signed [9:0] m46_14;
   assign m46_14 ={ {2{in46[5]}} , in46 , {2{1'b0}} };

   // m46_15 = W*in
   wire signed [9:0] m46_15;
   assign m46_15 =10'b0;

   // m46_16 = W*in
   wire signed [9:0] m46_16;
   assign m46_16 =10'b0;

   // m46_17 = W*in
   wire signed [9:0] m46_17;
   assign m46_17 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_18 = W*in
   wire signed [9:0] m46_18;
   assign m46_18 =10'b0;

   // m46_19 = W*in
   wire signed [9:0] m46_19;
   assign m46_19 =10'b0;

   // m46_20 = W*in
   wire signed [9:0] m46_20;
   assign m46_20 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_21 = W*in
   wire signed [9:0] m46_21;
   assign m46_21 =10'b0;

   // m46_22 = W*in
   wire signed [9:0] m46_22;
   assign m46_22 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_23 = W*in
   wire signed [9:0] m46_23;
   assign m46_23 =10'b0;

   // m46_24 = W*in
   wire signed [9:0] m46_24;
   assign m46_24 =10'b0;

   // m46_25 = W*in
   wire signed [9:0] m46_25;
   assign m46_25 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_26 = W*in
   wire signed [9:0] m46_26;
   assign m46_26 =10'b0;

   // m46_27 = W*in
   wire signed [9:0] m46_27;
   assign m46_27 =10'b0;

   // m46_28 = W*in
   wire signed [9:0] m46_28;
   assign m46_28 =10'b0;

   // m46_29 = W*in
   wire signed [9:0] m46_29;
   assign m46_29 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_30 = W*in
   wire signed [9:0] m46_30;
   assign m46_30 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_31 = W*in
   wire signed [9:0] m46_31;
   assign m46_31 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_32 = W*in
   wire signed [9:0] m46_32;
   assign m46_32 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_33 = W*in
   wire signed [9:0] m46_33;
   assign m46_33 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_34 = W*in
   wire signed [9:0] m46_34;
   assign m46_34 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_35 = W*in
   wire signed [9:0] m46_35;
   assign m46_35 =10'b0;

   // m46_36 = W*in
   wire signed [9:0] m46_36;
   assign m46_36 =10'b0;

   // m46_37 = W*in
   wire signed [9:0] m46_37;
   assign m46_37 ={ {2{in46[5]}} , in46 , {2{1'b0}} };

   // m46_38 = W*in
   wire signed [9:0] m46_38;
   assign m46_38 =10'b0;

   // m46_39 = W*in
   wire signed [9:0] m46_39;
   assign m46_39 =10'b0;

   // m46_40 = W*in
   wire signed [9:0] m46_40;
   assign m46_40 =10'b0;

   // m46_41 = W*in
   wire signed [9:0] m46_41;
   assign m46_41 =10'b0;

   // m46_42 = W*in
   wire signed [9:0] m46_42;
   assign m46_42 =10'b0;

   // m46_43 = W*in
   wire signed [9:0] m46_43;
   assign m46_43 ={ {2{in46[5]}} , in46 , {2{1'b0}} };

   // m46_44 = W*in
   wire signed [9:0] m46_44;
   assign m46_44 =10'b0;

   // m46_45 = W*in
   wire signed [9:0] m46_45;
   assign m46_45 =10'b0;

   // m46_46 = W*in
   wire signed [9:0] m46_46;
   assign m46_46 =10'b0;

   // m46_47 = W*in
   wire signed [9:0] m46_47;
   assign m46_47 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_48 = W*in
   wire signed [9:0] m46_48;
   assign m46_48 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_49 = W*in
   wire signed [9:0] m46_49;
   assign m46_49 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_50 = W*in
   wire signed [9:0] m46_50;
   assign m46_50 =10'b0;

   // m46_51 = W*in
   wire signed [9:0] m46_51;
   assign m46_51 =10'b0;

   // m46_52 = W*in
   wire signed [9:0] m46_52;
   assign m46_52 =10'b0;

   // m46_53 = W*in
   wire signed [9:0] m46_53;
   assign m46_53 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_54 = W*in
   wire signed [9:0] m46_54;
   assign m46_54 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_55 = W*in
   wire signed [9:0] m46_55;
   assign m46_55 =10'b0;

   // m46_56 = W*in
   wire signed [9:0] m46_56;
   assign m46_56 =10'b0;

   // m46_57 = W*in
   wire signed [9:0] m46_57;
   assign m46_57 =10'b0;

   // m46_58 = W*in
   wire signed [9:0] m46_58;
   assign m46_58 =10'b0;

   // m46_59 = W*in
   wire signed [9:0] m46_59;
   assign m46_59 =10'b0;

   // m46_60 = W*in
   wire signed [9:0] m46_60;
   assign m46_60 =10'b0;

   // m46_61 = W*in
   wire signed [9:0] m46_61;
   assign m46_61 =10'b0;

   // m46_62 = W*in
   wire signed [9:0] m46_62;
   assign m46_62 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_63 = W*in
   wire signed [9:0] m46_63;
   assign m46_63 ={ {2{in46[5]}} , in46 , {2{1'b0}} };

   // m46_64 = W*in
   wire signed [9:0] m46_64;
   assign m46_64 =10'b0;

   // m46_65 = W*in
   wire signed [9:0] m46_65;
   assign m46_65 =10'b0;

   // m46_66 = W*in
   wire signed [9:0] m46_66;
   assign m46_66 =10'b0;

   // m46_67 = W*in
   wire signed [9:0] m46_67;
   assign m46_67 =10'b0;

   // m46_68 = W*in
   wire signed [9:0] m46_68;
   assign m46_68 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_69 = W*in
   wire signed [9:0] m46_69;
   assign m46_69 =10'b0;

   // m46_70 = W*in
   wire signed [9:0] m46_70;
   assign m46_70 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_71 = W*in
   wire signed [9:0] m46_71;
   assign m46_71 =10'b0;

   // m46_72 = W*in
   wire signed [9:0] m46_72;
   assign m46_72 =10'b0;

   // m46_73 = W*in
   wire signed [9:0] m46_73;
   assign m46_73 =10'b0;

   // m46_74 = W*in
   wire signed [9:0] m46_74;
   assign m46_74 =10'b0;

   // m46_75 = W*in
   wire signed [9:0] m46_75;
   assign m46_75 =10'b0;

   // m46_76 = W*in
   wire signed [9:0] m46_76;
   assign m46_76 =10'b0;

   // m46_77 = W*in
   wire signed [9:0] m46_77;
   assign m46_77 ={ {3{neg46[5]}} , neg46 , {1{1'b0}} };

   // m46_78 = W*in
   wire signed [9:0] m46_78;
   assign m46_78 =10'b0;

   // m46_79 = W*in
   wire signed [9:0] m46_79;
   assign m46_79 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_80 = W*in
   wire signed [9:0] m46_80;
   assign m46_80 =10'b0;

   // m46_81 = W*in
   wire signed [9:0] m46_81;
   assign m46_81 =10'b0;

   // m47_1 = W*in
   wire signed [9:0] m47_1;
   assign m47_1 =10'b0;

   // m47_2 = W*in
   wire signed [9:0] m47_2;
   assign m47_2 =10'b0;

   // m47_3 = W*in
   wire signed [9:0] m47_3;
   assign m47_3 =10'b0;

   // m47_4 = W*in
   wire signed [9:0] m47_4;
   assign m47_4 =10'b0;

   // m47_5 = W*in
   wire signed [9:0] m47_5;
   assign m47_5 =10'b0;

   // m47_6 = W*in
   wire signed [9:0] m47_6;
   assign m47_6 =10'b0;

   // m47_7 = W*in
   wire signed [9:0] m47_7;
   assign m47_7 =10'b0;

   // m47_8 = W*in
   wire signed [9:0] m47_8;
   assign m47_8 =10'b0;

   // m47_9 = W*in
   wire signed [9:0] m47_9;
   assign m47_9 =10'b0;

   // m47_10 = W*in
   wire signed [9:0] m47_10;
   assign m47_10 =10'b0;

   // m47_11 = W*in
   wire signed [9:0] m47_11;
   assign m47_11 =10'b0;

   // m47_12 = W*in
   wire signed [9:0] m47_12;
   assign m47_12 =10'b0;

   // m47_13 = W*in
   wire signed [9:0] m47_13;
   assign m47_13 =10'b0;

   // m47_14 = W*in
   wire signed [9:0] m47_14;
   assign m47_14 =10'b0;

   // m47_15 = W*in
   wire signed [9:0] m47_15;
   assign m47_15 =10'b0;

   // m47_16 = W*in
   wire signed [9:0] m47_16;
   assign m47_16 =10'b0;

   // m47_17 = W*in
   wire signed [9:0] m47_17;
   assign m47_17 =10'b0;

   // m47_18 = W*in
   wire signed [9:0] m47_18;
   assign m47_18 =10'b0;

   // m47_19 = W*in
   wire signed [9:0] m47_19;
   assign m47_19 =10'b0;

   // m47_20 = W*in
   wire signed [9:0] m47_20;
   assign m47_20 =10'b0;

   // m47_21 = W*in
   wire signed [9:0] m47_21;
   assign m47_21 =10'b0;

   // m47_22 = W*in
   wire signed [9:0] m47_22;
   assign m47_22 ={ {3{neg47[5]}} , neg47 , {1{1'b0}} };

   // m47_23 = W*in
   wire signed [9:0] m47_23;
   assign m47_23 ={ {2{in47[5]}} , in47 , {2{1'b0}} };

   // m47_24 = W*in
   wire signed [9:0] m47_24;
   assign m47_24 ={ {3{in47[5]}} , in47 , {1{1'b0}} };

   // m47_25 = W*in
   wire signed [9:0] m47_25;
   assign m47_25 ={ {3{in47[5]}} , in47 , {1{1'b0}} };

   // m47_26 = W*in
   wire signed [9:0] m47_26;
   assign m47_26 =10'b0;

   // m47_27 = W*in
   wire signed [9:0] m47_27;
   assign m47_27 =10'b0;

   // m47_28 = W*in
   wire signed [9:0] m47_28;
   assign m47_28 ={ {3{in47[5]}} , in47 , {1{1'b0}} };

   // m47_29 = W*in
   wire signed [9:0] m47_29;
   assign m47_29 =10'b0;

   // m47_30 = W*in
   wire signed [9:0] m47_30;
   assign m47_30 ={ {3{in47[5]}} , in47 , {1{1'b0}} };

   // m47_31 = W*in
   wire signed [9:0] m47_31;
   assign m47_31 =10'b0;

   // m47_32 = W*in
   wire signed [9:0] m47_32;
   assign m47_32 =10'b0;

   // m47_33 = W*in
   wire signed [9:0] m47_33;
   assign m47_33 =10'b0;

   // m47_34 = W*in
   wire signed [9:0] m47_34;
   assign m47_34 =10'b0;

   // m47_35 = W*in
   wire signed [9:0] m47_35;
   assign m47_35 =10'b0;

   // m47_36 = W*in
   wire signed [9:0] m47_36;
   assign m47_36 =10'b0;

   // m47_37 = W*in
   wire signed [9:0] m47_37;
   assign m47_37 =10'b0;

   // m47_38 = W*in
   wire signed [9:0] m47_38;
   assign m47_38 =10'b0;

   // m47_39 = W*in
   wire signed [9:0] m47_39;
   assign m47_39 ={ {2{in47[5]}} , in47 , {2{1'b0}} };

   // m47_40 = W*in
   wire signed [9:0] m47_40;
   assign m47_40 =10'b0;

   // m47_41 = W*in
   wire signed [9:0] m47_41;
   assign m47_41 =10'b0;

   // m47_42 = W*in
   wire signed [9:0] m47_42;
   assign m47_42 =10'b0;

   // m47_43 = W*in
   wire signed [9:0] m47_43;
   assign m47_43 ={ {3{in47[5]}} , in47 , {1{1'b0}} };

   // m47_44 = W*in
   wire signed [9:0] m47_44;
   assign m47_44 =10'b0;

   // m47_45 = W*in
   wire signed [9:0] m47_45;
   assign m47_45 =10'b0;

   // m47_46 = W*in
   wire signed [9:0] m47_46;
   assign m47_46 =10'b0;

   // m47_47 = W*in
   wire signed [9:0] m47_47;
   assign m47_47 =10'b0;

   // m47_48 = W*in
   wire signed [9:0] m47_48;
   assign m47_48 =10'b0;

   // m47_49 = W*in
   wire signed [9:0] m47_49;
   assign m47_49 =10'b0;

   // m47_50 = W*in
   wire signed [9:0] m47_50;
   assign m47_50 =10'b0;

   // m47_51 = W*in
   wire signed [9:0] m47_51;
   assign m47_51 =10'b0;

   // m47_52 = W*in
   wire signed [9:0] m47_52;
   assign m47_52 =10'b0;

   // m47_53 = W*in
   wire signed [9:0] m47_53;
   assign m47_53 =10'b0;

   // m47_54 = W*in
   wire signed [9:0] m47_54;
   assign m47_54 =10'b0;

   // m47_55 = W*in
   wire signed [9:0] m47_55;
   assign m47_55 =10'b0;

   // m47_56 = W*in
   wire signed [9:0] m47_56;
   assign m47_56 =10'b0;

   // m47_57 = W*in
   wire signed [9:0] m47_57;
   assign m47_57 =10'b0;

   // m47_58 = W*in
   wire signed [9:0] m47_58;
   assign m47_58 =10'b0;

   // m47_59 = W*in
   wire signed [9:0] m47_59;
   assign m47_59 =10'b0;

   // m47_60 = W*in
   wire signed [9:0] m47_60;
   assign m47_60 ={ {3{neg47[5]}} , neg47 , {1{1'b0}} };

   // m47_61 = W*in
   wire signed [9:0] m47_61;
   assign m47_61 =10'b0;

   // m47_62 = W*in
   wire signed [9:0] m47_62;
   assign m47_62 =10'b0;

   // m47_63 = W*in
   wire signed [9:0] m47_63;
   assign m47_63 =10'b0;

   // m47_64 = W*in
   wire signed [9:0] m47_64;
   assign m47_64 ={ {3{in47[5]}} , in47 , {1{1'b0}} };

   // m47_65 = W*in
   wire signed [9:0] m47_65;
   assign m47_65 =10'b0;

   // m47_66 = W*in
   wire signed [9:0] m47_66;
   assign m47_66 =10'b0;

   // m47_67 = W*in
   wire signed [9:0] m47_67;
   assign m47_67 =10'b0;

   // m47_68 = W*in
   wire signed [9:0] m47_68;
   assign m47_68 =10'b0;

   // m47_69 = W*in
   wire signed [9:0] m47_69;
   assign m47_69 ={ {3{neg47[5]}} , neg47 , {1{1'b0}} };

   // m47_70 = W*in
   wire signed [9:0] m47_70;
   assign m47_70 =10'b0;

   // m47_71 = W*in
   wire signed [9:0] m47_71;
   assign m47_71 =10'b0;

   // m47_72 = W*in
   wire signed [9:0] m47_72;
   assign m47_72 =10'b0;

   // m47_73 = W*in
   wire signed [9:0] m47_73;
   assign m47_73 =10'b0;

   // m47_74 = W*in
   wire signed [9:0] m47_74;
   assign m47_74 =10'b0;

   // m47_75 = W*in
   wire signed [9:0] m47_75;
   assign m47_75 =10'b0;

   // m47_76 = W*in
   wire signed [9:0] m47_76;
   assign m47_76 =10'b0;

   // m47_77 = W*in
   wire signed [9:0] m47_77;
   assign m47_77 =10'b0;

   // m47_78 = W*in
   wire signed [9:0] m47_78;
   assign m47_78 =10'b0;

   // m47_79 = W*in
   wire signed [9:0] m47_79;
   assign m47_79 =10'b0;

   // m47_80 = W*in
   wire signed [9:0] m47_80;
   assign m47_80 =10'b0;

   // m47_81 = W*in
   wire signed [9:0] m47_81;
   assign m47_81 =10'b0;

   // m48_1 = W*in
   wire signed [9:0] m48_1;
   assign m48_1 =10'b0;

   // m48_2 = W*in
   wire signed [9:0] m48_2;
   assign m48_2 =10'b0;

   // m48_3 = W*in
   wire signed [9:0] m48_3;
   assign m48_3 =10'b0;

   // m48_4 = W*in
   wire signed [9:0] m48_4;
   assign m48_4 =10'b0;

   // m48_5 = W*in
   wire signed [9:0] m48_5;
   assign m48_5 =10'b0;

   // m48_6 = W*in
   wire signed [9:0] m48_6;
   assign m48_6 =10'b0;

   // m48_7 = W*in
   wire signed [9:0] m48_7;
   assign m48_7 =10'b0;

   // m48_8 = W*in
   wire signed [9:0] m48_8;
   assign m48_8 =10'b0;

   // m48_9 = W*in
   wire signed [9:0] m48_9;
   assign m48_9 =10'b0;

   // m48_10 = W*in
   wire signed [9:0] m48_10;
   assign m48_10 =10'b0;

   // m48_11 = W*in
   wire signed [9:0] m48_11;
   assign m48_11 =10'b0;

   // m48_12 = W*in
   wire signed [9:0] m48_12;
   assign m48_12 ={ {2{in48[5]}} , in48 , {2{1'b0}} };

   // m48_13 = W*in
   wire signed [9:0] m48_13;
   assign m48_13 =10'b0;

   // m48_14 = W*in
   wire signed [9:0] m48_14;
   assign m48_14 =10'b0;

   // m48_15 = W*in
   wire signed [9:0] m48_15;
   assign m48_15 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_16 = W*in
   wire signed [9:0] m48_16;
   assign m48_16 =10'b0;

   // m48_17 = W*in
   wire signed [9:0] m48_17;
   assign m48_17 =10'b0;

   // m48_18 = W*in
   wire signed [9:0] m48_18;
   assign m48_18 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_19 = W*in
   wire signed [9:0] m48_19;
   assign m48_19 =10'b0;

   // m48_20 = W*in
   wire signed [9:0] m48_20;
   assign m48_20 =10'b0;

   // m48_21 = W*in
   wire signed [9:0] m48_21;
   assign m48_21 =10'b0;

   // m48_22 = W*in
   wire signed [9:0] m48_22;
   assign m48_22 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_23 = W*in
   wire signed [9:0] m48_23;
   assign m48_23 ={ {2{in48[5]}} , in48 , {2{1'b0}} };

   // m48_24 = W*in
   wire signed [9:0] m48_24;
   assign m48_24 =10'b0;

   // m48_25 = W*in
   wire signed [9:0] m48_25;
   assign m48_25 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_26 = W*in
   wire signed [9:0] m48_26;
   assign m48_26 =10'b0;

   // m48_27 = W*in
   wire signed [9:0] m48_27;
   assign m48_27 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_28 = W*in
   wire signed [9:0] m48_28;
   assign m48_28 =10'b0;

   // m48_29 = W*in
   wire signed [9:0] m48_29;
   assign m48_29 =10'b0;

   // m48_30 = W*in
   wire signed [9:0] m48_30;
   assign m48_30 =10'b0;

   // m48_31 = W*in
   wire signed [9:0] m48_31;
   assign m48_31 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_32 = W*in
   wire signed [9:0] m48_32;
   assign m48_32 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_33 = W*in
   wire signed [9:0] m48_33;
   assign m48_33 =10'b0;

   // m48_34 = W*in
   wire signed [9:0] m48_34;
   assign m48_34 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_35 = W*in
   wire signed [9:0] m48_35;
   assign m48_35 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_36 = W*in
   wire signed [9:0] m48_36;
   assign m48_36 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_37 = W*in
   wire signed [9:0] m48_37;
   assign m48_37 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_38 = W*in
   wire signed [9:0] m48_38;
   assign m48_38 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_39 = W*in
   wire signed [9:0] m48_39;
   assign m48_39 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_40 = W*in
   wire signed [9:0] m48_40;
   assign m48_40 =10'b0;

   // m48_41 = W*in
   wire signed [9:0] m48_41;
   assign m48_41 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_42 = W*in
   wire signed [9:0] m48_42;
   assign m48_42 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_43 = W*in
   wire signed [9:0] m48_43;
   assign m48_43 =10'b0;

   // m48_44 = W*in
   wire signed [9:0] m48_44;
   assign m48_44 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_45 = W*in
   wire signed [9:0] m48_45;
   assign m48_45 =10'b0;

   // m48_46 = W*in
   wire signed [9:0] m48_46;
   assign m48_46 =10'b0;

   // m48_47 = W*in
   wire signed [9:0] m48_47;
   assign m48_47 =10'b0;

   // m48_48 = W*in
   wire signed [9:0] m48_48;
   assign m48_48 =10'b0;

   // m48_49 = W*in
   wire signed [9:0] m48_49;
   assign m48_49 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_50 = W*in
   wire signed [9:0] m48_50;
   assign m48_50 =10'b0;

   // m48_51 = W*in
   wire signed [9:0] m48_51;
   assign m48_51 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_52 = W*in
   wire signed [9:0] m48_52;
   assign m48_52 =10'b0;

   // m48_53 = W*in
   wire signed [9:0] m48_53;
   assign m48_53 =10'b0;

   // m48_54 = W*in
   wire signed [9:0] m48_54;
   assign m48_54 =10'b0;

   // m48_55 = W*in
   wire signed [9:0] m48_55;
   assign m48_55 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_56 = W*in
   wire signed [9:0] m48_56;
   assign m48_56 =10'b0;

   // m48_57 = W*in
   wire signed [9:0] m48_57;
   assign m48_57 =10'b0;

   // m48_58 = W*in
   wire signed [9:0] m48_58;
   assign m48_58 =10'b0;

   // m48_59 = W*in
   wire signed [9:0] m48_59;
   assign m48_59 =10'b0;

   // m48_60 = W*in
   wire signed [9:0] m48_60;
   assign m48_60 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_61 = W*in
   wire signed [9:0] m48_61;
   assign m48_61 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_62 = W*in
   wire signed [9:0] m48_62;
   assign m48_62 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_63 = W*in
   wire signed [9:0] m48_63;
   assign m48_63 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_64 = W*in
   wire signed [9:0] m48_64;
   assign m48_64 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_65 = W*in
   wire signed [9:0] m48_65;
   assign m48_65 =10'b0;

   // m48_66 = W*in
   wire signed [9:0] m48_66;
   assign m48_66 =10'b0;

   // m48_67 = W*in
   wire signed [9:0] m48_67;
   assign m48_67 ={ {2{in48[5]}} , in48 , {2{1'b0}} };

   // m48_68 = W*in
   wire signed [9:0] m48_68;
   assign m48_68 =10'b0;

   // m48_69 = W*in
   wire signed [9:0] m48_69;
   assign m48_69 =10'b0;

   // m48_70 = W*in
   wire signed [9:0] m48_70;
   assign m48_70 =10'b0;

   // m48_71 = W*in
   wire signed [9:0] m48_71;
   assign m48_71 ={ {2{in48[5]}} , in48 , {2{1'b0}} };

   // m48_72 = W*in
   wire signed [9:0] m48_72;
   assign m48_72 =10'b0;

   // m48_73 = W*in
   wire signed [9:0] m48_73;
   assign m48_73 =10'b0;

   // m48_74 = W*in
   wire signed [9:0] m48_74;
   assign m48_74 =10'b0;

   // m48_75 = W*in
   wire signed [9:0] m48_75;
   assign m48_75 =10'b0;

   // m48_76 = W*in
   wire signed [9:0] m48_76;
   assign m48_76 =10'b0;

   // m48_77 = W*in
   wire signed [9:0] m48_77;
   assign m48_77 =10'b0;

   // m48_78 = W*in
   wire signed [9:0] m48_78;
   assign m48_78 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_79 = W*in
   wire signed [9:0] m48_79;
   assign m48_79 =10'b0;

   // m48_80 = W*in
   wire signed [9:0] m48_80;
   assign m48_80 =10'b0;

   // m48_81 = W*in
   wire signed [9:0] m48_81;
   assign m48_81 =10'b0;

   // m49_1 = W*in
   wire signed [9:0] m49_1;
   assign m49_1 =10'b0;

   // m49_2 = W*in
   wire signed [9:0] m49_2;
   assign m49_2 =10'b0;

   // m49_3 = W*in
   wire signed [9:0] m49_3;
   assign m49_3 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_4 = W*in
   wire signed [9:0] m49_4;
   assign m49_4 =10'b0;

   // m49_5 = W*in
   wire signed [9:0] m49_5;
   assign m49_5 =10'b0;

   // m49_6 = W*in
   wire signed [9:0] m49_6;
   assign m49_6 =10'b0;

   // m49_7 = W*in
   wire signed [9:0] m49_7;
   assign m49_7 ={ {2{in49[5]}} , in49 , {2{1'b0}} };

   // m49_8 = W*in
   wire signed [9:0] m49_8;
   assign m49_8 =10'b0;

   // m49_9 = W*in
   wire signed [9:0] m49_9;
   assign m49_9 =10'b0;

   // m49_10 = W*in
   wire signed [9:0] m49_10;
   assign m49_10 =10'b0;

   // m49_11 = W*in
   wire signed [9:0] m49_11;
   assign m49_11 =10'b0;

   // m49_12 = W*in
   wire signed [9:0] m49_12;
   assign m49_12 =10'b0;

   // m49_13 = W*in
   wire signed [9:0] m49_13;
   assign m49_13 =10'b0;

   // m49_14 = W*in
   wire signed [9:0] m49_14;
   assign m49_14 =10'b0;

   // m49_15 = W*in
   wire signed [9:0] m49_15;
   assign m49_15 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_16 = W*in
   wire signed [9:0] m49_16;
   assign m49_16 =10'b0;

   // m49_17 = W*in
   wire signed [9:0] m49_17;
   assign m49_17 =10'b0;

   // m49_18 = W*in
   wire signed [9:0] m49_18;
   assign m49_18 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_19 = W*in
   wire signed [9:0] m49_19;
   assign m49_19 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_20 = W*in
   wire signed [9:0] m49_20;
   assign m49_20 =10'b0;

   // m49_21 = W*in
   wire signed [9:0] m49_21;
   assign m49_21 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_22 = W*in
   wire signed [9:0] m49_22;
   assign m49_22 =10'b0;

   // m49_23 = W*in
   wire signed [9:0] m49_23;
   assign m49_23 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_24 = W*in
   wire signed [9:0] m49_24;
   assign m49_24 =10'b0;

   // m49_25 = W*in
   wire signed [9:0] m49_25;
   assign m49_25 =10'b0;

   // m49_26 = W*in
   wire signed [9:0] m49_26;
   assign m49_26 =10'b0;

   // m49_27 = W*in
   wire signed [9:0] m49_27;
   assign m49_27 =10'b0;

   // m49_28 = W*in
   wire signed [9:0] m49_28;
   assign m49_28 =10'b0;

   // m49_29 = W*in
   wire signed [9:0] m49_29;
   assign m49_29 =10'b0;

   // m49_30 = W*in
   wire signed [9:0] m49_30;
   assign m49_30 =10'b0;

   // m49_31 = W*in
   wire signed [9:0] m49_31;
   assign m49_31 =10'b0;

   // m49_32 = W*in
   wire signed [9:0] m49_32;
   assign m49_32 =10'b0;

   // m49_33 = W*in
   wire signed [9:0] m49_33;
   assign m49_33 =10'b0;

   // m49_34 = W*in
   wire signed [9:0] m49_34;
   assign m49_34 =10'b0;

   // m49_35 = W*in
   wire signed [9:0] m49_35;
   assign m49_35 =10'b0;

   // m49_36 = W*in
   wire signed [9:0] m49_36;
   assign m49_36 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_37 = W*in
   wire signed [9:0] m49_37;
   assign m49_37 =10'b0;

   // m49_38 = W*in
   wire signed [9:0] m49_38;
   assign m49_38 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_39 = W*in
   wire signed [9:0] m49_39;
   assign m49_39 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_40 = W*in
   wire signed [9:0] m49_40;
   assign m49_40 =10'b0;

   // m49_41 = W*in
   wire signed [9:0] m49_41;
   assign m49_41 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_42 = W*in
   wire signed [9:0] m49_42;
   assign m49_42 ={ {2{neg49[5]}} , neg49 , {2{1'b0}} };

   // m49_43 = W*in
   wire signed [9:0] m49_43;
   assign m49_43 =10'b0;

   // m49_44 = W*in
   wire signed [9:0] m49_44;
   assign m49_44 =10'b0;

   // m49_45 = W*in
   wire signed [9:0] m49_45;
   assign m49_45 =10'b0;

   // m49_46 = W*in
   wire signed [9:0] m49_46;
   assign m49_46 =10'b0;

   // m49_47 = W*in
   wire signed [9:0] m49_47;
   assign m49_47 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_48 = W*in
   wire signed [9:0] m49_48;
   assign m49_48 =10'b0;

   // m49_49 = W*in
   wire signed [9:0] m49_49;
   assign m49_49 =10'b0;

   // m49_50 = W*in
   wire signed [9:0] m49_50;
   assign m49_50 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_51 = W*in
   wire signed [9:0] m49_51;
   assign m49_51 ={ {2{in49[5]}} , in49 , {2{1'b0}} };

   // m49_52 = W*in
   wire signed [9:0] m49_52;
   assign m49_52 =10'b0;

   // m49_53 = W*in
   wire signed [9:0] m49_53;
   assign m49_53 =10'b0;

   // m49_54 = W*in
   wire signed [9:0] m49_54;
   assign m49_54 =10'b0;

   // m49_55 = W*in
   wire signed [9:0] m49_55;
   assign m49_55 =10'b0;

   // m49_56 = W*in
   wire signed [9:0] m49_56;
   assign m49_56 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_57 = W*in
   wire signed [9:0] m49_57;
   assign m49_57 =10'b0;

   // m49_58 = W*in
   wire signed [9:0] m49_58;
   assign m49_58 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_59 = W*in
   wire signed [9:0] m49_59;
   assign m49_59 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_60 = W*in
   wire signed [9:0] m49_60;
   assign m49_60 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_61 = W*in
   wire signed [9:0] m49_61;
   assign m49_61 =10'b0;

   // m49_62 = W*in
   wire signed [9:0] m49_62;
   assign m49_62 =10'b0;

   // m49_63 = W*in
   wire signed [9:0] m49_63;
   assign m49_63 =10'b0;

   // m49_64 = W*in
   wire signed [9:0] m49_64;
   assign m49_64 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_65 = W*in
   wire signed [9:0] m49_65;
   assign m49_65 =10'b0;

   // m49_66 = W*in
   wire signed [9:0] m49_66;
   assign m49_66 =10'b0;

   // m49_67 = W*in
   wire signed [9:0] m49_67;
   assign m49_67 =10'b0;

   // m49_68 = W*in
   wire signed [9:0] m49_68;
   assign m49_68 =10'b0;

   // m49_69 = W*in
   wire signed [9:0] m49_69;
   assign m49_69 ={ {2{in49[5]}} , in49 , {2{1'b0}} };

   // m49_70 = W*in
   wire signed [9:0] m49_70;
   assign m49_70 =10'b0;

   // m49_71 = W*in
   wire signed [9:0] m49_71;
   assign m49_71 =10'b0;

   // m49_72 = W*in
   wire signed [9:0] m49_72;
   assign m49_72 =10'b0;

   // m49_73 = W*in
   wire signed [9:0] m49_73;
   assign m49_73 =10'b0;

   // m49_74 = W*in
   wire signed [9:0] m49_74;
   assign m49_74 =10'b0;

   // m49_75 = W*in
   wire signed [9:0] m49_75;
   assign m49_75 =10'b0;

   // m49_76 = W*in
   wire signed [9:0] m49_76;
   assign m49_76 =10'b0;

   // m49_77 = W*in
   wire signed [9:0] m49_77;
   assign m49_77 =10'b0;

   // m49_78 = W*in
   wire signed [9:0] m49_78;
   assign m49_78 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_79 = W*in
   wire signed [9:0] m49_79;
   assign m49_79 =10'b0;

   // m49_80 = W*in
   wire signed [9:0] m49_80;
   assign m49_80 =10'b0;

   // m49_81 = W*in
   wire signed [9:0] m49_81;
   assign m49_81 =10'b0;

   // m50_1 = W*in
   wire signed [9:0] m50_1;
   assign m50_1 =10'b0;

   // m50_2 = W*in
   wire signed [9:0] m50_2;
   assign m50_2 =10'b0;

   // m50_3 = W*in
   wire signed [9:0] m50_3;
   assign m50_3 =10'b0;

   // m50_4 = W*in
   wire signed [9:0] m50_4;
   assign m50_4 =10'b0;

   // m50_5 = W*in
   wire signed [9:0] m50_5;
   assign m50_5 =10'b0;

   // m50_6 = W*in
   wire signed [9:0] m50_6;
   assign m50_6 =10'b0;

   // m50_7 = W*in
   wire signed [9:0] m50_7;
   assign m50_7 =10'b0;

   // m50_8 = W*in
   wire signed [9:0] m50_8;
   assign m50_8 =10'b0;

   // m50_9 = W*in
   wire signed [9:0] m50_9;
   assign m50_9 =10'b0;

   // m50_10 = W*in
   wire signed [9:0] m50_10;
   assign m50_10 =10'b0;

   // m50_11 = W*in
   wire signed [9:0] m50_11;
   assign m50_11 =10'b0;

   // m50_12 = W*in
   wire signed [9:0] m50_12;
   assign m50_12 =10'b0;

   // m50_13 = W*in
   wire signed [9:0] m50_13;
   assign m50_13 =10'b0;

   // m50_14 = W*in
   wire signed [9:0] m50_14;
   assign m50_14 =10'b0;

   // m50_15 = W*in
   wire signed [9:0] m50_15;
   assign m50_15 =10'b0;

   // m50_16 = W*in
   wire signed [9:0] m50_16;
   assign m50_16 =10'b0;

   // m50_17 = W*in
   wire signed [9:0] m50_17;
   assign m50_17 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_18 = W*in
   wire signed [9:0] m50_18;
   assign m50_18 =10'b0;

   // m50_19 = W*in
   wire signed [9:0] m50_19;
   assign m50_19 =10'b0;

   // m50_20 = W*in
   wire signed [9:0] m50_20;
   assign m50_20 ={ {2{in50[5]}} , in50 , {2{1'b0}} };

   // m50_21 = W*in
   wire signed [9:0] m50_21;
   assign m50_21 =10'b0;

   // m50_22 = W*in
   wire signed [9:0] m50_22;
   assign m50_22 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_23 = W*in
   wire signed [9:0] m50_23;
   assign m50_23 =10'b0;

   // m50_24 = W*in
   wire signed [9:0] m50_24;
   assign m50_24 =10'b0;

   // m50_25 = W*in
   wire signed [9:0] m50_25;
   assign m50_25 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_26 = W*in
   wire signed [9:0] m50_26;
   assign m50_26 =10'b0;

   // m50_27 = W*in
   wire signed [9:0] m50_27;
   assign m50_27 =10'b0;

   // m50_28 = W*in
   wire signed [9:0] m50_28;
   assign m50_28 =10'b0;

   // m50_29 = W*in
   wire signed [9:0] m50_29;
   assign m50_29 ={ {2{in50[5]}} , in50 , {2{1'b0}} };

   // m50_30 = W*in
   wire signed [9:0] m50_30;
   assign m50_30 =10'b0;

   // m50_31 = W*in
   wire signed [9:0] m50_31;
   assign m50_31 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_32 = W*in
   wire signed [9:0] m50_32;
   assign m50_32 =10'b0;

   // m50_33 = W*in
   wire signed [9:0] m50_33;
   assign m50_33 =10'b0;

   // m50_34 = W*in
   wire signed [9:0] m50_34;
   assign m50_34 =10'b0;

   // m50_35 = W*in
   wire signed [9:0] m50_35;
   assign m50_35 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_36 = W*in
   wire signed [9:0] m50_36;
   assign m50_36 =10'b0;

   // m50_37 = W*in
   wire signed [9:0] m50_37;
   assign m50_37 =10'b0;

   // m50_38 = W*in
   wire signed [9:0] m50_38;
   assign m50_38 =10'b0;

   // m50_39 = W*in
   wire signed [9:0] m50_39;
   assign m50_39 =10'b0;

   // m50_40 = W*in
   wire signed [9:0] m50_40;
   assign m50_40 =10'b0;

   // m50_41 = W*in
   wire signed [9:0] m50_41;
   assign m50_41 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_42 = W*in
   wire signed [9:0] m50_42;
   assign m50_42 =10'b0;

   // m50_43 = W*in
   wire signed [9:0] m50_43;
   assign m50_43 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_44 = W*in
   wire signed [9:0] m50_44;
   assign m50_44 =10'b0;

   // m50_45 = W*in
   wire signed [9:0] m50_45;
   assign m50_45 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_46 = W*in
   wire signed [9:0] m50_46;
   assign m50_46 =10'b0;

   // m50_47 = W*in
   wire signed [9:0] m50_47;
   assign m50_47 =10'b0;

   // m50_48 = W*in
   wire signed [9:0] m50_48;
   assign m50_48 ={ {2{in50[5]}} , in50 , {2{1'b0}} };

   // m50_49 = W*in
   wire signed [9:0] m50_49;
   assign m50_49 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_50 = W*in
   wire signed [9:0] m50_50;
   assign m50_50 =10'b0;

   // m50_51 = W*in
   wire signed [9:0] m50_51;
   assign m50_51 =10'b0;

   // m50_52 = W*in
   wire signed [9:0] m50_52;
   assign m50_52 =10'b0;

   // m50_53 = W*in
   wire signed [9:0] m50_53;
   assign m50_53 =10'b0;

   // m50_54 = W*in
   wire signed [9:0] m50_54;
   assign m50_54 =10'b0;

   // m50_55 = W*in
   wire signed [9:0] m50_55;
   assign m50_55 =10'b0;

   // m50_56 = W*in
   wire signed [9:0] m50_56;
   assign m50_56 =10'b0;

   // m50_57 = W*in
   wire signed [9:0] m50_57;
   assign m50_57 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_58 = W*in
   wire signed [9:0] m50_58;
   assign m50_58 =10'b0;

   // m50_59 = W*in
   wire signed [9:0] m50_59;
   assign m50_59 =10'b0;

   // m50_60 = W*in
   wire signed [9:0] m50_60;
   assign m50_60 =10'b0;

   // m50_61 = W*in
   wire signed [9:0] m50_61;
   assign m50_61 =10'b0;

   // m50_62 = W*in
   wire signed [9:0] m50_62;
   assign m50_62 =10'b0;

   // m50_63 = W*in
   wire signed [9:0] m50_63;
   assign m50_63 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_64 = W*in
   wire signed [9:0] m50_64;
   assign m50_64 ={ {2{in50[5]}} , in50 , {2{1'b0}} };

   // m50_65 = W*in
   wire signed [9:0] m50_65;
   assign m50_65 =10'b0;

   // m50_66 = W*in
   wire signed [9:0] m50_66;
   assign m50_66 =10'b0;

   // m50_67 = W*in
   wire signed [9:0] m50_67;
   assign m50_67 =10'b0;

   // m50_68 = W*in
   wire signed [9:0] m50_68;
   assign m50_68 =10'b0;

   // m50_69 = W*in
   wire signed [9:0] m50_69;
   assign m50_69 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_70 = W*in
   wire signed [9:0] m50_70;
   assign m50_70 =10'b0;

   // m50_71 = W*in
   wire signed [9:0] m50_71;
   assign m50_71 =10'b0;

   // m50_72 = W*in
   wire signed [9:0] m50_72;
   assign m50_72 =10'b0;

   // m50_73 = W*in
   wire signed [9:0] m50_73;
   assign m50_73 =10'b0;

   // m50_74 = W*in
   wire signed [9:0] m50_74;
   assign m50_74 =10'b0;

   // m50_75 = W*in
   wire signed [9:0] m50_75;
   assign m50_75 =10'b0;

   // m50_76 = W*in
   wire signed [9:0] m50_76;
   assign m50_76 =10'b0;

   // m50_77 = W*in
   wire signed [9:0] m50_77;
   assign m50_77 =10'b0;

   // m50_78 = W*in
   wire signed [9:0] m50_78;
   assign m50_78 =10'b0;

   // m50_79 = W*in
   wire signed [9:0] m50_79;
   assign m50_79 =10'b0;

   // m50_80 = W*in
   wire signed [9:0] m50_80;
   assign m50_80 =10'b0;

   // m50_81 = W*in
   wire signed [9:0] m50_81;
   assign m50_81 =10'b0;

   // m51_1 = W*in
   wire signed [9:0] m51_1;
   assign m51_1 =10'b0;

   // m51_2 = W*in
   wire signed [9:0] m51_2;
   assign m51_2 =10'b0;

   // m51_3 = W*in
   wire signed [9:0] m51_3;
   assign m51_3 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_4 = W*in
   wire signed [9:0] m51_4;
   assign m51_4 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_5 = W*in
   wire signed [9:0] m51_5;
   assign m51_5 =10'b0;

   // m51_6 = W*in
   wire signed [9:0] m51_6;
   assign m51_6 =10'b0;

   // m51_7 = W*in
   wire signed [9:0] m51_7;
   assign m51_7 =10'b0;

   // m51_8 = W*in
   wire signed [9:0] m51_8;
   assign m51_8 =10'b0;

   // m51_9 = W*in
   wire signed [9:0] m51_9;
   assign m51_9 =10'b0;

   // m51_10 = W*in
   wire signed [9:0] m51_10;
   assign m51_10 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_11 = W*in
   wire signed [9:0] m51_11;
   assign m51_11 =10'b0;

   // m51_12 = W*in
   wire signed [9:0] m51_12;
   assign m51_12 =10'b0;

   // m51_13 = W*in
   wire signed [9:0] m51_13;
   assign m51_13 =10'b0;

   // m51_14 = W*in
   wire signed [9:0] m51_14;
   assign m51_14 =10'b0;

   // m51_15 = W*in
   wire signed [9:0] m51_15;
   assign m51_15 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_16 = W*in
   wire signed [9:0] m51_16;
   assign m51_16 =10'b0;

   // m51_17 = W*in
   wire signed [9:0] m51_17;
   assign m51_17 =10'b0;

   // m51_18 = W*in
   wire signed [9:0] m51_18;
   assign m51_18 =10'b0;

   // m51_19 = W*in
   wire signed [9:0] m51_19;
   assign m51_19 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_20 = W*in
   wire signed [9:0] m51_20;
   assign m51_20 =10'b0;

   // m51_21 = W*in
   wire signed [9:0] m51_21;
   assign m51_21 =10'b0;

   // m51_22 = W*in
   wire signed [9:0] m51_22;
   assign m51_22 =10'b0;

   // m51_23 = W*in
   wire signed [9:0] m51_23;
   assign m51_23 =10'b0;

   // m51_24 = W*in
   wire signed [9:0] m51_24;
   assign m51_24 =10'b0;

   // m51_25 = W*in
   wire signed [9:0] m51_25;
   assign m51_25 =10'b0;

   // m51_26 = W*in
   wire signed [9:0] m51_26;
   assign m51_26 =10'b0;

   // m51_27 = W*in
   wire signed [9:0] m51_27;
   assign m51_27 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_28 = W*in
   wire signed [9:0] m51_28;
   assign m51_28 =10'b0;

   // m51_29 = W*in
   wire signed [9:0] m51_29;
   assign m51_29 =10'b0;

   // m51_30 = W*in
   wire signed [9:0] m51_30;
   assign m51_30 =10'b0;

   // m51_31 = W*in
   wire signed [9:0] m51_31;
   assign m51_31 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_32 = W*in
   wire signed [9:0] m51_32;
   assign m51_32 =10'b0;

   // m51_33 = W*in
   wire signed [9:0] m51_33;
   assign m51_33 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_34 = W*in
   wire signed [9:0] m51_34;
   assign m51_34 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_35 = W*in
   wire signed [9:0] m51_35;
   assign m51_35 =10'b0;

   // m51_36 = W*in
   wire signed [9:0] m51_36;
   assign m51_36 =10'b0;

   // m51_37 = W*in
   wire signed [9:0] m51_37;
   assign m51_37 =10'b0;

   // m51_38 = W*in
   wire signed [9:0] m51_38;
   assign m51_38 =10'b0;

   // m51_39 = W*in
   wire signed [9:0] m51_39;
   assign m51_39 =10'b0;

   // m51_40 = W*in
   wire signed [9:0] m51_40;
   assign m51_40 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_41 = W*in
   wire signed [9:0] m51_41;
   assign m51_41 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_42 = W*in
   wire signed [9:0] m51_42;
   assign m51_42 =10'b0;

   // m51_43 = W*in
   wire signed [9:0] m51_43;
   assign m51_43 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_44 = W*in
   wire signed [9:0] m51_44;
   assign m51_44 ={ {2{in51[5]}} , in51 , {2{1'b0}} };

   // m51_45 = W*in
   wire signed [9:0] m51_45;
   assign m51_45 =10'b0;

   // m51_46 = W*in
   wire signed [9:0] m51_46;
   assign m51_46 =10'b0;

   // m51_47 = W*in
   wire signed [9:0] m51_47;
   assign m51_47 =10'b0;

   // m51_48 = W*in
   wire signed [9:0] m51_48;
   assign m51_48 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_49 = W*in
   wire signed [9:0] m51_49;
   assign m51_49 ={ {2{in51[5]}} , in51 , {2{1'b0}} };

   // m51_50 = W*in
   wire signed [9:0] m51_50;
   assign m51_50 =10'b0;

   // m51_51 = W*in
   wire signed [9:0] m51_51;
   assign m51_51 =10'b0;

   // m51_52 = W*in
   wire signed [9:0] m51_52;
   assign m51_52 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_53 = W*in
   wire signed [9:0] m51_53;
   assign m51_53 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_54 = W*in
   wire signed [9:0] m51_54;
   assign m51_54 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_55 = W*in
   wire signed [9:0] m51_55;
   assign m51_55 ={ {2{in51[5]}} , in51 , {2{1'b0}} };

   // m51_56 = W*in
   wire signed [9:0] m51_56;
   assign m51_56 ={ {2{neg51[5]}} , neg51 , {2{1'b0}} };

   // m51_57 = W*in
   wire signed [9:0] m51_57;
   assign m51_57 =10'b0;

   // m51_58 = W*in
   wire signed [9:0] m51_58;
   assign m51_58 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_59 = W*in
   wire signed [9:0] m51_59;
   assign m51_59 =10'b0;

   // m51_60 = W*in
   wire signed [9:0] m51_60;
   assign m51_60 =10'b0;

   // m51_61 = W*in
   wire signed [9:0] m51_61;
   assign m51_61 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_62 = W*in
   wire signed [9:0] m51_62;
   assign m51_62 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_63 = W*in
   wire signed [9:0] m51_63;
   assign m51_63 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_64 = W*in
   wire signed [9:0] m51_64;
   assign m51_64 =10'b0;

   // m51_65 = W*in
   wire signed [9:0] m51_65;
   assign m51_65 =10'b0;

   // m51_66 = W*in
   wire signed [9:0] m51_66;
   assign m51_66 ={ {2{in51[5]}} , in51 , {2{1'b0}} };

   // m51_67 = W*in
   wire signed [9:0] m51_67;
   assign m51_67 ={ {3{in51[5]}} , in51 , {1{1'b0}} };

   // m51_68 = W*in
   wire signed [9:0] m51_68;
   assign m51_68 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_69 = W*in
   wire signed [9:0] m51_69;
   assign m51_69 =10'b0;

   // m51_70 = W*in
   wire signed [9:0] m51_70;
   assign m51_70 ={ {2{in51[5]}} , in51 , {2{1'b0}} };

   // m51_71 = W*in
   wire signed [9:0] m51_71;
   assign m51_71 =10'b0;

   // m51_72 = W*in
   wire signed [9:0] m51_72;
   assign m51_72 =10'b0;

   // m51_73 = W*in
   wire signed [9:0] m51_73;
   assign m51_73 =10'b0;

   // m51_74 = W*in
   wire signed [9:0] m51_74;
   assign m51_74 =10'b0;

   // m51_75 = W*in
   wire signed [9:0] m51_75;
   assign m51_75 =10'b0;

   // m51_76 = W*in
   wire signed [9:0] m51_76;
   assign m51_76 =10'b0;

   // m51_77 = W*in
   wire signed [9:0] m51_77;
   assign m51_77 ={ {3{neg51[5]}} , neg51 , {1{1'b0}} };

   // m51_78 = W*in
   wire signed [9:0] m51_78;
   assign m51_78 =10'b0;

   // m51_79 = W*in
   wire signed [9:0] m51_79;
   assign m51_79 =10'b0;

   // m51_80 = W*in
   wire signed [9:0] m51_80;
   assign m51_80 =10'b0;

   // m51_81 = W*in
   wire signed [9:0] m51_81;
   assign m51_81 =10'b0;

   // m52_1 = W*in
   wire signed [9:0] m52_1;
   assign m52_1 =10'b0;

   // m52_2 = W*in
   wire signed [9:0] m52_2;
   assign m52_2 =10'b0;

   // m52_3 = W*in
   wire signed [9:0] m52_3;
   assign m52_3 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_4 = W*in
   wire signed [9:0] m52_4;
   assign m52_4 =10'b0;

   // m52_5 = W*in
   wire signed [9:0] m52_5;
   assign m52_5 =10'b0;

   // m52_6 = W*in
   wire signed [9:0] m52_6;
   assign m52_6 =10'b0;

   // m52_7 = W*in
   wire signed [9:0] m52_7;
   assign m52_7 =10'b0;

   // m52_8 = W*in
   wire signed [9:0] m52_8;
   assign m52_8 =10'b0;

   // m52_9 = W*in
   wire signed [9:0] m52_9;
   assign m52_9 =10'b0;

   // m52_10 = W*in
   wire signed [9:0] m52_10;
   assign m52_10 =10'b0;

   // m52_11 = W*in
   wire signed [9:0] m52_11;
   assign m52_11 =10'b0;

   // m52_12 = W*in
   wire signed [9:0] m52_12;
   assign m52_12 =10'b0;

   // m52_13 = W*in
   wire signed [9:0] m52_13;
   assign m52_13 =10'b0;

   // m52_14 = W*in
   wire signed [9:0] m52_14;
   assign m52_14 =10'b0;

   // m52_15 = W*in
   wire signed [9:0] m52_15;
   assign m52_15 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_16 = W*in
   wire signed [9:0] m52_16;
   assign m52_16 =10'b0;

   // m52_17 = W*in
   wire signed [9:0] m52_17;
   assign m52_17 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_18 = W*in
   wire signed [9:0] m52_18;
   assign m52_18 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_19 = W*in
   wire signed [9:0] m52_19;
   assign m52_19 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_20 = W*in
   wire signed [9:0] m52_20;
   assign m52_20 =10'b0;

   // m52_21 = W*in
   wire signed [9:0] m52_21;
   assign m52_21 =10'b0;

   // m52_22 = W*in
   wire signed [9:0] m52_22;
   assign m52_22 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_23 = W*in
   wire signed [9:0] m52_23;
   assign m52_23 ={ {3{neg52[5]}} , neg52 , {1{1'b0}} };

   // m52_24 = W*in
   wire signed [9:0] m52_24;
   assign m52_24 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_25 = W*in
   wire signed [9:0] m52_25;
   assign m52_25 =10'b0;

   // m52_26 = W*in
   wire signed [9:0] m52_26;
   assign m52_26 =10'b0;

   // m52_27 = W*in
   wire signed [9:0] m52_27;
   assign m52_27 =10'b0;

   // m52_28 = W*in
   wire signed [9:0] m52_28;
   assign m52_28 =10'b0;

   // m52_29 = W*in
   wire signed [9:0] m52_29;
   assign m52_29 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_30 = W*in
   wire signed [9:0] m52_30;
   assign m52_30 ={ {3{neg52[5]}} , neg52 , {1{1'b0}} };

   // m52_31 = W*in
   wire signed [9:0] m52_31;
   assign m52_31 =10'b0;

   // m52_32 = W*in
   wire signed [9:0] m52_32;
   assign m52_32 =10'b0;

   // m52_33 = W*in
   wire signed [9:0] m52_33;
   assign m52_33 =10'b0;

   // m52_34 = W*in
   wire signed [9:0] m52_34;
   assign m52_34 =10'b0;

   // m52_35 = W*in
   wire signed [9:0] m52_35;
   assign m52_35 =10'b0;

   // m52_36 = W*in
   wire signed [9:0] m52_36;
   assign m52_36 ={ {3{neg52[5]}} , neg52 , {1{1'b0}} };

   // m52_37 = W*in
   wire signed [9:0] m52_37;
   assign m52_37 =10'b0;

   // m52_38 = W*in
   wire signed [9:0] m52_38;
   assign m52_38 =10'b0;

   // m52_39 = W*in
   wire signed [9:0] m52_39;
   assign m52_39 =10'b0;

   // m52_40 = W*in
   wire signed [9:0] m52_40;
   assign m52_40 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_41 = W*in
   wire signed [9:0] m52_41;
   assign m52_41 =10'b0;

   // m52_42 = W*in
   wire signed [9:0] m52_42;
   assign m52_42 =10'b0;

   // m52_43 = W*in
   wire signed [9:0] m52_43;
   assign m52_43 =10'b0;

   // m52_44 = W*in
   wire signed [9:0] m52_44;
   assign m52_44 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_45 = W*in
   wire signed [9:0] m52_45;
   assign m52_45 =10'b0;

   // m52_46 = W*in
   wire signed [9:0] m52_46;
   assign m52_46 =10'b0;

   // m52_47 = W*in
   wire signed [9:0] m52_47;
   assign m52_47 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_48 = W*in
   wire signed [9:0] m52_48;
   assign m52_48 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_49 = W*in
   wire signed [9:0] m52_49;
   assign m52_49 =10'b0;

   // m52_50 = W*in
   wire signed [9:0] m52_50;
   assign m52_50 ={ {3{neg52[5]}} , neg52 , {1{1'b0}} };

   // m52_51 = W*in
   wire signed [9:0] m52_51;
   assign m52_51 =10'b0;

   // m52_52 = W*in
   wire signed [9:0] m52_52;
   assign m52_52 =10'b0;

   // m52_53 = W*in
   wire signed [9:0] m52_53;
   assign m52_53 =10'b0;

   // m52_54 = W*in
   wire signed [9:0] m52_54;
   assign m52_54 =10'b0;

   // m52_55 = W*in
   wire signed [9:0] m52_55;
   assign m52_55 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_56 = W*in
   wire signed [9:0] m52_56;
   assign m52_56 =10'b0;

   // m52_57 = W*in
   wire signed [9:0] m52_57;
   assign m52_57 =10'b0;

   // m52_58 = W*in
   wire signed [9:0] m52_58;
   assign m52_58 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_59 = W*in
   wire signed [9:0] m52_59;
   assign m52_59 =10'b0;

   // m52_60 = W*in
   wire signed [9:0] m52_60;
   assign m52_60 =10'b0;

   // m52_61 = W*in
   wire signed [9:0] m52_61;
   assign m52_61 =10'b0;

   // m52_62 = W*in
   wire signed [9:0] m52_62;
   assign m52_62 =10'b0;

   // m52_63 = W*in
   wire signed [9:0] m52_63;
   assign m52_63 =10'b0;

   // m52_64 = W*in
   wire signed [9:0] m52_64;
   assign m52_64 =10'b0;

   // m52_65 = W*in
   wire signed [9:0] m52_65;
   assign m52_65 =10'b0;

   // m52_66 = W*in
   wire signed [9:0] m52_66;
   assign m52_66 =10'b0;

   // m52_67 = W*in
   wire signed [9:0] m52_67;
   assign m52_67 =10'b0;

   // m52_68 = W*in
   wire signed [9:0] m52_68;
   assign m52_68 =10'b0;

   // m52_69 = W*in
   wire signed [9:0] m52_69;
   assign m52_69 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_70 = W*in
   wire signed [9:0] m52_70;
   assign m52_70 ={ {2{in52[5]}} , in52 , {2{1'b0}} };

   // m52_71 = W*in
   wire signed [9:0] m52_71;
   assign m52_71 =10'b0;

   // m52_72 = W*in
   wire signed [9:0] m52_72;
   assign m52_72 =10'b0;

   // m52_73 = W*in
   wire signed [9:0] m52_73;
   assign m52_73 =10'b0;

   // m52_74 = W*in
   wire signed [9:0] m52_74;
   assign m52_74 =10'b0;

   // m52_75 = W*in
   wire signed [9:0] m52_75;
   assign m52_75 =10'b0;

   // m52_76 = W*in
   wire signed [9:0] m52_76;
   assign m52_76 =10'b0;

   // m52_77 = W*in
   wire signed [9:0] m52_77;
   assign m52_77 =10'b0;

   // m52_78 = W*in
   wire signed [9:0] m52_78;
   assign m52_78 ={ {3{in52[5]}} , in52 , {1{1'b0}} };

   // m52_79 = W*in
   wire signed [9:0] m52_79;
   assign m52_79 =10'b0;

   // m52_80 = W*in
   wire signed [9:0] m52_80;
   assign m52_80 =10'b0;

   // m52_81 = W*in
   wire signed [9:0] m52_81;
   assign m52_81 =10'b0;

   // m53_1 = W*in
   wire signed [9:0] m53_1;
   assign m53_1 =10'b0;

   // m53_2 = W*in
   wire signed [9:0] m53_2;
   assign m53_2 =10'b0;

   // m53_3 = W*in
   wire signed [9:0] m53_3;
   assign m53_3 =10'b0;

   // m53_4 = W*in
   wire signed [9:0] m53_4;
   assign m53_4 =10'b0;

   // m53_5 = W*in
   wire signed [9:0] m53_5;
   assign m53_5 =10'b0;

   // m53_6 = W*in
   wire signed [9:0] m53_6;
   assign m53_6 =10'b0;

   // m53_7 = W*in
   wire signed [9:0] m53_7;
   assign m53_7 ={ {2{in53[5]}} , in53 , {2{1'b0}} };

   // m53_8 = W*in
   wire signed [9:0] m53_8;
   assign m53_8 =10'b0;

   // m53_9 = W*in
   wire signed [9:0] m53_9;
   assign m53_9 =10'b0;

   // m53_10 = W*in
   wire signed [9:0] m53_10;
   assign m53_10 =10'b0;

   // m53_11 = W*in
   wire signed [9:0] m53_11;
   assign m53_11 =10'b0;

   // m53_12 = W*in
   wire signed [9:0] m53_12;
   assign m53_12 =10'b0;

   // m53_13 = W*in
   wire signed [9:0] m53_13;
   assign m53_13 =10'b0;

   // m53_14 = W*in
   wire signed [9:0] m53_14;
   assign m53_14 =10'b0;

   // m53_15 = W*in
   wire signed [9:0] m53_15;
   assign m53_15 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_16 = W*in
   wire signed [9:0] m53_16;
   assign m53_16 =10'b0;

   // m53_17 = W*in
   wire signed [9:0] m53_17;
   assign m53_17 =10'b0;

   // m53_18 = W*in
   wire signed [9:0] m53_18;
   assign m53_18 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_19 = W*in
   wire signed [9:0] m53_19;
   assign m53_19 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_20 = W*in
   wire signed [9:0] m53_20;
   assign m53_20 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_21 = W*in
   wire signed [9:0] m53_21;
   assign m53_21 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_22 = W*in
   wire signed [9:0] m53_22;
   assign m53_22 =10'b0;

   // m53_23 = W*in
   wire signed [9:0] m53_23;
   assign m53_23 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_24 = W*in
   wire signed [9:0] m53_24;
   assign m53_24 =10'b0;

   // m53_25 = W*in
   wire signed [9:0] m53_25;
   assign m53_25 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_26 = W*in
   wire signed [9:0] m53_26;
   assign m53_26 =10'b0;

   // m53_27 = W*in
   wire signed [9:0] m53_27;
   assign m53_27 =10'b0;

   // m53_28 = W*in
   wire signed [9:0] m53_28;
   assign m53_28 =10'b0;

   // m53_29 = W*in
   wire signed [9:0] m53_29;
   assign m53_29 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_30 = W*in
   wire signed [9:0] m53_30;
   assign m53_30 =10'b0;

   // m53_31 = W*in
   wire signed [9:0] m53_31;
   assign m53_31 =10'b0;

   // m53_32 = W*in
   wire signed [9:0] m53_32;
   assign m53_32 =10'b0;

   // m53_33 = W*in
   wire signed [9:0] m53_33;
   assign m53_33 =10'b0;

   // m53_34 = W*in
   wire signed [9:0] m53_34;
   assign m53_34 =10'b0;

   // m53_35 = W*in
   wire signed [9:0] m53_35;
   assign m53_35 =10'b0;

   // m53_36 = W*in
   wire signed [9:0] m53_36;
   assign m53_36 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_37 = W*in
   wire signed [9:0] m53_37;
   assign m53_37 =10'b0;

   // m53_38 = W*in
   wire signed [9:0] m53_38;
   assign m53_38 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_39 = W*in
   wire signed [9:0] m53_39;
   assign m53_39 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_40 = W*in
   wire signed [9:0] m53_40;
   assign m53_40 =10'b0;

   // m53_41 = W*in
   wire signed [9:0] m53_41;
   assign m53_41 =10'b0;

   // m53_42 = W*in
   wire signed [9:0] m53_42;
   assign m53_42 ={ {2{neg53[5]}} , neg53 , {2{1'b0}} };

   // m53_43 = W*in
   wire signed [9:0] m53_43;
   assign m53_43 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_44 = W*in
   wire signed [9:0] m53_44;
   assign m53_44 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_45 = W*in
   wire signed [9:0] m53_45;
   assign m53_45 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_46 = W*in
   wire signed [9:0] m53_46;
   assign m53_46 =10'b0;

   // m53_47 = W*in
   wire signed [9:0] m53_47;
   assign m53_47 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_48 = W*in
   wire signed [9:0] m53_48;
   assign m53_48 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_49 = W*in
   wire signed [9:0] m53_49;
   assign m53_49 =10'b0;

   // m53_50 = W*in
   wire signed [9:0] m53_50;
   assign m53_50 ={ {3{neg53[5]}} , neg53 , {1{1'b0}} };

   // m53_51 = W*in
   wire signed [9:0] m53_51;
   assign m53_51 ={ {2{in53[5]}} , in53 , {2{1'b0}} };

   // m53_52 = W*in
   wire signed [9:0] m53_52;
   assign m53_52 =10'b0;

   // m53_53 = W*in
   wire signed [9:0] m53_53;
   assign m53_53 =10'b0;

   // m53_54 = W*in
   wire signed [9:0] m53_54;
   assign m53_54 =10'b0;

   // m53_55 = W*in
   wire signed [9:0] m53_55;
   assign m53_55 =10'b0;

   // m53_56 = W*in
   wire signed [9:0] m53_56;
   assign m53_56 =10'b0;

   // m53_57 = W*in
   wire signed [9:0] m53_57;
   assign m53_57 =10'b0;

   // m53_58 = W*in
   wire signed [9:0] m53_58;
   assign m53_58 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_59 = W*in
   wire signed [9:0] m53_59;
   assign m53_59 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_60 = W*in
   wire signed [9:0] m53_60;
   assign m53_60 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_61 = W*in
   wire signed [9:0] m53_61;
   assign m53_61 =10'b0;

   // m53_62 = W*in
   wire signed [9:0] m53_62;
   assign m53_62 =10'b0;

   // m53_63 = W*in
   wire signed [9:0] m53_63;
   assign m53_63 =10'b0;

   // m53_64 = W*in
   wire signed [9:0] m53_64;
   assign m53_64 =10'b0;

   // m53_65 = W*in
   wire signed [9:0] m53_65;
   assign m53_65 =10'b0;

   // m53_66 = W*in
   wire signed [9:0] m53_66;
   assign m53_66 =10'b0;

   // m53_67 = W*in
   wire signed [9:0] m53_67;
   assign m53_67 =10'b0;

   // m53_68 = W*in
   wire signed [9:0] m53_68;
   assign m53_68 =10'b0;

   // m53_69 = W*in
   wire signed [9:0] m53_69;
   assign m53_69 ={ {2{in53[5]}} , in53 , {2{1'b0}} };

   // m53_70 = W*in
   wire signed [9:0] m53_70;
   assign m53_70 =10'b0;

   // m53_71 = W*in
   wire signed [9:0] m53_71;
   assign m53_71 =10'b0;

   // m53_72 = W*in
   wire signed [9:0] m53_72;
   assign m53_72 =10'b0;

   // m53_73 = W*in
   wire signed [9:0] m53_73;
   assign m53_73 =10'b0;

   // m53_74 = W*in
   wire signed [9:0] m53_74;
   assign m53_74 =10'b0;

   // m53_75 = W*in
   wire signed [9:0] m53_75;
   assign m53_75 =10'b0;

   // m53_76 = W*in
   wire signed [9:0] m53_76;
   assign m53_76 =10'b0;

   // m53_77 = W*in
   wire signed [9:0] m53_77;
   assign m53_77 =10'b0;

   // m53_78 = W*in
   wire signed [9:0] m53_78;
   assign m53_78 =10'b0;

   // m53_79 = W*in
   wire signed [9:0] m53_79;
   assign m53_79 ={ {3{in53[5]}} , in53 , {1{1'b0}} };

   // m53_80 = W*in
   wire signed [9:0] m53_80;
   assign m53_80 =10'b0;

   // m53_81 = W*in
   wire signed [9:0] m53_81;
   assign m53_81 =10'b0;

   // m54_1 = W*in
   wire signed [9:0] m54_1;
   assign m54_1 =10'b0;

   // m54_2 = W*in
   wire signed [9:0] m54_2;
   assign m54_2 =10'b0;

   // m54_3 = W*in
   wire signed [9:0] m54_3;
   assign m54_3 =10'b0;

   // m54_4 = W*in
   wire signed [9:0] m54_4;
   assign m54_4 =10'b0;

   // m54_5 = W*in
   wire signed [9:0] m54_5;
   assign m54_5 =10'b0;

   // m54_6 = W*in
   wire signed [9:0] m54_6;
   assign m54_6 =10'b0;

   // m54_7 = W*in
   wire signed [9:0] m54_7;
   assign m54_7 =10'b0;

   // m54_8 = W*in
   wire signed [9:0] m54_8;
   assign m54_8 =10'b0;

   // m54_9 = W*in
   wire signed [9:0] m54_9;
   assign m54_9 =10'b0;

   // m54_10 = W*in
   wire signed [9:0] m54_10;
   assign m54_10 =10'b0;

   // m54_11 = W*in
   wire signed [9:0] m54_11;
   assign m54_11 =10'b0;

   // m54_12 = W*in
   wire signed [9:0] m54_12;
   assign m54_12 =10'b0;

   // m54_13 = W*in
   wire signed [9:0] m54_13;
   assign m54_13 =10'b0;

   // m54_14 = W*in
   wire signed [9:0] m54_14;
   assign m54_14 =10'b0;

   // m54_15 = W*in
   wire signed [9:0] m54_15;
   assign m54_15 ={ {2{in54[5]}} , in54 , {2{1'b0}} };

   // m54_16 = W*in
   wire signed [9:0] m54_16;
   assign m54_16 =10'b0;

   // m54_17 = W*in
   wire signed [9:0] m54_17;
   assign m54_17 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_18 = W*in
   wire signed [9:0] m54_18;
   assign m54_18 =10'b0;

   // m54_19 = W*in
   wire signed [9:0] m54_19;
   assign m54_19 =10'b0;

   // m54_20 = W*in
   wire signed [9:0] m54_20;
   assign m54_20 =10'b0;

   // m54_21 = W*in
   wire signed [9:0] m54_21;
   assign m54_21 =10'b0;

   // m54_22 = W*in
   wire signed [9:0] m54_22;
   assign m54_22 =10'b0;

   // m54_23 = W*in
   wire signed [9:0] m54_23;
   assign m54_23 =10'b0;

   // m54_24 = W*in
   wire signed [9:0] m54_24;
   assign m54_24 =10'b0;

   // m54_25 = W*in
   wire signed [9:0] m54_25;
   assign m54_25 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_26 = W*in
   wire signed [9:0] m54_26;
   assign m54_26 =10'b0;

   // m54_27 = W*in
   wire signed [9:0] m54_27;
   assign m54_27 =10'b0;

   // m54_28 = W*in
   wire signed [9:0] m54_28;
   assign m54_28 =10'b0;

   // m54_29 = W*in
   wire signed [9:0] m54_29;
   assign m54_29 =10'b0;

   // m54_30 = W*in
   wire signed [9:0] m54_30;
   assign m54_30 =10'b0;

   // m54_31 = W*in
   wire signed [9:0] m54_31;
   assign m54_31 =10'b0;

   // m54_32 = W*in
   wire signed [9:0] m54_32;
   assign m54_32 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_33 = W*in
   wire signed [9:0] m54_33;
   assign m54_33 =10'b0;

   // m54_34 = W*in
   wire signed [9:0] m54_34;
   assign m54_34 =10'b0;

   // m54_35 = W*in
   wire signed [9:0] m54_35;
   assign m54_35 =10'b0;

   // m54_36 = W*in
   wire signed [9:0] m54_36;
   assign m54_36 ={ {3{neg54[5]}} , neg54 , {1{1'b0}} };

   // m54_37 = W*in
   wire signed [9:0] m54_37;
   assign m54_37 =10'b0;

   // m54_38 = W*in
   wire signed [9:0] m54_38;
   assign m54_38 ={ {3{neg54[5]}} , neg54 , {1{1'b0}} };

   // m54_39 = W*in
   wire signed [9:0] m54_39;
   assign m54_39 ={ {3{neg54[5]}} , neg54 , {1{1'b0}} };

   // m54_40 = W*in
   wire signed [9:0] m54_40;
   assign m54_40 =10'b0;

   // m54_41 = W*in
   wire signed [9:0] m54_41;
   assign m54_41 =10'b0;

   // m54_42 = W*in
   wire signed [9:0] m54_42;
   assign m54_42 =10'b0;

   // m54_43 = W*in
   wire signed [9:0] m54_43;
   assign m54_43 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_44 = W*in
   wire signed [9:0] m54_44;
   assign m54_44 =10'b0;

   // m54_45 = W*in
   wire signed [9:0] m54_45;
   assign m54_45 =10'b0;

   // m54_46 = W*in
   wire signed [9:0] m54_46;
   assign m54_46 =10'b0;

   // m54_47 = W*in
   wire signed [9:0] m54_47;
   assign m54_47 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_48 = W*in
   wire signed [9:0] m54_48;
   assign m54_48 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_49 = W*in
   wire signed [9:0] m54_49;
   assign m54_49 =10'b0;

   // m54_50 = W*in
   wire signed [9:0] m54_50;
   assign m54_50 ={ {3{neg54[5]}} , neg54 , {1{1'b0}} };

   // m54_51 = W*in
   wire signed [9:0] m54_51;
   assign m54_51 =10'b0;

   // m54_52 = W*in
   wire signed [9:0] m54_52;
   assign m54_52 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_53 = W*in
   wire signed [9:0] m54_53;
   assign m54_53 =10'b0;

   // m54_54 = W*in
   wire signed [9:0] m54_54;
   assign m54_54 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_55 = W*in
   wire signed [9:0] m54_55;
   assign m54_55 =10'b0;

   // m54_56 = W*in
   wire signed [9:0] m54_56;
   assign m54_56 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_57 = W*in
   wire signed [9:0] m54_57;
   assign m54_57 ={ {2{in54[5]}} , in54 , {2{1'b0}} };

   // m54_58 = W*in
   wire signed [9:0] m54_58;
   assign m54_58 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_59 = W*in
   wire signed [9:0] m54_59;
   assign m54_59 =10'b0;

   // m54_60 = W*in
   wire signed [9:0] m54_60;
   assign m54_60 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_61 = W*in
   wire signed [9:0] m54_61;
   assign m54_61 =10'b0;

   // m54_62 = W*in
   wire signed [9:0] m54_62;
   assign m54_62 ={ {3{in54[5]}} , in54 , {1{1'b0}} };

   // m54_63 = W*in
   wire signed [9:0] m54_63;
   assign m54_63 =10'b0;

   // m54_64 = W*in
   wire signed [9:0] m54_64;
   assign m54_64 ={ {3{neg54[5]}} , neg54 , {1{1'b0}} };

   // m54_65 = W*in
   wire signed [9:0] m54_65;
   assign m54_65 =10'b0;

   // m54_66 = W*in
   wire signed [9:0] m54_66;
   assign m54_66 =10'b0;

   // m54_67 = W*in
   wire signed [9:0] m54_67;
   assign m54_67 =10'b0;

   // m54_68 = W*in
   wire signed [9:0] m54_68;
   assign m54_68 =10'b0;

   // m54_69 = W*in
   wire signed [9:0] m54_69;
   assign m54_69 =10'b0;

   // m54_70 = W*in
   wire signed [9:0] m54_70;
   assign m54_70 =10'b0;

   // m54_71 = W*in
   wire signed [9:0] m54_71;
   assign m54_71 =10'b0;

   // m54_72 = W*in
   wire signed [9:0] m54_72;
   assign m54_72 =10'b0;

   // m54_73 = W*in
   wire signed [9:0] m54_73;
   assign m54_73 =10'b0;

   // m54_74 = W*in
   wire signed [9:0] m54_74;
   assign m54_74 =10'b0;

   // m54_75 = W*in
   wire signed [9:0] m54_75;
   assign m54_75 =10'b0;

   // m54_76 = W*in
   wire signed [9:0] m54_76;
   assign m54_76 =10'b0;

   // m54_77 = W*in
   wire signed [9:0] m54_77;
   assign m54_77 =10'b0;

   // m54_78 = W*in
   wire signed [9:0] m54_78;
   assign m54_78 ={ {3{neg54[5]}} , neg54 , {1{1'b0}} };

   // m54_79 = W*in
   wire signed [9:0] m54_79;
   assign m54_79 =10'b0;

   // m54_80 = W*in
   wire signed [9:0] m54_80;
   assign m54_80 =10'b0;

   // m54_81 = W*in
   wire signed [9:0] m54_81;
   assign m54_81 =10'b0;

   // m55_1 = W*in
   wire signed [9:0] m55_1;
   assign m55_1 =10'b0;

   // m55_2 = W*in
   wire signed [9:0] m55_2;
   assign m55_2 =10'b0;

   // m55_3 = W*in
   wire signed [9:0] m55_3;
   assign m55_3 ={ {3{in55[5]}} , in55 , {1{1'b0}} };

   // m55_4 = W*in
   wire signed [9:0] m55_4;
   assign m55_4 =10'b0;

   // m55_5 = W*in
   wire signed [9:0] m55_5;
   assign m55_5 =10'b0;

   // m55_6 = W*in
   wire signed [9:0] m55_6;
   assign m55_6 =10'b0;

   // m55_7 = W*in
   wire signed [9:0] m55_7;
   assign m55_7 =10'b0;

   // m55_8 = W*in
   wire signed [9:0] m55_8;
   assign m55_8 =10'b0;

   // m55_9 = W*in
   wire signed [9:0] m55_9;
   assign m55_9 =10'b0;

   // m55_10 = W*in
   wire signed [9:0] m55_10;
   assign m55_10 =10'b0;

   // m55_11 = W*in
   wire signed [9:0] m55_11;
   assign m55_11 =10'b0;

   // m55_12 = W*in
   wire signed [9:0] m55_12;
   assign m55_12 =10'b0;

   // m55_13 = W*in
   wire signed [9:0] m55_13;
   assign m55_13 =10'b0;

   // m55_14 = W*in
   wire signed [9:0] m55_14;
   assign m55_14 =10'b0;

   // m55_15 = W*in
   wire signed [9:0] m55_15;
   assign m55_15 =10'b0;

   // m55_16 = W*in
   wire signed [9:0] m55_16;
   assign m55_16 =10'b0;

   // m55_17 = W*in
   wire signed [9:0] m55_17;
   assign m55_17 =10'b0;

   // m55_18 = W*in
   wire signed [9:0] m55_18;
   assign m55_18 =10'b0;

   // m55_19 = W*in
   wire signed [9:0] m55_19;
   assign m55_19 =10'b0;

   // m55_20 = W*in
   wire signed [9:0] m55_20;
   assign m55_20 =10'b0;

   // m55_21 = W*in
   wire signed [9:0] m55_21;
   assign m55_21 =10'b0;

   // m55_22 = W*in
   wire signed [9:0] m55_22;
   assign m55_22 =10'b0;

   // m55_23 = W*in
   wire signed [9:0] m55_23;
   assign m55_23 =10'b0;

   // m55_24 = W*in
   wire signed [9:0] m55_24;
   assign m55_24 =10'b0;

   // m55_25 = W*in
   wire signed [9:0] m55_25;
   assign m55_25 =10'b0;

   // m55_26 = W*in
   wire signed [9:0] m55_26;
   assign m55_26 =10'b0;

   // m55_27 = W*in
   wire signed [9:0] m55_27;
   assign m55_27 =10'b0;

   // m55_28 = W*in
   wire signed [9:0] m55_28;
   assign m55_28 =10'b0;

   // m55_29 = W*in
   wire signed [9:0] m55_29;
   assign m55_29 =10'b0;

   // m55_30 = W*in
   wire signed [9:0] m55_30;
   assign m55_30 =10'b0;

   // m55_31 = W*in
   wire signed [9:0] m55_31;
   assign m55_31 =10'b0;

   // m55_32 = W*in
   wire signed [9:0] m55_32;
   assign m55_32 =10'b0;

   // m55_33 = W*in
   wire signed [9:0] m55_33;
   assign m55_33 =10'b0;

   // m55_34 = W*in
   wire signed [9:0] m55_34;
   assign m55_34 =10'b0;

   // m55_35 = W*in
   wire signed [9:0] m55_35;
   assign m55_35 =10'b0;

   // m55_36 = W*in
   wire signed [9:0] m55_36;
   assign m55_36 ={ {2{in55[5]}} , in55 , {2{1'b0}} };

   // m55_37 = W*in
   wire signed [9:0] m55_37;
   assign m55_37 =10'b0;

   // m55_38 = W*in
   wire signed [9:0] m55_38;
   assign m55_38 ={ {2{in55[5]}} , in55 , {2{1'b0}} };

   // m55_39 = W*in
   wire signed [9:0] m55_39;
   assign m55_39 =10'b0;

   // m55_40 = W*in
   wire signed [9:0] m55_40;
   assign m55_40 =10'b0;

   // m55_41 = W*in
   wire signed [9:0] m55_41;
   assign m55_41 ={ {3{in55[5]}} , in55 , {1{1'b0}} };

   // m55_42 = W*in
   wire signed [9:0] m55_42;
   assign m55_42 ={ {3{in55[5]}} , in55 , {1{1'b0}} };

   // m55_43 = W*in
   wire signed [9:0] m55_43;
   assign m55_43 =10'b0;

   // m55_44 = W*in
   wire signed [9:0] m55_44;
   assign m55_44 =10'b0;

   // m55_45 = W*in
   wire signed [9:0] m55_45;
   assign m55_45 =10'b0;

   // m55_46 = W*in
   wire signed [9:0] m55_46;
   assign m55_46 =10'b0;

   // m55_47 = W*in
   wire signed [9:0] m55_47;
   assign m55_47 =10'b0;

   // m55_48 = W*in
   wire signed [9:0] m55_48;
   assign m55_48 =10'b0;

   // m55_49 = W*in
   wire signed [9:0] m55_49;
   assign m55_49 =10'b0;

   // m55_50 = W*in
   wire signed [9:0] m55_50;
   assign m55_50 ={ {3{in55[5]}} , in55 , {1{1'b0}} };

   // m55_51 = W*in
   wire signed [9:0] m55_51;
   assign m55_51 =10'b0;

   // m55_52 = W*in
   wire signed [9:0] m55_52;
   assign m55_52 =10'b0;

   // m55_53 = W*in
   wire signed [9:0] m55_53;
   assign m55_53 =10'b0;

   // m55_54 = W*in
   wire signed [9:0] m55_54;
   assign m55_54 =10'b0;

   // m55_55 = W*in
   wire signed [9:0] m55_55;
   assign m55_55 =10'b0;

   // m55_56 = W*in
   wire signed [9:0] m55_56;
   assign m55_56 =10'b0;

   // m55_57 = W*in
   wire signed [9:0] m55_57;
   assign m55_57 =10'b0;

   // m55_58 = W*in
   wire signed [9:0] m55_58;
   assign m55_58 =10'b0;

   // m55_59 = W*in
   wire signed [9:0] m55_59;
   assign m55_59 =10'b0;

   // m55_60 = W*in
   wire signed [9:0] m55_60;
   assign m55_60 =10'b0;

   // m55_61 = W*in
   wire signed [9:0] m55_61;
   assign m55_61 =10'b0;

   // m55_62 = W*in
   wire signed [9:0] m55_62;
   assign m55_62 =10'b0;

   // m55_63 = W*in
   wire signed [9:0] m55_63;
   assign m55_63 =10'b0;

   // m55_64 = W*in
   wire signed [9:0] m55_64;
   assign m55_64 =10'b0;

   // m55_65 = W*in
   wire signed [9:0] m55_65;
   assign m55_65 =10'b0;

   // m55_66 = W*in
   wire signed [9:0] m55_66;
   assign m55_66 =10'b0;

   // m55_67 = W*in
   wire signed [9:0] m55_67;
   assign m55_67 =10'b0;

   // m55_68 = W*in
   wire signed [9:0] m55_68;
   assign m55_68 =10'b0;

   // m55_69 = W*in
   wire signed [9:0] m55_69;
   assign m55_69 =10'b0;

   // m55_70 = W*in
   wire signed [9:0] m55_70;
   assign m55_70 =10'b0;

   // m55_71 = W*in
   wire signed [9:0] m55_71;
   assign m55_71 =10'b0;

   // m55_72 = W*in
   wire signed [9:0] m55_72;
   assign m55_72 =10'b0;

   // m55_73 = W*in
   wire signed [9:0] m55_73;
   assign m55_73 ={ {3{in55[5]}} , in55 , {1{1'b0}} };

   // m55_74 = W*in
   wire signed [9:0] m55_74;
   assign m55_74 =10'b0;

   // m55_75 = W*in
   wire signed [9:0] m55_75;
   assign m55_75 =10'b0;

   // m55_76 = W*in
   wire signed [9:0] m55_76;
   assign m55_76 =10'b0;

   // m55_77 = W*in
   wire signed [9:0] m55_77;
   assign m55_77 =10'b0;

   // m55_78 = W*in
   wire signed [9:0] m55_78;
   assign m55_78 =10'b0;

   // m55_79 = W*in
   wire signed [9:0] m55_79;
   assign m55_79 =10'b0;

   // m55_80 = W*in
   wire signed [9:0] m55_80;
   assign m55_80 =10'b0;

   // m55_81 = W*in
   wire signed [9:0] m55_81;
   assign m55_81 =10'b0;

   // m56_1 = W*in
   wire signed [9:0] m56_1;
   assign m56_1 =10'b0;

   // m56_2 = W*in
   wire signed [9:0] m56_2;
   assign m56_2 =10'b0;

   // m56_3 = W*in
   wire signed [9:0] m56_3;
   assign m56_3 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_4 = W*in
   wire signed [9:0] m56_4;
   assign m56_4 =10'b0;

   // m56_5 = W*in
   wire signed [9:0] m56_5;
   assign m56_5 =10'b0;

   // m56_6 = W*in
   wire signed [9:0] m56_6;
   assign m56_6 =10'b0;

   // m56_7 = W*in
   wire signed [9:0] m56_7;
   assign m56_7 =10'b0;

   // m56_8 = W*in
   wire signed [9:0] m56_8;
   assign m56_8 =10'b0;

   // m56_9 = W*in
   wire signed [9:0] m56_9;
   assign m56_9 ={ {2{in56[5]}} , in56 , {2{1'b0}} };

   // m56_10 = W*in
   wire signed [9:0] m56_10;
   assign m56_10 =10'b0;

   // m56_11 = W*in
   wire signed [9:0] m56_11;
   assign m56_11 =10'b0;

   // m56_12 = W*in
   wire signed [9:0] m56_12;
   assign m56_12 =10'b0;

   // m56_13 = W*in
   wire signed [9:0] m56_13;
   assign m56_13 =10'b0;

   // m56_14 = W*in
   wire signed [9:0] m56_14;
   assign m56_14 =10'b0;

   // m56_15 = W*in
   wire signed [9:0] m56_15;
   assign m56_15 ={ {2{in56[5]}} , in56 , {2{1'b0}} };

   // m56_16 = W*in
   wire signed [9:0] m56_16;
   assign m56_16 =10'b0;

   // m56_17 = W*in
   wire signed [9:0] m56_17;
   assign m56_17 =10'b0;

   // m56_18 = W*in
   wire signed [9:0] m56_18;
   assign m56_18 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_19 = W*in
   wire signed [9:0] m56_19;
   assign m56_19 =10'b0;

   // m56_20 = W*in
   wire signed [9:0] m56_20;
   assign m56_20 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_21 = W*in
   wire signed [9:0] m56_21;
   assign m56_21 =10'b0;

   // m56_22 = W*in
   wire signed [9:0] m56_22;
   assign m56_22 =10'b0;

   // m56_23 = W*in
   wire signed [9:0] m56_23;
   assign m56_23 =10'b0;

   // m56_24 = W*in
   wire signed [9:0] m56_24;
   assign m56_24 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_25 = W*in
   wire signed [9:0] m56_25;
   assign m56_25 =10'b0;

   // m56_26 = W*in
   wire signed [9:0] m56_26;
   assign m56_26 =10'b0;

   // m56_27 = W*in
   wire signed [9:0] m56_27;
   assign m56_27 =10'b0;

   // m56_28 = W*in
   wire signed [9:0] m56_28;
   assign m56_28 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_29 = W*in
   wire signed [9:0] m56_29;
   assign m56_29 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_30 = W*in
   wire signed [9:0] m56_30;
   assign m56_30 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_31 = W*in
   wire signed [9:0] m56_31;
   assign m56_31 =10'b0;

   // m56_32 = W*in
   wire signed [9:0] m56_32;
   assign m56_32 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_33 = W*in
   wire signed [9:0] m56_33;
   assign m56_33 =10'b0;

   // m56_34 = W*in
   wire signed [9:0] m56_34;
   assign m56_34 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_35 = W*in
   wire signed [9:0] m56_35;
   assign m56_35 =10'b0;

   // m56_36 = W*in
   wire signed [9:0] m56_36;
   assign m56_36 =10'b0;

   // m56_37 = W*in
   wire signed [9:0] m56_37;
   assign m56_37 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_38 = W*in
   wire signed [9:0] m56_38;
   assign m56_38 =10'b0;

   // m56_39 = W*in
   wire signed [9:0] m56_39;
   assign m56_39 =10'b0;

   // m56_40 = W*in
   wire signed [9:0] m56_40;
   assign m56_40 =10'b0;

   // m56_41 = W*in
   wire signed [9:0] m56_41;
   assign m56_41 =10'b0;

   // m56_42 = W*in
   wire signed [9:0] m56_42;
   assign m56_42 ={ {2{in56[5]}} , in56 , {2{1'b0}} };

   // m56_43 = W*in
   wire signed [9:0] m56_43;
   assign m56_43 =10'b0;

   // m56_44 = W*in
   wire signed [9:0] m56_44;
   assign m56_44 =10'b0;

   // m56_45 = W*in
   wire signed [9:0] m56_45;
   assign m56_45 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_46 = W*in
   wire signed [9:0] m56_46;
   assign m56_46 =10'b0;

   // m56_47 = W*in
   wire signed [9:0] m56_47;
   assign m56_47 =10'b0;

   // m56_48 = W*in
   wire signed [9:0] m56_48;
   assign m56_48 =10'b0;

   // m56_49 = W*in
   wire signed [9:0] m56_49;
   assign m56_49 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_50 = W*in
   wire signed [9:0] m56_50;
   assign m56_50 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_51 = W*in
   wire signed [9:0] m56_51;
   assign m56_51 =10'b0;

   // m56_52 = W*in
   wire signed [9:0] m56_52;
   assign m56_52 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_53 = W*in
   wire signed [9:0] m56_53;
   assign m56_53 =10'b0;

   // m56_54 = W*in
   wire signed [9:0] m56_54;
   assign m56_54 =10'b0;

   // m56_55 = W*in
   wire signed [9:0] m56_55;
   assign m56_55 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_56 = W*in
   wire signed [9:0] m56_56;
   assign m56_56 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_57 = W*in
   wire signed [9:0] m56_57;
   assign m56_57 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_58 = W*in
   wire signed [9:0] m56_58;
   assign m56_58 =10'b0;

   // m56_59 = W*in
   wire signed [9:0] m56_59;
   assign m56_59 =10'b0;

   // m56_60 = W*in
   wire signed [9:0] m56_60;
   assign m56_60 =10'b0;

   // m56_61 = W*in
   wire signed [9:0] m56_61;
   assign m56_61 =10'b0;

   // m56_62 = W*in
   wire signed [9:0] m56_62;
   assign m56_62 ={ {2{in56[5]}} , in56 , {2{1'b0}} };

   // m56_63 = W*in
   wire signed [9:0] m56_63;
   assign m56_63 =10'b0;

   // m56_64 = W*in
   wire signed [9:0] m56_64;
   assign m56_64 =10'b0;

   // m56_65 = W*in
   wire signed [9:0] m56_65;
   assign m56_65 =10'b0;

   // m56_66 = W*in
   wire signed [9:0] m56_66;
   assign m56_66 ={ {2{in56[5]}} , in56 , {2{1'b0}} };

   // m56_67 = W*in
   wire signed [9:0] m56_67;
   assign m56_67 =10'b0;

   // m56_68 = W*in
   wire signed [9:0] m56_68;
   assign m56_68 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_69 = W*in
   wire signed [9:0] m56_69;
   assign m56_69 =10'b0;

   // m56_70 = W*in
   wire signed [9:0] m56_70;
   assign m56_70 =10'b0;

   // m56_71 = W*in
   wire signed [9:0] m56_71;
   assign m56_71 =10'b0;

   // m56_72 = W*in
   wire signed [9:0] m56_72;
   assign m56_72 =10'b0;

   // m56_73 = W*in
   wire signed [9:0] m56_73;
   assign m56_73 =10'b0;

   // m56_74 = W*in
   wire signed [9:0] m56_74;
   assign m56_74 =10'b0;

   // m56_75 = W*in
   wire signed [9:0] m56_75;
   assign m56_75 =10'b0;

   // m56_76 = W*in
   wire signed [9:0] m56_76;
   assign m56_76 =10'b0;

   // m56_77 = W*in
   wire signed [9:0] m56_77;
   assign m56_77 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_78 = W*in
   wire signed [9:0] m56_78;
   assign m56_78 =10'b0;

   // m56_79 = W*in
   wire signed [9:0] m56_79;
   assign m56_79 =10'b0;

   // m56_80 = W*in
   wire signed [9:0] m56_80;
   assign m56_80 =10'b0;

   // m56_81 = W*in
   wire signed [9:0] m56_81;
   assign m56_81 =10'b0;

   // m57_1 = W*in
   wire signed [9:0] m57_1;
   assign m57_1 =10'b0;

   // m57_2 = W*in
   wire signed [9:0] m57_2;
   assign m57_2 =10'b0;

   // m57_3 = W*in
   wire signed [9:0] m57_3;
   assign m57_3 =10'b0;

   // m57_4 = W*in
   wire signed [9:0] m57_4;
   assign m57_4 =10'b0;

   // m57_5 = W*in
   wire signed [9:0] m57_5;
   assign m57_5 =10'b0;

   // m57_6 = W*in
   wire signed [9:0] m57_6;
   assign m57_6 =10'b0;

   // m57_7 = W*in
   wire signed [9:0] m57_7;
   assign m57_7 =10'b0;

   // m57_8 = W*in
   wire signed [9:0] m57_8;
   assign m57_8 =10'b0;

   // m57_9 = W*in
   wire signed [9:0] m57_9;
   assign m57_9 =10'b0;

   // m57_10 = W*in
   wire signed [9:0] m57_10;
   assign m57_10 =10'b0;

   // m57_11 = W*in
   wire signed [9:0] m57_11;
   assign m57_11 =10'b0;

   // m57_12 = W*in
   wire signed [9:0] m57_12;
   assign m57_12 =10'b0;

   // m57_13 = W*in
   wire signed [9:0] m57_13;
   assign m57_13 =10'b0;

   // m57_14 = W*in
   wire signed [9:0] m57_14;
   assign m57_14 =10'b0;

   // m57_15 = W*in
   wire signed [9:0] m57_15;
   assign m57_15 =10'b0;

   // m57_16 = W*in
   wire signed [9:0] m57_16;
   assign m57_16 =10'b0;

   // m57_17 = W*in
   wire signed [9:0] m57_17;
   assign m57_17 =10'b0;

   // m57_18 = W*in
   wire signed [9:0] m57_18;
   assign m57_18 =10'b0;

   // m57_19 = W*in
   wire signed [9:0] m57_19;
   assign m57_19 =10'b0;

   // m57_20 = W*in
   wire signed [9:0] m57_20;
   assign m57_20 =10'b0;

   // m57_21 = W*in
   wire signed [9:0] m57_21;
   assign m57_21 =10'b0;

   // m57_22 = W*in
   wire signed [9:0] m57_22;
   assign m57_22 =10'b0;

   // m57_23 = W*in
   wire signed [9:0] m57_23;
   assign m57_23 =10'b0;

   // m57_24 = W*in
   wire signed [9:0] m57_24;
   assign m57_24 =10'b0;

   // m57_25 = W*in
   wire signed [9:0] m57_25;
   assign m57_25 =10'b0;

   // m57_26 = W*in
   wire signed [9:0] m57_26;
   assign m57_26 =10'b0;

   // m57_27 = W*in
   wire signed [9:0] m57_27;
   assign m57_27 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_28 = W*in
   wire signed [9:0] m57_28;
   assign m57_28 =10'b0;

   // m57_29 = W*in
   wire signed [9:0] m57_29;
   assign m57_29 =10'b0;

   // m57_30 = W*in
   wire signed [9:0] m57_30;
   assign m57_30 =10'b0;

   // m57_31 = W*in
   wire signed [9:0] m57_31;
   assign m57_31 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_32 = W*in
   wire signed [9:0] m57_32;
   assign m57_32 =10'b0;

   // m57_33 = W*in
   wire signed [9:0] m57_33;
   assign m57_33 =10'b0;

   // m57_34 = W*in
   wire signed [9:0] m57_34;
   assign m57_34 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_35 = W*in
   wire signed [9:0] m57_35;
   assign m57_35 =10'b0;

   // m57_36 = W*in
   wire signed [9:0] m57_36;
   assign m57_36 =10'b0;

   // m57_37 = W*in
   wire signed [9:0] m57_37;
   assign m57_37 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_38 = W*in
   wire signed [9:0] m57_38;
   assign m57_38 =10'b0;

   // m57_39 = W*in
   wire signed [9:0] m57_39;
   assign m57_39 =10'b0;

   // m57_40 = W*in
   wire signed [9:0] m57_40;
   assign m57_40 =10'b0;

   // m57_41 = W*in
   wire signed [9:0] m57_41;
   assign m57_41 =10'b0;

   // m57_42 = W*in
   wire signed [9:0] m57_42;
   assign m57_42 =10'b0;

   // m57_43 = W*in
   wire signed [9:0] m57_43;
   assign m57_43 =10'b0;

   // m57_44 = W*in
   wire signed [9:0] m57_44;
   assign m57_44 =10'b0;

   // m57_45 = W*in
   wire signed [9:0] m57_45;
   assign m57_45 =10'b0;

   // m57_46 = W*in
   wire signed [9:0] m57_46;
   assign m57_46 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_47 = W*in
   wire signed [9:0] m57_47;
   assign m57_47 =10'b0;

   // m57_48 = W*in
   wire signed [9:0] m57_48;
   assign m57_48 =10'b0;

   // m57_49 = W*in
   wire signed [9:0] m57_49;
   assign m57_49 =10'b0;

   // m57_50 = W*in
   wire signed [9:0] m57_50;
   assign m57_50 =10'b0;

   // m57_51 = W*in
   wire signed [9:0] m57_51;
   assign m57_51 =10'b0;

   // m57_52 = W*in
   wire signed [9:0] m57_52;
   assign m57_52 =10'b0;

   // m57_53 = W*in
   wire signed [9:0] m57_53;
   assign m57_53 =10'b0;

   // m57_54 = W*in
   wire signed [9:0] m57_54;
   assign m57_54 =10'b0;

   // m57_55 = W*in
   wire signed [9:0] m57_55;
   assign m57_55 =10'b0;

   // m57_56 = W*in
   wire signed [9:0] m57_56;
   assign m57_56 =10'b0;

   // m57_57 = W*in
   wire signed [9:0] m57_57;
   assign m57_57 =10'b0;

   // m57_58 = W*in
   wire signed [9:0] m57_58;
   assign m57_58 =10'b0;

   // m57_59 = W*in
   wire signed [9:0] m57_59;
   assign m57_59 =10'b0;

   // m57_60 = W*in
   wire signed [9:0] m57_60;
   assign m57_60 =10'b0;

   // m57_61 = W*in
   wire signed [9:0] m57_61;
   assign m57_61 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_62 = W*in
   wire signed [9:0] m57_62;
   assign m57_62 =10'b0;

   // m57_63 = W*in
   wire signed [9:0] m57_63;
   assign m57_63 =10'b0;

   // m57_64 = W*in
   wire signed [9:0] m57_64;
   assign m57_64 =10'b0;

   // m57_65 = W*in
   wire signed [9:0] m57_65;
   assign m57_65 =10'b0;

   // m57_66 = W*in
   wire signed [9:0] m57_66;
   assign m57_66 =10'b0;

   // m57_67 = W*in
   wire signed [9:0] m57_67;
   assign m57_67 =10'b0;

   // m57_68 = W*in
   wire signed [9:0] m57_68;
   assign m57_68 =10'b0;

   // m57_69 = W*in
   wire signed [9:0] m57_69;
   assign m57_69 =10'b0;

   // m57_70 = W*in
   wire signed [9:0] m57_70;
   assign m57_70 =10'b0;

   // m57_71 = W*in
   wire signed [9:0] m57_71;
   assign m57_71 =10'b0;

   // m57_72 = W*in
   wire signed [9:0] m57_72;
   assign m57_72 =10'b0;

   // m57_73 = W*in
   wire signed [9:0] m57_73;
   assign m57_73 =10'b0;

   // m57_74 = W*in
   wire signed [9:0] m57_74;
   assign m57_74 =10'b0;

   // m57_75 = W*in
   wire signed [9:0] m57_75;
   assign m57_75 =10'b0;

   // m57_76 = W*in
   wire signed [9:0] m57_76;
   assign m57_76 =10'b0;

   // m57_77 = W*in
   wire signed [9:0] m57_77;
   assign m57_77 =10'b0;

   // m57_78 = W*in
   wire signed [9:0] m57_78;
   assign m57_78 ={ {3{in57[5]}} , in57 , {1{1'b0}} };

   // m57_79 = W*in
   wire signed [9:0] m57_79;
   assign m57_79 =10'b0;

   // m57_80 = W*in
   wire signed [9:0] m57_80;
   assign m57_80 =10'b0;

   // m57_81 = W*in
   wire signed [9:0] m57_81;
   assign m57_81 =10'b0;

   // m58_1 = W*in
   wire signed [9:0] m58_1;
   assign m58_1 =10'b0;

   // m58_2 = W*in
   wire signed [9:0] m58_2;
   assign m58_2 =10'b0;

   // m58_3 = W*in
   wire signed [9:0] m58_3;
   assign m58_3 =10'b0;

   // m58_4 = W*in
   wire signed [9:0] m58_4;
   assign m58_4 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_5 = W*in
   wire signed [9:0] m58_5;
   assign m58_5 =10'b0;

   // m58_6 = W*in
   wire signed [9:0] m58_6;
   assign m58_6 =10'b0;

   // m58_7 = W*in
   wire signed [9:0] m58_7;
   assign m58_7 =10'b0;

   // m58_8 = W*in
   wire signed [9:0] m58_8;
   assign m58_8 =10'b0;

   // m58_9 = W*in
   wire signed [9:0] m58_9;
   assign m58_9 =10'b0;

   // m58_10 = W*in
   wire signed [9:0] m58_10;
   assign m58_10 =10'b0;

   // m58_11 = W*in
   wire signed [9:0] m58_11;
   assign m58_11 =10'b0;

   // m58_12 = W*in
   wire signed [9:0] m58_12;
   assign m58_12 =10'b0;

   // m58_13 = W*in
   wire signed [9:0] m58_13;
   assign m58_13 =10'b0;

   // m58_14 = W*in
   wire signed [9:0] m58_14;
   assign m58_14 =10'b0;

   // m58_15 = W*in
   wire signed [9:0] m58_15;
   assign m58_15 =10'b0;

   // m58_16 = W*in
   wire signed [9:0] m58_16;
   assign m58_16 =10'b0;

   // m58_17 = W*in
   wire signed [9:0] m58_17;
   assign m58_17 =10'b0;

   // m58_18 = W*in
   wire signed [9:0] m58_18;
   assign m58_18 =10'b0;

   // m58_19 = W*in
   wire signed [9:0] m58_19;
   assign m58_19 =10'b0;

   // m58_20 = W*in
   wire signed [9:0] m58_20;
   assign m58_20 =10'b0;

   // m58_21 = W*in
   wire signed [9:0] m58_21;
   assign m58_21 =10'b0;

   // m58_22 = W*in
   wire signed [9:0] m58_22;
   assign m58_22 =10'b0;

   // m58_23 = W*in
   wire signed [9:0] m58_23;
   assign m58_23 =10'b0;

   // m58_24 = W*in
   wire signed [9:0] m58_24;
   assign m58_24 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_25 = W*in
   wire signed [9:0] m58_25;
   assign m58_25 =10'b0;

   // m58_26 = W*in
   wire signed [9:0] m58_26;
   assign m58_26 =10'b0;

   // m58_27 = W*in
   wire signed [9:0] m58_27;
   assign m58_27 =10'b0;

   // m58_28 = W*in
   wire signed [9:0] m58_28;
   assign m58_28 =10'b0;

   // m58_29 = W*in
   wire signed [9:0] m58_29;
   assign m58_29 =10'b0;

   // m58_30 = W*in
   wire signed [9:0] m58_30;
   assign m58_30 =10'b0;

   // m58_31 = W*in
   wire signed [9:0] m58_31;
   assign m58_31 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_32 = W*in
   wire signed [9:0] m58_32;
   assign m58_32 =10'b0;

   // m58_33 = W*in
   wire signed [9:0] m58_33;
   assign m58_33 =10'b0;

   // m58_34 = W*in
   wire signed [9:0] m58_34;
   assign m58_34 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_35 = W*in
   wire signed [9:0] m58_35;
   assign m58_35 =10'b0;

   // m58_36 = W*in
   wire signed [9:0] m58_36;
   assign m58_36 =10'b0;

   // m58_37 = W*in
   wire signed [9:0] m58_37;
   assign m58_37 =10'b0;

   // m58_38 = W*in
   wire signed [9:0] m58_38;
   assign m58_38 =10'b0;

   // m58_39 = W*in
   wire signed [9:0] m58_39;
   assign m58_39 =10'b0;

   // m58_40 = W*in
   wire signed [9:0] m58_40;
   assign m58_40 =10'b0;

   // m58_41 = W*in
   wire signed [9:0] m58_41;
   assign m58_41 =10'b0;

   // m58_42 = W*in
   wire signed [9:0] m58_42;
   assign m58_42 ={ {3{neg58[5]}} , neg58 , {1{1'b0}} };

   // m58_43 = W*in
   wire signed [9:0] m58_43;
   assign m58_43 =10'b0;

   // m58_44 = W*in
   wire signed [9:0] m58_44;
   assign m58_44 =10'b0;

   // m58_45 = W*in
   wire signed [9:0] m58_45;
   assign m58_45 =10'b0;

   // m58_46 = W*in
   wire signed [9:0] m58_46;
   assign m58_46 =10'b0;

   // m58_47 = W*in
   wire signed [9:0] m58_47;
   assign m58_47 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_48 = W*in
   wire signed [9:0] m58_48;
   assign m58_48 =10'b0;

   // m58_49 = W*in
   wire signed [9:0] m58_49;
   assign m58_49 =10'b0;

   // m58_50 = W*in
   wire signed [9:0] m58_50;
   assign m58_50 =10'b0;

   // m58_51 = W*in
   wire signed [9:0] m58_51;
   assign m58_51 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_52 = W*in
   wire signed [9:0] m58_52;
   assign m58_52 =10'b0;

   // m58_53 = W*in
   wire signed [9:0] m58_53;
   assign m58_53 =10'b0;

   // m58_54 = W*in
   wire signed [9:0] m58_54;
   assign m58_54 =10'b0;

   // m58_55 = W*in
   wire signed [9:0] m58_55;
   assign m58_55 =10'b0;

   // m58_56 = W*in
   wire signed [9:0] m58_56;
   assign m58_56 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_57 = W*in
   wire signed [9:0] m58_57;
   assign m58_57 =10'b0;

   // m58_58 = W*in
   wire signed [9:0] m58_58;
   assign m58_58 =10'b0;

   // m58_59 = W*in
   wire signed [9:0] m58_59;
   assign m58_59 =10'b0;

   // m58_60 = W*in
   wire signed [9:0] m58_60;
   assign m58_60 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_61 = W*in
   wire signed [9:0] m58_61;
   assign m58_61 =10'b0;

   // m58_62 = W*in
   wire signed [9:0] m58_62;
   assign m58_62 =10'b0;

   // m58_63 = W*in
   wire signed [9:0] m58_63;
   assign m58_63 =10'b0;

   // m58_64 = W*in
   wire signed [9:0] m58_64;
   assign m58_64 =10'b0;

   // m58_65 = W*in
   wire signed [9:0] m58_65;
   assign m58_65 =10'b0;

   // m58_66 = W*in
   wire signed [9:0] m58_66;
   assign m58_66 =10'b0;

   // m58_67 = W*in
   wire signed [9:0] m58_67;
   assign m58_67 =10'b0;

   // m58_68 = W*in
   wire signed [9:0] m58_68;
   assign m58_68 =10'b0;

   // m58_69 = W*in
   wire signed [9:0] m58_69;
   assign m58_69 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_70 = W*in
   wire signed [9:0] m58_70;
   assign m58_70 =10'b0;

   // m58_71 = W*in
   wire signed [9:0] m58_71;
   assign m58_71 =10'b0;

   // m58_72 = W*in
   wire signed [9:0] m58_72;
   assign m58_72 =10'b0;

   // m58_73 = W*in
   wire signed [9:0] m58_73;
   assign m58_73 =10'b0;

   // m58_74 = W*in
   wire signed [9:0] m58_74;
   assign m58_74 =10'b0;

   // m58_75 = W*in
   wire signed [9:0] m58_75;
   assign m58_75 =10'b0;

   // m58_76 = W*in
   wire signed [9:0] m58_76;
   assign m58_76 =10'b0;

   // m58_77 = W*in
   wire signed [9:0] m58_77;
   assign m58_77 =10'b0;

   // m58_78 = W*in
   wire signed [9:0] m58_78;
   assign m58_78 =10'b0;

   // m58_79 = W*in
   wire signed [9:0] m58_79;
   assign m58_79 =10'b0;

   // m58_80 = W*in
   wire signed [9:0] m58_80;
   assign m58_80 =10'b0;

   // m58_81 = W*in
   wire signed [9:0] m58_81;
   assign m58_81 =10'b0;

   // m59_1 = W*in
   wire signed [9:0] m59_1;
   assign m59_1 =10'b0;

   // m59_2 = W*in
   wire signed [9:0] m59_2;
   assign m59_2 =10'b0;

   // m59_3 = W*in
   wire signed [9:0] m59_3;
   assign m59_3 ={ {3{in59[5]}} , in59 , {1{1'b0}} };

   // m59_4 = W*in
   wire signed [9:0] m59_4;
   assign m59_4 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_5 = W*in
   wire signed [9:0] m59_5;
   assign m59_5 =10'b0;

   // m59_6 = W*in
   wire signed [9:0] m59_6;
   assign m59_6 =10'b0;

   // m59_7 = W*in
   wire signed [9:0] m59_7;
   assign m59_7 =10'b0;

   // m59_8 = W*in
   wire signed [9:0] m59_8;
   assign m59_8 =10'b0;

   // m59_9 = W*in
   wire signed [9:0] m59_9;
   assign m59_9 =10'b0;

   // m59_10 = W*in
   wire signed [9:0] m59_10;
   assign m59_10 =10'b0;

   // m59_11 = W*in
   wire signed [9:0] m59_11;
   assign m59_11 =10'b0;

   // m59_12 = W*in
   wire signed [9:0] m59_12;
   assign m59_12 =10'b0;

   // m59_13 = W*in
   wire signed [9:0] m59_13;
   assign m59_13 =10'b0;

   // m59_14 = W*in
   wire signed [9:0] m59_14;
   assign m59_14 =10'b0;

   // m59_15 = W*in
   wire signed [9:0] m59_15;
   assign m59_15 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m59_16 = W*in
   wire signed [9:0] m59_16;
   assign m59_16 =10'b0;

   // m59_17 = W*in
   wire signed [9:0] m59_17;
   assign m59_17 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_18 = W*in
   wire signed [9:0] m59_18;
   assign m59_18 =10'b0;

   // m59_19 = W*in
   wire signed [9:0] m59_19;
   assign m59_19 =10'b0;

   // m59_20 = W*in
   wire signed [9:0] m59_20;
   assign m59_20 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_21 = W*in
   wire signed [9:0] m59_21;
   assign m59_21 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_22 = W*in
   wire signed [9:0] m59_22;
   assign m59_22 =10'b0;

   // m59_23 = W*in
   wire signed [9:0] m59_23;
   assign m59_23 =10'b0;

   // m59_24 = W*in
   wire signed [9:0] m59_24;
   assign m59_24 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_25 = W*in
   wire signed [9:0] m59_25;
   assign m59_25 =10'b0;

   // m59_26 = W*in
   wire signed [9:0] m59_26;
   assign m59_26 =10'b0;

   // m59_27 = W*in
   wire signed [9:0] m59_27;
   assign m59_27 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_28 = W*in
   wire signed [9:0] m59_28;
   assign m59_28 =10'b0;

   // m59_29 = W*in
   wire signed [9:0] m59_29;
   assign m59_29 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_30 = W*in
   wire signed [9:0] m59_30;
   assign m59_30 ={ {3{in59[5]}} , in59 , {1{1'b0}} };

   // m59_31 = W*in
   wire signed [9:0] m59_31;
   assign m59_31 =10'b0;

   // m59_32 = W*in
   wire signed [9:0] m59_32;
   assign m59_32 =10'b0;

   // m59_33 = W*in
   wire signed [9:0] m59_33;
   assign m59_33 =10'b0;

   // m59_34 = W*in
   wire signed [9:0] m59_34;
   assign m59_34 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_35 = W*in
   wire signed [9:0] m59_35;
   assign m59_35 =10'b0;

   // m59_36 = W*in
   wire signed [9:0] m59_36;
   assign m59_36 =10'b0;

   // m59_37 = W*in
   wire signed [9:0] m59_37;
   assign m59_37 =10'b0;

   // m59_38 = W*in
   wire signed [9:0] m59_38;
   assign m59_38 =10'b0;

   // m59_39 = W*in
   wire signed [9:0] m59_39;
   assign m59_39 ={ {3{in59[5]}} , in59 , {1{1'b0}} };

   // m59_40 = W*in
   wire signed [9:0] m59_40;
   assign m59_40 =10'b0;

   // m59_41 = W*in
   wire signed [9:0] m59_41;
   assign m59_41 =10'b0;

   // m59_42 = W*in
   wire signed [9:0] m59_42;
   assign m59_42 =10'b0;

   // m59_43 = W*in
   wire signed [9:0] m59_43;
   assign m59_43 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m59_44 = W*in
   wire signed [9:0] m59_44;
   assign m59_44 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m59_45 = W*in
   wire signed [9:0] m59_45;
   assign m59_45 =10'b0;

   // m59_46 = W*in
   wire signed [9:0] m59_46;
   assign m59_46 =10'b0;

   // m59_47 = W*in
   wire signed [9:0] m59_47;
   assign m59_47 =10'b0;

   // m59_48 = W*in
   wire signed [9:0] m59_48;
   assign m59_48 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_49 = W*in
   wire signed [9:0] m59_49;
   assign m59_49 =10'b0;

   // m59_50 = W*in
   wire signed [9:0] m59_50;
   assign m59_50 =10'b0;

   // m59_51 = W*in
   wire signed [9:0] m59_51;
   assign m59_51 =10'b0;

   // m59_52 = W*in
   wire signed [9:0] m59_52;
   assign m59_52 =10'b0;

   // m59_53 = W*in
   wire signed [9:0] m59_53;
   assign m59_53 =10'b0;

   // m59_54 = W*in
   wire signed [9:0] m59_54;
   assign m59_54 =10'b0;

   // m59_55 = W*in
   wire signed [9:0] m59_55;
   assign m59_55 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m59_56 = W*in
   wire signed [9:0] m59_56;
   assign m59_56 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_57 = W*in
   wire signed [9:0] m59_57;
   assign m59_57 ={ {3{in59[5]}} , in59 , {1{1'b0}} };

   // m59_58 = W*in
   wire signed [9:0] m59_58;
   assign m59_58 ={ {3{in59[5]}} , in59 , {1{1'b0}} };

   // m59_59 = W*in
   wire signed [9:0] m59_59;
   assign m59_59 =10'b0;

   // m59_60 = W*in
   wire signed [9:0] m59_60;
   assign m59_60 =10'b0;

   // m59_61 = W*in
   wire signed [9:0] m59_61;
   assign m59_61 =10'b0;

   // m59_62 = W*in
   wire signed [9:0] m59_62;
   assign m59_62 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m59_63 = W*in
   wire signed [9:0] m59_63;
   assign m59_63 =10'b0;

   // m59_64 = W*in
   wire signed [9:0] m59_64;
   assign m59_64 =10'b0;

   // m59_65 = W*in
   wire signed [9:0] m59_65;
   assign m59_65 =10'b0;

   // m59_66 = W*in
   wire signed [9:0] m59_66;
   assign m59_66 =10'b0;

   // m59_67 = W*in
   wire signed [9:0] m59_67;
   assign m59_67 =10'b0;

   // m59_68 = W*in
   wire signed [9:0] m59_68;
   assign m59_68 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_69 = W*in
   wire signed [9:0] m59_69;
   assign m59_69 =10'b0;

   // m59_70 = W*in
   wire signed [9:0] m59_70;
   assign m59_70 =10'b0;

   // m59_71 = W*in
   wire signed [9:0] m59_71;
   assign m59_71 =10'b0;

   // m59_72 = W*in
   wire signed [9:0] m59_72;
   assign m59_72 =10'b0;

   // m59_73 = W*in
   wire signed [9:0] m59_73;
   assign m59_73 =10'b0;

   // m59_74 = W*in
   wire signed [9:0] m59_74;
   assign m59_74 =10'b0;

   // m59_75 = W*in
   wire signed [9:0] m59_75;
   assign m59_75 =10'b0;

   // m59_76 = W*in
   wire signed [9:0] m59_76;
   assign m59_76 =10'b0;

   // m59_77 = W*in
   wire signed [9:0] m59_77;
   assign m59_77 ={ {3{neg59[5]}} , neg59 , {1{1'b0}} };

   // m59_78 = W*in
   wire signed [9:0] m59_78;
   assign m59_78 =10'b0;

   // m59_79 = W*in
   wire signed [9:0] m59_79;
   assign m59_79 =10'b0;

   // m59_80 = W*in
   wire signed [9:0] m59_80;
   assign m59_80 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m59_81 = W*in
   wire signed [9:0] m59_81;
   assign m59_81 ={ {2{in59[5]}} , in59 , {2{1'b0}} };

   // m60_1 = W*in
   wire signed [9:0] m60_1;
   assign m60_1 =10'b0;

   // m60_2 = W*in
   wire signed [9:0] m60_2;
   assign m60_2 =10'b0;

   // m60_3 = W*in
   wire signed [9:0] m60_3;
   assign m60_3 =10'b0;

   // m60_4 = W*in
   wire signed [9:0] m60_4;
   assign m60_4 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_5 = W*in
   wire signed [9:0] m60_5;
   assign m60_5 =10'b0;

   // m60_6 = W*in
   wire signed [9:0] m60_6;
   assign m60_6 =10'b0;

   // m60_7 = W*in
   wire signed [9:0] m60_7;
   assign m60_7 =10'b0;

   // m60_8 = W*in
   wire signed [9:0] m60_8;
   assign m60_8 =10'b0;

   // m60_9 = W*in
   wire signed [9:0] m60_9;
   assign m60_9 =10'b0;

   // m60_10 = W*in
   wire signed [9:0] m60_10;
   assign m60_10 =10'b0;

   // m60_11 = W*in
   wire signed [9:0] m60_11;
   assign m60_11 =10'b0;

   // m60_12 = W*in
   wire signed [9:0] m60_12;
   assign m60_12 =10'b0;

   // m60_13 = W*in
   wire signed [9:0] m60_13;
   assign m60_13 =10'b0;

   // m60_14 = W*in
   wire signed [9:0] m60_14;
   assign m60_14 =10'b0;

   // m60_15 = W*in
   wire signed [9:0] m60_15;
   assign m60_15 =10'b0;

   // m60_16 = W*in
   wire signed [9:0] m60_16;
   assign m60_16 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_17 = W*in
   wire signed [9:0] m60_17;
   assign m60_17 =10'b0;

   // m60_18 = W*in
   wire signed [9:0] m60_18;
   assign m60_18 =10'b0;

   // m60_19 = W*in
   wire signed [9:0] m60_19;
   assign m60_19 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_20 = W*in
   wire signed [9:0] m60_20;
   assign m60_20 =10'b0;

   // m60_21 = W*in
   wire signed [9:0] m60_21;
   assign m60_21 =10'b0;

   // m60_22 = W*in
   wire signed [9:0] m60_22;
   assign m60_22 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_23 = W*in
   wire signed [9:0] m60_23;
   assign m60_23 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_24 = W*in
   wire signed [9:0] m60_24;
   assign m60_24 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_25 = W*in
   wire signed [9:0] m60_25;
   assign m60_25 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_26 = W*in
   wire signed [9:0] m60_26;
   assign m60_26 =10'b0;

   // m60_27 = W*in
   wire signed [9:0] m60_27;
   assign m60_27 =10'b0;

   // m60_28 = W*in
   wire signed [9:0] m60_28;
   assign m60_28 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_29 = W*in
   wire signed [9:0] m60_29;
   assign m60_29 =10'b0;

   // m60_30 = W*in
   wire signed [9:0] m60_30;
   assign m60_30 ={ {2{in60[5]}} , in60 , {2{1'b0}} };

   // m60_31 = W*in
   wire signed [9:0] m60_31;
   assign m60_31 =10'b0;

   // m60_32 = W*in
   wire signed [9:0] m60_32;
   assign m60_32 ={ {2{in60[5]}} , in60 , {2{1'b0}} };

   // m60_33 = W*in
   wire signed [9:0] m60_33;
   assign m60_33 =10'b0;

   // m60_34 = W*in
   wire signed [9:0] m60_34;
   assign m60_34 =10'b0;

   // m60_35 = W*in
   wire signed [9:0] m60_35;
   assign m60_35 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_36 = W*in
   wire signed [9:0] m60_36;
   assign m60_36 =10'b0;

   // m60_37 = W*in
   wire signed [9:0] m60_37;
   assign m60_37 =10'b0;

   // m60_38 = W*in
   wire signed [9:0] m60_38;
   assign m60_38 =10'b0;

   // m60_39 = W*in
   wire signed [9:0] m60_39;
   assign m60_39 =10'b0;

   // m60_40 = W*in
   wire signed [9:0] m60_40;
   assign m60_40 =10'b0;

   // m60_41 = W*in
   wire signed [9:0] m60_41;
   assign m60_41 =10'b0;

   // m60_42 = W*in
   wire signed [9:0] m60_42;
   assign m60_42 =10'b0;

   // m60_43 = W*in
   wire signed [9:0] m60_43;
   assign m60_43 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_44 = W*in
   wire signed [9:0] m60_44;
   assign m60_44 =10'b0;

   // m60_45 = W*in
   wire signed [9:0] m60_45;
   assign m60_45 =10'b0;

   // m60_46 = W*in
   wire signed [9:0] m60_46;
   assign m60_46 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_47 = W*in
   wire signed [9:0] m60_47;
   assign m60_47 =10'b0;

   // m60_48 = W*in
   wire signed [9:0] m60_48;
   assign m60_48 =10'b0;

   // m60_49 = W*in
   wire signed [9:0] m60_49;
   assign m60_49 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_50 = W*in
   wire signed [9:0] m60_50;
   assign m60_50 =10'b0;

   // m60_51 = W*in
   wire signed [9:0] m60_51;
   assign m60_51 =10'b0;

   // m60_52 = W*in
   wire signed [9:0] m60_52;
   assign m60_52 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_53 = W*in
   wire signed [9:0] m60_53;
   assign m60_53 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_54 = W*in
   wire signed [9:0] m60_54;
   assign m60_54 =10'b0;

   // m60_55 = W*in
   wire signed [9:0] m60_55;
   assign m60_55 =10'b0;

   // m60_56 = W*in
   wire signed [9:0] m60_56;
   assign m60_56 =10'b0;

   // m60_57 = W*in
   wire signed [9:0] m60_57;
   assign m60_57 =10'b0;

   // m60_58 = W*in
   wire signed [9:0] m60_58;
   assign m60_58 =10'b0;

   // m60_59 = W*in
   wire signed [9:0] m60_59;
   assign m60_59 =10'b0;

   // m60_60 = W*in
   wire signed [9:0] m60_60;
   assign m60_60 =10'b0;

   // m60_61 = W*in
   wire signed [9:0] m60_61;
   assign m60_61 =10'b0;

   // m60_62 = W*in
   wire signed [9:0] m60_62;
   assign m60_62 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_63 = W*in
   wire signed [9:0] m60_63;
   assign m60_63 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_64 = W*in
   wire signed [9:0] m60_64;
   assign m60_64 =10'b0;

   // m60_65 = W*in
   wire signed [9:0] m60_65;
   assign m60_65 =10'b0;

   // m60_66 = W*in
   wire signed [9:0] m60_66;
   assign m60_66 =10'b0;

   // m60_67 = W*in
   wire signed [9:0] m60_67;
   assign m60_67 =10'b0;

   // m60_68 = W*in
   wire signed [9:0] m60_68;
   assign m60_68 =10'b0;

   // m60_69 = W*in
   wire signed [9:0] m60_69;
   assign m60_69 =10'b0;

   // m60_70 = W*in
   wire signed [9:0] m60_70;
   assign m60_70 =10'b0;

   // m60_71 = W*in
   wire signed [9:0] m60_71;
   assign m60_71 =10'b0;

   // m60_72 = W*in
   wire signed [9:0] m60_72;
   assign m60_72 =10'b0;

   // m60_73 = W*in
   wire signed [9:0] m60_73;
   assign m60_73 =10'b0;

   // m60_74 = W*in
   wire signed [9:0] m60_74;
   assign m60_74 =10'b0;

   // m60_75 = W*in
   wire signed [9:0] m60_75;
   assign m60_75 =10'b0;

   // m60_76 = W*in
   wire signed [9:0] m60_76;
   assign m60_76 =10'b0;

   // m60_77 = W*in
   wire signed [9:0] m60_77;
   assign m60_77 ={ {3{neg60[5]}} , neg60 , {1{1'b0}} };

   // m60_78 = W*in
   wire signed [9:0] m60_78;
   assign m60_78 =10'b0;

   // m60_79 = W*in
   wire signed [9:0] m60_79;
   assign m60_79 ={ {2{in60[5]}} , in60 , {2{1'b0}} };

   // m60_80 = W*in
   wire signed [9:0] m60_80;
   assign m60_80 =10'b0;

   // m60_81 = W*in
   wire signed [9:0] m60_81;
   assign m60_81 =10'b0;

   // m61_1 = W*in
   wire signed [9:0] m61_1;
   assign m61_1 =10'b0;

   // m61_2 = W*in
   wire signed [9:0] m61_2;
   assign m61_2 =10'b0;

   // m61_3 = W*in
   wire signed [9:0] m61_3;
   assign m61_3 =10'b0;

   // m61_4 = W*in
   wire signed [9:0] m61_4;
   assign m61_4 =10'b0;

   // m61_5 = W*in
   wire signed [9:0] m61_5;
   assign m61_5 =10'b0;

   // m61_6 = W*in
   wire signed [9:0] m61_6;
   assign m61_6 =10'b0;

   // m61_7 = W*in
   wire signed [9:0] m61_7;
   assign m61_7 =10'b0;

   // m61_8 = W*in
   wire signed [9:0] m61_8;
   assign m61_8 =10'b0;

   // m61_9 = W*in
   wire signed [9:0] m61_9;
   assign m61_9 =10'b0;

   // m61_10 = W*in
   wire signed [9:0] m61_10;
   assign m61_10 =10'b0;

   // m61_11 = W*in
   wire signed [9:0] m61_11;
   assign m61_11 =10'b0;

   // m61_12 = W*in
   wire signed [9:0] m61_12;
   assign m61_12 =10'b0;

   // m61_13 = W*in
   wire signed [9:0] m61_13;
   assign m61_13 =10'b0;

   // m61_14 = W*in
   wire signed [9:0] m61_14;
   assign m61_14 =10'b0;

   // m61_15 = W*in
   wire signed [9:0] m61_15;
   assign m61_15 ={ {2{in61[5]}} , in61 , {2{1'b0}} };

   // m61_16 = W*in
   wire signed [9:0] m61_16;
   assign m61_16 ={ {2{in61[5]}} , in61 , {2{1'b0}} };

   // m61_17 = W*in
   wire signed [9:0] m61_17;
   assign m61_17 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_18 = W*in
   wire signed [9:0] m61_18;
   assign m61_18 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_19 = W*in
   wire signed [9:0] m61_19;
   assign m61_19 =10'b0;

   // m61_20 = W*in
   wire signed [9:0] m61_20;
   assign m61_20 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_21 = W*in
   wire signed [9:0] m61_21;
   assign m61_21 =10'b0;

   // m61_22 = W*in
   wire signed [9:0] m61_22;
   assign m61_22 =10'b0;

   // m61_23 = W*in
   wire signed [9:0] m61_23;
   assign m61_23 =10'b0;

   // m61_24 = W*in
   wire signed [9:0] m61_24;
   assign m61_24 =10'b0;

   // m61_25 = W*in
   wire signed [9:0] m61_25;
   assign m61_25 =10'b0;

   // m61_26 = W*in
   wire signed [9:0] m61_26;
   assign m61_26 =10'b0;

   // m61_27 = W*in
   wire signed [9:0] m61_27;
   assign m61_27 =10'b0;

   // m61_28 = W*in
   wire signed [9:0] m61_28;
   assign m61_28 =10'b0;

   // m61_29 = W*in
   wire signed [9:0] m61_29;
   assign m61_29 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_30 = W*in
   wire signed [9:0] m61_30;
   assign m61_30 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_31 = W*in
   wire signed [9:0] m61_31;
   assign m61_31 =10'b0;

   // m61_32 = W*in
   wire signed [9:0] m61_32;
   assign m61_32 ={ {2{in61[5]}} , in61 , {2{1'b0}} };

   // m61_33 = W*in
   wire signed [9:0] m61_33;
   assign m61_33 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_34 = W*in
   wire signed [9:0] m61_34;
   assign m61_34 =10'b0;

   // m61_35 = W*in
   wire signed [9:0] m61_35;
   assign m61_35 =10'b0;

   // m61_36 = W*in
   wire signed [9:0] m61_36;
   assign m61_36 =10'b0;

   // m61_37 = W*in
   wire signed [9:0] m61_37;
   assign m61_37 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_38 = W*in
   wire signed [9:0] m61_38;
   assign m61_38 =10'b0;

   // m61_39 = W*in
   wire signed [9:0] m61_39;
   assign m61_39 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_40 = W*in
   wire signed [9:0] m61_40;
   assign m61_40 ={ {2{in61[5]}} , in61 , {2{1'b0}} };

   // m61_41 = W*in
   wire signed [9:0] m61_41;
   assign m61_41 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_42 = W*in
   wire signed [9:0] m61_42;
   assign m61_42 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_43 = W*in
   wire signed [9:0] m61_43;
   assign m61_43 =10'b0;

   // m61_44 = W*in
   wire signed [9:0] m61_44;
   assign m61_44 =10'b0;

   // m61_45 = W*in
   wire signed [9:0] m61_45;
   assign m61_45 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_46 = W*in
   wire signed [9:0] m61_46;
   assign m61_46 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_47 = W*in
   wire signed [9:0] m61_47;
   assign m61_47 =10'b0;

   // m61_48 = W*in
   wire signed [9:0] m61_48;
   assign m61_48 =10'b0;

   // m61_49 = W*in
   wire signed [9:0] m61_49;
   assign m61_49 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_50 = W*in
   wire signed [9:0] m61_50;
   assign m61_50 =10'b0;

   // m61_51 = W*in
   wire signed [9:0] m61_51;
   assign m61_51 =10'b0;

   // m61_52 = W*in
   wire signed [9:0] m61_52;
   assign m61_52 =10'b0;

   // m61_53 = W*in
   wire signed [9:0] m61_53;
   assign m61_53 =10'b0;

   // m61_54 = W*in
   wire signed [9:0] m61_54;
   assign m61_54 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_55 = W*in
   wire signed [9:0] m61_55;
   assign m61_55 =10'b0;

   // m61_56 = W*in
   wire signed [9:0] m61_56;
   assign m61_56 =10'b0;

   // m61_57 = W*in
   wire signed [9:0] m61_57;
   assign m61_57 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_58 = W*in
   wire signed [9:0] m61_58;
   assign m61_58 =10'b0;

   // m61_59 = W*in
   wire signed [9:0] m61_59;
   assign m61_59 =10'b0;

   // m61_60 = W*in
   wire signed [9:0] m61_60;
   assign m61_60 =10'b0;

   // m61_61 = W*in
   wire signed [9:0] m61_61;
   assign m61_61 =10'b0;

   // m61_62 = W*in
   wire signed [9:0] m61_62;
   assign m61_62 ={ {2{in61[5]}} , in61 , {2{1'b0}} };

   // m61_63 = W*in
   wire signed [9:0] m61_63;
   assign m61_63 =10'b0;

   // m61_64 = W*in
   wire signed [9:0] m61_64;
   assign m61_64 =10'b0;

   // m61_65 = W*in
   wire signed [9:0] m61_65;
   assign m61_65 =10'b0;

   // m61_66 = W*in
   wire signed [9:0] m61_66;
   assign m61_66 =10'b0;

   // m61_67 = W*in
   wire signed [9:0] m61_67;
   assign m61_67 =10'b0;

   // m61_68 = W*in
   wire signed [9:0] m61_68;
   assign m61_68 =10'b0;

   // m61_69 = W*in
   wire signed [9:0] m61_69;
   assign m61_69 =10'b0;

   // m61_70 = W*in
   wire signed [9:0] m61_70;
   assign m61_70 =10'b0;

   // m61_71 = W*in
   wire signed [9:0] m61_71;
   assign m61_71 =10'b0;

   // m61_72 = W*in
   wire signed [9:0] m61_72;
   assign m61_72 =10'b0;

   // m61_73 = W*in
   wire signed [9:0] m61_73;
   assign m61_73 ={ {3{neg61[5]}} , neg61 , {1{1'b0}} };

   // m61_74 = W*in
   wire signed [9:0] m61_74;
   assign m61_74 =10'b0;

   // m61_75 = W*in
   wire signed [9:0] m61_75;
   assign m61_75 =10'b0;

   // m61_76 = W*in
   wire signed [9:0] m61_76;
   assign m61_76 =10'b0;

   // m61_77 = W*in
   wire signed [9:0] m61_77;
   assign m61_77 =10'b0;

   // m61_78 = W*in
   wire signed [9:0] m61_78;
   assign m61_78 =10'b0;

   // m61_79 = W*in
   wire signed [9:0] m61_79;
   assign m61_79 ={ {3{in61[5]}} , in61 , {1{1'b0}} };

   // m61_80 = W*in
   wire signed [9:0] m61_80;
   assign m61_80 =10'b0;

   // m61_81 = W*in
   wire signed [9:0] m61_81;
   assign m61_81 =10'b0;

   // m62_1 = W*in
   wire signed [9:0] m62_1;
   assign m62_1 =10'b0;

   // m62_2 = W*in
   wire signed [9:0] m62_2;
   assign m62_2 =10'b0;

   // m62_3 = W*in
   wire signed [9:0] m62_3;
   assign m62_3 ={ {3{neg62[5]}} , neg62 , {1{1'b0}} };

   // m62_4 = W*in
   wire signed [9:0] m62_4;
   assign m62_4 =10'b0;

   // m62_5 = W*in
   wire signed [9:0] m62_5;
   assign m62_5 =10'b0;

   // m62_6 = W*in
   wire signed [9:0] m62_6;
   assign m62_6 =10'b0;

   // m62_7 = W*in
   wire signed [9:0] m62_7;
   assign m62_7 =10'b0;

   // m62_8 = W*in
   wire signed [9:0] m62_8;
   assign m62_8 =10'b0;

   // m62_9 = W*in
   wire signed [9:0] m62_9;
   assign m62_9 =10'b0;

   // m62_10 = W*in
   wire signed [9:0] m62_10;
   assign m62_10 =10'b0;

   // m62_11 = W*in
   wire signed [9:0] m62_11;
   assign m62_11 =10'b0;

   // m62_12 = W*in
   wire signed [9:0] m62_12;
   assign m62_12 =10'b0;

   // m62_13 = W*in
   wire signed [9:0] m62_13;
   assign m62_13 =10'b0;

   // m62_14 = W*in
   wire signed [9:0] m62_14;
   assign m62_14 =10'b0;

   // m62_15 = W*in
   wire signed [9:0] m62_15;
   assign m62_15 =10'b0;

   // m62_16 = W*in
   wire signed [9:0] m62_16;
   assign m62_16 =10'b0;

   // m62_17 = W*in
   wire signed [9:0] m62_17;
   assign m62_17 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_18 = W*in
   wire signed [9:0] m62_18;
   assign m62_18 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_19 = W*in
   wire signed [9:0] m62_19;
   assign m62_19 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_20 = W*in
   wire signed [9:0] m62_20;
   assign m62_20 =10'b0;

   // m62_21 = W*in
   wire signed [9:0] m62_21;
   assign m62_21 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_22 = W*in
   wire signed [9:0] m62_22;
   assign m62_22 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_23 = W*in
   wire signed [9:0] m62_23;
   assign m62_23 =10'b0;

   // m62_24 = W*in
   wire signed [9:0] m62_24;
   assign m62_24 =10'b0;

   // m62_25 = W*in
   wire signed [9:0] m62_25;
   assign m62_25 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_26 = W*in
   wire signed [9:0] m62_26;
   assign m62_26 =10'b0;

   // m62_27 = W*in
   wire signed [9:0] m62_27;
   assign m62_27 =10'b0;

   // m62_28 = W*in
   wire signed [9:0] m62_28;
   assign m62_28 =10'b0;

   // m62_29 = W*in
   wire signed [9:0] m62_29;
   assign m62_29 =10'b0;

   // m62_30 = W*in
   wire signed [9:0] m62_30;
   assign m62_30 ={ {3{neg62[5]}} , neg62 , {1{1'b0}} };

   // m62_31 = W*in
   wire signed [9:0] m62_31;
   assign m62_31 =10'b0;

   // m62_32 = W*in
   wire signed [9:0] m62_32;
   assign m62_32 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_33 = W*in
   wire signed [9:0] m62_33;
   assign m62_33 =10'b0;

   // m62_34 = W*in
   wire signed [9:0] m62_34;
   assign m62_34 =10'b0;

   // m62_35 = W*in
   wire signed [9:0] m62_35;
   assign m62_35 =10'b0;

   // m62_36 = W*in
   wire signed [9:0] m62_36;
   assign m62_36 ={ {3{neg62[5]}} , neg62 , {1{1'b0}} };

   // m62_37 = W*in
   wire signed [9:0] m62_37;
   assign m62_37 =10'b0;

   // m62_38 = W*in
   wire signed [9:0] m62_38;
   assign m62_38 =10'b0;

   // m62_39 = W*in
   wire signed [9:0] m62_39;
   assign m62_39 =10'b0;

   // m62_40 = W*in
   wire signed [9:0] m62_40;
   assign m62_40 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_41 = W*in
   wire signed [9:0] m62_41;
   assign m62_41 =10'b0;

   // m62_42 = W*in
   wire signed [9:0] m62_42;
   assign m62_42 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_43 = W*in
   wire signed [9:0] m62_43;
   assign m62_43 =10'b0;

   // m62_44 = W*in
   wire signed [9:0] m62_44;
   assign m62_44 =10'b0;

   // m62_45 = W*in
   wire signed [9:0] m62_45;
   assign m62_45 =10'b0;

   // m62_46 = W*in
   wire signed [9:0] m62_46;
   assign m62_46 =10'b0;

   // m62_47 = W*in
   wire signed [9:0] m62_47;
   assign m62_47 =10'b0;

   // m62_48 = W*in
   wire signed [9:0] m62_48;
   assign m62_48 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_49 = W*in
   wire signed [9:0] m62_49;
   assign m62_49 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_50 = W*in
   wire signed [9:0] m62_50;
   assign m62_50 =10'b0;

   // m62_51 = W*in
   wire signed [9:0] m62_51;
   assign m62_51 =10'b0;

   // m62_52 = W*in
   wire signed [9:0] m62_52;
   assign m62_52 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_53 = W*in
   wire signed [9:0] m62_53;
   assign m62_53 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_54 = W*in
   wire signed [9:0] m62_54;
   assign m62_54 =10'b0;

   // m62_55 = W*in
   wire signed [9:0] m62_55;
   assign m62_55 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_56 = W*in
   wire signed [9:0] m62_56;
   assign m62_56 =10'b0;

   // m62_57 = W*in
   wire signed [9:0] m62_57;
   assign m62_57 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_58 = W*in
   wire signed [9:0] m62_58;
   assign m62_58 =10'b0;

   // m62_59 = W*in
   wire signed [9:0] m62_59;
   assign m62_59 =10'b0;

   // m62_60 = W*in
   wire signed [9:0] m62_60;
   assign m62_60 =10'b0;

   // m62_61 = W*in
   wire signed [9:0] m62_61;
   assign m62_61 =10'b0;

   // m62_62 = W*in
   wire signed [9:0] m62_62;
   assign m62_62 =10'b0;

   // m62_63 = W*in
   wire signed [9:0] m62_63;
   assign m62_63 =10'b0;

   // m62_64 = W*in
   wire signed [9:0] m62_64;
   assign m62_64 =10'b0;

   // m62_65 = W*in
   wire signed [9:0] m62_65;
   assign m62_65 =10'b0;

   // m62_66 = W*in
   wire signed [9:0] m62_66;
   assign m62_66 =10'b0;

   // m62_67 = W*in
   wire signed [9:0] m62_67;
   assign m62_67 =10'b0;

   // m62_68 = W*in
   wire signed [9:0] m62_68;
   assign m62_68 =10'b0;

   // m62_69 = W*in
   wire signed [9:0] m62_69;
   assign m62_69 =10'b0;

   // m62_70 = W*in
   wire signed [9:0] m62_70;
   assign m62_70 ={ {3{in62[5]}} , in62 , {1{1'b0}} };

   // m62_71 = W*in
   wire signed [9:0] m62_71;
   assign m62_71 =10'b0;

   // m62_72 = W*in
   wire signed [9:0] m62_72;
   assign m62_72 =10'b0;

   // m62_73 = W*in
   wire signed [9:0] m62_73;
   assign m62_73 =10'b0;

   // m62_74 = W*in
   wire signed [9:0] m62_74;
   assign m62_74 =10'b0;

   // m62_75 = W*in
   wire signed [9:0] m62_75;
   assign m62_75 =10'b0;

   // m62_76 = W*in
   wire signed [9:0] m62_76;
   assign m62_76 =10'b0;

   // m62_77 = W*in
   wire signed [9:0] m62_77;
   assign m62_77 =10'b0;

   // m62_78 = W*in
   wire signed [9:0] m62_78;
   assign m62_78 =10'b0;

   // m62_79 = W*in
   wire signed [9:0] m62_79;
   assign m62_79 =10'b0;

   // m62_80 = W*in
   wire signed [9:0] m62_80;
   assign m62_80 =10'b0;

   // m62_81 = W*in
   wire signed [9:0] m62_81;
   assign m62_81 =10'b0;

   // m63_1 = W*in
   wire signed [9:0] m63_1;
   assign m63_1 =10'b0;

   // m63_2 = W*in
   wire signed [9:0] m63_2;
   assign m63_2 =10'b0;

   // m63_3 = W*in
   wire signed [9:0] m63_3;
   assign m63_3 =10'b0;

   // m63_4 = W*in
   wire signed [9:0] m63_4;
   assign m63_4 ={ {2{in63[5]}} , in63 , {2{1'b0}} };

   // m63_5 = W*in
   wire signed [9:0] m63_5;
   assign m63_5 =10'b0;

   // m63_6 = W*in
   wire signed [9:0] m63_6;
   assign m63_6 =10'b0;

   // m63_7 = W*in
   wire signed [9:0] m63_7;
   assign m63_7 =10'b0;

   // m63_8 = W*in
   wire signed [9:0] m63_8;
   assign m63_8 =10'b0;

   // m63_9 = W*in
   wire signed [9:0] m63_9;
   assign m63_9 =10'b0;

   // m63_10 = W*in
   wire signed [9:0] m63_10;
   assign m63_10 ={ {2{in63[5]}} , in63 , {2{1'b0}} };

   // m63_11 = W*in
   wire signed [9:0] m63_11;
   assign m63_11 =10'b0;

   // m63_12 = W*in
   wire signed [9:0] m63_12;
   assign m63_12 ={ {2{in63[5]}} , in63 , {2{1'b0}} };

   // m63_13 = W*in
   wire signed [9:0] m63_13;
   assign m63_13 =10'b0;

   // m63_14 = W*in
   wire signed [9:0] m63_14;
   assign m63_14 =10'b0;

   // m63_15 = W*in
   wire signed [9:0] m63_15;
   assign m63_15 =10'b0;

   // m63_16 = W*in
   wire signed [9:0] m63_16;
   assign m63_16 =10'b0;

   // m63_17 = W*in
   wire signed [9:0] m63_17;
   assign m63_17 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_18 = W*in
   wire signed [9:0] m63_18;
   assign m63_18 =10'b0;

   // m63_19 = W*in
   wire signed [9:0] m63_19;
   assign m63_19 =10'b0;

   // m63_20 = W*in
   wire signed [9:0] m63_20;
   assign m63_20 ={ {2{in63[5]}} , in63 , {2{1'b0}} };

   // m63_21 = W*in
   wire signed [9:0] m63_21;
   assign m63_21 =10'b0;

   // m63_22 = W*in
   wire signed [9:0] m63_22;
   assign m63_22 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_23 = W*in
   wire signed [9:0] m63_23;
   assign m63_23 =10'b0;

   // m63_24 = W*in
   wire signed [9:0] m63_24;
   assign m63_24 =10'b0;

   // m63_25 = W*in
   wire signed [9:0] m63_25;
   assign m63_25 =10'b0;

   // m63_26 = W*in
   wire signed [9:0] m63_26;
   assign m63_26 =10'b0;

   // m63_27 = W*in
   wire signed [9:0] m63_27;
   assign m63_27 =10'b0;

   // m63_28 = W*in
   wire signed [9:0] m63_28;
   assign m63_28 =10'b0;

   // m63_29 = W*in
   wire signed [9:0] m63_29;
   assign m63_29 ={ {2{in63[5]}} , in63 , {2{1'b0}} };

   // m63_30 = W*in
   wire signed [9:0] m63_30;
   assign m63_30 =10'b0;

   // m63_31 = W*in
   wire signed [9:0] m63_31;
   assign m63_31 =10'b0;

   // m63_32 = W*in
   wire signed [9:0] m63_32;
   assign m63_32 =10'b0;

   // m63_33 = W*in
   wire signed [9:0] m63_33;
   assign m63_33 =10'b0;

   // m63_34 = W*in
   wire signed [9:0] m63_34;
   assign m63_34 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_35 = W*in
   wire signed [9:0] m63_35;
   assign m63_35 =10'b0;

   // m63_36 = W*in
   wire signed [9:0] m63_36;
   assign m63_36 =10'b0;

   // m63_37 = W*in
   wire signed [9:0] m63_37;
   assign m63_37 ={ {3{neg63[5]}} , neg63 , {1{1'b0}} };

   // m63_38 = W*in
   wire signed [9:0] m63_38;
   assign m63_38 =10'b0;

   // m63_39 = W*in
   wire signed [9:0] m63_39;
   assign m63_39 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_40 = W*in
   wire signed [9:0] m63_40;
   assign m63_40 ={ {3{neg63[5]}} , neg63 , {1{1'b0}} };

   // m63_41 = W*in
   wire signed [9:0] m63_41;
   assign m63_41 =10'b0;

   // m63_42 = W*in
   wire signed [9:0] m63_42;
   assign m63_42 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_43 = W*in
   wire signed [9:0] m63_43;
   assign m63_43 =10'b0;

   // m63_44 = W*in
   wire signed [9:0] m63_44;
   assign m63_44 ={ {3{neg63[5]}} , neg63 , {1{1'b0}} };

   // m63_45 = W*in
   wire signed [9:0] m63_45;
   assign m63_45 =10'b0;

   // m63_46 = W*in
   wire signed [9:0] m63_46;
   assign m63_46 =10'b0;

   // m63_47 = W*in
   wire signed [9:0] m63_47;
   assign m63_47 =10'b0;

   // m63_48 = W*in
   wire signed [9:0] m63_48;
   assign m63_48 =10'b0;

   // m63_49 = W*in
   wire signed [9:0] m63_49;
   assign m63_49 =10'b0;

   // m63_50 = W*in
   wire signed [9:0] m63_50;
   assign m63_50 =10'b0;

   // m63_51 = W*in
   wire signed [9:0] m63_51;
   assign m63_51 =10'b0;

   // m63_52 = W*in
   wire signed [9:0] m63_52;
   assign m63_52 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_53 = W*in
   wire signed [9:0] m63_53;
   assign m63_53 =10'b0;

   // m63_54 = W*in
   wire signed [9:0] m63_54;
   assign m63_54 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_55 = W*in
   wire signed [9:0] m63_55;
   assign m63_55 ={ {3{neg63[5]}} , neg63 , {1{1'b0}} };

   // m63_56 = W*in
   wire signed [9:0] m63_56;
   assign m63_56 =10'b0;

   // m63_57 = W*in
   wire signed [9:0] m63_57;
   assign m63_57 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_58 = W*in
   wire signed [9:0] m63_58;
   assign m63_58 =10'b0;

   // m63_59 = W*in
   wire signed [9:0] m63_59;
   assign m63_59 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_60 = W*in
   wire signed [9:0] m63_60;
   assign m63_60 =10'b0;

   // m63_61 = W*in
   wire signed [9:0] m63_61;
   assign m63_61 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_62 = W*in
   wire signed [9:0] m63_62;
   assign m63_62 =10'b0;

   // m63_63 = W*in
   wire signed [9:0] m63_63;
   assign m63_63 =10'b0;

   // m63_64 = W*in
   wire signed [9:0] m63_64;
   assign m63_64 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_65 = W*in
   wire signed [9:0] m63_65;
   assign m63_65 =10'b0;

   // m63_66 = W*in
   wire signed [9:0] m63_66;
   assign m63_66 =10'b0;

   // m63_67 = W*in
   wire signed [9:0] m63_67;
   assign m63_67 =10'b0;

   // m63_68 = W*in
   wire signed [9:0] m63_68;
   assign m63_68 =10'b0;

   // m63_69 = W*in
   wire signed [9:0] m63_69;
   assign m63_69 =10'b0;

   // m63_70 = W*in
   wire signed [9:0] m63_70;
   assign m63_70 ={ {3{neg63[5]}} , neg63 , {1{1'b0}} };

   // m63_71 = W*in
   wire signed [9:0] m63_71;
   assign m63_71 =10'b0;

   // m63_72 = W*in
   wire signed [9:0] m63_72;
   assign m63_72 =10'b0;

   // m63_73 = W*in
   wire signed [9:0] m63_73;
   assign m63_73 =10'b0;

   // m63_74 = W*in
   wire signed [9:0] m63_74;
   assign m63_74 =10'b0;

   // m63_75 = W*in
   wire signed [9:0] m63_75;
   assign m63_75 =10'b0;

   // m63_76 = W*in
   wire signed [9:0] m63_76;
   assign m63_76 ={ {2{in63[5]}} , in63 , {2{1'b0}} };

   // m63_77 = W*in
   wire signed [9:0] m63_77;
   assign m63_77 ={ {3{in63[5]}} , in63 , {1{1'b0}} };

   // m63_78 = W*in
   wire signed [9:0] m63_78;
   assign m63_78 =10'b0;

   // m63_79 = W*in
   wire signed [9:0] m63_79;
   assign m63_79 =10'b0;

   // m63_80 = W*in
   wire signed [9:0] m63_80;
   assign m63_80 =10'b0;

   // m63_81 = W*in
   wire signed [9:0] m63_81;
   assign m63_81 =10'b0;

   // m64_1 = W*in
   wire signed [9:0] m64_1;
   assign m64_1 ={ {2{in64[5]}} , in64 , {2{1'b0}} };

   // m64_2 = W*in
   wire signed [9:0] m64_2;
   assign m64_2 =10'b0;

   // m64_3 = W*in
   wire signed [9:0] m64_3;
   assign m64_3 =10'b0;

   // m64_4 = W*in
   wire signed [9:0] m64_4;
   assign m64_4 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_5 = W*in
   wire signed [9:0] m64_5;
   assign m64_5 =10'b0;

   // m64_6 = W*in
   wire signed [9:0] m64_6;
   assign m64_6 =10'b0;

   // m64_7 = W*in
   wire signed [9:0] m64_7;
   assign m64_7 =10'b0;

   // m64_8 = W*in
   wire signed [9:0] m64_8;
   assign m64_8 =10'b0;

   // m64_9 = W*in
   wire signed [9:0] m64_9;
   assign m64_9 =10'b0;

   // m64_10 = W*in
   wire signed [9:0] m64_10;
   assign m64_10 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_11 = W*in
   wire signed [9:0] m64_11;
   assign m64_11 =10'b0;

   // m64_12 = W*in
   wire signed [9:0] m64_12;
   assign m64_12 =10'b0;

   // m64_13 = W*in
   wire signed [9:0] m64_13;
   assign m64_13 =10'b0;

   // m64_14 = W*in
   wire signed [9:0] m64_14;
   assign m64_14 =10'b0;

   // m64_15 = W*in
   wire signed [9:0] m64_15;
   assign m64_15 =10'b0;

   // m64_16 = W*in
   wire signed [9:0] m64_16;
   assign m64_16 =10'b0;

   // m64_17 = W*in
   wire signed [9:0] m64_17;
   assign m64_17 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_18 = W*in
   wire signed [9:0] m64_18;
   assign m64_18 =10'b0;

   // m64_19 = W*in
   wire signed [9:0] m64_19;
   assign m64_19 =10'b0;

   // m64_20 = W*in
   wire signed [9:0] m64_20;
   assign m64_20 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_21 = W*in
   wire signed [9:0] m64_21;
   assign m64_21 =10'b0;

   // m64_22 = W*in
   wire signed [9:0] m64_22;
   assign m64_22 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_23 = W*in
   wire signed [9:0] m64_23;
   assign m64_23 =10'b0;

   // m64_24 = W*in
   wire signed [9:0] m64_24;
   assign m64_24 =10'b0;

   // m64_25 = W*in
   wire signed [9:0] m64_25;
   assign m64_25 =10'b0;

   // m64_26 = W*in
   wire signed [9:0] m64_26;
   assign m64_26 =10'b0;

   // m64_27 = W*in
   wire signed [9:0] m64_27;
   assign m64_27 ={ {2{in64[5]}} , in64 , {2{1'b0}} };

   // m64_28 = W*in
   wire signed [9:0] m64_28;
   assign m64_28 =10'b0;

   // m64_29 = W*in
   wire signed [9:0] m64_29;
   assign m64_29 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_30 = W*in
   wire signed [9:0] m64_30;
   assign m64_30 =10'b0;

   // m64_31 = W*in
   wire signed [9:0] m64_31;
   assign m64_31 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_32 = W*in
   wire signed [9:0] m64_32;
   assign m64_32 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_33 = W*in
   wire signed [9:0] m64_33;
   assign m64_33 =10'b0;

   // m64_34 = W*in
   wire signed [9:0] m64_34;
   assign m64_34 =10'b0;

   // m64_35 = W*in
   wire signed [9:0] m64_35;
   assign m64_35 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_36 = W*in
   wire signed [9:0] m64_36;
   assign m64_36 =10'b0;

   // m64_37 = W*in
   wire signed [9:0] m64_37;
   assign m64_37 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_38 = W*in
   wire signed [9:0] m64_38;
   assign m64_38 =10'b0;

   // m64_39 = W*in
   wire signed [9:0] m64_39;
   assign m64_39 =10'b0;

   // m64_40 = W*in
   wire signed [9:0] m64_40;
   assign m64_40 =10'b0;

   // m64_41 = W*in
   wire signed [9:0] m64_41;
   assign m64_41 =10'b0;

   // m64_42 = W*in
   wire signed [9:0] m64_42;
   assign m64_42 =10'b0;

   // m64_43 = W*in
   wire signed [9:0] m64_43;
   assign m64_43 =10'b0;

   // m64_44 = W*in
   wire signed [9:0] m64_44;
   assign m64_44 =10'b0;

   // m64_45 = W*in
   wire signed [9:0] m64_45;
   assign m64_45 =10'b0;

   // m64_46 = W*in
   wire signed [9:0] m64_46;
   assign m64_46 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_47 = W*in
   wire signed [9:0] m64_47;
   assign m64_47 =10'b0;

   // m64_48 = W*in
   wire signed [9:0] m64_48;
   assign m64_48 =10'b0;

   // m64_49 = W*in
   wire signed [9:0] m64_49;
   assign m64_49 =10'b0;

   // m64_50 = W*in
   wire signed [9:0] m64_50;
   assign m64_50 =10'b0;

   // m64_51 = W*in
   wire signed [9:0] m64_51;
   assign m64_51 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_52 = W*in
   wire signed [9:0] m64_52;
   assign m64_52 =10'b0;

   // m64_53 = W*in
   wire signed [9:0] m64_53;
   assign m64_53 =10'b0;

   // m64_54 = W*in
   wire signed [9:0] m64_54;
   assign m64_54 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_55 = W*in
   wire signed [9:0] m64_55;
   assign m64_55 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_56 = W*in
   wire signed [9:0] m64_56;
   assign m64_56 =10'b0;

   // m64_57 = W*in
   wire signed [9:0] m64_57;
   assign m64_57 =10'b0;

   // m64_58 = W*in
   wire signed [9:0] m64_58;
   assign m64_58 =10'b0;

   // m64_59 = W*in
   wire signed [9:0] m64_59;
   assign m64_59 =10'b0;

   // m64_60 = W*in
   wire signed [9:0] m64_60;
   assign m64_60 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_61 = W*in
   wire signed [9:0] m64_61;
   assign m64_61 ={ {2{in64[5]}} , in64 , {2{1'b0}} };

   // m64_62 = W*in
   wire signed [9:0] m64_62;
   assign m64_62 =10'b0;

   // m64_63 = W*in
   wire signed [9:0] m64_63;
   assign m64_63 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_64 = W*in
   wire signed [9:0] m64_64;
   assign m64_64 =10'b0;

   // m64_65 = W*in
   wire signed [9:0] m64_65;
   assign m64_65 =10'b0;

   // m64_66 = W*in
   wire signed [9:0] m64_66;
   assign m64_66 =10'b0;

   // m64_67 = W*in
   wire signed [9:0] m64_67;
   assign m64_67 =10'b0;

   // m64_68 = W*in
   wire signed [9:0] m64_68;
   assign m64_68 =10'b0;

   // m64_69 = W*in
   wire signed [9:0] m64_69;
   assign m64_69 ={ {3{neg64[5]}} , neg64 , {1{1'b0}} };

   // m64_70 = W*in
   wire signed [9:0] m64_70;
   assign m64_70 =10'b0;

   // m64_71 = W*in
   wire signed [9:0] m64_71;
   assign m64_71 =10'b0;

   // m64_72 = W*in
   wire signed [9:0] m64_72;
   assign m64_72 =10'b0;

   // m64_73 = W*in
   wire signed [9:0] m64_73;
   assign m64_73 =10'b0;

   // m64_74 = W*in
   wire signed [9:0] m64_74;
   assign m64_74 =10'b0;

   // m64_75 = W*in
   wire signed [9:0] m64_75;
   assign m64_75 =10'b0;

   // m64_76 = W*in
   wire signed [9:0] m64_76;
   assign m64_76 =10'b0;

   // m64_77 = W*in
   wire signed [9:0] m64_77;
   assign m64_77 =10'b0;

   // m64_78 = W*in
   wire signed [9:0] m64_78;
   assign m64_78 ={ {3{in64[5]}} , in64 , {1{1'b0}} };

   // m64_79 = W*in
   wire signed [9:0] m64_79;
   assign m64_79 =10'b0;

   // m64_80 = W*in
   wire signed [9:0] m64_80;
   assign m64_80 =10'b0;

   // m64_81 = W*in
   wire signed [9:0] m64_81;
   assign m64_81 =10'b0;

   // m65_1 = W*in
   wire signed [9:0] m65_1;
   assign m65_1 ={ {2{in65[5]}} , in65 , {2{1'b0}} };

   // m65_2 = W*in
   wire signed [9:0] m65_2;
   assign m65_2 =10'b0;

   // m65_3 = W*in
   wire signed [9:0] m65_3;
   assign m65_3 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_4 = W*in
   wire signed [9:0] m65_4;
   assign m65_4 =10'b0;

   // m65_5 = W*in
   wire signed [9:0] m65_5;
   assign m65_5 =10'b0;

   // m65_6 = W*in
   wire signed [9:0] m65_6;
   assign m65_6 =10'b0;

   // m65_7 = W*in
   wire signed [9:0] m65_7;
   assign m65_7 =10'b0;

   // m65_8 = W*in
   wire signed [9:0] m65_8;
   assign m65_8 =10'b0;

   // m65_9 = W*in
   wire signed [9:0] m65_9;
   assign m65_9 =10'b0;

   // m65_10 = W*in
   wire signed [9:0] m65_10;
   assign m65_10 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_11 = W*in
   wire signed [9:0] m65_11;
   assign m65_11 =10'b0;

   // m65_12 = W*in
   wire signed [9:0] m65_12;
   assign m65_12 =10'b0;

   // m65_13 = W*in
   wire signed [9:0] m65_13;
   assign m65_13 =10'b0;

   // m65_14 = W*in
   wire signed [9:0] m65_14;
   assign m65_14 =10'b0;

   // m65_15 = W*in
   wire signed [9:0] m65_15;
   assign m65_15 =10'b0;

   // m65_16 = W*in
   wire signed [9:0] m65_16;
   assign m65_16 =10'b0;

   // m65_17 = W*in
   wire signed [9:0] m65_17;
   assign m65_17 =10'b0;

   // m65_18 = W*in
   wire signed [9:0] m65_18;
   assign m65_18 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_19 = W*in
   wire signed [9:0] m65_19;
   assign m65_19 =10'b0;

   // m65_20 = W*in
   wire signed [9:0] m65_20;
   assign m65_20 =10'b0;

   // m65_21 = W*in
   wire signed [9:0] m65_21;
   assign m65_21 =10'b0;

   // m65_22 = W*in
   wire signed [9:0] m65_22;
   assign m65_22 ={ {2{in65[5]}} , in65 , {2{1'b0}} };

   // m65_23 = W*in
   wire signed [9:0] m65_23;
   assign m65_23 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_24 = W*in
   wire signed [9:0] m65_24;
   assign m65_24 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_25 = W*in
   wire signed [9:0] m65_25;
   assign m65_25 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_26 = W*in
   wire signed [9:0] m65_26;
   assign m65_26 =10'b0;

   // m65_27 = W*in
   wire signed [9:0] m65_27;
   assign m65_27 =10'b0;

   // m65_28 = W*in
   wire signed [9:0] m65_28;
   assign m65_28 =10'b0;

   // m65_29 = W*in
   wire signed [9:0] m65_29;
   assign m65_29 =10'b0;

   // m65_30 = W*in
   wire signed [9:0] m65_30;
   assign m65_30 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_31 = W*in
   wire signed [9:0] m65_31;
   assign m65_31 ={ {2{in65[5]}} , in65 , {2{1'b0}} };

   // m65_32 = W*in
   wire signed [9:0] m65_32;
   assign m65_32 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_33 = W*in
   wire signed [9:0] m65_33;
   assign m65_33 =10'b0;

   // m65_34 = W*in
   wire signed [9:0] m65_34;
   assign m65_34 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_35 = W*in
   wire signed [9:0] m65_35;
   assign m65_35 =10'b0;

   // m65_36 = W*in
   wire signed [9:0] m65_36;
   assign m65_36 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_37 = W*in
   wire signed [9:0] m65_37;
   assign m65_37 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_38 = W*in
   wire signed [9:0] m65_38;
   assign m65_38 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_39 = W*in
   wire signed [9:0] m65_39;
   assign m65_39 =10'b0;

   // m65_40 = W*in
   wire signed [9:0] m65_40;
   assign m65_40 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_41 = W*in
   wire signed [9:0] m65_41;
   assign m65_41 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_42 = W*in
   wire signed [9:0] m65_42;
   assign m65_42 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_43 = W*in
   wire signed [9:0] m65_43;
   assign m65_43 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_44 = W*in
   wire signed [9:0] m65_44;
   assign m65_44 =10'b0;

   // m65_45 = W*in
   wire signed [9:0] m65_45;
   assign m65_45 =10'b0;

   // m65_46 = W*in
   wire signed [9:0] m65_46;
   assign m65_46 =10'b0;

   // m65_47 = W*in
   wire signed [9:0] m65_47;
   assign m65_47 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_48 = W*in
   wire signed [9:0] m65_48;
   assign m65_48 =10'b0;

   // m65_49 = W*in
   wire signed [9:0] m65_49;
   assign m65_49 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_50 = W*in
   wire signed [9:0] m65_50;
   assign m65_50 ={ {2{in65[5]}} , in65 , {2{1'b0}} };

   // m65_51 = W*in
   wire signed [9:0] m65_51;
   assign m65_51 =10'b0;

   // m65_52 = W*in
   wire signed [9:0] m65_52;
   assign m65_52 =10'b0;

   // m65_53 = W*in
   wire signed [9:0] m65_53;
   assign m65_53 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_54 = W*in
   wire signed [9:0] m65_54;
   assign m65_54 =10'b0;

   // m65_55 = W*in
   wire signed [9:0] m65_55;
   assign m65_55 ={ {2{neg65[5]}} , neg65 , {2{1'b0}} };

   // m65_56 = W*in
   wire signed [9:0] m65_56;
   assign m65_56 =10'b0;

   // m65_57 = W*in
   wire signed [9:0] m65_57;
   assign m65_57 =10'b0;

   // m65_58 = W*in
   wire signed [9:0] m65_58;
   assign m65_58 =10'b0;

   // m65_59 = W*in
   wire signed [9:0] m65_59;
   assign m65_59 =10'b0;

   // m65_60 = W*in
   wire signed [9:0] m65_60;
   assign m65_60 =10'b0;

   // m65_61 = W*in
   wire signed [9:0] m65_61;
   assign m65_61 ={ {2{in65[5]}} , in65 , {2{1'b0}} };

   // m65_62 = W*in
   wire signed [9:0] m65_62;
   assign m65_62 =10'b0;

   // m65_63 = W*in
   wire signed [9:0] m65_63;
   assign m65_63 =10'b0;

   // m65_64 = W*in
   wire signed [9:0] m65_64;
   assign m65_64 =10'b0;

   // m65_65 = W*in
   wire signed [9:0] m65_65;
   assign m65_65 =10'b0;

   // m65_66 = W*in
   wire signed [9:0] m65_66;
   assign m65_66 =10'b0;

   // m65_67 = W*in
   wire signed [9:0] m65_67;
   assign m65_67 =10'b0;

   // m65_68 = W*in
   wire signed [9:0] m65_68;
   assign m65_68 =10'b0;

   // m65_69 = W*in
   wire signed [9:0] m65_69;
   assign m65_69 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_70 = W*in
   wire signed [9:0] m65_70;
   assign m65_70 =10'b0;

   // m65_71 = W*in
   wire signed [9:0] m65_71;
   assign m65_71 =10'b0;

   // m65_72 = W*in
   wire signed [9:0] m65_72;
   assign m65_72 =10'b0;

   // m65_73 = W*in
   wire signed [9:0] m65_73;
   assign m65_73 =10'b0;

   // m65_74 = W*in
   wire signed [9:0] m65_74;
   assign m65_74 =10'b0;

   // m65_75 = W*in
   wire signed [9:0] m65_75;
   assign m65_75 =10'b0;

   // m65_76 = W*in
   wire signed [9:0] m65_76;
   assign m65_76 =10'b0;

   // m65_77 = W*in
   wire signed [9:0] m65_77;
   assign m65_77 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_78 = W*in
   wire signed [9:0] m65_78;
   assign m65_78 =10'b0;

   // m65_79 = W*in
   wire signed [9:0] m65_79;
   assign m65_79 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_80 = W*in
   wire signed [9:0] m65_80;
   assign m65_80 =10'b0;

   // m65_81 = W*in
   wire signed [9:0] m65_81;
   assign m65_81 =10'b0;

   // m66_1 = W*in
   wire signed [9:0] m66_1;
   assign m66_1 =10'b0;

   // m66_2 = W*in
   wire signed [9:0] m66_2;
   assign m66_2 =10'b0;

   // m66_3 = W*in
   wire signed [9:0] m66_3;
   assign m66_3 =10'b0;

   // m66_4 = W*in
   wire signed [9:0] m66_4;
   assign m66_4 =10'b0;

   // m66_5 = W*in
   wire signed [9:0] m66_5;
   assign m66_5 =10'b0;

   // m66_6 = W*in
   wire signed [9:0] m66_6;
   assign m66_6 =10'b0;

   // m66_7 = W*in
   wire signed [9:0] m66_7;
   assign m66_7 =10'b0;

   // m66_8 = W*in
   wire signed [9:0] m66_8;
   assign m66_8 =10'b0;

   // m66_9 = W*in
   wire signed [9:0] m66_9;
   assign m66_9 =10'b0;

   // m66_10 = W*in
   wire signed [9:0] m66_10;
   assign m66_10 =10'b0;

   // m66_11 = W*in
   wire signed [9:0] m66_11;
   assign m66_11 ={ {2{in66[5]}} , in66 , {2{1'b0}} };

   // m66_12 = W*in
   wire signed [9:0] m66_12;
   assign m66_12 =10'b0;

   // m66_13 = W*in
   wire signed [9:0] m66_13;
   assign m66_13 =10'b0;

   // m66_14 = W*in
   wire signed [9:0] m66_14;
   assign m66_14 =10'b0;

   // m66_15 = W*in
   wire signed [9:0] m66_15;
   assign m66_15 =10'b0;

   // m66_16 = W*in
   wire signed [9:0] m66_16;
   assign m66_16 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_17 = W*in
   wire signed [9:0] m66_17;
   assign m66_17 ={ {2{neg66[5]}} , neg66 , {2{1'b0}} };

   // m66_18 = W*in
   wire signed [9:0] m66_18;
   assign m66_18 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_19 = W*in
   wire signed [9:0] m66_19;
   assign m66_19 =10'b0;

   // m66_20 = W*in
   wire signed [9:0] m66_20;
   assign m66_20 =10'b0;

   // m66_21 = W*in
   wire signed [9:0] m66_21;
   assign m66_21 =10'b0;

   // m66_22 = W*in
   wire signed [9:0] m66_22;
   assign m66_22 =10'b0;

   // m66_23 = W*in
   wire signed [9:0] m66_23;
   assign m66_23 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_24 = W*in
   wire signed [9:0] m66_24;
   assign m66_24 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_25 = W*in
   wire signed [9:0] m66_25;
   assign m66_25 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_26 = W*in
   wire signed [9:0] m66_26;
   assign m66_26 =10'b0;

   // m66_27 = W*in
   wire signed [9:0] m66_27;
   assign m66_27 =10'b0;

   // m66_28 = W*in
   wire signed [9:0] m66_28;
   assign m66_28 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_29 = W*in
   wire signed [9:0] m66_29;
   assign m66_29 =10'b0;

   // m66_30 = W*in
   wire signed [9:0] m66_30;
   assign m66_30 =10'b0;

   // m66_31 = W*in
   wire signed [9:0] m66_31;
   assign m66_31 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_32 = W*in
   wire signed [9:0] m66_32;
   assign m66_32 =10'b0;

   // m66_33 = W*in
   wire signed [9:0] m66_33;
   assign m66_33 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_34 = W*in
   wire signed [9:0] m66_34;
   assign m66_34 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_35 = W*in
   wire signed [9:0] m66_35;
   assign m66_35 =10'b0;

   // m66_36 = W*in
   wire signed [9:0] m66_36;
   assign m66_36 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_37 = W*in
   wire signed [9:0] m66_37;
   assign m66_37 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_38 = W*in
   wire signed [9:0] m66_38;
   assign m66_38 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_39 = W*in
   wire signed [9:0] m66_39;
   assign m66_39 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_40 = W*in
   wire signed [9:0] m66_40;
   assign m66_40 =10'b0;

   // m66_41 = W*in
   wire signed [9:0] m66_41;
   assign m66_41 ={ {2{in66[5]}} , in66 , {2{1'b0}} };

   // m66_42 = W*in
   wire signed [9:0] m66_42;
   assign m66_42 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_43 = W*in
   wire signed [9:0] m66_43;
   assign m66_43 =10'b0;

   // m66_44 = W*in
   wire signed [9:0] m66_44;
   assign m66_44 =10'b0;

   // m66_45 = W*in
   wire signed [9:0] m66_45;
   assign m66_45 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_46 = W*in
   wire signed [9:0] m66_46;
   assign m66_46 =10'b0;

   // m66_47 = W*in
   wire signed [9:0] m66_47;
   assign m66_47 =10'b0;

   // m66_48 = W*in
   wire signed [9:0] m66_48;
   assign m66_48 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_49 = W*in
   wire signed [9:0] m66_49;
   assign m66_49 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_50 = W*in
   wire signed [9:0] m66_50;
   assign m66_50 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_51 = W*in
   wire signed [9:0] m66_51;
   assign m66_51 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_52 = W*in
   wire signed [9:0] m66_52;
   assign m66_52 =10'b0;

   // m66_53 = W*in
   wire signed [9:0] m66_53;
   assign m66_53 =10'b0;

   // m66_54 = W*in
   wire signed [9:0] m66_54;
   assign m66_54 =10'b0;

   // m66_55 = W*in
   wire signed [9:0] m66_55;
   assign m66_55 =10'b0;

   // m66_56 = W*in
   wire signed [9:0] m66_56;
   assign m66_56 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_57 = W*in
   wire signed [9:0] m66_57;
   assign m66_57 =10'b0;

   // m66_58 = W*in
   wire signed [9:0] m66_58;
   assign m66_58 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_59 = W*in
   wire signed [9:0] m66_59;
   assign m66_59 ={ {2{in66[5]}} , in66 , {2{1'b0}} };

   // m66_60 = W*in
   wire signed [9:0] m66_60;
   assign m66_60 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_61 = W*in
   wire signed [9:0] m66_61;
   assign m66_61 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_62 = W*in
   wire signed [9:0] m66_62;
   assign m66_62 =10'b0;

   // m66_63 = W*in
   wire signed [9:0] m66_63;
   assign m66_63 ={ {2{in66[5]}} , in66 , {2{1'b0}} };

   // m66_64 = W*in
   wire signed [9:0] m66_64;
   assign m66_64 =10'b0;

   // m66_65 = W*in
   wire signed [9:0] m66_65;
   assign m66_65 =10'b0;

   // m66_66 = W*in
   wire signed [9:0] m66_66;
   assign m66_66 =10'b0;

   // m66_67 = W*in
   wire signed [9:0] m66_67;
   assign m66_67 =10'b0;

   // m66_68 = W*in
   wire signed [9:0] m66_68;
   assign m66_68 =10'b0;

   // m66_69 = W*in
   wire signed [9:0] m66_69;
   assign m66_69 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_70 = W*in
   wire signed [9:0] m66_70;
   assign m66_70 =10'b0;

   // m66_71 = W*in
   wire signed [9:0] m66_71;
   assign m66_71 =10'b0;

   // m66_72 = W*in
   wire signed [9:0] m66_72;
   assign m66_72 =10'b0;

   // m66_73 = W*in
   wire signed [9:0] m66_73;
   assign m66_73 =10'b0;

   // m66_74 = W*in
   wire signed [9:0] m66_74;
   assign m66_74 =10'b0;

   // m66_75 = W*in
   wire signed [9:0] m66_75;
   assign m66_75 =10'b0;

   // m66_76 = W*in
   wire signed [9:0] m66_76;
   assign m66_76 =10'b0;

   // m66_77 = W*in
   wire signed [9:0] m66_77;
   assign m66_77 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_78 = W*in
   wire signed [9:0] m66_78;
   assign m66_78 =10'b0;

   // m66_79 = W*in
   wire signed [9:0] m66_79;
   assign m66_79 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_80 = W*in
   wire signed [9:0] m66_80;
   assign m66_80 =10'b0;

   // m66_81 = W*in
   wire signed [9:0] m66_81;
   assign m66_81 =10'b0;

   // m67_1 = W*in
   wire signed [9:0] m67_1;
   assign m67_1 =10'b0;

   // m67_2 = W*in
   wire signed [9:0] m67_2;
   assign m67_2 =10'b0;

   // m67_3 = W*in
   wire signed [9:0] m67_3;
   assign m67_3 =10'b0;

   // m67_4 = W*in
   wire signed [9:0] m67_4;
   assign m67_4 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_5 = W*in
   wire signed [9:0] m67_5;
   assign m67_5 =10'b0;

   // m67_6 = W*in
   wire signed [9:0] m67_6;
   assign m67_6 =10'b0;

   // m67_7 = W*in
   wire signed [9:0] m67_7;
   assign m67_7 ={ {2{in67[5]}} , in67 , {2{1'b0}} };

   // m67_8 = W*in
   wire signed [9:0] m67_8;
   assign m67_8 =10'b0;

   // m67_9 = W*in
   wire signed [9:0] m67_9;
   assign m67_9 =10'b0;

   // m67_10 = W*in
   wire signed [9:0] m67_10;
   assign m67_10 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_11 = W*in
   wire signed [9:0] m67_11;
   assign m67_11 =10'b0;

   // m67_12 = W*in
   wire signed [9:0] m67_12;
   assign m67_12 =10'b0;

   // m67_13 = W*in
   wire signed [9:0] m67_13;
   assign m67_13 =10'b0;

   // m67_14 = W*in
   wire signed [9:0] m67_14;
   assign m67_14 =10'b0;

   // m67_15 = W*in
   wire signed [9:0] m67_15;
   assign m67_15 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_16 = W*in
   wire signed [9:0] m67_16;
   assign m67_16 =10'b0;

   // m67_17 = W*in
   wire signed [9:0] m67_17;
   assign m67_17 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_18 = W*in
   wire signed [9:0] m67_18;
   assign m67_18 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_19 = W*in
   wire signed [9:0] m67_19;
   assign m67_19 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_20 = W*in
   wire signed [9:0] m67_20;
   assign m67_20 ={ {2{in67[5]}} , in67 , {2{1'b0}} };

   // m67_21 = W*in
   wire signed [9:0] m67_21;
   assign m67_21 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_22 = W*in
   wire signed [9:0] m67_22;
   assign m67_22 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_23 = W*in
   wire signed [9:0] m67_23;
   assign m67_23 =10'b0;

   // m67_24 = W*in
   wire signed [9:0] m67_24;
   assign m67_24 =10'b0;

   // m67_25 = W*in
   wire signed [9:0] m67_25;
   assign m67_25 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_26 = W*in
   wire signed [9:0] m67_26;
   assign m67_26 =10'b0;

   // m67_27 = W*in
   wire signed [9:0] m67_27;
   assign m67_27 =10'b0;

   // m67_28 = W*in
   wire signed [9:0] m67_28;
   assign m67_28 =10'b0;

   // m67_29 = W*in
   wire signed [9:0] m67_29;
   assign m67_29 ={ {2{in67[5]}} , in67 , {2{1'b0}} };

   // m67_30 = W*in
   wire signed [9:0] m67_30;
   assign m67_30 =10'b0;

   // m67_31 = W*in
   wire signed [9:0] m67_31;
   assign m67_31 =10'b0;

   // m67_32 = W*in
   wire signed [9:0] m67_32;
   assign m67_32 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_33 = W*in
   wire signed [9:0] m67_33;
   assign m67_33 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_34 = W*in
   wire signed [9:0] m67_34;
   assign m67_34 =10'b0;

   // m67_35 = W*in
   wire signed [9:0] m67_35;
   assign m67_35 =10'b0;

   // m67_36 = W*in
   wire signed [9:0] m67_36;
   assign m67_36 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_37 = W*in
   wire signed [9:0] m67_37;
   assign m67_37 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_38 = W*in
   wire signed [9:0] m67_38;
   assign m67_38 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_39 = W*in
   wire signed [9:0] m67_39;
   assign m67_39 =10'b0;

   // m67_40 = W*in
   wire signed [9:0] m67_40;
   assign m67_40 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_41 = W*in
   wire signed [9:0] m67_41;
   assign m67_41 =10'b0;

   // m67_42 = W*in
   wire signed [9:0] m67_42;
   assign m67_42 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_43 = W*in
   wire signed [9:0] m67_43;
   assign m67_43 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_44 = W*in
   wire signed [9:0] m67_44;
   assign m67_44 =10'b0;

   // m67_45 = W*in
   wire signed [9:0] m67_45;
   assign m67_45 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_46 = W*in
   wire signed [9:0] m67_46;
   assign m67_46 =10'b0;

   // m67_47 = W*in
   wire signed [9:0] m67_47;
   assign m67_47 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_48 = W*in
   wire signed [9:0] m67_48;
   assign m67_48 ={ {2{in67[5]}} , in67 , {2{1'b0}} };

   // m67_49 = W*in
   wire signed [9:0] m67_49;
   assign m67_49 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_50 = W*in
   wire signed [9:0] m67_50;
   assign m67_50 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_51 = W*in
   wire signed [9:0] m67_51;
   assign m67_51 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_52 = W*in
   wire signed [9:0] m67_52;
   assign m67_52 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_53 = W*in
   wire signed [9:0] m67_53;
   assign m67_53 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_54 = W*in
   wire signed [9:0] m67_54;
   assign m67_54 =10'b0;

   // m67_55 = W*in
   wire signed [9:0] m67_55;
   assign m67_55 =10'b0;

   // m67_56 = W*in
   wire signed [9:0] m67_56;
   assign m67_56 =10'b0;

   // m67_57 = W*in
   wire signed [9:0] m67_57;
   assign m67_57 =10'b0;

   // m67_58 = W*in
   wire signed [9:0] m67_58;
   assign m67_58 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_59 = W*in
   wire signed [9:0] m67_59;
   assign m67_59 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_60 = W*in
   wire signed [9:0] m67_60;
   assign m67_60 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_61 = W*in
   wire signed [9:0] m67_61;
   assign m67_61 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_62 = W*in
   wire signed [9:0] m67_62;
   assign m67_62 ={ {3{neg67[5]}} , neg67 , {1{1'b0}} };

   // m67_63 = W*in
   wire signed [9:0] m67_63;
   assign m67_63 =10'b0;

   // m67_64 = W*in
   wire signed [9:0] m67_64;
   assign m67_64 =10'b0;

   // m67_65 = W*in
   wire signed [9:0] m67_65;
   assign m67_65 =10'b0;

   // m67_66 = W*in
   wire signed [9:0] m67_66;
   assign m67_66 =10'b0;

   // m67_67 = W*in
   wire signed [9:0] m67_67;
   assign m67_67 =10'b0;

   // m67_68 = W*in
   wire signed [9:0] m67_68;
   assign m67_68 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_69 = W*in
   wire signed [9:0] m67_69;
   assign m67_69 ={ {2{in67[5]}} , in67 , {2{1'b0}} };

   // m67_70 = W*in
   wire signed [9:0] m67_70;
   assign m67_70 =10'b0;

   // m67_71 = W*in
   wire signed [9:0] m67_71;
   assign m67_71 =10'b0;

   // m67_72 = W*in
   wire signed [9:0] m67_72;
   assign m67_72 =10'b0;

   // m67_73 = W*in
   wire signed [9:0] m67_73;
   assign m67_73 =10'b0;

   // m67_74 = W*in
   wire signed [9:0] m67_74;
   assign m67_74 =10'b0;

   // m67_75 = W*in
   wire signed [9:0] m67_75;
   assign m67_75 =10'b0;

   // m67_76 = W*in
   wire signed [9:0] m67_76;
   assign m67_76 =10'b0;

   // m67_77 = W*in
   wire signed [9:0] m67_77;
   assign m67_77 ={ {3{in67[5]}} , in67 , {1{1'b0}} };

   // m67_78 = W*in
   wire signed [9:0] m67_78;
   assign m67_78 =10'b0;

   // m67_79 = W*in
   wire signed [9:0] m67_79;
   assign m67_79 =10'b0;

   // m67_80 = W*in
   wire signed [9:0] m67_80;
   assign m67_80 =10'b0;

   // m67_81 = W*in
   wire signed [9:0] m67_81;
   assign m67_81 =10'b0;

   // m68_1 = W*in
   wire signed [9:0] m68_1;
   assign m68_1 =10'b0;

   // m68_2 = W*in
   wire signed [9:0] m68_2;
   assign m68_2 ={ {2{in68[5]}} , in68 , {2{1'b0}} };

   // m68_3 = W*in
   wire signed [9:0] m68_3;
   assign m68_3 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_4 = W*in
   wire signed [9:0] m68_4;
   assign m68_4 =10'b0;

   // m68_5 = W*in
   wire signed [9:0] m68_5;
   assign m68_5 =10'b0;

   // m68_6 = W*in
   wire signed [9:0] m68_6;
   assign m68_6 =10'b0;

   // m68_7 = W*in
   wire signed [9:0] m68_7;
   assign m68_7 =10'b0;

   // m68_8 = W*in
   wire signed [9:0] m68_8;
   assign m68_8 ={ {2{in68[5]}} , in68 , {2{1'b0}} };

   // m68_9 = W*in
   wire signed [9:0] m68_9;
   assign m68_9 =10'b0;

   // m68_10 = W*in
   wire signed [9:0] m68_10;
   assign m68_10 =10'b0;

   // m68_11 = W*in
   wire signed [9:0] m68_11;
   assign m68_11 =10'b0;

   // m68_12 = W*in
   wire signed [9:0] m68_12;
   assign m68_12 =10'b0;

   // m68_13 = W*in
   wire signed [9:0] m68_13;
   assign m68_13 =10'b0;

   // m68_14 = W*in
   wire signed [9:0] m68_14;
   assign m68_14 =10'b0;

   // m68_15 = W*in
   wire signed [9:0] m68_15;
   assign m68_15 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_16 = W*in
   wire signed [9:0] m68_16;
   assign m68_16 =10'b0;

   // m68_17 = W*in
   wire signed [9:0] m68_17;
   assign m68_17 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_18 = W*in
   wire signed [9:0] m68_18;
   assign m68_18 =10'b0;

   // m68_19 = W*in
   wire signed [9:0] m68_19;
   assign m68_19 =10'b0;

   // m68_20 = W*in
   wire signed [9:0] m68_20;
   assign m68_20 =10'b0;

   // m68_21 = W*in
   wire signed [9:0] m68_21;
   assign m68_21 =10'b0;

   // m68_22 = W*in
   wire signed [9:0] m68_22;
   assign m68_22 =10'b0;

   // m68_23 = W*in
   wire signed [9:0] m68_23;
   assign m68_23 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_24 = W*in
   wire signed [9:0] m68_24;
   assign m68_24 =10'b0;

   // m68_25 = W*in
   wire signed [9:0] m68_25;
   assign m68_25 =10'b0;

   // m68_26 = W*in
   wire signed [9:0] m68_26;
   assign m68_26 =10'b0;

   // m68_27 = W*in
   wire signed [9:0] m68_27;
   assign m68_27 =10'b0;

   // m68_28 = W*in
   wire signed [9:0] m68_28;
   assign m68_28 =10'b0;

   // m68_29 = W*in
   wire signed [9:0] m68_29;
   assign m68_29 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_30 = W*in
   wire signed [9:0] m68_30;
   assign m68_30 =10'b0;

   // m68_31 = W*in
   wire signed [9:0] m68_31;
   assign m68_31 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_32 = W*in
   wire signed [9:0] m68_32;
   assign m68_32 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_33 = W*in
   wire signed [9:0] m68_33;
   assign m68_33 =10'b0;

   // m68_34 = W*in
   wire signed [9:0] m68_34;
   assign m68_34 =10'b0;

   // m68_35 = W*in
   wire signed [9:0] m68_35;
   assign m68_35 =10'b0;

   // m68_36 = W*in
   wire signed [9:0] m68_36;
   assign m68_36 =10'b0;

   // m68_37 = W*in
   wire signed [9:0] m68_37;
   assign m68_37 =10'b0;

   // m68_38 = W*in
   wire signed [9:0] m68_38;
   assign m68_38 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_39 = W*in
   wire signed [9:0] m68_39;
   assign m68_39 =10'b0;

   // m68_40 = W*in
   wire signed [9:0] m68_40;
   assign m68_40 =10'b0;

   // m68_41 = W*in
   wire signed [9:0] m68_41;
   assign m68_41 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_42 = W*in
   wire signed [9:0] m68_42;
   assign m68_42 =10'b0;

   // m68_43 = W*in
   wire signed [9:0] m68_43;
   assign m68_43 =10'b0;

   // m68_44 = W*in
   wire signed [9:0] m68_44;
   assign m68_44 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_45 = W*in
   wire signed [9:0] m68_45;
   assign m68_45 ={ {2{in68[5]}} , in68 , {2{1'b0}} };

   // m68_46 = W*in
   wire signed [9:0] m68_46;
   assign m68_46 =10'b0;

   // m68_47 = W*in
   wire signed [9:0] m68_47;
   assign m68_47 =10'b0;

   // m68_48 = W*in
   wire signed [9:0] m68_48;
   assign m68_48 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_49 = W*in
   wire signed [9:0] m68_49;
   assign m68_49 ={ {2{in68[5]}} , in68 , {2{1'b0}} };

   // m68_50 = W*in
   wire signed [9:0] m68_50;
   assign m68_50 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_51 = W*in
   wire signed [9:0] m68_51;
   assign m68_51 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_52 = W*in
   wire signed [9:0] m68_52;
   assign m68_52 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_53 = W*in
   wire signed [9:0] m68_53;
   assign m68_53 =10'b0;

   // m68_54 = W*in
   wire signed [9:0] m68_54;
   assign m68_54 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_55 = W*in
   wire signed [9:0] m68_55;
   assign m68_55 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_56 = W*in
   wire signed [9:0] m68_56;
   assign m68_56 =10'b0;

   // m68_57 = W*in
   wire signed [9:0] m68_57;
   assign m68_57 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_58 = W*in
   wire signed [9:0] m68_58;
   assign m68_58 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_59 = W*in
   wire signed [9:0] m68_59;
   assign m68_59 =10'b0;

   // m68_60 = W*in
   wire signed [9:0] m68_60;
   assign m68_60 =10'b0;

   // m68_61 = W*in
   wire signed [9:0] m68_61;
   assign m68_61 ={ {3{neg68[5]}} , neg68 , {1{1'b0}} };

   // m68_62 = W*in
   wire signed [9:0] m68_62;
   assign m68_62 =10'b0;

   // m68_63 = W*in
   wire signed [9:0] m68_63;
   assign m68_63 =10'b0;

   // m68_64 = W*in
   wire signed [9:0] m68_64;
   assign m68_64 =10'b0;

   // m68_65 = W*in
   wire signed [9:0] m68_65;
   assign m68_65 =10'b0;

   // m68_66 = W*in
   wire signed [9:0] m68_66;
   assign m68_66 =10'b0;

   // m68_67 = W*in
   wire signed [9:0] m68_67;
   assign m68_67 ={ {2{in68[5]}} , in68 , {2{1'b0}} };

   // m68_68 = W*in
   wire signed [9:0] m68_68;
   assign m68_68 =10'b0;

   // m68_69 = W*in
   wire signed [9:0] m68_69;
   assign m68_69 =10'b0;

   // m68_70 = W*in
   wire signed [9:0] m68_70;
   assign m68_70 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_71 = W*in
   wire signed [9:0] m68_71;
   assign m68_71 =10'b0;

   // m68_72 = W*in
   wire signed [9:0] m68_72;
   assign m68_72 =10'b0;

   // m68_73 = W*in
   wire signed [9:0] m68_73;
   assign m68_73 ={ {2{in68[5]}} , in68 , {2{1'b0}} };

   // m68_74 = W*in
   wire signed [9:0] m68_74;
   assign m68_74 =10'b0;

   // m68_75 = W*in
   wire signed [9:0] m68_75;
   assign m68_75 =10'b0;

   // m68_76 = W*in
   wire signed [9:0] m68_76;
   assign m68_76 =10'b0;

   // m68_77 = W*in
   wire signed [9:0] m68_77;
   assign m68_77 =10'b0;

   // m68_78 = W*in
   wire signed [9:0] m68_78;
   assign m68_78 =10'b0;

   // m68_79 = W*in
   wire signed [9:0] m68_79;
   assign m68_79 ={ {3{in68[5]}} , in68 , {1{1'b0}} };

   // m68_80 = W*in
   wire signed [9:0] m68_80;
   assign m68_80 =10'b0;

   // m68_81 = W*in
   wire signed [9:0] m68_81;
   assign m68_81 =10'b0;

   // m69_1 = W*in
   wire signed [9:0] m69_1;
   assign m69_1 =10'b0;

   // m69_2 = W*in
   wire signed [9:0] m69_2;
   assign m69_2 =10'b0;

   // m69_3 = W*in
   wire signed [9:0] m69_3;
   assign m69_3 =10'b0;

   // m69_4 = W*in
   wire signed [9:0] m69_4;
   assign m69_4 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_5 = W*in
   wire signed [9:0] m69_5;
   assign m69_5 =10'b0;

   // m69_6 = W*in
   wire signed [9:0] m69_6;
   assign m69_6 =10'b0;

   // m69_7 = W*in
   wire signed [9:0] m69_7;
   assign m69_7 =10'b0;

   // m69_8 = W*in
   wire signed [9:0] m69_8;
   assign m69_8 =10'b0;

   // m69_9 = W*in
   wire signed [9:0] m69_9;
   assign m69_9 =10'b0;

   // m69_10 = W*in
   wire signed [9:0] m69_10;
   assign m69_10 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_11 = W*in
   wire signed [9:0] m69_11;
   assign m69_11 =10'b0;

   // m69_12 = W*in
   wire signed [9:0] m69_12;
   assign m69_12 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_13 = W*in
   wire signed [9:0] m69_13;
   assign m69_13 =10'b0;

   // m69_14 = W*in
   wire signed [9:0] m69_14;
   assign m69_14 =10'b0;

   // m69_15 = W*in
   wire signed [9:0] m69_15;
   assign m69_15 =10'b0;

   // m69_16 = W*in
   wire signed [9:0] m69_16;
   assign m69_16 =10'b0;

   // m69_17 = W*in
   wire signed [9:0] m69_17;
   assign m69_17 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_18 = W*in
   wire signed [9:0] m69_18;
   assign m69_18 =10'b0;

   // m69_19 = W*in
   wire signed [9:0] m69_19;
   assign m69_19 =10'b0;

   // m69_20 = W*in
   wire signed [9:0] m69_20;
   assign m69_20 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_21 = W*in
   wire signed [9:0] m69_21;
   assign m69_21 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_22 = W*in
   wire signed [9:0] m69_22;
   assign m69_22 =10'b0;

   // m69_23 = W*in
   wire signed [9:0] m69_23;
   assign m69_23 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_24 = W*in
   wire signed [9:0] m69_24;
   assign m69_24 =10'b0;

   // m69_25 = W*in
   wire signed [9:0] m69_25;
   assign m69_25 =10'b0;

   // m69_26 = W*in
   wire signed [9:0] m69_26;
   assign m69_26 =10'b0;

   // m69_27 = W*in
   wire signed [9:0] m69_27;
   assign m69_27 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_28 = W*in
   wire signed [9:0] m69_28;
   assign m69_28 =10'b0;

   // m69_29 = W*in
   wire signed [9:0] m69_29;
   assign m69_29 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_30 = W*in
   wire signed [9:0] m69_30;
   assign m69_30 =10'b0;

   // m69_31 = W*in
   wire signed [9:0] m69_31;
   assign m69_31 =10'b0;

   // m69_32 = W*in
   wire signed [9:0] m69_32;
   assign m69_32 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_33 = W*in
   wire signed [9:0] m69_33;
   assign m69_33 =10'b0;

   // m69_34 = W*in
   wire signed [9:0] m69_34;
   assign m69_34 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_35 = W*in
   wire signed [9:0] m69_35;
   assign m69_35 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_36 = W*in
   wire signed [9:0] m69_36;
   assign m69_36 =10'b0;

   // m69_37 = W*in
   wire signed [9:0] m69_37;
   assign m69_37 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_38 = W*in
   wire signed [9:0] m69_38;
   assign m69_38 =10'b0;

   // m69_39 = W*in
   wire signed [9:0] m69_39;
   assign m69_39 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_40 = W*in
   wire signed [9:0] m69_40;
   assign m69_40 =10'b0;

   // m69_41 = W*in
   wire signed [9:0] m69_41;
   assign m69_41 =10'b0;

   // m69_42 = W*in
   wire signed [9:0] m69_42;
   assign m69_42 =10'b0;

   // m69_43 = W*in
   wire signed [9:0] m69_43;
   assign m69_43 =10'b0;

   // m69_44 = W*in
   wire signed [9:0] m69_44;
   assign m69_44 =10'b0;

   // m69_45 = W*in
   wire signed [9:0] m69_45;
   assign m69_45 =10'b0;

   // m69_46 = W*in
   wire signed [9:0] m69_46;
   assign m69_46 =10'b0;

   // m69_47 = W*in
   wire signed [9:0] m69_47;
   assign m69_47 =10'b0;

   // m69_48 = W*in
   wire signed [9:0] m69_48;
   assign m69_48 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_49 = W*in
   wire signed [9:0] m69_49;
   assign m69_49 =10'b0;

   // m69_50 = W*in
   wire signed [9:0] m69_50;
   assign m69_50 =10'b0;

   // m69_51 = W*in
   wire signed [9:0] m69_51;
   assign m69_51 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_52 = W*in
   wire signed [9:0] m69_52;
   assign m69_52 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_53 = W*in
   wire signed [9:0] m69_53;
   assign m69_53 =10'b0;

   // m69_54 = W*in
   wire signed [9:0] m69_54;
   assign m69_54 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_55 = W*in
   wire signed [9:0] m69_55;
   assign m69_55 =10'b0;

   // m69_56 = W*in
   wire signed [9:0] m69_56;
   assign m69_56 =10'b0;

   // m69_57 = W*in
   wire signed [9:0] m69_57;
   assign m69_57 =10'b0;

   // m69_58 = W*in
   wire signed [9:0] m69_58;
   assign m69_58 =10'b0;

   // m69_59 = W*in
   wire signed [9:0] m69_59;
   assign m69_59 =10'b0;

   // m69_60 = W*in
   wire signed [9:0] m69_60;
   assign m69_60 =10'b0;

   // m69_61 = W*in
   wire signed [9:0] m69_61;
   assign m69_61 =10'b0;

   // m69_62 = W*in
   wire signed [9:0] m69_62;
   assign m69_62 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_63 = W*in
   wire signed [9:0] m69_63;
   assign m69_63 ={ {3{neg69[5]}} , neg69 , {1{1'b0}} };

   // m69_64 = W*in
   wire signed [9:0] m69_64;
   assign m69_64 =10'b0;

   // m69_65 = W*in
   wire signed [9:0] m69_65;
   assign m69_65 =10'b0;

   // m69_66 = W*in
   wire signed [9:0] m69_66;
   assign m69_66 =10'b0;

   // m69_67 = W*in
   wire signed [9:0] m69_67;
   assign m69_67 =10'b0;

   // m69_68 = W*in
   wire signed [9:0] m69_68;
   assign m69_68 =10'b0;

   // m69_69 = W*in
   wire signed [9:0] m69_69;
   assign m69_69 =10'b0;

   // m69_70 = W*in
   wire signed [9:0] m69_70;
   assign m69_70 =10'b0;

   // m69_71 = W*in
   wire signed [9:0] m69_71;
   assign m69_71 =10'b0;

   // m69_72 = W*in
   wire signed [9:0] m69_72;
   assign m69_72 =10'b0;

   // m69_73 = W*in
   wire signed [9:0] m69_73;
   assign m69_73 =10'b0;

   // m69_74 = W*in
   wire signed [9:0] m69_74;
   assign m69_74 =10'b0;

   // m69_75 = W*in
   wire signed [9:0] m69_75;
   assign m69_75 =10'b0;

   // m69_76 = W*in
   wire signed [9:0] m69_76;
   assign m69_76 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_77 = W*in
   wire signed [9:0] m69_77;
   assign m69_77 ={ {2{in69[5]}} , in69 , {2{1'b0}} };

   // m69_78 = W*in
   wire signed [9:0] m69_78;
   assign m69_78 ={ {3{in69[5]}} , in69 , {1{1'b0}} };

   // m69_79 = W*in
   wire signed [9:0] m69_79;
   assign m69_79 =10'b0;

   // m69_80 = W*in
   wire signed [9:0] m69_80;
   assign m69_80 =10'b0;

   // m69_81 = W*in
   wire signed [9:0] m69_81;
   assign m69_81 =10'b0;

   // m70_1 = W*in
   wire signed [9:0] m70_1;
   assign m70_1 =10'b0;

   // m70_2 = W*in
   wire signed [9:0] m70_2;
   assign m70_2 =10'b0;

   // m70_3 = W*in
   wire signed [9:0] m70_3;
   assign m70_3 =10'b0;

   // m70_4 = W*in
   wire signed [9:0] m70_4;
   assign m70_4 ={ {2{in70[5]}} , in70 , {2{1'b0}} };

   // m70_5 = W*in
   wire signed [9:0] m70_5;
   assign m70_5 =10'b0;

   // m70_6 = W*in
   wire signed [9:0] m70_6;
   assign m70_6 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_7 = W*in
   wire signed [9:0] m70_7;
   assign m70_7 =10'b0;

   // m70_8 = W*in
   wire signed [9:0] m70_8;
   assign m70_8 =10'b0;

   // m70_9 = W*in
   wire signed [9:0] m70_9;
   assign m70_9 =10'b0;

   // m70_10 = W*in
   wire signed [9:0] m70_10;
   assign m70_10 ={ {2{in70[5]}} , in70 , {2{1'b0}} };

   // m70_11 = W*in
   wire signed [9:0] m70_11;
   assign m70_11 =10'b0;

   // m70_12 = W*in
   wire signed [9:0] m70_12;
   assign m70_12 =10'b0;

   // m70_13 = W*in
   wire signed [9:0] m70_13;
   assign m70_13 =10'b0;

   // m70_14 = W*in
   wire signed [9:0] m70_14;
   assign m70_14 =10'b0;

   // m70_15 = W*in
   wire signed [9:0] m70_15;
   assign m70_15 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_16 = W*in
   wire signed [9:0] m70_16;
   assign m70_16 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_17 = W*in
   wire signed [9:0] m70_17;
   assign m70_17 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_18 = W*in
   wire signed [9:0] m70_18;
   assign m70_18 =10'b0;

   // m70_19 = W*in
   wire signed [9:0] m70_19;
   assign m70_19 =10'b0;

   // m70_20 = W*in
   wire signed [9:0] m70_20;
   assign m70_20 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_21 = W*in
   wire signed [9:0] m70_21;
   assign m70_21 ={ {2{in70[5]}} , in70 , {2{1'b0}} };

   // m70_22 = W*in
   wire signed [9:0] m70_22;
   assign m70_22 =10'b0;

   // m70_23 = W*in
   wire signed [9:0] m70_23;
   assign m70_23 =10'b0;

   // m70_24 = W*in
   wire signed [9:0] m70_24;
   assign m70_24 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_25 = W*in
   wire signed [9:0] m70_25;
   assign m70_25 =10'b0;

   // m70_26 = W*in
   wire signed [9:0] m70_26;
   assign m70_26 =10'b0;

   // m70_27 = W*in
   wire signed [9:0] m70_27;
   assign m70_27 =10'b0;

   // m70_28 = W*in
   wire signed [9:0] m70_28;
   assign m70_28 =10'b0;

   // m70_29 = W*in
   wire signed [9:0] m70_29;
   assign m70_29 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_30 = W*in
   wire signed [9:0] m70_30;
   assign m70_30 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_31 = W*in
   wire signed [9:0] m70_31;
   assign m70_31 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_32 = W*in
   wire signed [9:0] m70_32;
   assign m70_32 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_33 = W*in
   wire signed [9:0] m70_33;
   assign m70_33 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_34 = W*in
   wire signed [9:0] m70_34;
   assign m70_34 ={ {2{in70[5]}} , in70 , {2{1'b0}} };

   // m70_35 = W*in
   wire signed [9:0] m70_35;
   assign m70_35 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_36 = W*in
   wire signed [9:0] m70_36;
   assign m70_36 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_37 = W*in
   wire signed [9:0] m70_37;
   assign m70_37 =10'b0;

   // m70_38 = W*in
   wire signed [9:0] m70_38;
   assign m70_38 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_39 = W*in
   wire signed [9:0] m70_39;
   assign m70_39 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_40 = W*in
   wire signed [9:0] m70_40;
   assign m70_40 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_41 = W*in
   wire signed [9:0] m70_41;
   assign m70_41 =10'b0;

   // m70_42 = W*in
   wire signed [9:0] m70_42;
   assign m70_42 =10'b0;

   // m70_43 = W*in
   wire signed [9:0] m70_43;
   assign m70_43 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_44 = W*in
   wire signed [9:0] m70_44;
   assign m70_44 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_45 = W*in
   wire signed [9:0] m70_45;
   assign m70_45 =10'b0;

   // m70_46 = W*in
   wire signed [9:0] m70_46;
   assign m70_46 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_47 = W*in
   wire signed [9:0] m70_47;
   assign m70_47 =10'b0;

   // m70_48 = W*in
   wire signed [9:0] m70_48;
   assign m70_48 =10'b0;

   // m70_49 = W*in
   wire signed [9:0] m70_49;
   assign m70_49 =10'b0;

   // m70_50 = W*in
   wire signed [9:0] m70_50;
   assign m70_50 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_51 = W*in
   wire signed [9:0] m70_51;
   assign m70_51 =10'b0;

   // m70_52 = W*in
   wire signed [9:0] m70_52;
   assign m70_52 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_53 = W*in
   wire signed [9:0] m70_53;
   assign m70_53 =10'b0;

   // m70_54 = W*in
   wire signed [9:0] m70_54;
   assign m70_54 =10'b0;

   // m70_55 = W*in
   wire signed [9:0] m70_55;
   assign m70_55 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_56 = W*in
   wire signed [9:0] m70_56;
   assign m70_56 =10'b0;

   // m70_57 = W*in
   wire signed [9:0] m70_57;
   assign m70_57 =10'b0;

   // m70_58 = W*in
   wire signed [9:0] m70_58;
   assign m70_58 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_59 = W*in
   wire signed [9:0] m70_59;
   assign m70_59 =10'b0;

   // m70_60 = W*in
   wire signed [9:0] m70_60;
   assign m70_60 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_61 = W*in
   wire signed [9:0] m70_61;
   assign m70_61 =10'b0;

   // m70_62 = W*in
   wire signed [9:0] m70_62;
   assign m70_62 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_63 = W*in
   wire signed [9:0] m70_63;
   assign m70_63 =10'b0;

   // m70_64 = W*in
   wire signed [9:0] m70_64;
   assign m70_64 =10'b0;

   // m70_65 = W*in
   wire signed [9:0] m70_65;
   assign m70_65 =10'b0;

   // m70_66 = W*in
   wire signed [9:0] m70_66;
   assign m70_66 =10'b0;

   // m70_67 = W*in
   wire signed [9:0] m70_67;
   assign m70_67 =10'b0;

   // m70_68 = W*in
   wire signed [9:0] m70_68;
   assign m70_68 ={ {3{in70[5]}} , in70 , {1{1'b0}} };

   // m70_69 = W*in
   wire signed [9:0] m70_69;
   assign m70_69 =10'b0;

   // m70_70 = W*in
   wire signed [9:0] m70_70;
   assign m70_70 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_71 = W*in
   wire signed [9:0] m70_71;
   assign m70_71 =10'b0;

   // m70_72 = W*in
   wire signed [9:0] m70_72;
   assign m70_72 =10'b0;

   // m70_73 = W*in
   wire signed [9:0] m70_73;
   assign m70_73 =10'b0;

   // m70_74 = W*in
   wire signed [9:0] m70_74;
   assign m70_74 =10'b0;

   // m70_75 = W*in
   wire signed [9:0] m70_75;
   assign m70_75 =10'b0;

   // m70_76 = W*in
   wire signed [9:0] m70_76;
   assign m70_76 =10'b0;

   // m70_77 = W*in
   wire signed [9:0] m70_77;
   assign m70_77 ={ {2{in70[5]}} , in70 , {2{1'b0}} };

   // m70_78 = W*in
   wire signed [9:0] m70_78;
   assign m70_78 =10'b0;

   // m70_79 = W*in
   wire signed [9:0] m70_79;
   assign m70_79 ={ {3{neg70[5]}} , neg70 , {1{1'b0}} };

   // m70_80 = W*in
   wire signed [9:0] m70_80;
   assign m70_80 =10'b0;

   // m70_81 = W*in
   wire signed [9:0] m70_81;
   assign m70_81 =10'b0;

   // m71_1 = W*in
   wire signed [9:0] m71_1;
   assign m71_1 =10'b0;

   // m71_2 = W*in
   wire signed [9:0] m71_2;
   assign m71_2 =10'b0;

   // m71_3 = W*in
   wire signed [9:0] m71_3;
   assign m71_3 =10'b0;

   // m71_4 = W*in
   wire signed [9:0] m71_4;
   assign m71_4 =10'b0;

   // m71_5 = W*in
   wire signed [9:0] m71_5;
   assign m71_5 =10'b0;

   // m71_6 = W*in
   wire signed [9:0] m71_6;
   assign m71_6 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_7 = W*in
   wire signed [9:0] m71_7;
   assign m71_7 =10'b0;

   // m71_8 = W*in
   wire signed [9:0] m71_8;
   assign m71_8 ={ {2{in71[5]}} , in71 , {2{1'b0}} };

   // m71_9 = W*in
   wire signed [9:0] m71_9;
   assign m71_9 =10'b0;

   // m71_10 = W*in
   wire signed [9:0] m71_10;
   assign m71_10 =10'b0;

   // m71_11 = W*in
   wire signed [9:0] m71_11;
   assign m71_11 =10'b0;

   // m71_12 = W*in
   wire signed [9:0] m71_12;
   assign m71_12 =10'b0;

   // m71_13 = W*in
   wire signed [9:0] m71_13;
   assign m71_13 =10'b0;

   // m71_14 = W*in
   wire signed [9:0] m71_14;
   assign m71_14 =10'b0;

   // m71_15 = W*in
   wire signed [9:0] m71_15;
   assign m71_15 =10'b0;

   // m71_16 = W*in
   wire signed [9:0] m71_16;
   assign m71_16 =10'b0;

   // m71_17 = W*in
   wire signed [9:0] m71_17;
   assign m71_17 =10'b0;

   // m71_18 = W*in
   wire signed [9:0] m71_18;
   assign m71_18 =10'b0;

   // m71_19 = W*in
   wire signed [9:0] m71_19;
   assign m71_19 =10'b0;

   // m71_20 = W*in
   wire signed [9:0] m71_20;
   assign m71_20 =10'b0;

   // m71_21 = W*in
   wire signed [9:0] m71_21;
   assign m71_21 =10'b0;

   // m71_22 = W*in
   wire signed [9:0] m71_22;
   assign m71_22 ={ {3{neg71[5]}} , neg71 , {1{1'b0}} };

   // m71_23 = W*in
   wire signed [9:0] m71_23;
   assign m71_23 =10'b0;

   // m71_24 = W*in
   wire signed [9:0] m71_24;
   assign m71_24 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_25 = W*in
   wire signed [9:0] m71_25;
   assign m71_25 ={ {2{in71[5]}} , in71 , {2{1'b0}} };

   // m71_26 = W*in
   wire signed [9:0] m71_26;
   assign m71_26 =10'b0;

   // m71_27 = W*in
   wire signed [9:0] m71_27;
   assign m71_27 =10'b0;

   // m71_28 = W*in
   wire signed [9:0] m71_28;
   assign m71_28 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_29 = W*in
   wire signed [9:0] m71_29;
   assign m71_29 =10'b0;

   // m71_30 = W*in
   wire signed [9:0] m71_30;
   assign m71_30 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_31 = W*in
   wire signed [9:0] m71_31;
   assign m71_31 =10'b0;

   // m71_32 = W*in
   wire signed [9:0] m71_32;
   assign m71_32 =10'b0;

   // m71_33 = W*in
   wire signed [9:0] m71_33;
   assign m71_33 ={ {2{in71[5]}} , in71 , {2{1'b0}} };

   // m71_34 = W*in
   wire signed [9:0] m71_34;
   assign m71_34 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_35 = W*in
   wire signed [9:0] m71_35;
   assign m71_35 =10'b0;

   // m71_36 = W*in
   wire signed [9:0] m71_36;
   assign m71_36 =10'b0;

   // m71_37 = W*in
   wire signed [9:0] m71_37;
   assign m71_37 ={ {2{in71[5]}} , in71 , {2{1'b0}} };

   // m71_38 = W*in
   wire signed [9:0] m71_38;
   assign m71_38 =10'b0;

   // m71_39 = W*in
   wire signed [9:0] m71_39;
   assign m71_39 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_40 = W*in
   wire signed [9:0] m71_40;
   assign m71_40 =10'b0;

   // m71_41 = W*in
   wire signed [9:0] m71_41;
   assign m71_41 =10'b0;

   // m71_42 = W*in
   wire signed [9:0] m71_42;
   assign m71_42 =10'b0;

   // m71_43 = W*in
   wire signed [9:0] m71_43;
   assign m71_43 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_44 = W*in
   wire signed [9:0] m71_44;
   assign m71_44 =10'b0;

   // m71_45 = W*in
   wire signed [9:0] m71_45;
   assign m71_45 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_46 = W*in
   wire signed [9:0] m71_46;
   assign m71_46 =10'b0;

   // m71_47 = W*in
   wire signed [9:0] m71_47;
   assign m71_47 =10'b0;

   // m71_48 = W*in
   wire signed [9:0] m71_48;
   assign m71_48 =10'b0;

   // m71_49 = W*in
   wire signed [9:0] m71_49;
   assign m71_49 =10'b0;

   // m71_50 = W*in
   wire signed [9:0] m71_50;
   assign m71_50 =10'b0;

   // m71_51 = W*in
   wire signed [9:0] m71_51;
   assign m71_51 =10'b0;

   // m71_52 = W*in
   wire signed [9:0] m71_52;
   assign m71_52 ={ {3{neg71[5]}} , neg71 , {1{1'b0}} };

   // m71_53 = W*in
   wire signed [9:0] m71_53;
   assign m71_53 =10'b0;

   // m71_54 = W*in
   wire signed [9:0] m71_54;
   assign m71_54 =10'b0;

   // m71_55 = W*in
   wire signed [9:0] m71_55;
   assign m71_55 =10'b0;

   // m71_56 = W*in
   wire signed [9:0] m71_56;
   assign m71_56 =10'b0;

   // m71_57 = W*in
   wire signed [9:0] m71_57;
   assign m71_57 =10'b0;

   // m71_58 = W*in
   wire signed [9:0] m71_58;
   assign m71_58 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_59 = W*in
   wire signed [9:0] m71_59;
   assign m71_59 =10'b0;

   // m71_60 = W*in
   wire signed [9:0] m71_60;
   assign m71_60 =10'b0;

   // m71_61 = W*in
   wire signed [9:0] m71_61;
   assign m71_61 =10'b0;

   // m71_62 = W*in
   wire signed [9:0] m71_62;
   assign m71_62 =10'b0;

   // m71_63 = W*in
   wire signed [9:0] m71_63;
   assign m71_63 ={ {3{in71[5]}} , in71 , {1{1'b0}} };

   // m71_64 = W*in
   wire signed [9:0] m71_64;
   assign m71_64 =10'b0;

   // m71_65 = W*in
   wire signed [9:0] m71_65;
   assign m71_65 =10'b0;

   // m71_66 = W*in
   wire signed [9:0] m71_66;
   assign m71_66 =10'b0;

   // m71_67 = W*in
   wire signed [9:0] m71_67;
   assign m71_67 =10'b0;

   // m71_68 = W*in
   wire signed [9:0] m71_68;
   assign m71_68 =10'b0;

   // m71_69 = W*in
   wire signed [9:0] m71_69;
   assign m71_69 =10'b0;

   // m71_70 = W*in
   wire signed [9:0] m71_70;
   assign m71_70 =10'b0;

   // m71_71 = W*in
   wire signed [9:0] m71_71;
   assign m71_71 =10'b0;

   // m71_72 = W*in
   wire signed [9:0] m71_72;
   assign m71_72 =10'b0;

   // m71_73 = W*in
   wire signed [9:0] m71_73;
   assign m71_73 =10'b0;

   // m71_74 = W*in
   wire signed [9:0] m71_74;
   assign m71_74 =10'b0;

   // m71_75 = W*in
   wire signed [9:0] m71_75;
   assign m71_75 =10'b0;

   // m71_76 = W*in
   wire signed [9:0] m71_76;
   assign m71_76 =10'b0;

   // m71_77 = W*in
   wire signed [9:0] m71_77;
   assign m71_77 =10'b0;

   // m71_78 = W*in
   wire signed [9:0] m71_78;
   assign m71_78 =10'b0;

   // m71_79 = W*in
   wire signed [9:0] m71_79;
   assign m71_79 =10'b0;

   // m71_80 = W*in
   wire signed [9:0] m71_80;
   assign m71_80 =10'b0;

   // m71_81 = W*in
   wire signed [9:0] m71_81;
   assign m71_81 =10'b0;

   // m72_1 = W*in
   wire signed [9:0] m72_1;
   assign m72_1 =10'b0;

   // m72_2 = W*in
   wire signed [9:0] m72_2;
   assign m72_2 =10'b0;

   // m72_3 = W*in
   wire signed [9:0] m72_3;
   assign m72_3 =10'b0;

   // m72_4 = W*in
   wire signed [9:0] m72_4;
   assign m72_4 =10'b0;

   // m72_5 = W*in
   wire signed [9:0] m72_5;
   assign m72_5 =10'b0;

   // m72_6 = W*in
   wire signed [9:0] m72_6;
   assign m72_6 =10'b0;

   // m72_7 = W*in
   wire signed [9:0] m72_7;
   assign m72_7 =10'b0;

   // m72_8 = W*in
   wire signed [9:0] m72_8;
   assign m72_8 =10'b0;

   // m72_9 = W*in
   wire signed [9:0] m72_9;
   assign m72_9 =10'b0;

   // m72_10 = W*in
   wire signed [9:0] m72_10;
   assign m72_10 =10'b0;

   // m72_11 = W*in
   wire signed [9:0] m72_11;
   assign m72_11 =10'b0;

   // m72_12 = W*in
   wire signed [9:0] m72_12;
   assign m72_12 =10'b0;

   // m72_13 = W*in
   wire signed [9:0] m72_13;
   assign m72_13 =10'b0;

   // m72_14 = W*in
   wire signed [9:0] m72_14;
   assign m72_14 =10'b0;

   // m72_15 = W*in
   wire signed [9:0] m72_15;
   assign m72_15 =10'b0;

   // m72_16 = W*in
   wire signed [9:0] m72_16;
   assign m72_16 =10'b0;

   // m72_17 = W*in
   wire signed [9:0] m72_17;
   assign m72_17 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_18 = W*in
   wire signed [9:0] m72_18;
   assign m72_18 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_19 = W*in
   wire signed [9:0] m72_19;
   assign m72_19 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_20 = W*in
   wire signed [9:0] m72_20;
   assign m72_20 =10'b0;

   // m72_21 = W*in
   wire signed [9:0] m72_21;
   assign m72_21 =10'b0;

   // m72_22 = W*in
   wire signed [9:0] m72_22;
   assign m72_22 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_23 = W*in
   wire signed [9:0] m72_23;
   assign m72_23 ={ {2{in72[5]}} , in72 , {2{1'b0}} };

   // m72_24 = W*in
   wire signed [9:0] m72_24;
   assign m72_24 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_25 = W*in
   wire signed [9:0] m72_25;
   assign m72_25 ={ {2{in72[5]}} , in72 , {2{1'b0}} };

   // m72_26 = W*in
   wire signed [9:0] m72_26;
   assign m72_26 =10'b0;

   // m72_27 = W*in
   wire signed [9:0] m72_27;
   assign m72_27 =10'b0;

   // m72_28 = W*in
   wire signed [9:0] m72_28;
   assign m72_28 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_29 = W*in
   wire signed [9:0] m72_29;
   assign m72_29 =10'b0;

   // m72_30 = W*in
   wire signed [9:0] m72_30;
   assign m72_30 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_31 = W*in
   wire signed [9:0] m72_31;
   assign m72_31 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_32 = W*in
   wire signed [9:0] m72_32;
   assign m72_32 =10'b0;

   // m72_33 = W*in
   wire signed [9:0] m72_33;
   assign m72_33 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_34 = W*in
   wire signed [9:0] m72_34;
   assign m72_34 =10'b0;

   // m72_35 = W*in
   wire signed [9:0] m72_35;
   assign m72_35 =10'b0;

   // m72_36 = W*in
   wire signed [9:0] m72_36;
   assign m72_36 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_37 = W*in
   wire signed [9:0] m72_37;
   assign m72_37 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_38 = W*in
   wire signed [9:0] m72_38;
   assign m72_38 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_39 = W*in
   wire signed [9:0] m72_39;
   assign m72_39 ={ {2{in72[5]}} , in72 , {2{1'b0}} };

   // m72_40 = W*in
   wire signed [9:0] m72_40;
   assign m72_40 =10'b0;

   // m72_41 = W*in
   wire signed [9:0] m72_41;
   assign m72_41 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_42 = W*in
   wire signed [9:0] m72_42;
   assign m72_42 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_43 = W*in
   wire signed [9:0] m72_43;
   assign m72_43 =10'b0;

   // m72_44 = W*in
   wire signed [9:0] m72_44;
   assign m72_44 =10'b0;

   // m72_45 = W*in
   wire signed [9:0] m72_45;
   assign m72_45 =10'b0;

   // m72_46 = W*in
   wire signed [9:0] m72_46;
   assign m72_46 =10'b0;

   // m72_47 = W*in
   wire signed [9:0] m72_47;
   assign m72_47 =10'b0;

   // m72_48 = W*in
   wire signed [9:0] m72_48;
   assign m72_48 =10'b0;

   // m72_49 = W*in
   wire signed [9:0] m72_49;
   assign m72_49 =10'b0;

   // m72_50 = W*in
   wire signed [9:0] m72_50;
   assign m72_50 =10'b0;

   // m72_51 = W*in
   wire signed [9:0] m72_51;
   assign m72_51 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_52 = W*in
   wire signed [9:0] m72_52;
   assign m72_52 =10'b0;

   // m72_53 = W*in
   wire signed [9:0] m72_53;
   assign m72_53 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_54 = W*in
   wire signed [9:0] m72_54;
   assign m72_54 =10'b0;

   // m72_55 = W*in
   wire signed [9:0] m72_55;
   assign m72_55 =10'b0;

   // m72_56 = W*in
   wire signed [9:0] m72_56;
   assign m72_56 =10'b0;

   // m72_57 = W*in
   wire signed [9:0] m72_57;
   assign m72_57 =10'b0;

   // m72_58 = W*in
   wire signed [9:0] m72_58;
   assign m72_58 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_59 = W*in
   wire signed [9:0] m72_59;
   assign m72_59 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_60 = W*in
   wire signed [9:0] m72_60;
   assign m72_60 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_61 = W*in
   wire signed [9:0] m72_61;
   assign m72_61 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_62 = W*in
   wire signed [9:0] m72_62;
   assign m72_62 =10'b0;

   // m72_63 = W*in
   wire signed [9:0] m72_63;
   assign m72_63 =10'b0;

   // m72_64 = W*in
   wire signed [9:0] m72_64;
   assign m72_64 =10'b0;

   // m72_65 = W*in
   wire signed [9:0] m72_65;
   assign m72_65 =10'b0;

   // m72_66 = W*in
   wire signed [9:0] m72_66;
   assign m72_66 =10'b0;

   // m72_67 = W*in
   wire signed [9:0] m72_67;
   assign m72_67 ={ {4{in72[5]}} , in72[5:0] };

   // m72_68 = W*in
   wire signed [9:0] m72_68;
   assign m72_68 =10'b0;

   // m72_69 = W*in
   wire signed [9:0] m72_69;
   assign m72_69 =10'b0;

   // m72_70 = W*in
   wire signed [9:0] m72_70;
   assign m72_70 =10'b0;

   // m72_71 = W*in
   wire signed [9:0] m72_71;
   assign m72_71 ={ {2{in72[5]}} , in72 , {2{1'b0}} };

   // m72_72 = W*in
   wire signed [9:0] m72_72;
   assign m72_72 =10'b0;

   // m72_73 = W*in
   wire signed [9:0] m72_73;
   assign m72_73 =10'b0;

   // m72_74 = W*in
   wire signed [9:0] m72_74;
   assign m72_74 =10'b0;

   // m72_75 = W*in
   wire signed [9:0] m72_75;
   assign m72_75 ={ {3{in72[5]}} , in72 , {1{1'b0}} };

   // m72_76 = W*in
   wire signed [9:0] m72_76;
   assign m72_76 =10'b0;

   // m72_77 = W*in
   wire signed [9:0] m72_77;
   assign m72_77 =10'b0;

   // m72_78 = W*in
   wire signed [9:0] m72_78;
   assign m72_78 =10'b0;

   // m72_79 = W*in
   wire signed [9:0] m72_79;
   assign m72_79 =10'b0;

   // m72_80 = W*in
   wire signed [9:0] m72_80;
   assign m72_80 =10'b0;

   // m72_81 = W*in
   wire signed [9:0] m72_81;
   assign m72_81 =10'b0;

   // m73_1 = W*in
   wire signed [9:0] m73_1;
   assign m73_1 =10'b0;

   // m73_2 = W*in
   wire signed [9:0] m73_2;
   assign m73_2 =10'b0;

   // m73_3 = W*in
   wire signed [9:0] m73_3;
   assign m73_3 ={ {2{in73[5]}} , in73 , {2{1'b0}} };

   // m73_4 = W*in
   wire signed [9:0] m73_4;
   assign m73_4 =10'b0;

   // m73_5 = W*in
   wire signed [9:0] m73_5;
   assign m73_5 =10'b0;

   // m73_6 = W*in
   wire signed [9:0] m73_6;
   assign m73_6 ={ {3{neg73[5]}} , neg73 , {1{1'b0}} };

   // m73_7 = W*in
   wire signed [9:0] m73_7;
   assign m73_7 =10'b0;

   // m73_8 = W*in
   wire signed [9:0] m73_8;
   assign m73_8 =10'b0;

   // m73_9 = W*in
   wire signed [9:0] m73_9;
   assign m73_9 =10'b0;

   // m73_10 = W*in
   wire signed [9:0] m73_10;
   assign m73_10 =10'b0;

   // m73_11 = W*in
   wire signed [9:0] m73_11;
   assign m73_11 =10'b0;

   // m73_12 = W*in
   wire signed [9:0] m73_12;
   assign m73_12 =10'b0;

   // m73_13 = W*in
   wire signed [9:0] m73_13;
   assign m73_13 =10'b0;

   // m73_14 = W*in
   wire signed [9:0] m73_14;
   assign m73_14 =10'b0;

   // m73_15 = W*in
   wire signed [9:0] m73_15;
   assign m73_15 ={ {2{in73[5]}} , in73 , {2{1'b0}} };

   // m73_16 = W*in
   wire signed [9:0] m73_16;
   assign m73_16 =10'b0;

   // m73_17 = W*in
   wire signed [9:0] m73_17;
   assign m73_17 ={ {3{neg73[5]}} , neg73 , {1{1'b0}} };

   // m73_18 = W*in
   wire signed [9:0] m73_18;
   assign m73_18 =10'b0;

   // m73_19 = W*in
   wire signed [9:0] m73_19;
   assign m73_19 =10'b0;

   // m73_20 = W*in
   wire signed [9:0] m73_20;
   assign m73_20 =10'b0;

   // m73_21 = W*in
   wire signed [9:0] m73_21;
   assign m73_21 ={ {3{neg73[5]}} , neg73 , {1{1'b0}} };

   // m73_22 = W*in
   wire signed [9:0] m73_22;
   assign m73_22 =10'b0;

   // m73_23 = W*in
   wire signed [9:0] m73_23;
   assign m73_23 =10'b0;

   // m73_24 = W*in
   wire signed [9:0] m73_24;
   assign m73_24 =10'b0;

   // m73_25 = W*in
   wire signed [9:0] m73_25;
   assign m73_25 =10'b0;

   // m73_26 = W*in
   wire signed [9:0] m73_26;
   assign m73_26 =10'b0;

   // m73_27 = W*in
   wire signed [9:0] m73_27;
   assign m73_27 =10'b0;

   // m73_28 = W*in
   wire signed [9:0] m73_28;
   assign m73_28 =10'b0;

   // m73_29 = W*in
   wire signed [9:0] m73_29;
   assign m73_29 =10'b0;

   // m73_30 = W*in
   wire signed [9:0] m73_30;
   assign m73_30 =10'b0;

   // m73_31 = W*in
   wire signed [9:0] m73_31;
   assign m73_31 =10'b0;

   // m73_32 = W*in
   wire signed [9:0] m73_32;
   assign m73_32 =10'b0;

   // m73_33 = W*in
   wire signed [9:0] m73_33;
   assign m73_33 =10'b0;

   // m73_34 = W*in
   wire signed [9:0] m73_34;
   assign m73_34 =10'b0;

   // m73_35 = W*in
   wire signed [9:0] m73_35;
   assign m73_35 =10'b0;

   // m73_36 = W*in
   wire signed [9:0] m73_36;
   assign m73_36 =10'b0;

   // m73_37 = W*in
   wire signed [9:0] m73_37;
   assign m73_37 =10'b0;

   // m73_38 = W*in
   wire signed [9:0] m73_38;
   assign m73_38 =10'b0;

   // m73_39 = W*in
   wire signed [9:0] m73_39;
   assign m73_39 =10'b0;

   // m73_40 = W*in
   wire signed [9:0] m73_40;
   assign m73_40 =10'b0;

   // m73_41 = W*in
   wire signed [9:0] m73_41;
   assign m73_41 =10'b0;

   // m73_42 = W*in
   wire signed [9:0] m73_42;
   assign m73_42 =10'b0;

   // m73_43 = W*in
   wire signed [9:0] m73_43;
   assign m73_43 ={ {3{in73[5]}} , in73 , {1{1'b0}} };

   // m73_44 = W*in
   wire signed [9:0] m73_44;
   assign m73_44 ={ {2{in73[5]}} , in73 , {2{1'b0}} };

   // m73_45 = W*in
   wire signed [9:0] m73_45;
   assign m73_45 =10'b0;

   // m73_46 = W*in
   wire signed [9:0] m73_46;
   assign m73_46 =10'b0;

   // m73_47 = W*in
   wire signed [9:0] m73_47;
   assign m73_47 ={ {3{in73[5]}} , in73 , {1{1'b0}} };

   // m73_48 = W*in
   wire signed [9:0] m73_48;
   assign m73_48 =10'b0;

   // m73_49 = W*in
   wire signed [9:0] m73_49;
   assign m73_49 =10'b0;

   // m73_50 = W*in
   wire signed [9:0] m73_50;
   assign m73_50 =10'b0;

   // m73_51 = W*in
   wire signed [9:0] m73_51;
   assign m73_51 =10'b0;

   // m73_52 = W*in
   wire signed [9:0] m73_52;
   assign m73_52 =10'b0;

   // m73_53 = W*in
   wire signed [9:0] m73_53;
   assign m73_53 =10'b0;

   // m73_54 = W*in
   wire signed [9:0] m73_54;
   assign m73_54 =10'b0;

   // m73_55 = W*in
   wire signed [9:0] m73_55;
   assign m73_55 ={ {2{in73[5]}} , in73 , {2{1'b0}} };

   // m73_56 = W*in
   wire signed [9:0] m73_56;
   assign m73_56 =10'b0;

   // m73_57 = W*in
   wire signed [9:0] m73_57;
   assign m73_57 =10'b0;

   // m73_58 = W*in
   wire signed [9:0] m73_58;
   assign m73_58 ={ {3{in73[5]}} , in73 , {1{1'b0}} };

   // m73_59 = W*in
   wire signed [9:0] m73_59;
   assign m73_59 ={ {3{in73[5]}} , in73 , {1{1'b0}} };

   // m73_60 = W*in
   wire signed [9:0] m73_60;
   assign m73_60 =10'b0;

   // m73_61 = W*in
   wire signed [9:0] m73_61;
   assign m73_61 =10'b0;

   // m73_62 = W*in
   wire signed [9:0] m73_62;
   assign m73_62 =10'b0;

   // m73_63 = W*in
   wire signed [9:0] m73_63;
   assign m73_63 =10'b0;

   // m73_64 = W*in
   wire signed [9:0] m73_64;
   assign m73_64 =10'b0;

   // m73_65 = W*in
   wire signed [9:0] m73_65;
   assign m73_65 =10'b0;

   // m73_66 = W*in
   wire signed [9:0] m73_66;
   assign m73_66 =10'b0;

   // m73_67 = W*in
   wire signed [9:0] m73_67;
   assign m73_67 =10'b0;

   // m73_68 = W*in
   wire signed [9:0] m73_68;
   assign m73_68 ={ {3{neg73[5]}} , neg73 , {1{1'b0}} };

   // m73_69 = W*in
   wire signed [9:0] m73_69;
   assign m73_69 ={ {3{in73[5]}} , in73 , {1{1'b0}} };

   // m73_70 = W*in
   wire signed [9:0] m73_70;
   assign m73_70 =10'b0;

   // m73_71 = W*in
   wire signed [9:0] m73_71;
   assign m73_71 =10'b0;

   // m73_72 = W*in
   wire signed [9:0] m73_72;
   assign m73_72 =10'b0;

   // m73_73 = W*in
   wire signed [9:0] m73_73;
   assign m73_73 =10'b0;

   // m73_74 = W*in
   wire signed [9:0] m73_74;
   assign m73_74 =10'b0;

   // m73_75 = W*in
   wire signed [9:0] m73_75;
   assign m73_75 =10'b0;

   // m73_76 = W*in
   wire signed [9:0] m73_76;
   assign m73_76 =10'b0;

   // m73_77 = W*in
   wire signed [9:0] m73_77;
   assign m73_77 ={ {3{neg73[5]}} , neg73 , {1{1'b0}} };

   // m73_78 = W*in
   wire signed [9:0] m73_78;
   assign m73_78 =10'b0;

   // m73_79 = W*in
   wire signed [9:0] m73_79;
   assign m73_79 ={ {3{in73[5]}} , in73 , {1{1'b0}} };

   // m73_80 = W*in
   wire signed [9:0] m73_80;
   assign m73_80 =10'b0;

   // m73_81 = W*in
   wire signed [9:0] m73_81;
   assign m73_81 =10'b0;

   // m74_1 = W*in
   wire signed [9:0] m74_1;
   assign m74_1 =10'b0;

   // m74_2 = W*in
   wire signed [9:0] m74_2;
   assign m74_2 =10'b0;

   // m74_3 = W*in
   wire signed [9:0] m74_3;
   assign m74_3 ={ {3{neg74[5]}} , neg74 , {1{1'b0}} };

   // m74_4 = W*in
   wire signed [9:0] m74_4;
   assign m74_4 =10'b0;

   // m74_5 = W*in
   wire signed [9:0] m74_5;
   assign m74_5 =10'b0;

   // m74_6 = W*in
   wire signed [9:0] m74_6;
   assign m74_6 =10'b0;

   // m74_7 = W*in
   wire signed [9:0] m74_7;
   assign m74_7 =10'b0;

   // m74_8 = W*in
   wire signed [9:0] m74_8;
   assign m74_8 =10'b0;

   // m74_9 = W*in
   wire signed [9:0] m74_9;
   assign m74_9 =10'b0;

   // m74_10 = W*in
   wire signed [9:0] m74_10;
   assign m74_10 =10'b0;

   // m74_11 = W*in
   wire signed [9:0] m74_11;
   assign m74_11 =10'b0;

   // m74_12 = W*in
   wire signed [9:0] m74_12;
   assign m74_12 =10'b0;

   // m74_13 = W*in
   wire signed [9:0] m74_13;
   assign m74_13 ={ {2{in74[5]}} , in74 , {2{1'b0}} };

   // m74_14 = W*in
   wire signed [9:0] m74_14;
   assign m74_14 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_15 = W*in
   wire signed [9:0] m74_15;
   assign m74_15 ={ {3{neg74[5]}} , neg74 , {1{1'b0}} };

   // m74_16 = W*in
   wire signed [9:0] m74_16;
   assign m74_16 =10'b0;

   // m74_17 = W*in
   wire signed [9:0] m74_17;
   assign m74_17 =10'b0;

   // m74_18 = W*in
   wire signed [9:0] m74_18;
   assign m74_18 =10'b0;

   // m74_19 = W*in
   wire signed [9:0] m74_19;
   assign m74_19 =10'b0;

   // m74_20 = W*in
   wire signed [9:0] m74_20;
   assign m74_20 =10'b0;

   // m74_21 = W*in
   wire signed [9:0] m74_21;
   assign m74_21 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_22 = W*in
   wire signed [9:0] m74_22;
   assign m74_22 =10'b0;

   // m74_23 = W*in
   wire signed [9:0] m74_23;
   assign m74_23 =10'b0;

   // m74_24 = W*in
   wire signed [9:0] m74_24;
   assign m74_24 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_25 = W*in
   wire signed [9:0] m74_25;
   assign m74_25 =10'b0;

   // m74_26 = W*in
   wire signed [9:0] m74_26;
   assign m74_26 =10'b0;

   // m74_27 = W*in
   wire signed [9:0] m74_27;
   assign m74_27 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_28 = W*in
   wire signed [9:0] m74_28;
   assign m74_28 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_29 = W*in
   wire signed [9:0] m74_29;
   assign m74_29 =10'b0;

   // m74_30 = W*in
   wire signed [9:0] m74_30;
   assign m74_30 =10'b0;

   // m74_31 = W*in
   wire signed [9:0] m74_31;
   assign m74_31 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_32 = W*in
   wire signed [9:0] m74_32;
   assign m74_32 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_33 = W*in
   wire signed [9:0] m74_33;
   assign m74_33 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_34 = W*in
   wire signed [9:0] m74_34;
   assign m74_34 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_35 = W*in
   wire signed [9:0] m74_35;
   assign m74_35 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_36 = W*in
   wire signed [9:0] m74_36;
   assign m74_36 =10'b0;

   // m74_37 = W*in
   wire signed [9:0] m74_37;
   assign m74_37 =10'b0;

   // m74_38 = W*in
   wire signed [9:0] m74_38;
   assign m74_38 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_39 = W*in
   wire signed [9:0] m74_39;
   assign m74_39 =10'b0;

   // m74_40 = W*in
   wire signed [9:0] m74_40;
   assign m74_40 =10'b0;

   // m74_41 = W*in
   wire signed [9:0] m74_41;
   assign m74_41 =10'b0;

   // m74_42 = W*in
   wire signed [9:0] m74_42;
   assign m74_42 =10'b0;

   // m74_43 = W*in
   wire signed [9:0] m74_43;
   assign m74_43 ={ {3{neg74[5]}} , neg74 , {1{1'b0}} };

   // m74_44 = W*in
   wire signed [9:0] m74_44;
   assign m74_44 ={ {3{neg74[5]}} , neg74 , {1{1'b0}} };

   // m74_45 = W*in
   wire signed [9:0] m74_45;
   assign m74_45 =10'b0;

   // m74_46 = W*in
   wire signed [9:0] m74_46;
   assign m74_46 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_47 = W*in
   wire signed [9:0] m74_47;
   assign m74_47 =10'b0;

   // m74_48 = W*in
   wire signed [9:0] m74_48;
   assign m74_48 =10'b0;

   // m74_49 = W*in
   wire signed [9:0] m74_49;
   assign m74_49 =10'b0;

   // m74_50 = W*in
   wire signed [9:0] m74_50;
   assign m74_50 =10'b0;

   // m74_51 = W*in
   wire signed [9:0] m74_51;
   assign m74_51 =10'b0;

   // m74_52 = W*in
   wire signed [9:0] m74_52;
   assign m74_52 =10'b0;

   // m74_53 = W*in
   wire signed [9:0] m74_53;
   assign m74_53 =10'b0;

   // m74_54 = W*in
   wire signed [9:0] m74_54;
   assign m74_54 =10'b0;

   // m74_55 = W*in
   wire signed [9:0] m74_55;
   assign m74_55 =10'b0;

   // m74_56 = W*in
   wire signed [9:0] m74_56;
   assign m74_56 =10'b0;

   // m74_57 = W*in
   wire signed [9:0] m74_57;
   assign m74_57 =10'b0;

   // m74_58 = W*in
   wire signed [9:0] m74_58;
   assign m74_58 =10'b0;

   // m74_59 = W*in
   wire signed [9:0] m74_59;
   assign m74_59 =10'b0;

   // m74_60 = W*in
   wire signed [9:0] m74_60;
   assign m74_60 =10'b0;

   // m74_61 = W*in
   wire signed [9:0] m74_61;
   assign m74_61 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_62 = W*in
   wire signed [9:0] m74_62;
   assign m74_62 =10'b0;

   // m74_63 = W*in
   wire signed [9:0] m74_63;
   assign m74_63 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_64 = W*in
   wire signed [9:0] m74_64;
   assign m74_64 =10'b0;

   // m74_65 = W*in
   wire signed [9:0] m74_65;
   assign m74_65 =10'b0;

   // m74_66 = W*in
   wire signed [9:0] m74_66;
   assign m74_66 =10'b0;

   // m74_67 = W*in
   wire signed [9:0] m74_67;
   assign m74_67 =10'b0;

   // m74_68 = W*in
   wire signed [9:0] m74_68;
   assign m74_68 ={ {3{in74[5]}} , in74 , {1{1'b0}} };

   // m74_69 = W*in
   wire signed [9:0] m74_69;
   assign m74_69 =10'b0;

   // m74_70 = W*in
   wire signed [9:0] m74_70;
   assign m74_70 =10'b0;

   // m74_71 = W*in
   wire signed [9:0] m74_71;
   assign m74_71 =10'b0;

   // m74_72 = W*in
   wire signed [9:0] m74_72;
   assign m74_72 =10'b0;

   // m74_73 = W*in
   wire signed [9:0] m74_73;
   assign m74_73 =10'b0;

   // m74_74 = W*in
   wire signed [9:0] m74_74;
   assign m74_74 =10'b0;

   // m74_75 = W*in
   wire signed [9:0] m74_75;
   assign m74_75 =10'b0;

   // m74_76 = W*in
   wire signed [9:0] m74_76;
   assign m74_76 =10'b0;

   // m74_77 = W*in
   wire signed [9:0] m74_77;
   assign m74_77 =10'b0;

   // m74_78 = W*in
   wire signed [9:0] m74_78;
   assign m74_78 =10'b0;

   // m74_79 = W*in
   wire signed [9:0] m74_79;
   assign m74_79 =10'b0;

   // m74_80 = W*in
   wire signed [9:0] m74_80;
   assign m74_80 =10'b0;

   // m74_81 = W*in
   wire signed [9:0] m74_81;
   assign m74_81 =10'b0;

   // m75_1 = W*in
   wire signed [9:0] m75_1;
   assign m75_1 =10'b0;

   // m75_2 = W*in
   wire signed [9:0] m75_2;
   assign m75_2 =10'b0;

   // m75_3 = W*in
   wire signed [9:0] m75_3;
   assign m75_3 =10'b0;

   // m75_4 = W*in
   wire signed [9:0] m75_4;
   assign m75_4 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_5 = W*in
   wire signed [9:0] m75_5;
   assign m75_5 =10'b0;

   // m75_6 = W*in
   wire signed [9:0] m75_6;
   assign m75_6 =10'b0;

   // m75_7 = W*in
   wire signed [9:0] m75_7;
   assign m75_7 =10'b0;

   // m75_8 = W*in
   wire signed [9:0] m75_8;
   assign m75_8 =10'b0;

   // m75_9 = W*in
   wire signed [9:0] m75_9;
   assign m75_9 =10'b0;

   // m75_10 = W*in
   wire signed [9:0] m75_10;
   assign m75_10 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_11 = W*in
   wire signed [9:0] m75_11;
   assign m75_11 =10'b0;

   // m75_12 = W*in
   wire signed [9:0] m75_12;
   assign m75_12 =10'b0;

   // m75_13 = W*in
   wire signed [9:0] m75_13;
   assign m75_13 =10'b0;

   // m75_14 = W*in
   wire signed [9:0] m75_14;
   assign m75_14 =10'b0;

   // m75_15 = W*in
   wire signed [9:0] m75_15;
   assign m75_15 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_16 = W*in
   wire signed [9:0] m75_16;
   assign m75_16 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_17 = W*in
   wire signed [9:0] m75_17;
   assign m75_17 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_18 = W*in
   wire signed [9:0] m75_18;
   assign m75_18 ={ {2{in75[5]}} , in75 , {2{1'b0}} };

   // m75_19 = W*in
   wire signed [9:0] m75_19;
   assign m75_19 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_20 = W*in
   wire signed [9:0] m75_20;
   assign m75_20 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_21 = W*in
   wire signed [9:0] m75_21;
   assign m75_21 =10'b0;

   // m75_22 = W*in
   wire signed [9:0] m75_22;
   assign m75_22 =10'b0;

   // m75_23 = W*in
   wire signed [9:0] m75_23;
   assign m75_23 =10'b0;

   // m75_24 = W*in
   wire signed [9:0] m75_24;
   assign m75_24 =10'b0;

   // m75_25 = W*in
   wire signed [9:0] m75_25;
   assign m75_25 =10'b0;

   // m75_26 = W*in
   wire signed [9:0] m75_26;
   assign m75_26 =10'b0;

   // m75_27 = W*in
   wire signed [9:0] m75_27;
   assign m75_27 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_28 = W*in
   wire signed [9:0] m75_28;
   assign m75_28 =10'b0;

   // m75_29 = W*in
   wire signed [9:0] m75_29;
   assign m75_29 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_30 = W*in
   wire signed [9:0] m75_30;
   assign m75_30 =10'b0;

   // m75_31 = W*in
   wire signed [9:0] m75_31;
   assign m75_31 =10'b0;

   // m75_32 = W*in
   wire signed [9:0] m75_32;
   assign m75_32 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_33 = W*in
   wire signed [9:0] m75_33;
   assign m75_33 =10'b0;

   // m75_34 = W*in
   wire signed [9:0] m75_34;
   assign m75_34 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_35 = W*in
   wire signed [9:0] m75_35;
   assign m75_35 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_36 = W*in
   wire signed [9:0] m75_36;
   assign m75_36 =10'b0;

   // m75_37 = W*in
   wire signed [9:0] m75_37;
   assign m75_37 =10'b0;

   // m75_38 = W*in
   wire signed [9:0] m75_38;
   assign m75_38 =10'b0;

   // m75_39 = W*in
   wire signed [9:0] m75_39;
   assign m75_39 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_40 = W*in
   wire signed [9:0] m75_40;
   assign m75_40 =10'b0;

   // m75_41 = W*in
   wire signed [9:0] m75_41;
   assign m75_41 =10'b0;

   // m75_42 = W*in
   wire signed [9:0] m75_42;
   assign m75_42 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_43 = W*in
   wire signed [9:0] m75_43;
   assign m75_43 =10'b0;

   // m75_44 = W*in
   wire signed [9:0] m75_44;
   assign m75_44 =10'b0;

   // m75_45 = W*in
   wire signed [9:0] m75_45;
   assign m75_45 =10'b0;

   // m75_46 = W*in
   wire signed [9:0] m75_46;
   assign m75_46 ={ {3{in75[5]}} , in75 , {1{1'b0}} };

   // m75_47 = W*in
   wire signed [9:0] m75_47;
   assign m75_47 =10'b0;

   // m75_48 = W*in
   wire signed [9:0] m75_48;
   assign m75_48 =10'b0;

   // m75_49 = W*in
   wire signed [9:0] m75_49;
   assign m75_49 =10'b0;

   // m75_50 = W*in
   wire signed [9:0] m75_50;
   assign m75_50 =10'b0;

   // m75_51 = W*in
   wire signed [9:0] m75_51;
   assign m75_51 =10'b0;

   // m75_52 = W*in
   wire signed [9:0] m75_52;
   assign m75_52 =10'b0;

   // m75_53 = W*in
   wire signed [9:0] m75_53;
   assign m75_53 =10'b0;

   // m75_54 = W*in
   wire signed [9:0] m75_54;
   assign m75_54 =10'b0;

   // m75_55 = W*in
   wire signed [9:0] m75_55;
   assign m75_55 =10'b0;

   // m75_56 = W*in
   wire signed [9:0] m75_56;
   assign m75_56 =10'b0;

   // m75_57 = W*in
   wire signed [9:0] m75_57;
   assign m75_57 =10'b0;

   // m75_58 = W*in
   wire signed [9:0] m75_58;
   assign m75_58 =10'b0;

   // m75_59 = W*in
   wire signed [9:0] m75_59;
   assign m75_59 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_60 = W*in
   wire signed [9:0] m75_60;
   assign m75_60 =10'b0;

   // m75_61 = W*in
   wire signed [9:0] m75_61;
   assign m75_61 =10'b0;

   // m75_62 = W*in
   wire signed [9:0] m75_62;
   assign m75_62 ={ {2{in75[5]}} , in75 , {2{1'b0}} };

   // m75_63 = W*in
   wire signed [9:0] m75_63;
   assign m75_63 =10'b0;

   // m75_64 = W*in
   wire signed [9:0] m75_64;
   assign m75_64 =10'b0;

   // m75_65 = W*in
   wire signed [9:0] m75_65;
   assign m75_65 =10'b0;

   // m75_66 = W*in
   wire signed [9:0] m75_66;
   assign m75_66 =10'b0;

   // m75_67 = W*in
   wire signed [9:0] m75_67;
   assign m75_67 =10'b0;

   // m75_68 = W*in
   wire signed [9:0] m75_68;
   assign m75_68 =10'b0;

   // m75_69 = W*in
   wire signed [9:0] m75_69;
   assign m75_69 =10'b0;

   // m75_70 = W*in
   wire signed [9:0] m75_70;
   assign m75_70 =10'b0;

   // m75_71 = W*in
   wire signed [9:0] m75_71;
   assign m75_71 =10'b0;

   // m75_72 = W*in
   wire signed [9:0] m75_72;
   assign m75_72 =10'b0;

   // m75_73 = W*in
   wire signed [9:0] m75_73;
   assign m75_73 =10'b0;

   // m75_74 = W*in
   wire signed [9:0] m75_74;
   assign m75_74 =10'b0;

   // m75_75 = W*in
   wire signed [9:0] m75_75;
   assign m75_75 =10'b0;

   // m75_76 = W*in
   wire signed [9:0] m75_76;
   assign m75_76 =10'b0;

   // m75_77 = W*in
   wire signed [9:0] m75_77;
   assign m75_77 ={ {3{neg75[5]}} , neg75 , {1{1'b0}} };

   // m75_78 = W*in
   wire signed [9:0] m75_78;
   assign m75_78 =10'b0;

   // m75_79 = W*in
   wire signed [9:0] m75_79;
   assign m75_79 =10'b0;

   // m75_80 = W*in
   wire signed [9:0] m75_80;
   assign m75_80 =10'b0;

   // m75_81 = W*in
   wire signed [9:0] m75_81;
   assign m75_81 =10'b0;

   // m76_1 = W*in
   wire signed [9:0] m76_1;
   assign m76_1 =10'b0;

   // m76_2 = W*in
   wire signed [9:0] m76_2;
   assign m76_2 =10'b0;

   // m76_3 = W*in
   wire signed [9:0] m76_3;
   assign m76_3 =10'b0;

   // m76_4 = W*in
   wire signed [9:0] m76_4;
   assign m76_4 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_5 = W*in
   wire signed [9:0] m76_5;
   assign m76_5 ={ {2{in76[5]}} , in76 , {2{1'b0}} };

   // m76_6 = W*in
   wire signed [9:0] m76_6;
   assign m76_6 =10'b0;

   // m76_7 = W*in
   wire signed [9:0] m76_7;
   assign m76_7 =10'b0;

   // m76_8 = W*in
   wire signed [9:0] m76_8;
   assign m76_8 =10'b0;

   // m76_9 = W*in
   wire signed [9:0] m76_9;
   assign m76_9 =10'b0;

   // m76_10 = W*in
   wire signed [9:0] m76_10;
   assign m76_10 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_11 = W*in
   wire signed [9:0] m76_11;
   assign m76_11 =10'b0;

   // m76_12 = W*in
   wire signed [9:0] m76_12;
   assign m76_12 =10'b0;

   // m76_13 = W*in
   wire signed [9:0] m76_13;
   assign m76_13 =10'b0;

   // m76_14 = W*in
   wire signed [9:0] m76_14;
   assign m76_14 =10'b0;

   // m76_15 = W*in
   wire signed [9:0] m76_15;
   assign m76_15 ={ {3{neg76[5]}} , neg76 , {1{1'b0}} };

   // m76_16 = W*in
   wire signed [9:0] m76_16;
   assign m76_16 =10'b0;

   // m76_17 = W*in
   wire signed [9:0] m76_17;
   assign m76_17 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_18 = W*in
   wire signed [9:0] m76_18;
   assign m76_18 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_19 = W*in
   wire signed [9:0] m76_19;
   assign m76_19 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_20 = W*in
   wire signed [9:0] m76_20;
   assign m76_20 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_21 = W*in
   wire signed [9:0] m76_21;
   assign m76_21 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_22 = W*in
   wire signed [9:0] m76_22;
   assign m76_22 ={ {2{in76[5]}} , in76 , {2{1'b0}} };

   // m76_23 = W*in
   wire signed [9:0] m76_23;
   assign m76_23 =10'b0;

   // m76_24 = W*in
   wire signed [9:0] m76_24;
   assign m76_24 ={ {2{in76[5]}} , in76 , {2{1'b0}} };

   // m76_25 = W*in
   wire signed [9:0] m76_25;
   assign m76_25 =10'b0;

   // m76_26 = W*in
   wire signed [9:0] m76_26;
   assign m76_26 =10'b0;

   // m76_27 = W*in
   wire signed [9:0] m76_27;
   assign m76_27 =10'b0;

   // m76_28 = W*in
   wire signed [9:0] m76_28;
   assign m76_28 ={ {2{in76[5]}} , in76 , {2{1'b0}} };

   // m76_29 = W*in
   wire signed [9:0] m76_29;
   assign m76_29 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_30 = W*in
   wire signed [9:0] m76_30;
   assign m76_30 ={ {3{neg76[5]}} , neg76 , {1{1'b0}} };

   // m76_31 = W*in
   wire signed [9:0] m76_31;
   assign m76_31 =10'b0;

   // m76_32 = W*in
   wire signed [9:0] m76_32;
   assign m76_32 =10'b0;

   // m76_33 = W*in
   wire signed [9:0] m76_33;
   assign m76_33 ={ {3{neg76[5]}} , neg76 , {1{1'b0}} };

   // m76_34 = W*in
   wire signed [9:0] m76_34;
   assign m76_34 =10'b0;

   // m76_35 = W*in
   wire signed [9:0] m76_35;
   assign m76_35 =10'b0;

   // m76_36 = W*in
   wire signed [9:0] m76_36;
   assign m76_36 =10'b0;

   // m76_37 = W*in
   wire signed [9:0] m76_37;
   assign m76_37 =10'b0;

   // m76_38 = W*in
   wire signed [9:0] m76_38;
   assign m76_38 =10'b0;

   // m76_39 = W*in
   wire signed [9:0] m76_39;
   assign m76_39 =10'b0;

   // m76_40 = W*in
   wire signed [9:0] m76_40;
   assign m76_40 =10'b0;

   // m76_41 = W*in
   wire signed [9:0] m76_41;
   assign m76_41 =10'b0;

   // m76_42 = W*in
   wire signed [9:0] m76_42;
   assign m76_42 =10'b0;

   // m76_43 = W*in
   wire signed [9:0] m76_43;
   assign m76_43 ={ {3{neg76[5]}} , neg76 , {1{1'b0}} };

   // m76_44 = W*in
   wire signed [9:0] m76_44;
   assign m76_44 ={ {3{neg76[5]}} , neg76 , {1{1'b0}} };

   // m76_45 = W*in
   wire signed [9:0] m76_45;
   assign m76_45 ={ {2{in76[5]}} , in76 , {2{1'b0}} };

   // m76_46 = W*in
   wire signed [9:0] m76_46;
   assign m76_46 =10'b0;

   // m76_47 = W*in
   wire signed [9:0] m76_47;
   assign m76_47 =10'b0;

   // m76_48 = W*in
   wire signed [9:0] m76_48;
   assign m76_48 ={ {2{in76[5]}} , in76 , {2{1'b0}} };

   // m76_49 = W*in
   wire signed [9:0] m76_49;
   assign m76_49 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_50 = W*in
   wire signed [9:0] m76_50;
   assign m76_50 =10'b0;

   // m76_51 = W*in
   wire signed [9:0] m76_51;
   assign m76_51 =10'b0;

   // m76_52 = W*in
   wire signed [9:0] m76_52;
   assign m76_52 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_53 = W*in
   wire signed [9:0] m76_53;
   assign m76_53 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_54 = W*in
   wire signed [9:0] m76_54;
   assign m76_54 =10'b0;

   // m76_55 = W*in
   wire signed [9:0] m76_55;
   assign m76_55 =10'b0;

   // m76_56 = W*in
   wire signed [9:0] m76_56;
   assign m76_56 =10'b0;

   // m76_57 = W*in
   wire signed [9:0] m76_57;
   assign m76_57 =10'b0;

   // m76_58 = W*in
   wire signed [9:0] m76_58;
   assign m76_58 =10'b0;

   // m76_59 = W*in
   wire signed [9:0] m76_59;
   assign m76_59 =10'b0;

   // m76_60 = W*in
   wire signed [9:0] m76_60;
   assign m76_60 =10'b0;

   // m76_61 = W*in
   wire signed [9:0] m76_61;
   assign m76_61 =10'b0;

   // m76_62 = W*in
   wire signed [9:0] m76_62;
   assign m76_62 ={ {3{neg76[5]}} , neg76 , {1{1'b0}} };

   // m76_63 = W*in
   wire signed [9:0] m76_63;
   assign m76_63 =10'b0;

   // m76_64 = W*in
   wire signed [9:0] m76_64;
   assign m76_64 =10'b0;

   // m76_65 = W*in
   wire signed [9:0] m76_65;
   assign m76_65 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_66 = W*in
   wire signed [9:0] m76_66;
   assign m76_66 =10'b0;

   // m76_67 = W*in
   wire signed [9:0] m76_67;
   assign m76_67 =10'b0;

   // m76_68 = W*in
   wire signed [9:0] m76_68;
   assign m76_68 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_69 = W*in
   wire signed [9:0] m76_69;
   assign m76_69 =10'b0;

   // m76_70 = W*in
   wire signed [9:0] m76_70;
   assign m76_70 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_71 = W*in
   wire signed [9:0] m76_71;
   assign m76_71 =10'b0;

   // m76_72 = W*in
   wire signed [9:0] m76_72;
   assign m76_72 =10'b0;

   // m76_73 = W*in
   wire signed [9:0] m76_73;
   assign m76_73 =10'b0;

   // m76_74 = W*in
   wire signed [9:0] m76_74;
   assign m76_74 =10'b0;

   // m76_75 = W*in
   wire signed [9:0] m76_75;
   assign m76_75 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_76 = W*in
   wire signed [9:0] m76_76;
   assign m76_76 =10'b0;

   // m76_77 = W*in
   wire signed [9:0] m76_77;
   assign m76_77 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_78 = W*in
   wire signed [9:0] m76_78;
   assign m76_78 ={ {3{in76[5]}} , in76 , {1{1'b0}} };

   // m76_79 = W*in
   wire signed [9:0] m76_79;
   assign m76_79 =10'b0;

   // m76_80 = W*in
   wire signed [9:0] m76_80;
   assign m76_80 =10'b0;

   // m76_81 = W*in
   wire signed [9:0] m76_81;
   assign m76_81 ={ {2{neg76[5]}} , neg76 , {2{1'b0}} };

   // m77_1 = W*in
   wire signed [9:0] m77_1;
   assign m77_1 =10'b0;

   // m77_2 = W*in
   wire signed [9:0] m77_2;
   assign m77_2 =10'b0;

   // m77_3 = W*in
   wire signed [9:0] m77_3;
   assign m77_3 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_4 = W*in
   wire signed [9:0] m77_4;
   assign m77_4 =10'b0;

   // m77_5 = W*in
   wire signed [9:0] m77_5;
   assign m77_5 ={ {2{in77[5]}} , in77 , {2{1'b0}} };

   // m77_6 = W*in
   wire signed [9:0] m77_6;
   assign m77_6 =10'b0;

   // m77_7 = W*in
   wire signed [9:0] m77_7;
   assign m77_7 =10'b0;

   // m77_8 = W*in
   wire signed [9:0] m77_8;
   assign m77_8 =10'b0;

   // m77_9 = W*in
   wire signed [9:0] m77_9;
   assign m77_9 =10'b0;

   // m77_10 = W*in
   wire signed [9:0] m77_10;
   assign m77_10 =10'b0;

   // m77_11 = W*in
   wire signed [9:0] m77_11;
   assign m77_11 =10'b0;

   // m77_12 = W*in
   wire signed [9:0] m77_12;
   assign m77_12 =10'b0;

   // m77_13 = W*in
   wire signed [9:0] m77_13;
   assign m77_13 =10'b0;

   // m77_14 = W*in
   wire signed [9:0] m77_14;
   assign m77_14 =10'b0;

   // m77_15 = W*in
   wire signed [9:0] m77_15;
   assign m77_15 =10'b0;

   // m77_16 = W*in
   wire signed [9:0] m77_16;
   assign m77_16 =10'b0;

   // m77_17 = W*in
   wire signed [9:0] m77_17;
   assign m77_17 =10'b0;

   // m77_18 = W*in
   wire signed [9:0] m77_18;
   assign m77_18 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_19 = W*in
   wire signed [9:0] m77_19;
   assign m77_19 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_20 = W*in
   wire signed [9:0] m77_20;
   assign m77_20 =10'b0;

   // m77_21 = W*in
   wire signed [9:0] m77_21;
   assign m77_21 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_22 = W*in
   wire signed [9:0] m77_22;
   assign m77_22 =10'b0;

   // m77_23 = W*in
   wire signed [9:0] m77_23;
   assign m77_23 =10'b0;

   // m77_24 = W*in
   wire signed [9:0] m77_24;
   assign m77_24 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_25 = W*in
   wire signed [9:0] m77_25;
   assign m77_25 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_26 = W*in
   wire signed [9:0] m77_26;
   assign m77_26 =10'b0;

   // m77_27 = W*in
   wire signed [9:0] m77_27;
   assign m77_27 =10'b0;

   // m77_28 = W*in
   wire signed [9:0] m77_28;
   assign m77_28 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_29 = W*in
   wire signed [9:0] m77_29;
   assign m77_29 =10'b0;

   // m77_30 = W*in
   wire signed [9:0] m77_30;
   assign m77_30 =10'b0;

   // m77_31 = W*in
   wire signed [9:0] m77_31;
   assign m77_31 =10'b0;

   // m77_32 = W*in
   wire signed [9:0] m77_32;
   assign m77_32 =10'b0;

   // m77_33 = W*in
   wire signed [9:0] m77_33;
   assign m77_33 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_34 = W*in
   wire signed [9:0] m77_34;
   assign m77_34 =10'b0;

   // m77_35 = W*in
   wire signed [9:0] m77_35;
   assign m77_35 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_36 = W*in
   wire signed [9:0] m77_36;
   assign m77_36 =10'b0;

   // m77_37 = W*in
   wire signed [9:0] m77_37;
   assign m77_37 =10'b0;

   // m77_38 = W*in
   wire signed [9:0] m77_38;
   assign m77_38 =10'b0;

   // m77_39 = W*in
   wire signed [9:0] m77_39;
   assign m77_39 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_40 = W*in
   wire signed [9:0] m77_40;
   assign m77_40 =10'b0;

   // m77_41 = W*in
   wire signed [9:0] m77_41;
   assign m77_41 =10'b0;

   // m77_42 = W*in
   wire signed [9:0] m77_42;
   assign m77_42 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_43 = W*in
   wire signed [9:0] m77_43;
   assign m77_43 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_44 = W*in
   wire signed [9:0] m77_44;
   assign m77_44 =10'b0;

   // m77_45 = W*in
   wire signed [9:0] m77_45;
   assign m77_45 =10'b0;

   // m77_46 = W*in
   wire signed [9:0] m77_46;
   assign m77_46 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_47 = W*in
   wire signed [9:0] m77_47;
   assign m77_47 =10'b0;

   // m77_48 = W*in
   wire signed [9:0] m77_48;
   assign m77_48 =10'b0;

   // m77_49 = W*in
   wire signed [9:0] m77_49;
   assign m77_49 =10'b0;

   // m77_50 = W*in
   wire signed [9:0] m77_50;
   assign m77_50 =10'b0;

   // m77_51 = W*in
   wire signed [9:0] m77_51;
   assign m77_51 =10'b0;

   // m77_52 = W*in
   wire signed [9:0] m77_52;
   assign m77_52 =10'b0;

   // m77_53 = W*in
   wire signed [9:0] m77_53;
   assign m77_53 =10'b0;

   // m77_54 = W*in
   wire signed [9:0] m77_54;
   assign m77_54 =10'b0;

   // m77_55 = W*in
   wire signed [9:0] m77_55;
   assign m77_55 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_56 = W*in
   wire signed [9:0] m77_56;
   assign m77_56 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_57 = W*in
   wire signed [9:0] m77_57;
   assign m77_57 =10'b0;

   // m77_58 = W*in
   wire signed [9:0] m77_58;
   assign m77_58 ={ {2{in77[5]}} , in77 , {2{1'b0}} };

   // m77_59 = W*in
   wire signed [9:0] m77_59;
   assign m77_59 =10'b0;

   // m77_60 = W*in
   wire signed [9:0] m77_60;
   assign m77_60 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_61 = W*in
   wire signed [9:0] m77_61;
   assign m77_61 =10'b0;

   // m77_62 = W*in
   wire signed [9:0] m77_62;
   assign m77_62 =10'b0;

   // m77_63 = W*in
   wire signed [9:0] m77_63;
   assign m77_63 =10'b0;

   // m77_64 = W*in
   wire signed [9:0] m77_64;
   assign m77_64 =10'b0;

   // m77_65 = W*in
   wire signed [9:0] m77_65;
   assign m77_65 =10'b0;

   // m77_66 = W*in
   wire signed [9:0] m77_66;
   assign m77_66 =10'b0;

   // m77_67 = W*in
   wire signed [9:0] m77_67;
   assign m77_67 =10'b0;

   // m77_68 = W*in
   wire signed [9:0] m77_68;
   assign m77_68 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_69 = W*in
   wire signed [9:0] m77_69;
   assign m77_69 =10'b0;

   // m77_70 = W*in
   wire signed [9:0] m77_70;
   assign m77_70 =10'b0;

   // m77_71 = W*in
   wire signed [9:0] m77_71;
   assign m77_71 =10'b0;

   // m77_72 = W*in
   wire signed [9:0] m77_72;
   assign m77_72 =10'b0;

   // m77_73 = W*in
   wire signed [9:0] m77_73;
   assign m77_73 =10'b0;

   // m77_74 = W*in
   wire signed [9:0] m77_74;
   assign m77_74 =10'b0;

   // m77_75 = W*in
   wire signed [9:0] m77_75;
   assign m77_75 =10'b0;

   // m77_76 = W*in
   wire signed [9:0] m77_76;
   assign m77_76 =10'b0;

   // m77_77 = W*in
   wire signed [9:0] m77_77;
   assign m77_77 =10'b0;

   // m77_78 = W*in
   wire signed [9:0] m77_78;
   assign m77_78 ={ {3{neg77[5]}} , neg77 , {1{1'b0}} };

   // m77_79 = W*in
   wire signed [9:0] m77_79;
   assign m77_79 =10'b0;

   // m77_80 = W*in
   wire signed [9:0] m77_80;
   assign m77_80 ={ {2{in77[5]}} , in77 , {2{1'b0}} };

   // m77_81 = W*in
   wire signed [9:0] m77_81;
   assign m77_81 =10'b0;

   // m78_1 = W*in
   wire signed [9:0] m78_1;
   assign m78_1 =10'b0;

   // m78_2 = W*in
   wire signed [9:0] m78_2;
   assign m78_2 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_3 = W*in
   wire signed [9:0] m78_3;
   assign m78_3 =10'b0;

   // m78_4 = W*in
   wire signed [9:0] m78_4;
   assign m78_4 =10'b0;

   // m78_5 = W*in
   wire signed [9:0] m78_5;
   assign m78_5 =10'b0;

   // m78_6 = W*in
   wire signed [9:0] m78_6;
   assign m78_6 =10'b0;

   // m78_7 = W*in
   wire signed [9:0] m78_7;
   assign m78_7 =10'b0;

   // m78_8 = W*in
   wire signed [9:0] m78_8;
   assign m78_8 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_9 = W*in
   wire signed [9:0] m78_9;
   assign m78_9 =10'b0;

   // m78_10 = W*in
   wire signed [9:0] m78_10;
   assign m78_10 =10'b0;

   // m78_11 = W*in
   wire signed [9:0] m78_11;
   assign m78_11 =10'b0;

   // m78_12 = W*in
   wire signed [9:0] m78_12;
   assign m78_12 =10'b0;

   // m78_13 = W*in
   wire signed [9:0] m78_13;
   assign m78_13 =10'b0;

   // m78_14 = W*in
   wire signed [9:0] m78_14;
   assign m78_14 =10'b0;

   // m78_15 = W*in
   wire signed [9:0] m78_15;
   assign m78_15 =10'b0;

   // m78_16 = W*in
   wire signed [9:0] m78_16;
   assign m78_16 =10'b0;

   // m78_17 = W*in
   wire signed [9:0] m78_17;
   assign m78_17 =10'b0;

   // m78_18 = W*in
   wire signed [9:0] m78_18;
   assign m78_18 =10'b0;

   // m78_19 = W*in
   wire signed [9:0] m78_19;
   assign m78_19 =10'b0;

   // m78_20 = W*in
   wire signed [9:0] m78_20;
   assign m78_20 =10'b0;

   // m78_21 = W*in
   wire signed [9:0] m78_21;
   assign m78_21 =10'b0;

   // m78_22 = W*in
   wire signed [9:0] m78_22;
   assign m78_22 =10'b0;

   // m78_23 = W*in
   wire signed [9:0] m78_23;
   assign m78_23 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_24 = W*in
   wire signed [9:0] m78_24;
   assign m78_24 =10'b0;

   // m78_25 = W*in
   wire signed [9:0] m78_25;
   assign m78_25 ={ {3{in78[5]}} , in78 , {1{1'b0}} };

   // m78_26 = W*in
   wire signed [9:0] m78_26;
   assign m78_26 =10'b0;

   // m78_27 = W*in
   wire signed [9:0] m78_27;
   assign m78_27 =10'b0;

   // m78_28 = W*in
   wire signed [9:0] m78_28;
   assign m78_28 =10'b0;

   // m78_29 = W*in
   wire signed [9:0] m78_29;
   assign m78_29 =10'b0;

   // m78_30 = W*in
   wire signed [9:0] m78_30;
   assign m78_30 =10'b0;

   // m78_31 = W*in
   wire signed [9:0] m78_31;
   assign m78_31 =10'b0;

   // m78_32 = W*in
   wire signed [9:0] m78_32;
   assign m78_32 =10'b0;

   // m78_33 = W*in
   wire signed [9:0] m78_33;
   assign m78_33 =10'b0;

   // m78_34 = W*in
   wire signed [9:0] m78_34;
   assign m78_34 =10'b0;

   // m78_35 = W*in
   wire signed [9:0] m78_35;
   assign m78_35 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_36 = W*in
   wire signed [9:0] m78_36;
   assign m78_36 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_37 = W*in
   wire signed [9:0] m78_37;
   assign m78_37 =10'b0;

   // m78_38 = W*in
   wire signed [9:0] m78_38;
   assign m78_38 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_39 = W*in
   wire signed [9:0] m78_39;
   assign m78_39 ={ {3{in78[5]}} , in78 , {1{1'b0}} };

   // m78_40 = W*in
   wire signed [9:0] m78_40;
   assign m78_40 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_41 = W*in
   wire signed [9:0] m78_41;
   assign m78_41 =10'b0;

   // m78_42 = W*in
   wire signed [9:0] m78_42;
   assign m78_42 ={ {3{in78[5]}} , in78 , {1{1'b0}} };

   // m78_43 = W*in
   wire signed [9:0] m78_43;
   assign m78_43 =10'b0;

   // m78_44 = W*in
   wire signed [9:0] m78_44;
   assign m78_44 =10'b0;

   // m78_45 = W*in
   wire signed [9:0] m78_45;
   assign m78_45 =10'b0;

   // m78_46 = W*in
   wire signed [9:0] m78_46;
   assign m78_46 =10'b0;

   // m78_47 = W*in
   wire signed [9:0] m78_47;
   assign m78_47 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_48 = W*in
   wire signed [9:0] m78_48;
   assign m78_48 =10'b0;

   // m78_49 = W*in
   wire signed [9:0] m78_49;
   assign m78_49 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_50 = W*in
   wire signed [9:0] m78_50;
   assign m78_50 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_51 = W*in
   wire signed [9:0] m78_51;
   assign m78_51 =10'b0;

   // m78_52 = W*in
   wire signed [9:0] m78_52;
   assign m78_52 =10'b0;

   // m78_53 = W*in
   wire signed [9:0] m78_53;
   assign m78_53 =10'b0;

   // m78_54 = W*in
   wire signed [9:0] m78_54;
   assign m78_54 =10'b0;

   // m78_55 = W*in
   wire signed [9:0] m78_55;
   assign m78_55 =10'b0;

   // m78_56 = W*in
   wire signed [9:0] m78_56;
   assign m78_56 =10'b0;

   // m78_57 = W*in
   wire signed [9:0] m78_57;
   assign m78_57 =10'b0;

   // m78_58 = W*in
   wire signed [9:0] m78_58;
   assign m78_58 =10'b0;

   // m78_59 = W*in
   wire signed [9:0] m78_59;
   assign m78_59 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_60 = W*in
   wire signed [9:0] m78_60;
   assign m78_60 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_61 = W*in
   wire signed [9:0] m78_61;
   assign m78_61 =10'b0;

   // m78_62 = W*in
   wire signed [9:0] m78_62;
   assign m78_62 =10'b0;

   // m78_63 = W*in
   wire signed [9:0] m78_63;
   assign m78_63 =10'b0;

   // m78_64 = W*in
   wire signed [9:0] m78_64;
   assign m78_64 =10'b0;

   // m78_65 = W*in
   wire signed [9:0] m78_65;
   assign m78_65 =10'b0;

   // m78_66 = W*in
   wire signed [9:0] m78_66;
   assign m78_66 =10'b0;

   // m78_67 = W*in
   wire signed [9:0] m78_67;
   assign m78_67 =10'b0;

   // m78_68 = W*in
   wire signed [9:0] m78_68;
   assign m78_68 =10'b0;

   // m78_69 = W*in
   wire signed [9:0] m78_69;
   assign m78_69 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_70 = W*in
   wire signed [9:0] m78_70;
   assign m78_70 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_71 = W*in
   wire signed [9:0] m78_71;
   assign m78_71 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_72 = W*in
   wire signed [9:0] m78_72;
   assign m78_72 =10'b0;

   // m78_73 = W*in
   wire signed [9:0] m78_73;
   assign m78_73 ={ {2{in78[5]}} , in78 , {2{1'b0}} };

   // m78_74 = W*in
   wire signed [9:0] m78_74;
   assign m78_74 =10'b0;

   // m78_75 = W*in
   wire signed [9:0] m78_75;
   assign m78_75 =10'b0;

   // m78_76 = W*in
   wire signed [9:0] m78_76;
   assign m78_76 =10'b0;

   // m78_77 = W*in
   wire signed [9:0] m78_77;
   assign m78_77 =10'b0;

   // m78_78 = W*in
   wire signed [9:0] m78_78;
   assign m78_78 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_79 = W*in
   wire signed [9:0] m78_79;
   assign m78_79 ={ {3{neg78[5]}} , neg78 , {1{1'b0}} };

   // m78_80 = W*in
   wire signed [9:0] m78_80;
   assign m78_80 =10'b0;

   // m78_81 = W*in
   wire signed [9:0] m78_81;
   assign m78_81 =10'b0;

   // m79_1 = W*in
   wire signed [9:0] m79_1;
   assign m79_1 =10'b0;

   // m79_2 = W*in
   wire signed [9:0] m79_2;
   assign m79_2 =10'b0;

   // m79_3 = W*in
   wire signed [9:0] m79_3;
   assign m79_3 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_4 = W*in
   wire signed [9:0] m79_4;
   assign m79_4 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_5 = W*in
   wire signed [9:0] m79_5;
   assign m79_5 =10'b0;

   // m79_6 = W*in
   wire signed [9:0] m79_6;
   assign m79_6 =10'b0;

   // m79_7 = W*in
   wire signed [9:0] m79_7;
   assign m79_7 =10'b0;

   // m79_8 = W*in
   wire signed [9:0] m79_8;
   assign m79_8 =10'b0;

   // m79_9 = W*in
   wire signed [9:0] m79_9;
   assign m79_9 =10'b0;

   // m79_10 = W*in
   wire signed [9:0] m79_10;
   assign m79_10 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_11 = W*in
   wire signed [9:0] m79_11;
   assign m79_11 =10'b0;

   // m79_12 = W*in
   wire signed [9:0] m79_12;
   assign m79_12 =10'b0;

   // m79_13 = W*in
   wire signed [9:0] m79_13;
   assign m79_13 =10'b0;

   // m79_14 = W*in
   wire signed [9:0] m79_14;
   assign m79_14 =10'b0;

   // m79_15 = W*in
   wire signed [9:0] m79_15;
   assign m79_15 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_16 = W*in
   wire signed [9:0] m79_16;
   assign m79_16 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_17 = W*in
   wire signed [9:0] m79_17;
   assign m79_17 =10'b0;

   // m79_18 = W*in
   wire signed [9:0] m79_18;
   assign m79_18 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_19 = W*in
   wire signed [9:0] m79_19;
   assign m79_19 =10'b0;

   // m79_20 = W*in
   wire signed [9:0] m79_20;
   assign m79_20 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_21 = W*in
   wire signed [9:0] m79_21;
   assign m79_21 =10'b0;

   // m79_22 = W*in
   wire signed [9:0] m79_22;
   assign m79_22 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_23 = W*in
   wire signed [9:0] m79_23;
   assign m79_23 ={ {3{neg79[5]}} , neg79 , {1{1'b0}} };

   // m79_24 = W*in
   wire signed [9:0] m79_24;
   assign m79_24 =10'b0;

   // m79_25 = W*in
   wire signed [9:0] m79_25;
   assign m79_25 ={ {3{neg79[5]}} , neg79 , {1{1'b0}} };

   // m79_26 = W*in
   wire signed [9:0] m79_26;
   assign m79_26 =10'b0;

   // m79_27 = W*in
   wire signed [9:0] m79_27;
   assign m79_27 =10'b0;

   // m79_28 = W*in
   wire signed [9:0] m79_28;
   assign m79_28 =10'b0;

   // m79_29 = W*in
   wire signed [9:0] m79_29;
   assign m79_29 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_30 = W*in
   wire signed [9:0] m79_30;
   assign m79_30 =10'b0;

   // m79_31 = W*in
   wire signed [9:0] m79_31;
   assign m79_31 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_32 = W*in
   wire signed [9:0] m79_32;
   assign m79_32 =10'b0;

   // m79_33 = W*in
   wire signed [9:0] m79_33;
   assign m79_33 ={ {3{neg79[5]}} , neg79 , {1{1'b0}} };

   // m79_34 = W*in
   wire signed [9:0] m79_34;
   assign m79_34 =10'b0;

   // m79_35 = W*in
   wire signed [9:0] m79_35;
   assign m79_35 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_36 = W*in
   wire signed [9:0] m79_36;
   assign m79_36 =10'b0;

   // m79_37 = W*in
   wire signed [9:0] m79_37;
   assign m79_37 ={ {3{neg79[5]}} , neg79 , {1{1'b0}} };

   // m79_38 = W*in
   wire signed [9:0] m79_38;
   assign m79_38 =10'b0;

   // m79_39 = W*in
   wire signed [9:0] m79_39;
   assign m79_39 =10'b0;

   // m79_40 = W*in
   wire signed [9:0] m79_40;
   assign m79_40 =10'b0;

   // m79_41 = W*in
   wire signed [9:0] m79_41;
   assign m79_41 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_42 = W*in
   wire signed [9:0] m79_42;
   assign m79_42 =10'b0;

   // m79_43 = W*in
   wire signed [9:0] m79_43;
   assign m79_43 ={ {3{neg79[5]}} , neg79 , {1{1'b0}} };

   // m79_44 = W*in
   wire signed [9:0] m79_44;
   assign m79_44 =10'b0;

   // m79_45 = W*in
   wire signed [9:0] m79_45;
   assign m79_45 =10'b0;

   // m79_46 = W*in
   wire signed [9:0] m79_46;
   assign m79_46 =10'b0;

   // m79_47 = W*in
   wire signed [9:0] m79_47;
   assign m79_47 =10'b0;

   // m79_48 = W*in
   wire signed [9:0] m79_48;
   assign m79_48 =10'b0;

   // m79_49 = W*in
   wire signed [9:0] m79_49;
   assign m79_49 =10'b0;

   // m79_50 = W*in
   wire signed [9:0] m79_50;
   assign m79_50 =10'b0;

   // m79_51 = W*in
   wire signed [9:0] m79_51;
   assign m79_51 =10'b0;

   // m79_52 = W*in
   wire signed [9:0] m79_52;
   assign m79_52 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_53 = W*in
   wire signed [9:0] m79_53;
   assign m79_53 =10'b0;

   // m79_54 = W*in
   wire signed [9:0] m79_54;
   assign m79_54 =10'b0;

   // m79_55 = W*in
   wire signed [9:0] m79_55;
   assign m79_55 =10'b0;

   // m79_56 = W*in
   wire signed [9:0] m79_56;
   assign m79_56 =10'b0;

   // m79_57 = W*in
   wire signed [9:0] m79_57;
   assign m79_57 =10'b0;

   // m79_58 = W*in
   wire signed [9:0] m79_58;
   assign m79_58 =10'b0;

   // m79_59 = W*in
   wire signed [9:0] m79_59;
   assign m79_59 =10'b0;

   // m79_60 = W*in
   wire signed [9:0] m79_60;
   assign m79_60 =10'b0;

   // m79_61 = W*in
   wire signed [9:0] m79_61;
   assign m79_61 ={ {2{in79[5]}} , in79 , {2{1'b0}} };

   // m79_62 = W*in
   wire signed [9:0] m79_62;
   assign m79_62 =10'b0;

   // m79_63 = W*in
   wire signed [9:0] m79_63;
   assign m79_63 =10'b0;

   // m79_64 = W*in
   wire signed [9:0] m79_64;
   assign m79_64 =10'b0;

   // m79_65 = W*in
   wire signed [9:0] m79_65;
   assign m79_65 =10'b0;

   // m79_66 = W*in
   wire signed [9:0] m79_66;
   assign m79_66 =10'b0;

   // m79_67 = W*in
   wire signed [9:0] m79_67;
   assign m79_67 =10'b0;

   // m79_68 = W*in
   wire signed [9:0] m79_68;
   assign m79_68 =10'b0;

   // m79_69 = W*in
   wire signed [9:0] m79_69;
   assign m79_69 =10'b0;

   // m79_70 = W*in
   wire signed [9:0] m79_70;
   assign m79_70 =10'b0;

   // m79_71 = W*in
   wire signed [9:0] m79_71;
   assign m79_71 =10'b0;

   // m79_72 = W*in
   wire signed [9:0] m79_72;
   assign m79_72 =10'b0;

   // m79_73 = W*in
   wire signed [9:0] m79_73;
   assign m79_73 =10'b0;

   // m79_74 = W*in
   wire signed [9:0] m79_74;
   assign m79_74 =10'b0;

   // m79_75 = W*in
   wire signed [9:0] m79_75;
   assign m79_75 =10'b0;

   // m79_76 = W*in
   wire signed [9:0] m79_76;
   assign m79_76 =10'b0;

   // m79_77 = W*in
   wire signed [9:0] m79_77;
   assign m79_77 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_78 = W*in
   wire signed [9:0] m79_78;
   assign m79_78 =10'b0;

   // m79_79 = W*in
   wire signed [9:0] m79_79;
   assign m79_79 ={ {3{in79[5]}} , in79 , {1{1'b0}} };

   // m79_80 = W*in
   wire signed [9:0] m79_80;
   assign m79_80 =10'b0;

   // m79_81 = W*in
   wire signed [9:0] m79_81;
   assign m79_81 =10'b0;

   // m80_1 = W*in
   wire signed [9:0] m80_1;
   assign m80_1 =10'b0;

   // m80_2 = W*in
   wire signed [9:0] m80_2;
   assign m80_2 =10'b0;

   // m80_3 = W*in
   wire signed [9:0] m80_3;
   assign m80_3 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_4 = W*in
   wire signed [9:0] m80_4;
   assign m80_4 =10'b0;

   // m80_5 = W*in
   wire signed [9:0] m80_5;
   assign m80_5 =10'b0;

   // m80_6 = W*in
   wire signed [9:0] m80_6;
   assign m80_6 =10'b0;

   // m80_7 = W*in
   wire signed [9:0] m80_7;
   assign m80_7 =10'b0;

   // m80_8 = W*in
   wire signed [9:0] m80_8;
   assign m80_8 =10'b0;

   // m80_9 = W*in
   wire signed [9:0] m80_9;
   assign m80_9 =10'b0;

   // m80_10 = W*in
   wire signed [9:0] m80_10;
   assign m80_10 =10'b0;

   // m80_11 = W*in
   wire signed [9:0] m80_11;
   assign m80_11 =10'b0;

   // m80_12 = W*in
   wire signed [9:0] m80_12;
   assign m80_12 =10'b0;

   // m80_13 = W*in
   wire signed [9:0] m80_13;
   assign m80_13 =10'b0;

   // m80_14 = W*in
   wire signed [9:0] m80_14;
   assign m80_14 =10'b0;

   // m80_15 = W*in
   wire signed [9:0] m80_15;
   assign m80_15 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_16 = W*in
   wire signed [9:0] m80_16;
   assign m80_16 =10'b0;

   // m80_17 = W*in
   wire signed [9:0] m80_17;
   assign m80_17 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_18 = W*in
   wire signed [9:0] m80_18;
   assign m80_18 =10'b0;

   // m80_19 = W*in
   wire signed [9:0] m80_19;
   assign m80_19 =10'b0;

   // m80_20 = W*in
   wire signed [9:0] m80_20;
   assign m80_20 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_21 = W*in
   wire signed [9:0] m80_21;
   assign m80_21 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_22 = W*in
   wire signed [9:0] m80_22;
   assign m80_22 =10'b0;

   // m80_23 = W*in
   wire signed [9:0] m80_23;
   assign m80_23 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_24 = W*in
   wire signed [9:0] m80_24;
   assign m80_24 =10'b0;

   // m80_25 = W*in
   wire signed [9:0] m80_25;
   assign m80_25 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_26 = W*in
   wire signed [9:0] m80_26;
   assign m80_26 =10'b0;

   // m80_27 = W*in
   wire signed [9:0] m80_27;
   assign m80_27 =10'b0;

   // m80_28 = W*in
   wire signed [9:0] m80_28;
   assign m80_28 =10'b0;

   // m80_29 = W*in
   wire signed [9:0] m80_29;
   assign m80_29 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_30 = W*in
   wire signed [9:0] m80_30;
   assign m80_30 =10'b0;

   // m80_31 = W*in
   wire signed [9:0] m80_31;
   assign m80_31 =10'b0;

   // m80_32 = W*in
   wire signed [9:0] m80_32;
   assign m80_32 =10'b0;

   // m80_33 = W*in
   wire signed [9:0] m80_33;
   assign m80_33 =10'b0;

   // m80_34 = W*in
   wire signed [9:0] m80_34;
   assign m80_34 =10'b0;

   // m80_35 = W*in
   wire signed [9:0] m80_35;
   assign m80_35 =10'b0;

   // m80_36 = W*in
   wire signed [9:0] m80_36;
   assign m80_36 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_37 = W*in
   wire signed [9:0] m80_37;
   assign m80_37 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_38 = W*in
   wire signed [9:0] m80_38;
   assign m80_38 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_39 = W*in
   wire signed [9:0] m80_39;
   assign m80_39 =10'b0;

   // m80_40 = W*in
   wire signed [9:0] m80_40;
   assign m80_40 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_41 = W*in
   wire signed [9:0] m80_41;
   assign m80_41 =10'b0;

   // m80_42 = W*in
   wire signed [9:0] m80_42;
   assign m80_42 ={ {3{neg80[5]}} , neg80 , {1{1'b0}} };

   // m80_43 = W*in
   wire signed [9:0] m80_43;
   assign m80_43 =10'b0;

   // m80_44 = W*in
   wire signed [9:0] m80_44;
   assign m80_44 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_45 = W*in
   wire signed [9:0] m80_45;
   assign m80_45 =10'b0;

   // m80_46 = W*in
   wire signed [9:0] m80_46;
   assign m80_46 =10'b0;

   // m80_47 = W*in
   wire signed [9:0] m80_47;
   assign m80_47 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_48 = W*in
   wire signed [9:0] m80_48;
   assign m80_48 =10'b0;

   // m80_49 = W*in
   wire signed [9:0] m80_49;
   assign m80_49 =10'b0;

   // m80_50 = W*in
   wire signed [9:0] m80_50;
   assign m80_50 =10'b0;

   // m80_51 = W*in
   wire signed [9:0] m80_51;
   assign m80_51 ={ {2{in80[5]}} , in80 , {2{1'b0}} };

   // m80_52 = W*in
   wire signed [9:0] m80_52;
   assign m80_52 =10'b0;

   // m80_53 = W*in
   wire signed [9:0] m80_53;
   assign m80_53 =10'b0;

   // m80_54 = W*in
   wire signed [9:0] m80_54;
   assign m80_54 =10'b0;

   // m80_55 = W*in
   wire signed [9:0] m80_55;
   assign m80_55 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_56 = W*in
   wire signed [9:0] m80_56;
   assign m80_56 =10'b0;

   // m80_57 = W*in
   wire signed [9:0] m80_57;
   assign m80_57 =10'b0;

   // m80_58 = W*in
   wire signed [9:0] m80_58;
   assign m80_58 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_59 = W*in
   wire signed [9:0] m80_59;
   assign m80_59 ={ {2{in80[5]}} , in80 , {2{1'b0}} };

   // m80_60 = W*in
   wire signed [9:0] m80_60;
   assign m80_60 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_61 = W*in
   wire signed [9:0] m80_61;
   assign m80_61 =10'b0;

   // m80_62 = W*in
   wire signed [9:0] m80_62;
   assign m80_62 =10'b0;

   // m80_63 = W*in
   wire signed [9:0] m80_63;
   assign m80_63 =10'b0;

   // m80_64 = W*in
   wire signed [9:0] m80_64;
   assign m80_64 =10'b0;

   // m80_65 = W*in
   wire signed [9:0] m80_65;
   assign m80_65 =10'b0;

   // m80_66 = W*in
   wire signed [9:0] m80_66;
   assign m80_66 =10'b0;

   // m80_67 = W*in
   wire signed [9:0] m80_67;
   assign m80_67 =10'b0;

   // m80_68 = W*in
   wire signed [9:0] m80_68;
   assign m80_68 =10'b0;

   // m80_69 = W*in
   wire signed [9:0] m80_69;
   assign m80_69 ={ {2{in80[5]}} , in80 , {2{1'b0}} };

   // m80_70 = W*in
   wire signed [9:0] m80_70;
   assign m80_70 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_71 = W*in
   wire signed [9:0] m80_71;
   assign m80_71 =10'b0;

   // m80_72 = W*in
   wire signed [9:0] m80_72;
   assign m80_72 =10'b0;

   // m80_73 = W*in
   wire signed [9:0] m80_73;
   assign m80_73 =10'b0;

   // m80_74 = W*in
   wire signed [9:0] m80_74;
   assign m80_74 =10'b0;

   // m80_75 = W*in
   wire signed [9:0] m80_75;
   assign m80_75 =10'b0;

   // m80_76 = W*in
   wire signed [9:0] m80_76;
   assign m80_76 =10'b0;

   // m80_77 = W*in
   wire signed [9:0] m80_77;
   assign m80_77 =10'b0;

   // m80_78 = W*in
   wire signed [9:0] m80_78;
   assign m80_78 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_79 = W*in
   wire signed [9:0] m80_79;
   assign m80_79 ={ {3{in80[5]}} , in80 , {1{1'b0}} };

   // m80_80 = W*in
   wire signed [9:0] m80_80;
   assign m80_80 =10'b0;

   // m80_81 = W*in
   wire signed [9:0] m80_81;
   assign m80_81 =10'b0;

   // m81_1 = W*in
   wire signed [9:0] m81_1;
   assign m81_1 ={ {2{in81[5]}} , in81 , {2{1'b0}} };

   // m81_2 = W*in
   wire signed [9:0] m81_2;
   assign m81_2 =10'b0;

   // m81_3 = W*in
   wire signed [9:0] m81_3;
   assign m81_3 =10'b0;

   // m81_4 = W*in
   wire signed [9:0] m81_4;
   assign m81_4 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_5 = W*in
   wire signed [9:0] m81_5;
   assign m81_5 =10'b0;

   // m81_6 = W*in
   wire signed [9:0] m81_6;
   assign m81_6 =10'b0;

   // m81_7 = W*in
   wire signed [9:0] m81_7;
   assign m81_7 =10'b0;

   // m81_8 = W*in
   wire signed [9:0] m81_8;
   assign m81_8 =10'b0;

   // m81_9 = W*in
   wire signed [9:0] m81_9;
   assign m81_9 =10'b0;

   // m81_10 = W*in
   wire signed [9:0] m81_10;
   assign m81_10 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_11 = W*in
   wire signed [9:0] m81_11;
   assign m81_11 =10'b0;

   // m81_12 = W*in
   wire signed [9:0] m81_12;
   assign m81_12 =10'b0;

   // m81_13 = W*in
   wire signed [9:0] m81_13;
   assign m81_13 ={ {2{in81[5]}} , in81 , {2{1'b0}} };

   // m81_14 = W*in
   wire signed [9:0] m81_14;
   assign m81_14 =10'b0;

   // m81_15 = W*in
   wire signed [9:0] m81_15;
   assign m81_15 =10'b0;

   // m81_16 = W*in
   wire signed [9:0] m81_16;
   assign m81_16 =10'b0;

   // m81_17 = W*in
   wire signed [9:0] m81_17;
   assign m81_17 =10'b0;

   // m81_18 = W*in
   wire signed [9:0] m81_18;
   assign m81_18 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_19 = W*in
   wire signed [9:0] m81_19;
   assign m81_19 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_20 = W*in
   wire signed [9:0] m81_20;
   assign m81_20 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_21 = W*in
   wire signed [9:0] m81_21;
   assign m81_21 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_22 = W*in
   wire signed [9:0] m81_22;
   assign m81_22 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_23 = W*in
   wire signed [9:0] m81_23;
   assign m81_23 =10'b0;

   // m81_24 = W*in
   wire signed [9:0] m81_24;
   assign m81_24 =10'b0;

   // m81_25 = W*in
   wire signed [9:0] m81_25;
   assign m81_25 =10'b0;

   // m81_26 = W*in
   wire signed [9:0] m81_26;
   assign m81_26 =10'b0;

   // m81_27 = W*in
   wire signed [9:0] m81_27;
   assign m81_27 ={ {2{in81[5]}} , in81 , {2{1'b0}} };

   // m81_28 = W*in
   wire signed [9:0] m81_28;
   assign m81_28 =10'b0;

   // m81_29 = W*in
   wire signed [9:0] m81_29;
   assign m81_29 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_30 = W*in
   wire signed [9:0] m81_30;
   assign m81_30 =10'b0;

   // m81_31 = W*in
   wire signed [9:0] m81_31;
   assign m81_31 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_32 = W*in
   wire signed [9:0] m81_32;
   assign m81_32 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_33 = W*in
   wire signed [9:0] m81_33;
   assign m81_33 =10'b0;

   // m81_34 = W*in
   wire signed [9:0] m81_34;
   assign m81_34 =10'b0;

   // m81_35 = W*in
   wire signed [9:0] m81_35;
   assign m81_35 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_36 = W*in
   wire signed [9:0] m81_36;
   assign m81_36 =10'b0;

   // m81_37 = W*in
   wire signed [9:0] m81_37;
   assign m81_37 =10'b0;

   // m81_38 = W*in
   wire signed [9:0] m81_38;
   assign m81_38 =10'b0;

   // m81_39 = W*in
   wire signed [9:0] m81_39;
   assign m81_39 =10'b0;

   // m81_40 = W*in
   wire signed [9:0] m81_40;
   assign m81_40 =10'b0;

   // m81_41 = W*in
   wire signed [9:0] m81_41;
   assign m81_41 =10'b0;

   // m81_42 = W*in
   wire signed [9:0] m81_42;
   assign m81_42 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_43 = W*in
   wire signed [9:0] m81_43;
   assign m81_43 =10'b0;

   // m81_44 = W*in
   wire signed [9:0] m81_44;
   assign m81_44 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_45 = W*in
   wire signed [9:0] m81_45;
   assign m81_45 =10'b0;

   // m81_46 = W*in
   wire signed [9:0] m81_46;
   assign m81_46 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_47 = W*in
   wire signed [9:0] m81_47;
   assign m81_47 =10'b0;

   // m81_48 = W*in
   wire signed [9:0] m81_48;
   assign m81_48 =10'b0;

   // m81_49 = W*in
   wire signed [9:0] m81_49;
   assign m81_49 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_50 = W*in
   wire signed [9:0] m81_50;
   assign m81_50 =10'b0;

   // m81_51 = W*in
   wire signed [9:0] m81_51;
   assign m81_51 =10'b0;

   // m81_52 = W*in
   wire signed [9:0] m81_52;
   assign m81_52 =10'b0;

   // m81_53 = W*in
   wire signed [9:0] m81_53;
   assign m81_53 ={ {2{in81[5]}} , in81 , {2{1'b0}} };

   // m81_54 = W*in
   wire signed [9:0] m81_54;
   assign m81_54 =10'b0;

   // m81_55 = W*in
   wire signed [9:0] m81_55;
   assign m81_55 =10'b0;

   // m81_56 = W*in
   wire signed [9:0] m81_56;
   assign m81_56 =10'b0;

   // m81_57 = W*in
   wire signed [9:0] m81_57;
   assign m81_57 =10'b0;

   // m81_58 = W*in
   wire signed [9:0] m81_58;
   assign m81_58 =10'b0;

   // m81_59 = W*in
   wire signed [9:0] m81_59;
   assign m81_59 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_60 = W*in
   wire signed [9:0] m81_60;
   assign m81_60 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_61 = W*in
   wire signed [9:0] m81_61;
   assign m81_61 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_62 = W*in
   wire signed [9:0] m81_62;
   assign m81_62 =10'b0;

   // m81_63 = W*in
   wire signed [9:0] m81_63;
   assign m81_63 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_64 = W*in
   wire signed [9:0] m81_64;
   assign m81_64 =10'b0;

   // m81_65 = W*in
   wire signed [9:0] m81_65;
   assign m81_65 =10'b0;

   // m81_66 = W*in
   wire signed [9:0] m81_66;
   assign m81_66 =10'b0;

   // m81_67 = W*in
   wire signed [9:0] m81_67;
   assign m81_67 =10'b0;

   // m81_68 = W*in
   wire signed [9:0] m81_68;
   assign m81_68 =10'b0;

   // m81_69 = W*in
   wire signed [9:0] m81_69;
   assign m81_69 =10'b0;

   // m81_70 = W*in
   wire signed [9:0] m81_70;
   assign m81_70 ={ {3{in81[5]}} , in81 , {1{1'b0}} };

   // m81_71 = W*in
   wire signed [9:0] m81_71;
   assign m81_71 =10'b0;

   // m81_72 = W*in
   wire signed [9:0] m81_72;
   assign m81_72 ={ {2{in81[5]}} , in81 , {2{1'b0}} };

   // m81_73 = W*in
   wire signed [9:0] m81_73;
   assign m81_73 =10'b0;

   // m81_74 = W*in
   wire signed [9:0] m81_74;
   assign m81_74 =10'b0;

   // m81_75 = W*in
   wire signed [9:0] m81_75;
   assign m81_75 =10'b0;

   // m81_76 = W*in
   wire signed [9:0] m81_76;
   assign m81_76 =10'b0;

   // m81_77 = W*in
   wire signed [9:0] m81_77;
   assign m81_77 =10'b0;

   // m81_78 = W*in
   wire signed [9:0] m81_78;
   assign m81_78 =10'b0;

   // m81_79 = W*in
   wire signed [9:0] m81_79;
   assign m81_79 =10'b0;

   // m81_80 = W*in
   wire signed [9:0] m81_80;
   assign m81_80 =10'b0;

   // m81_81 = W*in
   wire signed [9:0] m81_81;
   assign m81_81 =10'b0;

   // m82_1 = W*in
   wire signed [9:0] m82_1;
   assign m82_1 =10'b0;

   // m82_2 = W*in
   wire signed [9:0] m82_2;
   assign m82_2 =10'b0;

   // m82_3 = W*in
   wire signed [9:0] m82_3;
   assign m82_3 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_4 = W*in
   wire signed [9:0] m82_4;
   assign m82_4 ={ {2{in82[5]}} , in82 , {2{1'b0}} };

   // m82_5 = W*in
   wire signed [9:0] m82_5;
   assign m82_5 =10'b0;

   // m82_6 = W*in
   wire signed [9:0] m82_6;
   assign m82_6 =10'b0;

   // m82_7 = W*in
   wire signed [9:0] m82_7;
   assign m82_7 =10'b0;

   // m82_8 = W*in
   wire signed [9:0] m82_8;
   assign m82_8 =10'b0;

   // m82_9 = W*in
   wire signed [9:0] m82_9;
   assign m82_9 =10'b0;

   // m82_10 = W*in
   wire signed [9:0] m82_10;
   assign m82_10 ={ {2{in82[5]}} , in82 , {2{1'b0}} };

   // m82_11 = W*in
   wire signed [9:0] m82_11;
   assign m82_11 =10'b0;

   // m82_12 = W*in
   wire signed [9:0] m82_12;
   assign m82_12 ={ {2{in82[5]}} , in82 , {2{1'b0}} };

   // m82_13 = W*in
   wire signed [9:0] m82_13;
   assign m82_13 =10'b0;

   // m82_14 = W*in
   wire signed [9:0] m82_14;
   assign m82_14 =10'b0;

   // m82_15 = W*in
   wire signed [9:0] m82_15;
   assign m82_15 =10'b0;

   // m82_16 = W*in
   wire signed [9:0] m82_16;
   assign m82_16 =10'b0;

   // m82_17 = W*in
   wire signed [9:0] m82_17;
   assign m82_17 =10'b0;

   // m82_18 = W*in
   wire signed [9:0] m82_18;
   assign m82_18 =10'b0;

   // m82_19 = W*in
   wire signed [9:0] m82_19;
   assign m82_19 =10'b0;

   // m82_20 = W*in
   wire signed [9:0] m82_20;
   assign m82_20 ={ {2{in82[5]}} , in82 , {2{1'b0}} };

   // m82_21 = W*in
   wire signed [9:0] m82_21;
   assign m82_21 =10'b0;

   // m82_22 = W*in
   wire signed [9:0] m82_22;
   assign m82_22 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_23 = W*in
   wire signed [9:0] m82_23;
   assign m82_23 =10'b0;

   // m82_24 = W*in
   wire signed [9:0] m82_24;
   assign m82_24 =10'b0;

   // m82_25 = W*in
   wire signed [9:0] m82_25;
   assign m82_25 =10'b0;

   // m82_26 = W*in
   wire signed [9:0] m82_26;
   assign m82_26 =10'b0;

   // m82_27 = W*in
   wire signed [9:0] m82_27;
   assign m82_27 =10'b0;

   // m82_28 = W*in
   wire signed [9:0] m82_28;
   assign m82_28 =10'b0;

   // m82_29 = W*in
   wire signed [9:0] m82_29;
   assign m82_29 ={ {2{in82[5]}} , in82 , {2{1'b0}} };

   // m82_30 = W*in
   wire signed [9:0] m82_30;
   assign m82_30 ={ {3{neg82[5]}} , neg82 , {1{1'b0}} };

   // m82_31 = W*in
   wire signed [9:0] m82_31;
   assign m82_31 =10'b0;

   // m82_32 = W*in
   wire signed [9:0] m82_32;
   assign m82_32 ={ {3{neg82[5]}} , neg82 , {1{1'b0}} };

   // m82_33 = W*in
   wire signed [9:0] m82_33;
   assign m82_33 =10'b0;

   // m82_34 = W*in
   wire signed [9:0] m82_34;
   assign m82_34 =10'b0;

   // m82_35 = W*in
   wire signed [9:0] m82_35;
   assign m82_35 =10'b0;

   // m82_36 = W*in
   wire signed [9:0] m82_36;
   assign m82_36 =10'b0;

   // m82_37 = W*in
   wire signed [9:0] m82_37;
   assign m82_37 =10'b0;

   // m82_38 = W*in
   wire signed [9:0] m82_38;
   assign m82_38 =10'b0;

   // m82_39 = W*in
   wire signed [9:0] m82_39;
   assign m82_39 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_40 = W*in
   wire signed [9:0] m82_40;
   assign m82_40 =10'b0;

   // m82_41 = W*in
   wire signed [9:0] m82_41;
   assign m82_41 =10'b0;

   // m82_42 = W*in
   wire signed [9:0] m82_42;
   assign m82_42 =10'b0;

   // m82_43 = W*in
   wire signed [9:0] m82_43;
   assign m82_43 ={ {3{neg82[5]}} , neg82 , {1{1'b0}} };

   // m82_44 = W*in
   wire signed [9:0] m82_44;
   assign m82_44 =10'b0;

   // m82_45 = W*in
   wire signed [9:0] m82_45;
   assign m82_45 =10'b0;

   // m82_46 = W*in
   wire signed [9:0] m82_46;
   assign m82_46 =10'b0;

   // m82_47 = W*in
   wire signed [9:0] m82_47;
   assign m82_47 =10'b0;

   // m82_48 = W*in
   wire signed [9:0] m82_48;
   assign m82_48 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_49 = W*in
   wire signed [9:0] m82_49;
   assign m82_49 =10'b0;

   // m82_50 = W*in
   wire signed [9:0] m82_50;
   assign m82_50 =10'b0;

   // m82_51 = W*in
   wire signed [9:0] m82_51;
   assign m82_51 =10'b0;

   // m82_52 = W*in
   wire signed [9:0] m82_52;
   assign m82_52 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_53 = W*in
   wire signed [9:0] m82_53;
   assign m82_53 =10'b0;

   // m82_54 = W*in
   wire signed [9:0] m82_54;
   assign m82_54 =10'b0;

   // m82_55 = W*in
   wire signed [9:0] m82_55;
   assign m82_55 =10'b0;

   // m82_56 = W*in
   wire signed [9:0] m82_56;
   assign m82_56 =10'b0;

   // m82_57 = W*in
   wire signed [9:0] m82_57;
   assign m82_57 =10'b0;

   // m82_58 = W*in
   wire signed [9:0] m82_58;
   assign m82_58 =10'b0;

   // m82_59 = W*in
   wire signed [9:0] m82_59;
   assign m82_59 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_60 = W*in
   wire signed [9:0] m82_60;
   assign m82_60 =10'b0;

   // m82_61 = W*in
   wire signed [9:0] m82_61;
   assign m82_61 =10'b0;

   // m82_62 = W*in
   wire signed [9:0] m82_62;
   assign m82_62 ={ {3{neg82[5]}} , neg82 , {1{1'b0}} };

   // m82_63 = W*in
   wire signed [9:0] m82_63;
   assign m82_63 ={ {3{neg82[5]}} , neg82 , {1{1'b0}} };

   // m82_64 = W*in
   wire signed [9:0] m82_64;
   assign m82_64 =10'b0;

   // m82_65 = W*in
   wire signed [9:0] m82_65;
   assign m82_65 =10'b0;

   // m82_66 = W*in
   wire signed [9:0] m82_66;
   assign m82_66 =10'b0;

   // m82_67 = W*in
   wire signed [9:0] m82_67;
   assign m82_67 =10'b0;

   // m82_68 = W*in
   wire signed [9:0] m82_68;
   assign m82_68 =10'b0;

   // m82_69 = W*in
   wire signed [9:0] m82_69;
   assign m82_69 =10'b0;

   // m82_70 = W*in
   wire signed [9:0] m82_70;
   assign m82_70 =10'b0;

   // m82_71 = W*in
   wire signed [9:0] m82_71;
   assign m82_71 =10'b0;

   // m82_72 = W*in
   wire signed [9:0] m82_72;
   assign m82_72 =10'b0;

   // m82_73 = W*in
   wire signed [9:0] m82_73;
   assign m82_73 =10'b0;

   // m82_74 = W*in
   wire signed [9:0] m82_74;
   assign m82_74 =10'b0;

   // m82_75 = W*in
   wire signed [9:0] m82_75;
   assign m82_75 =10'b0;

   // m82_76 = W*in
   wire signed [9:0] m82_76;
   assign m82_76 =10'b0;

   // m82_77 = W*in
   wire signed [9:0] m82_77;
   assign m82_77 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_78 = W*in
   wire signed [9:0] m82_78;
   assign m82_78 ={ {3{in82[5]}} , in82 , {1{1'b0}} };

   // m82_79 = W*in
   wire signed [9:0] m82_79;
   assign m82_79 =10'b0;

   // m82_80 = W*in
   wire signed [9:0] m82_80;
   assign m82_80 =10'b0;

   // m82_81 = W*in
   wire signed [9:0] m82_81;
   assign m82_81 =10'b0;

   // m83_1 = W*in
   wire signed [9:0] m83_1;
   assign m83_1 =10'b0;

   // m83_2 = W*in
   wire signed [9:0] m83_2;
   assign m83_2 =10'b0;

   // m83_3 = W*in
   wire signed [9:0] m83_3;
   assign m83_3 =10'b0;

   // m83_4 = W*in
   wire signed [9:0] m83_4;
   assign m83_4 =10'b0;

   // m83_5 = W*in
   wire signed [9:0] m83_5;
   assign m83_5 =10'b0;

   // m83_6 = W*in
   wire signed [9:0] m83_6;
   assign m83_6 =10'b0;

   // m83_7 = W*in
   wire signed [9:0] m83_7;
   assign m83_7 =10'b0;

   // m83_8 = W*in
   wire signed [9:0] m83_8;
   assign m83_8 =10'b0;

   // m83_9 = W*in
   wire signed [9:0] m83_9;
   assign m83_9 =10'b0;

   // m83_10 = W*in
   wire signed [9:0] m83_10;
   assign m83_10 =10'b0;

   // m83_11 = W*in
   wire signed [9:0] m83_11;
   assign m83_11 =10'b0;

   // m83_12 = W*in
   wire signed [9:0] m83_12;
   assign m83_12 =10'b0;

   // m83_13 = W*in
   wire signed [9:0] m83_13;
   assign m83_13 =10'b0;

   // m83_14 = W*in
   wire signed [9:0] m83_14;
   assign m83_14 =10'b0;

   // m83_15 = W*in
   wire signed [9:0] m83_15;
   assign m83_15 =10'b0;

   // m83_16 = W*in
   wire signed [9:0] m83_16;
   assign m83_16 =10'b0;

   // m83_17 = W*in
   wire signed [9:0] m83_17;
   assign m83_17 ={ {2{in83[5]}} , in83 , {2{1'b0}} };

   // m83_18 = W*in
   wire signed [9:0] m83_18;
   assign m83_18 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_19 = W*in
   wire signed [9:0] m83_19;
   assign m83_19 ={ {2{in83[5]}} , in83 , {2{1'b0}} };

   // m83_20 = W*in
   wire signed [9:0] m83_20;
   assign m83_20 =10'b0;

   // m83_21 = W*in
   wire signed [9:0] m83_21;
   assign m83_21 ={ {2{in83[5]}} , in83 , {2{1'b0}} };

   // m83_22 = W*in
   wire signed [9:0] m83_22;
   assign m83_22 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_23 = W*in
   wire signed [9:0] m83_23;
   assign m83_23 =10'b0;

   // m83_24 = W*in
   wire signed [9:0] m83_24;
   assign m83_24 =10'b0;

   // m83_25 = W*in
   wire signed [9:0] m83_25;
   assign m83_25 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_26 = W*in
   wire signed [9:0] m83_26;
   assign m83_26 =10'b0;

   // m83_27 = W*in
   wire signed [9:0] m83_27;
   assign m83_27 =10'b0;

   // m83_28 = W*in
   wire signed [9:0] m83_28;
   assign m83_28 =10'b0;

   // m83_29 = W*in
   wire signed [9:0] m83_29;
   assign m83_29 =10'b0;

   // m83_30 = W*in
   wire signed [9:0] m83_30;
   assign m83_30 =10'b0;

   // m83_31 = W*in
   wire signed [9:0] m83_31;
   assign m83_31 =10'b0;

   // m83_32 = W*in
   wire signed [9:0] m83_32;
   assign m83_32 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_33 = W*in
   wire signed [9:0] m83_33;
   assign m83_33 =10'b0;

   // m83_34 = W*in
   wire signed [9:0] m83_34;
   assign m83_34 =10'b0;

   // m83_35 = W*in
   wire signed [9:0] m83_35;
   assign m83_35 =10'b0;

   // m83_36 = W*in
   wire signed [9:0] m83_36;
   assign m83_36 =10'b0;

   // m83_37 = W*in
   wire signed [9:0] m83_37;
   assign m83_37 =10'b0;

   // m83_38 = W*in
   wire signed [9:0] m83_38;
   assign m83_38 =10'b0;

   // m83_39 = W*in
   wire signed [9:0] m83_39;
   assign m83_39 =10'b0;

   // m83_40 = W*in
   wire signed [9:0] m83_40;
   assign m83_40 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_41 = W*in
   wire signed [9:0] m83_41;
   assign m83_41 =10'b0;

   // m83_42 = W*in
   wire signed [9:0] m83_42;
   assign m83_42 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_43 = W*in
   wire signed [9:0] m83_43;
   assign m83_43 =10'b0;

   // m83_44 = W*in
   wire signed [9:0] m83_44;
   assign m83_44 =10'b0;

   // m83_45 = W*in
   wire signed [9:0] m83_45;
   assign m83_45 =10'b0;

   // m83_46 = W*in
   wire signed [9:0] m83_46;
   assign m83_46 =10'b0;

   // m83_47 = W*in
   wire signed [9:0] m83_47;
   assign m83_47 =10'b0;

   // m83_48 = W*in
   wire signed [9:0] m83_48;
   assign m83_48 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_49 = W*in
   wire signed [9:0] m83_49;
   assign m83_49 =10'b0;

   // m83_50 = W*in
   wire signed [9:0] m83_50;
   assign m83_50 =10'b0;

   // m83_51 = W*in
   wire signed [9:0] m83_51;
   assign m83_51 =10'b0;

   // m83_52 = W*in
   wire signed [9:0] m83_52;
   assign m83_52 ={ {2{in83[5]}} , in83 , {2{1'b0}} };

   // m83_53 = W*in
   wire signed [9:0] m83_53;
   assign m83_53 ={ {2{in83[5]}} , in83 , {2{1'b0}} };

   // m83_54 = W*in
   wire signed [9:0] m83_54;
   assign m83_54 =10'b0;

   // m83_55 = W*in
   wire signed [9:0] m83_55;
   assign m83_55 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_56 = W*in
   wire signed [9:0] m83_56;
   assign m83_56 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_57 = W*in
   wire signed [9:0] m83_57;
   assign m83_57 ={ {2{in83[5]}} , in83 , {2{1'b0}} };

   // m83_58 = W*in
   wire signed [9:0] m83_58;
   assign m83_58 =10'b0;

   // m83_59 = W*in
   wire signed [9:0] m83_59;
   assign m83_59 =10'b0;

   // m83_60 = W*in
   wire signed [9:0] m83_60;
   assign m83_60 =10'b0;

   // m83_61 = W*in
   wire signed [9:0] m83_61;
   assign m83_61 =10'b0;

   // m83_62 = W*in
   wire signed [9:0] m83_62;
   assign m83_62 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_63 = W*in
   wire signed [9:0] m83_63;
   assign m83_63 =10'b0;

   // m83_64 = W*in
   wire signed [9:0] m83_64;
   assign m83_64 =10'b0;

   // m83_65 = W*in
   wire signed [9:0] m83_65;
   assign m83_65 =10'b0;

   // m83_66 = W*in
   wire signed [9:0] m83_66;
   assign m83_66 =10'b0;

   // m83_67 = W*in
   wire signed [9:0] m83_67;
   assign m83_67 =10'b0;

   // m83_68 = W*in
   wire signed [9:0] m83_68;
   assign m83_68 =10'b0;

   // m83_69 = W*in
   wire signed [9:0] m83_69;
   assign m83_69 =10'b0;

   // m83_70 = W*in
   wire signed [9:0] m83_70;
   assign m83_70 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_71 = W*in
   wire signed [9:0] m83_71;
   assign m83_71 =10'b0;

   // m83_72 = W*in
   wire signed [9:0] m83_72;
   assign m83_72 =10'b0;

   // m83_73 = W*in
   wire signed [9:0] m83_73;
   assign m83_73 =10'b0;

   // m83_74 = W*in
   wire signed [9:0] m83_74;
   assign m83_74 =10'b0;

   // m83_75 = W*in
   wire signed [9:0] m83_75;
   assign m83_75 =10'b0;

   // m83_76 = W*in
   wire signed [9:0] m83_76;
   assign m83_76 =10'b0;

   // m83_77 = W*in
   wire signed [9:0] m83_77;
   assign m83_77 =10'b0;

   // m83_78 = W*in
   wire signed [9:0] m83_78;
   assign m83_78 =10'b0;

   // m83_79 = W*in
   wire signed [9:0] m83_79;
   assign m83_79 =10'b0;

   // m83_80 = W*in
   wire signed [9:0] m83_80;
   assign m83_80 =10'b0;

   // m83_81 = W*in
   wire signed [9:0] m83_81;
   assign m83_81 =10'b0;

   // m84_1 = W*in
   wire signed [9:0] m84_1;
   assign m84_1 =10'b0;

   // m84_2 = W*in
   wire signed [9:0] m84_2;
   assign m84_2 =10'b0;

   // m84_3 = W*in
   wire signed [9:0] m84_3;
   assign m84_3 =10'b0;

   // m84_4 = W*in
   wire signed [9:0] m84_4;
   assign m84_4 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_5 = W*in
   wire signed [9:0] m84_5;
   assign m84_5 =10'b0;

   // m84_6 = W*in
   wire signed [9:0] m84_6;
   assign m84_6 =10'b0;

   // m84_7 = W*in
   wire signed [9:0] m84_7;
   assign m84_7 =10'b0;

   // m84_8 = W*in
   wire signed [9:0] m84_8;
   assign m84_8 =10'b0;

   // m84_9 = W*in
   wire signed [9:0] m84_9;
   assign m84_9 =10'b0;

   // m84_10 = W*in
   wire signed [9:0] m84_10;
   assign m84_10 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_11 = W*in
   wire signed [9:0] m84_11;
   assign m84_11 =10'b0;

   // m84_12 = W*in
   wire signed [9:0] m84_12;
   assign m84_12 =10'b0;

   // m84_13 = W*in
   wire signed [9:0] m84_13;
   assign m84_13 =10'b0;

   // m84_14 = W*in
   wire signed [9:0] m84_14;
   assign m84_14 =10'b0;

   // m84_15 = W*in
   wire signed [9:0] m84_15;
   assign m84_15 =10'b0;

   // m84_16 = W*in
   wire signed [9:0] m84_16;
   assign m84_16 =10'b0;

   // m84_17 = W*in
   wire signed [9:0] m84_17;
   assign m84_17 =10'b0;

   // m84_18 = W*in
   wire signed [9:0] m84_18;
   assign m84_18 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_19 = W*in
   wire signed [9:0] m84_19;
   assign m84_19 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_20 = W*in
   wire signed [9:0] m84_20;
   assign m84_20 =10'b0;

   // m84_21 = W*in
   wire signed [9:0] m84_21;
   assign m84_21 =10'b0;

   // m84_22 = W*in
   wire signed [9:0] m84_22;
   assign m84_22 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_23 = W*in
   wire signed [9:0] m84_23;
   assign m84_23 ={ {2{in84[5]}} , in84 , {2{1'b0}} };

   // m84_24 = W*in
   wire signed [9:0] m84_24;
   assign m84_24 =10'b0;

   // m84_25 = W*in
   wire signed [9:0] m84_25;
   assign m84_25 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_26 = W*in
   wire signed [9:0] m84_26;
   assign m84_26 =10'b0;

   // m84_27 = W*in
   wire signed [9:0] m84_27;
   assign m84_27 =10'b0;

   // m84_28 = W*in
   wire signed [9:0] m84_28;
   assign m84_28 =10'b0;

   // m84_29 = W*in
   wire signed [9:0] m84_29;
   assign m84_29 =10'b0;

   // m84_30 = W*in
   wire signed [9:0] m84_30;
   assign m84_30 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_31 = W*in
   wire signed [9:0] m84_31;
   assign m84_31 =10'b0;

   // m84_32 = W*in
   wire signed [9:0] m84_32;
   assign m84_32 =10'b0;

   // m84_33 = W*in
   wire signed [9:0] m84_33;
   assign m84_33 =10'b0;

   // m84_34 = W*in
   wire signed [9:0] m84_34;
   assign m84_34 =10'b0;

   // m84_35 = W*in
   wire signed [9:0] m84_35;
   assign m84_35 =10'b0;

   // m84_36 = W*in
   wire signed [9:0] m84_36;
   assign m84_36 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_37 = W*in
   wire signed [9:0] m84_37;
   assign m84_37 =10'b0;

   // m84_38 = W*in
   wire signed [9:0] m84_38;
   assign m84_38 =10'b0;

   // m84_39 = W*in
   wire signed [9:0] m84_39;
   assign m84_39 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_40 = W*in
   wire signed [9:0] m84_40;
   assign m84_40 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_41 = W*in
   wire signed [9:0] m84_41;
   assign m84_41 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_42 = W*in
   wire signed [9:0] m84_42;
   assign m84_42 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_43 = W*in
   wire signed [9:0] m84_43;
   assign m84_43 =10'b0;

   // m84_44 = W*in
   wire signed [9:0] m84_44;
   assign m84_44 =10'b0;

   // m84_45 = W*in
   wire signed [9:0] m84_45;
   assign m84_45 =10'b0;

   // m84_46 = W*in
   wire signed [9:0] m84_46;
   assign m84_46 =10'b0;

   // m84_47 = W*in
   wire signed [9:0] m84_47;
   assign m84_47 =10'b0;

   // m84_48 = W*in
   wire signed [9:0] m84_48;
   assign m84_48 =10'b0;

   // m84_49 = W*in
   wire signed [9:0] m84_49;
   assign m84_49 =10'b0;

   // m84_50 = W*in
   wire signed [9:0] m84_50;
   assign m84_50 =10'b0;

   // m84_51 = W*in
   wire signed [9:0] m84_51;
   assign m84_51 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_52 = W*in
   wire signed [9:0] m84_52;
   assign m84_52 =10'b0;

   // m84_53 = W*in
   wire signed [9:0] m84_53;
   assign m84_53 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_54 = W*in
   wire signed [9:0] m84_54;
   assign m84_54 =10'b0;

   // m84_55 = W*in
   wire signed [9:0] m84_55;
   assign m84_55 =10'b0;

   // m84_56 = W*in
   wire signed [9:0] m84_56;
   assign m84_56 =10'b0;

   // m84_57 = W*in
   wire signed [9:0] m84_57;
   assign m84_57 =10'b0;

   // m84_58 = W*in
   wire signed [9:0] m84_58;
   assign m84_58 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_59 = W*in
   wire signed [9:0] m84_59;
   assign m84_59 =10'b0;

   // m84_60 = W*in
   wire signed [9:0] m84_60;
   assign m84_60 ={ {3{neg84[5]}} , neg84 , {1{1'b0}} };

   // m84_61 = W*in
   wire signed [9:0] m84_61;
   assign m84_61 =10'b0;

   // m84_62 = W*in
   wire signed [9:0] m84_62;
   assign m84_62 ={ {3{in84[5]}} , in84 , {1{1'b0}} };

   // m84_63 = W*in
   wire signed [9:0] m84_63;
   assign m84_63 =10'b0;

   // m84_64 = W*in
   wire signed [9:0] m84_64;
   assign m84_64 =10'b0;

   // m84_65 = W*in
   wire signed [9:0] m84_65;
   assign m84_65 =10'b0;

   // m84_66 = W*in
   wire signed [9:0] m84_66;
   assign m84_66 =10'b0;

   // m84_67 = W*in
   wire signed [9:0] m84_67;
   assign m84_67 =10'b0;

   // m84_68 = W*in
   wire signed [9:0] m84_68;
   assign m84_68 =10'b0;

   // m84_69 = W*in
   wire signed [9:0] m84_69;
   assign m84_69 =10'b0;

   // m84_70 = W*in
   wire signed [9:0] m84_70;
   assign m84_70 =10'b0;

   // m84_71 = W*in
   wire signed [9:0] m84_71;
   assign m84_71 ={ {2{in84[5]}} , in84 , {2{1'b0}} };

   // m84_72 = W*in
   wire signed [9:0] m84_72;
   assign m84_72 =10'b0;

   // m84_73 = W*in
   wire signed [9:0] m84_73;
   assign m84_73 =10'b0;

   // m84_74 = W*in
   wire signed [9:0] m84_74;
   assign m84_74 =10'b0;

   // m84_75 = W*in
   wire signed [9:0] m84_75;
   assign m84_75 =10'b0;

   // m84_76 = W*in
   wire signed [9:0] m84_76;
   assign m84_76 =10'b0;

   // m84_77 = W*in
   wire signed [9:0] m84_77;
   assign m84_77 =10'b0;

   // m84_78 = W*in
   wire signed [9:0] m84_78;
   assign m84_78 =10'b0;

   // m84_79 = W*in
   wire signed [9:0] m84_79;
   assign m84_79 =10'b0;

   // m84_80 = W*in
   wire signed [9:0] m84_80;
   assign m84_80 =10'b0;

   // m84_81 = W*in
   wire signed [9:0] m84_81;
   assign m84_81 =10'b0;

   // m85_1 = W*in
   wire signed [9:0] m85_1;
   assign m85_1 =10'b0;

   // m85_2 = W*in
   wire signed [9:0] m85_2;
   assign m85_2 =10'b0;

   // m85_3 = W*in
   wire signed [9:0] m85_3;
   assign m85_3 =10'b0;

   // m85_4 = W*in
   wire signed [9:0] m85_4;
   assign m85_4 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_5 = W*in
   wire signed [9:0] m85_5;
   assign m85_5 =10'b0;

   // m85_6 = W*in
   wire signed [9:0] m85_6;
   assign m85_6 =10'b0;

   // m85_7 = W*in
   wire signed [9:0] m85_7;
   assign m85_7 =10'b0;

   // m85_8 = W*in
   wire signed [9:0] m85_8;
   assign m85_8 =10'b0;

   // m85_9 = W*in
   wire signed [9:0] m85_9;
   assign m85_9 =10'b0;

   // m85_10 = W*in
   wire signed [9:0] m85_10;
   assign m85_10 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_11 = W*in
   wire signed [9:0] m85_11;
   assign m85_11 =10'b0;

   // m85_12 = W*in
   wire signed [9:0] m85_12;
   assign m85_12 =10'b0;

   // m85_13 = W*in
   wire signed [9:0] m85_13;
   assign m85_13 =10'b0;

   // m85_14 = W*in
   wire signed [9:0] m85_14;
   assign m85_14 =10'b0;

   // m85_15 = W*in
   wire signed [9:0] m85_15;
   assign m85_15 =10'b0;

   // m85_16 = W*in
   wire signed [9:0] m85_16;
   assign m85_16 =10'b0;

   // m85_17 = W*in
   wire signed [9:0] m85_17;
   assign m85_17 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_18 = W*in
   wire signed [9:0] m85_18;
   assign m85_18 =10'b0;

   // m85_19 = W*in
   wire signed [9:0] m85_19;
   assign m85_19 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_20 = W*in
   wire signed [9:0] m85_20;
   assign m85_20 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_21 = W*in
   wire signed [9:0] m85_21;
   assign m85_21 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_22 = W*in
   wire signed [9:0] m85_22;
   assign m85_22 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_23 = W*in
   wire signed [9:0] m85_23;
   assign m85_23 =10'b0;

   // m85_24 = W*in
   wire signed [9:0] m85_24;
   assign m85_24 =10'b0;

   // m85_25 = W*in
   wire signed [9:0] m85_25;
   assign m85_25 =10'b0;

   // m85_26 = W*in
   wire signed [9:0] m85_26;
   assign m85_26 =10'b0;

   // m85_27 = W*in
   wire signed [9:0] m85_27;
   assign m85_27 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_28 = W*in
   wire signed [9:0] m85_28;
   assign m85_28 =10'b0;

   // m85_29 = W*in
   wire signed [9:0] m85_29;
   assign m85_29 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_30 = W*in
   wire signed [9:0] m85_30;
   assign m85_30 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_31 = W*in
   wire signed [9:0] m85_31;
   assign m85_31 =10'b0;

   // m85_32 = W*in
   wire signed [9:0] m85_32;
   assign m85_32 =10'b0;

   // m85_33 = W*in
   wire signed [9:0] m85_33;
   assign m85_33 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_34 = W*in
   wire signed [9:0] m85_34;
   assign m85_34 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_35 = W*in
   wire signed [9:0] m85_35;
   assign m85_35 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_36 = W*in
   wire signed [9:0] m85_36;
   assign m85_36 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_37 = W*in
   wire signed [9:0] m85_37;
   assign m85_37 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_38 = W*in
   wire signed [9:0] m85_38;
   assign m85_38 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_39 = W*in
   wire signed [9:0] m85_39;
   assign m85_39 =10'b0;

   // m85_40 = W*in
   wire signed [9:0] m85_40;
   assign m85_40 =10'b0;

   // m85_41 = W*in
   wire signed [9:0] m85_41;
   assign m85_41 =10'b0;

   // m85_42 = W*in
   wire signed [9:0] m85_42;
   assign m85_42 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_43 = W*in
   wire signed [9:0] m85_43;
   assign m85_43 =10'b0;

   // m85_44 = W*in
   wire signed [9:0] m85_44;
   assign m85_44 =10'b0;

   // m85_45 = W*in
   wire signed [9:0] m85_45;
   assign m85_45 =10'b0;

   // m85_46 = W*in
   wire signed [9:0] m85_46;
   assign m85_46 =10'b0;

   // m85_47 = W*in
   wire signed [9:0] m85_47;
   assign m85_47 =10'b0;

   // m85_48 = W*in
   wire signed [9:0] m85_48;
   assign m85_48 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_49 = W*in
   wire signed [9:0] m85_49;
   assign m85_49 =10'b0;

   // m85_50 = W*in
   wire signed [9:0] m85_50;
   assign m85_50 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_51 = W*in
   wire signed [9:0] m85_51;
   assign m85_51 =10'b0;

   // m85_52 = W*in
   wire signed [9:0] m85_52;
   assign m85_52 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_53 = W*in
   wire signed [9:0] m85_53;
   assign m85_53 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_54 = W*in
   wire signed [9:0] m85_54;
   assign m85_54 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_55 = W*in
   wire signed [9:0] m85_55;
   assign m85_55 =10'b0;

   // m85_56 = W*in
   wire signed [9:0] m85_56;
   assign m85_56 =10'b0;

   // m85_57 = W*in
   wire signed [9:0] m85_57;
   assign m85_57 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_58 = W*in
   wire signed [9:0] m85_58;
   assign m85_58 =10'b0;

   // m85_59 = W*in
   wire signed [9:0] m85_59;
   assign m85_59 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_60 = W*in
   wire signed [9:0] m85_60;
   assign m85_60 =10'b0;

   // m85_61 = W*in
   wire signed [9:0] m85_61;
   assign m85_61 =10'b0;

   // m85_62 = W*in
   wire signed [9:0] m85_62;
   assign m85_62 =10'b0;

   // m85_63 = W*in
   wire signed [9:0] m85_63;
   assign m85_63 ={ {3{neg85[5]}} , neg85 , {1{1'b0}} };

   // m85_64 = W*in
   wire signed [9:0] m85_64;
   assign m85_64 =10'b0;

   // m85_65 = W*in
   wire signed [9:0] m85_65;
   assign m85_65 ={ {2{in85[5]}} , in85 , {2{1'b0}} };

   // m85_66 = W*in
   wire signed [9:0] m85_66;
   assign m85_66 =10'b0;

   // m85_67 = W*in
   wire signed [9:0] m85_67;
   assign m85_67 =10'b0;

   // m85_68 = W*in
   wire signed [9:0] m85_68;
   assign m85_68 =10'b0;

   // m85_69 = W*in
   wire signed [9:0] m85_69;
   assign m85_69 =10'b0;

   // m85_70 = W*in
   wire signed [9:0] m85_70;
   assign m85_70 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_71 = W*in
   wire signed [9:0] m85_71;
   assign m85_71 =10'b0;

   // m85_72 = W*in
   wire signed [9:0] m85_72;
   assign m85_72 =10'b0;

   // m85_73 = W*in
   wire signed [9:0] m85_73;
   assign m85_73 =10'b0;

   // m85_74 = W*in
   wire signed [9:0] m85_74;
   assign m85_74 =10'b0;

   // m85_75 = W*in
   wire signed [9:0] m85_75;
   assign m85_75 =10'b0;

   // m85_76 = W*in
   wire signed [9:0] m85_76;
   assign m85_76 =10'b0;

   // m85_77 = W*in
   wire signed [9:0] m85_77;
   assign m85_77 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_78 = W*in
   wire signed [9:0] m85_78;
   assign m85_78 ={ {3{in85[5]}} , in85 , {1{1'b0}} };

   // m85_79 = W*in
   wire signed [9:0] m85_79;
   assign m85_79 =10'b0;

   // m85_80 = W*in
   wire signed [9:0] m85_80;
   assign m85_80 =10'b0;

   // m85_81 = W*in
   wire signed [9:0] m85_81;
   assign m85_81 =10'b0;

   // m86_1 = W*in
   wire signed [9:0] m86_1;
   assign m86_1 =10'b0;

   // m86_2 = W*in
   wire signed [9:0] m86_2;
   assign m86_2 =10'b0;

   // m86_3 = W*in
   wire signed [9:0] m86_3;
   assign m86_3 =10'b0;

   // m86_4 = W*in
   wire signed [9:0] m86_4;
   assign m86_4 =10'b0;

   // m86_5 = W*in
   wire signed [9:0] m86_5;
   assign m86_5 =10'b0;

   // m86_6 = W*in
   wire signed [9:0] m86_6;
   assign m86_6 =10'b0;

   // m86_7 = W*in
   wire signed [9:0] m86_7;
   assign m86_7 =10'b0;

   // m86_8 = W*in
   wire signed [9:0] m86_8;
   assign m86_8 =10'b0;

   // m86_9 = W*in
   wire signed [9:0] m86_9;
   assign m86_9 =10'b0;

   // m86_10 = W*in
   wire signed [9:0] m86_10;
   assign m86_10 =10'b0;

   // m86_11 = W*in
   wire signed [9:0] m86_11;
   assign m86_11 =10'b0;

   // m86_12 = W*in
   wire signed [9:0] m86_12;
   assign m86_12 =10'b0;

   // m86_13 = W*in
   wire signed [9:0] m86_13;
   assign m86_13 =10'b0;

   // m86_14 = W*in
   wire signed [9:0] m86_14;
   assign m86_14 =10'b0;

   // m86_15 = W*in
   wire signed [9:0] m86_15;
   assign m86_15 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_16 = W*in
   wire signed [9:0] m86_16;
   assign m86_16 =10'b0;

   // m86_17 = W*in
   wire signed [9:0] m86_17;
   assign m86_17 =10'b0;

   // m86_18 = W*in
   wire signed [9:0] m86_18;
   assign m86_18 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_19 = W*in
   wire signed [9:0] m86_19;
   assign m86_19 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_20 = W*in
   wire signed [9:0] m86_20;
   assign m86_20 =10'b0;

   // m86_21 = W*in
   wire signed [9:0] m86_21;
   assign m86_21 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_22 = W*in
   wire signed [9:0] m86_22;
   assign m86_22 =10'b0;

   // m86_23 = W*in
   wire signed [9:0] m86_23;
   assign m86_23 =10'b0;

   // m86_24 = W*in
   wire signed [9:0] m86_24;
   assign m86_24 =10'b0;

   // m86_25 = W*in
   wire signed [9:0] m86_25;
   assign m86_25 =10'b0;

   // m86_26 = W*in
   wire signed [9:0] m86_26;
   assign m86_26 =10'b0;

   // m86_27 = W*in
   wire signed [9:0] m86_27;
   assign m86_27 =10'b0;

   // m86_28 = W*in
   wire signed [9:0] m86_28;
   assign m86_28 =10'b0;

   // m86_29 = W*in
   wire signed [9:0] m86_29;
   assign m86_29 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_30 = W*in
   wire signed [9:0] m86_30;
   assign m86_30 =10'b0;

   // m86_31 = W*in
   wire signed [9:0] m86_31;
   assign m86_31 =10'b0;

   // m86_32 = W*in
   wire signed [9:0] m86_32;
   assign m86_32 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_33 = W*in
   wire signed [9:0] m86_33;
   assign m86_33 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_34 = W*in
   wire signed [9:0] m86_34;
   assign m86_34 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_35 = W*in
   wire signed [9:0] m86_35;
   assign m86_35 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_36 = W*in
   wire signed [9:0] m86_36;
   assign m86_36 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_37 = W*in
   wire signed [9:0] m86_37;
   assign m86_37 =10'b0;

   // m86_38 = W*in
   wire signed [9:0] m86_38;
   assign m86_38 ={ {2{in86[5]}} , in86 , {2{1'b0}} };

   // m86_39 = W*in
   wire signed [9:0] m86_39;
   assign m86_39 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_40 = W*in
   wire signed [9:0] m86_40;
   assign m86_40 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_41 = W*in
   wire signed [9:0] m86_41;
   assign m86_41 =10'b0;

   // m86_42 = W*in
   wire signed [9:0] m86_42;
   assign m86_42 ={ {3{in86[5]}} , in86 , {1{1'b0}} };

   // m86_43 = W*in
   wire signed [9:0] m86_43;
   assign m86_43 =10'b0;

   // m86_44 = W*in
   wire signed [9:0] m86_44;
   assign m86_44 =10'b0;

   // m86_45 = W*in
   wire signed [9:0] m86_45;
   assign m86_45 =10'b0;

   // m86_46 = W*in
   wire signed [9:0] m86_46;
   assign m86_46 =10'b0;

   // m86_47 = W*in
   wire signed [9:0] m86_47;
   assign m86_47 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_48 = W*in
   wire signed [9:0] m86_48;
   assign m86_48 =10'b0;

   // m86_49 = W*in
   wire signed [9:0] m86_49;
   assign m86_49 =10'b0;

   // m86_50 = W*in
   wire signed [9:0] m86_50;
   assign m86_50 ={ {2{in86[5]}} , in86 , {2{1'b0}} };

   // m86_51 = W*in
   wire signed [9:0] m86_51;
   assign m86_51 =10'b0;

   // m86_52 = W*in
   wire signed [9:0] m86_52;
   assign m86_52 =10'b0;

   // m86_53 = W*in
   wire signed [9:0] m86_53;
   assign m86_53 =10'b0;

   // m86_54 = W*in
   wire signed [9:0] m86_54;
   assign m86_54 =10'b0;

   // m86_55 = W*in
   wire signed [9:0] m86_55;
   assign m86_55 =10'b0;

   // m86_56 = W*in
   wire signed [9:0] m86_56;
   assign m86_56 =10'b0;

   // m86_57 = W*in
   wire signed [9:0] m86_57;
   assign m86_57 =10'b0;

   // m86_58 = W*in
   wire signed [9:0] m86_58;
   assign m86_58 =10'b0;

   // m86_59 = W*in
   wire signed [9:0] m86_59;
   assign m86_59 =10'b0;

   // m86_60 = W*in
   wire signed [9:0] m86_60;
   assign m86_60 =10'b0;

   // m86_61 = W*in
   wire signed [9:0] m86_61;
   assign m86_61 =10'b0;

   // m86_62 = W*in
   wire signed [9:0] m86_62;
   assign m86_62 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_63 = W*in
   wire signed [9:0] m86_63;
   assign m86_63 =10'b0;

   // m86_64 = W*in
   wire signed [9:0] m86_64;
   assign m86_64 =10'b0;

   // m86_65 = W*in
   wire signed [9:0] m86_65;
   assign m86_65 =10'b0;

   // m86_66 = W*in
   wire signed [9:0] m86_66;
   assign m86_66 =10'b0;

   // m86_67 = W*in
   wire signed [9:0] m86_67;
   assign m86_67 =10'b0;

   // m86_68 = W*in
   wire signed [9:0] m86_68;
   assign m86_68 =10'b0;

   // m86_69 = W*in
   wire signed [9:0] m86_69;
   assign m86_69 =10'b0;

   // m86_70 = W*in
   wire signed [9:0] m86_70;
   assign m86_70 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_71 = W*in
   wire signed [9:0] m86_71;
   assign m86_71 =10'b0;

   // m86_72 = W*in
   wire signed [9:0] m86_72;
   assign m86_72 =10'b0;

   // m86_73 = W*in
   wire signed [9:0] m86_73;
   assign m86_73 =10'b0;

   // m86_74 = W*in
   wire signed [9:0] m86_74;
   assign m86_74 =10'b0;

   // m86_75 = W*in
   wire signed [9:0] m86_75;
   assign m86_75 =10'b0;

   // m86_76 = W*in
   wire signed [9:0] m86_76;
   assign m86_76 =10'b0;

   // m86_77 = W*in
   wire signed [9:0] m86_77;
   assign m86_77 ={ {2{in86[5]}} , in86 , {2{1'b0}} };

   // m86_78 = W*in
   wire signed [9:0] m86_78;
   assign m86_78 =10'b0;

   // m86_79 = W*in
   wire signed [9:0] m86_79;
   assign m86_79 ={ {3{neg86[5]}} , neg86 , {1{1'b0}} };

   // m86_80 = W*in
   wire signed [9:0] m86_80;
   assign m86_80 =10'b0;

   // m86_81 = W*in
   wire signed [9:0] m86_81;
   assign m86_81 =10'b0;

   // m87_1 = W*in
   wire signed [9:0] m87_1;
   assign m87_1 =10'b0;

   // m87_2 = W*in
   wire signed [9:0] m87_2;
   assign m87_2 =10'b0;

   // m87_3 = W*in
   wire signed [9:0] m87_3;
   assign m87_3 ={ {3{neg87[5]}} , neg87 , {1{1'b0}} };

   // m87_4 = W*in
   wire signed [9:0] m87_4;
   assign m87_4 =10'b0;

   // m87_5 = W*in
   wire signed [9:0] m87_5;
   assign m87_5 =10'b0;

   // m87_6 = W*in
   wire signed [9:0] m87_6;
   assign m87_6 =10'b0;

   // m87_7 = W*in
   wire signed [9:0] m87_7;
   assign m87_7 =10'b0;

   // m87_8 = W*in
   wire signed [9:0] m87_8;
   assign m87_8 =10'b0;

   // m87_9 = W*in
   wire signed [9:0] m87_9;
   assign m87_9 =10'b0;

   // m87_10 = W*in
   wire signed [9:0] m87_10;
   assign m87_10 =10'b0;

   // m87_11 = W*in
   wire signed [9:0] m87_11;
   assign m87_11 =10'b0;

   // m87_12 = W*in
   wire signed [9:0] m87_12;
   assign m87_12 =10'b0;

   // m87_13 = W*in
   wire signed [9:0] m87_13;
   assign m87_13 =10'b0;

   // m87_14 = W*in
   wire signed [9:0] m87_14;
   assign m87_14 =10'b0;

   // m87_15 = W*in
   wire signed [9:0] m87_15;
   assign m87_15 ={ {3{neg87[5]}} , neg87 , {1{1'b0}} };

   // m87_16 = W*in
   wire signed [9:0] m87_16;
   assign m87_16 =10'b0;

   // m87_17 = W*in
   wire signed [9:0] m87_17;
   assign m87_17 =10'b0;

   // m87_18 = W*in
   wire signed [9:0] m87_18;
   assign m87_18 =10'b0;

   // m87_19 = W*in
   wire signed [9:0] m87_19;
   assign m87_19 =10'b0;

   // m87_20 = W*in
   wire signed [9:0] m87_20;
   assign m87_20 =10'b0;

   // m87_21 = W*in
   wire signed [9:0] m87_21;
   assign m87_21 =10'b0;

   // m87_22 = W*in
   wire signed [9:0] m87_22;
   assign m87_22 =10'b0;

   // m87_23 = W*in
   wire signed [9:0] m87_23;
   assign m87_23 ={ {2{in87[5]}} , in87 , {2{1'b0}} };

   // m87_24 = W*in
   wire signed [9:0] m87_24;
   assign m87_24 ={ {3{in87[5]}} , in87 , {1{1'b0}} };

   // m87_25 = W*in
   wire signed [9:0] m87_25;
   assign m87_25 ={ {2{in87[5]}} , in87 , {2{1'b0}} };

   // m87_26 = W*in
   wire signed [9:0] m87_26;
   assign m87_26 =10'b0;

   // m87_27 = W*in
   wire signed [9:0] m87_27;
   assign m87_27 =10'b0;

   // m87_28 = W*in
   wire signed [9:0] m87_28;
   assign m87_28 ={ {3{in87[5]}} , in87 , {1{1'b0}} };

   // m87_29 = W*in
   wire signed [9:0] m87_29;
   assign m87_29 =10'b0;

   // m87_30 = W*in
   wire signed [9:0] m87_30;
   assign m87_30 =10'b0;

   // m87_31 = W*in
   wire signed [9:0] m87_31;
   assign m87_31 =10'b0;

   // m87_32 = W*in
   wire signed [9:0] m87_32;
   assign m87_32 =10'b0;

   // m87_33 = W*in
   wire signed [9:0] m87_33;
   assign m87_33 ={ {3{in87[5]}} , in87 , {1{1'b0}} };

   // m87_34 = W*in
   wire signed [9:0] m87_34;
   assign m87_34 ={ {3{in87[5]}} , in87 , {1{1'b0}} };

   // m87_35 = W*in
   wire signed [9:0] m87_35;
   assign m87_35 =10'b0;

   // m87_36 = W*in
   wire signed [9:0] m87_36;
   assign m87_36 =10'b0;

   // m87_37 = W*in
   wire signed [9:0] m87_37;
   assign m87_37 =10'b0;

   // m87_38 = W*in
   wire signed [9:0] m87_38;
   assign m87_38 =10'b0;

   // m87_39 = W*in
   wire signed [9:0] m87_39;
   assign m87_39 ={ {2{in87[5]}} , in87 , {2{1'b0}} };

   // m87_40 = W*in
   wire signed [9:0] m87_40;
   assign m87_40 =10'b0;

   // m87_41 = W*in
   wire signed [9:0] m87_41;
   assign m87_41 =10'b0;

   // m87_42 = W*in
   wire signed [9:0] m87_42;
   assign m87_42 =10'b0;

   // m87_43 = W*in
   wire signed [9:0] m87_43;
   assign m87_43 =10'b0;

   // m87_44 = W*in
   wire signed [9:0] m87_44;
   assign m87_44 =10'b0;

   // m87_45 = W*in
   wire signed [9:0] m87_45;
   assign m87_45 ={ {2{in87[5]}} , in87 , {2{1'b0}} };

   // m87_46 = W*in
   wire signed [9:0] m87_46;
   assign m87_46 =10'b0;

   // m87_47 = W*in
   wire signed [9:0] m87_47;
   assign m87_47 =10'b0;

   // m87_48 = W*in
   wire signed [9:0] m87_48;
   assign m87_48 =10'b0;

   // m87_49 = W*in
   wire signed [9:0] m87_49;
   assign m87_49 =10'b0;

   // m87_50 = W*in
   wire signed [9:0] m87_50;
   assign m87_50 =10'b0;

   // m87_51 = W*in
   wire signed [9:0] m87_51;
   assign m87_51 =10'b0;

   // m87_52 = W*in
   wire signed [9:0] m87_52;
   assign m87_52 =10'b0;

   // m87_53 = W*in
   wire signed [9:0] m87_53;
   assign m87_53 =10'b0;

   // m87_54 = W*in
   wire signed [9:0] m87_54;
   assign m87_54 =10'b0;

   // m87_55 = W*in
   wire signed [9:0] m87_55;
   assign m87_55 =10'b0;

   // m87_56 = W*in
   wire signed [9:0] m87_56;
   assign m87_56 =10'b0;

   // m87_57 = W*in
   wire signed [9:0] m87_57;
   assign m87_57 =10'b0;

   // m87_58 = W*in
   wire signed [9:0] m87_58;
   assign m87_58 ={ {3{neg87[5]}} , neg87 , {1{1'b0}} };

   // m87_59 = W*in
   wire signed [9:0] m87_59;
   assign m87_59 ={ {3{neg87[5]}} , neg87 , {1{1'b0}} };

   // m87_60 = W*in
   wire signed [9:0] m87_60;
   assign m87_60 =10'b0;

   // m87_61 = W*in
   wire signed [9:0] m87_61;
   assign m87_61 =10'b0;

   // m87_62 = W*in
   wire signed [9:0] m87_62;
   assign m87_62 =10'b0;

   // m87_63 = W*in
   wire signed [9:0] m87_63;
   assign m87_63 =10'b0;

   // m87_64 = W*in
   wire signed [9:0] m87_64;
   assign m87_64 ={ {3{in87[5]}} , in87 , {1{1'b0}} };

   // m87_65 = W*in
   wire signed [9:0] m87_65;
   assign m87_65 =10'b0;

   // m87_66 = W*in
   wire signed [9:0] m87_66;
   assign m87_66 =10'b0;

   // m87_67 = W*in
   wire signed [9:0] m87_67;
   assign m87_67 =10'b0;

   // m87_68 = W*in
   wire signed [9:0] m87_68;
   assign m87_68 =10'b0;

   // m87_69 = W*in
   wire signed [9:0] m87_69;
   assign m87_69 ={ {3{neg87[5]}} , neg87 , {1{1'b0}} };

   // m87_70 = W*in
   wire signed [9:0] m87_70;
   assign m87_70 =10'b0;

   // m87_71 = W*in
   wire signed [9:0] m87_71;
   assign m87_71 =10'b0;

   // m87_72 = W*in
   wire signed [9:0] m87_72;
   assign m87_72 =10'b0;

   // m87_73 = W*in
   wire signed [9:0] m87_73;
   assign m87_73 =10'b0;

   // m87_74 = W*in
   wire signed [9:0] m87_74;
   assign m87_74 =10'b0;

   // m87_75 = W*in
   wire signed [9:0] m87_75;
   assign m87_75 =10'b0;

   // m87_76 = W*in
   wire signed [9:0] m87_76;
   assign m87_76 =10'b0;

   // m87_77 = W*in
   wire signed [9:0] m87_77;
   assign m87_77 =10'b0;

   // m87_78 = W*in
   wire signed [9:0] m87_78;
   assign m87_78 =10'b0;

   // m87_79 = W*in
   wire signed [9:0] m87_79;
   assign m87_79 =10'b0;

   // m87_80 = W*in
   wire signed [9:0] m87_80;
   assign m87_80 =10'b0;

   // m87_81 = W*in
   wire signed [9:0] m87_81;
   assign m87_81 =10'b0;

   // m88_1 = W*in
   wire signed [9:0] m88_1;
   assign m88_1 =10'b0;

   // m88_2 = W*in
   wire signed [9:0] m88_2;
   assign m88_2 =10'b0;

   // m88_3 = W*in
   wire signed [9:0] m88_3;
   assign m88_3 =10'b0;

   // m88_4 = W*in
   wire signed [9:0] m88_4;
   assign m88_4 =10'b0;

   // m88_5 = W*in
   wire signed [9:0] m88_5;
   assign m88_5 =10'b0;

   // m88_6 = W*in
   wire signed [9:0] m88_6;
   assign m88_6 =10'b0;

   // m88_7 = W*in
   wire signed [9:0] m88_7;
   assign m88_7 =10'b0;

   // m88_8 = W*in
   wire signed [9:0] m88_8;
   assign m88_8 =10'b0;

   // m88_9 = W*in
   wire signed [9:0] m88_9;
   assign m88_9 =10'b0;

   // m88_10 = W*in
   wire signed [9:0] m88_10;
   assign m88_10 =10'b0;

   // m88_11 = W*in
   wire signed [9:0] m88_11;
   assign m88_11 =10'b0;

   // m88_12 = W*in
   wire signed [9:0] m88_12;
   assign m88_12 =10'b0;

   // m88_13 = W*in
   wire signed [9:0] m88_13;
   assign m88_13 =10'b0;

   // m88_14 = W*in
   wire signed [9:0] m88_14;
   assign m88_14 ={ {3{neg88[5]}} , neg88 , {1{1'b0}} };

   // m88_15 = W*in
   wire signed [9:0] m88_15;
   assign m88_15 =10'b0;

   // m88_16 = W*in
   wire signed [9:0] m88_16;
   assign m88_16 =10'b0;

   // m88_17 = W*in
   wire signed [9:0] m88_17;
   assign m88_17 =10'b0;

   // m88_18 = W*in
   wire signed [9:0] m88_18;
   assign m88_18 =10'b0;

   // m88_19 = W*in
   wire signed [9:0] m88_19;
   assign m88_19 =10'b0;

   // m88_20 = W*in
   wire signed [9:0] m88_20;
   assign m88_20 ={ {2{in88[5]}} , in88 , {2{1'b0}} };

   // m88_21 = W*in
   wire signed [9:0] m88_21;
   assign m88_21 =10'b0;

   // m88_22 = W*in
   wire signed [9:0] m88_22;
   assign m88_22 =10'b0;

   // m88_23 = W*in
   wire signed [9:0] m88_23;
   assign m88_23 =10'b0;

   // m88_24 = W*in
   wire signed [9:0] m88_24;
   assign m88_24 ={ {3{in88[5]}} , in88 , {1{1'b0}} };

   // m88_25 = W*in
   wire signed [9:0] m88_25;
   assign m88_25 ={ {3{neg88[5]}} , neg88 , {1{1'b0}} };

   // m88_26 = W*in
   wire signed [9:0] m88_26;
   assign m88_26 =10'b0;

   // m88_27 = W*in
   wire signed [9:0] m88_27;
   assign m88_27 =10'b0;

   // m88_28 = W*in
   wire signed [9:0] m88_28;
   assign m88_28 =10'b0;

   // m88_29 = W*in
   wire signed [9:0] m88_29;
   assign m88_29 ={ {3{in88[5]}} , in88 , {1{1'b0}} };

   // m88_30 = W*in
   wire signed [9:0] m88_30;
   assign m88_30 =10'b0;

   // m88_31 = W*in
   wire signed [9:0] m88_31;
   assign m88_31 ={ {3{neg88[5]}} , neg88 , {1{1'b0}} };

   // m88_32 = W*in
   wire signed [9:0] m88_32;
   assign m88_32 =10'b0;

   // m88_33 = W*in
   wire signed [9:0] m88_33;
   assign m88_33 =10'b0;

   // m88_34 = W*in
   wire signed [9:0] m88_34;
   assign m88_34 =10'b0;

   // m88_35 = W*in
   wire signed [9:0] m88_35;
   assign m88_35 =10'b0;

   // m88_36 = W*in
   wire signed [9:0] m88_36;
   assign m88_36 ={ {3{in88[5]}} , in88 , {1{1'b0}} };

   // m88_37 = W*in
   wire signed [9:0] m88_37;
   assign m88_37 =10'b0;

   // m88_38 = W*in
   wire signed [9:0] m88_38;
   assign m88_38 =10'b0;

   // m88_39 = W*in
   wire signed [9:0] m88_39;
   assign m88_39 =10'b0;

   // m88_40 = W*in
   wire signed [9:0] m88_40;
   assign m88_40 ={ {3{in88[5]}} , in88 , {1{1'b0}} };

   // m88_41 = W*in
   wire signed [9:0] m88_41;
   assign m88_41 =10'b0;

   // m88_42 = W*in
   wire signed [9:0] m88_42;
   assign m88_42 =10'b0;

   // m88_43 = W*in
   wire signed [9:0] m88_43;
   assign m88_43 ={ {3{neg88[5]}} , neg88 , {1{1'b0}} };

   // m88_44 = W*in
   wire signed [9:0] m88_44;
   assign m88_44 =10'b0;

   // m88_45 = W*in
   wire signed [9:0] m88_45;
   assign m88_45 ={ {3{in88[5]}} , in88 , {1{1'b0}} };

   // m88_46 = W*in
   wire signed [9:0] m88_46;
   assign m88_46 =10'b0;

   // m88_47 = W*in
   wire signed [9:0] m88_47;
   assign m88_47 =10'b0;

   // m88_48 = W*in
   wire signed [9:0] m88_48;
   assign m88_48 ={ {2{in88[5]}} , in88 , {2{1'b0}} };

   // m88_49 = W*in
   wire signed [9:0] m88_49;
   assign m88_49 ={ {3{in88[5]}} , in88 , {1{1'b0}} };

   // m88_50 = W*in
   wire signed [9:0] m88_50;
   assign m88_50 =10'b0;

   // m88_51 = W*in
   wire signed [9:0] m88_51;
   assign m88_51 =10'b0;

   // m88_52 = W*in
   wire signed [9:0] m88_52;
   assign m88_52 ={ {3{neg88[5]}} , neg88 , {1{1'b0}} };

   // m88_53 = W*in
   wire signed [9:0] m88_53;
   assign m88_53 =10'b0;

   // m88_54 = W*in
   wire signed [9:0] m88_54;
   assign m88_54 =10'b0;

   // m88_55 = W*in
   wire signed [9:0] m88_55;
   assign m88_55 =10'b0;

   // m88_56 = W*in
   wire signed [9:0] m88_56;
   assign m88_56 =10'b0;

   // m88_57 = W*in
   wire signed [9:0] m88_57;
   assign m88_57 =10'b0;

   // m88_58 = W*in
   wire signed [9:0] m88_58;
   assign m88_58 =10'b0;

   // m88_59 = W*in
   wire signed [9:0] m88_59;
   assign m88_59 =10'b0;

   // m88_60 = W*in
   wire signed [9:0] m88_60;
   assign m88_60 =10'b0;

   // m88_61 = W*in
   wire signed [9:0] m88_61;
   assign m88_61 ={ {3{neg88[5]}} , neg88 , {1{1'b0}} };

   // m88_62 = W*in
   wire signed [9:0] m88_62;
   assign m88_62 =10'b0;

   // m88_63 = W*in
   wire signed [9:0] m88_63;
   assign m88_63 =10'b0;

   // m88_64 = W*in
   wire signed [9:0] m88_64;
   assign m88_64 =10'b0;

   // m88_65 = W*in
   wire signed [9:0] m88_65;
   assign m88_65 =10'b0;

   // m88_66 = W*in
   wire signed [9:0] m88_66;
   assign m88_66 =10'b0;

   // m88_67 = W*in
   wire signed [9:0] m88_67;
   assign m88_67 =10'b0;

   // m88_68 = W*in
   wire signed [9:0] m88_68;
   assign m88_68 =10'b0;

   // m88_69 = W*in
   wire signed [9:0] m88_69;
   assign m88_69 =10'b0;

   // m88_70 = W*in
   wire signed [9:0] m88_70;
   assign m88_70 =10'b0;

   // m88_71 = W*in
   wire signed [9:0] m88_71;
   assign m88_71 =10'b0;

   // m88_72 = W*in
   wire signed [9:0] m88_72;
   assign m88_72 =10'b0;

   // m88_73 = W*in
   wire signed [9:0] m88_73;
   assign m88_73 =10'b0;

   // m88_74 = W*in
   wire signed [9:0] m88_74;
   assign m88_74 =10'b0;

   // m88_75 = W*in
   wire signed [9:0] m88_75;
   assign m88_75 ={ {2{in88[5]}} , in88 , {2{1'b0}} };

   // m88_76 = W*in
   wire signed [9:0] m88_76;
   assign m88_76 =10'b0;

   // m88_77 = W*in
   wire signed [9:0] m88_77;
   assign m88_77 =10'b0;

   // m88_78 = W*in
   wire signed [9:0] m88_78;
   assign m88_78 =10'b0;

   // m88_79 = W*in
   wire signed [9:0] m88_79;
   assign m88_79 =10'b0;

   // m88_80 = W*in
   wire signed [9:0] m88_80;
   assign m88_80 =10'b0;

   // m88_81 = W*in
   wire signed [9:0] m88_81;
   assign m88_81 =10'b0;

   // m89_1 = W*in
   wire signed [9:0] m89_1;
   assign m89_1 =10'b0;

   // m89_2 = W*in
   wire signed [9:0] m89_2;
   assign m89_2 =10'b0;

   // m89_3 = W*in
   wire signed [9:0] m89_3;
   assign m89_3 =10'b0;

   // m89_4 = W*in
   wire signed [9:0] m89_4;
   assign m89_4 =10'b0;

   // m89_5 = W*in
   wire signed [9:0] m89_5;
   assign m89_5 =10'b0;

   // m89_6 = W*in
   wire signed [9:0] m89_6;
   assign m89_6 =10'b0;

   // m89_7 = W*in
   wire signed [9:0] m89_7;
   assign m89_7 =10'b0;

   // m89_8 = W*in
   wire signed [9:0] m89_8;
   assign m89_8 =10'b0;

   // m89_9 = W*in
   wire signed [9:0] m89_9;
   assign m89_9 =10'b0;

   // m89_10 = W*in
   wire signed [9:0] m89_10;
   assign m89_10 =10'b0;

   // m89_11 = W*in
   wire signed [9:0] m89_11;
   assign m89_11 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_12 = W*in
   wire signed [9:0] m89_12;
   assign m89_12 =10'b0;

   // m89_13 = W*in
   wire signed [9:0] m89_13;
   assign m89_13 =10'b0;

   // m89_14 = W*in
   wire signed [9:0] m89_14;
   assign m89_14 =10'b0;

   // m89_15 = W*in
   wire signed [9:0] m89_15;
   assign m89_15 =10'b0;

   // m89_16 = W*in
   wire signed [9:0] m89_16;
   assign m89_16 =10'b0;

   // m89_17 = W*in
   wire signed [9:0] m89_17;
   assign m89_17 =10'b0;

   // m89_18 = W*in
   wire signed [9:0] m89_18;
   assign m89_18 =10'b0;

   // m89_19 = W*in
   wire signed [9:0] m89_19;
   assign m89_19 =10'b0;

   // m89_20 = W*in
   wire signed [9:0] m89_20;
   assign m89_20 =10'b0;

   // m89_21 = W*in
   wire signed [9:0] m89_21;
   assign m89_21 =10'b0;

   // m89_22 = W*in
   wire signed [9:0] m89_22;
   assign m89_22 =10'b0;

   // m89_23 = W*in
   wire signed [9:0] m89_23;
   assign m89_23 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_24 = W*in
   wire signed [9:0] m89_24;
   assign m89_24 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_25 = W*in
   wire signed [9:0] m89_25;
   assign m89_25 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_26 = W*in
   wire signed [9:0] m89_26;
   assign m89_26 =10'b0;

   // m89_27 = W*in
   wire signed [9:0] m89_27;
   assign m89_27 =10'b0;

   // m89_28 = W*in
   wire signed [9:0] m89_28;
   assign m89_28 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_29 = W*in
   wire signed [9:0] m89_29;
   assign m89_29 =10'b0;

   // m89_30 = W*in
   wire signed [9:0] m89_30;
   assign m89_30 =10'b0;

   // m89_31 = W*in
   wire signed [9:0] m89_31;
   assign m89_31 =10'b0;

   // m89_32 = W*in
   wire signed [9:0] m89_32;
   assign m89_32 =10'b0;

   // m89_33 = W*in
   wire signed [9:0] m89_33;
   assign m89_33 =10'b0;

   // m89_34 = W*in
   wire signed [9:0] m89_34;
   assign m89_34 =10'b0;

   // m89_35 = W*in
   wire signed [9:0] m89_35;
   assign m89_35 =10'b0;

   // m89_36 = W*in
   wire signed [9:0] m89_36;
   assign m89_36 =10'b0;

   // m89_37 = W*in
   wire signed [9:0] m89_37;
   assign m89_37 =10'b0;

   // m89_38 = W*in
   wire signed [9:0] m89_38;
   assign m89_38 =10'b0;

   // m89_39 = W*in
   wire signed [9:0] m89_39;
   assign m89_39 ={ {2{in89[5]}} , in89 , {2{1'b0}} };

   // m89_40 = W*in
   wire signed [9:0] m89_40;
   assign m89_40 =10'b0;

   // m89_41 = W*in
   wire signed [9:0] m89_41;
   assign m89_41 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_42 = W*in
   wire signed [9:0] m89_42;
   assign m89_42 =10'b0;

   // m89_43 = W*in
   wire signed [9:0] m89_43;
   assign m89_43 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_44 = W*in
   wire signed [9:0] m89_44;
   assign m89_44 =10'b0;

   // m89_45 = W*in
   wire signed [9:0] m89_45;
   assign m89_45 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_46 = W*in
   wire signed [9:0] m89_46;
   assign m89_46 =10'b0;

   // m89_47 = W*in
   wire signed [9:0] m89_47;
   assign m89_47 =10'b0;

   // m89_48 = W*in
   wire signed [9:0] m89_48;
   assign m89_48 =10'b0;

   // m89_49 = W*in
   wire signed [9:0] m89_49;
   assign m89_49 =10'b0;

   // m89_50 = W*in
   wire signed [9:0] m89_50;
   assign m89_50 =10'b0;

   // m89_51 = W*in
   wire signed [9:0] m89_51;
   assign m89_51 =10'b0;

   // m89_52 = W*in
   wire signed [9:0] m89_52;
   assign m89_52 =10'b0;

   // m89_53 = W*in
   wire signed [9:0] m89_53;
   assign m89_53 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_54 = W*in
   wire signed [9:0] m89_54;
   assign m89_54 =10'b0;

   // m89_55 = W*in
   wire signed [9:0] m89_55;
   assign m89_55 =10'b0;

   // m89_56 = W*in
   wire signed [9:0] m89_56;
   assign m89_56 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_57 = W*in
   wire signed [9:0] m89_57;
   assign m89_57 =10'b0;

   // m89_58 = W*in
   wire signed [9:0] m89_58;
   assign m89_58 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_59 = W*in
   wire signed [9:0] m89_59;
   assign m89_59 =10'b0;

   // m89_60 = W*in
   wire signed [9:0] m89_60;
   assign m89_60 =10'b0;

   // m89_61 = W*in
   wire signed [9:0] m89_61;
   assign m89_61 =10'b0;

   // m89_62 = W*in
   wire signed [9:0] m89_62;
   assign m89_62 =10'b0;

   // m89_63 = W*in
   wire signed [9:0] m89_63;
   assign m89_63 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_64 = W*in
   wire signed [9:0] m89_64;
   assign m89_64 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_65 = W*in
   wire signed [9:0] m89_65;
   assign m89_65 ={ {2{in89[5]}} , in89 , {2{1'b0}} };

   // m89_66 = W*in
   wire signed [9:0] m89_66;
   assign m89_66 =10'b0;

   // m89_67 = W*in
   wire signed [9:0] m89_67;
   assign m89_67 =10'b0;

   // m89_68 = W*in
   wire signed [9:0] m89_68;
   assign m89_68 ={ {3{neg89[5]}} , neg89 , {1{1'b0}} };

   // m89_69 = W*in
   wire signed [9:0] m89_69;
   assign m89_69 =10'b0;

   // m89_70 = W*in
   wire signed [9:0] m89_70;
   assign m89_70 =10'b0;

   // m89_71 = W*in
   wire signed [9:0] m89_71;
   assign m89_71 =10'b0;

   // m89_72 = W*in
   wire signed [9:0] m89_72;
   assign m89_72 =10'b0;

   // m89_73 = W*in
   wire signed [9:0] m89_73;
   assign m89_73 =10'b0;

   // m89_74 = W*in
   wire signed [9:0] m89_74;
   assign m89_74 =10'b0;

   // m89_75 = W*in
   wire signed [9:0] m89_75;
   assign m89_75 =10'b0;

   // m89_76 = W*in
   wire signed [9:0] m89_76;
   assign m89_76 =10'b0;

   // m89_77 = W*in
   wire signed [9:0] m89_77;
   assign m89_77 =10'b0;

   // m89_78 = W*in
   wire signed [9:0] m89_78;
   assign m89_78 ={ {3{in89[5]}} , in89 , {1{1'b0}} };

   // m89_79 = W*in
   wire signed [9:0] m89_79;
   assign m89_79 =10'b0;

   // m89_80 = W*in
   wire signed [9:0] m89_80;
   assign m89_80 =10'b0;

   // m89_81 = W*in
   wire signed [9:0] m89_81;
   assign m89_81 =10'b0;

   // m90_1 = W*in
   wire signed [9:0] m90_1;
   assign m90_1 =10'b0;

   // m90_2 = W*in
   wire signed [9:0] m90_2;
   assign m90_2 =10'b0;

   // m90_3 = W*in
   wire signed [9:0] m90_3;
   assign m90_3 =10'b0;

   // m90_4 = W*in
   wire signed [9:0] m90_4;
   assign m90_4 =10'b0;

   // m90_5 = W*in
   wire signed [9:0] m90_5;
   assign m90_5 =10'b0;

   // m90_6 = W*in
   wire signed [9:0] m90_6;
   assign m90_6 =10'b0;

   // m90_7 = W*in
   wire signed [9:0] m90_7;
   assign m90_7 =10'b0;

   // m90_8 = W*in
   wire signed [9:0] m90_8;
   assign m90_8 =10'b0;

   // m90_9 = W*in
   wire signed [9:0] m90_9;
   assign m90_9 =10'b0;

   // m90_10 = W*in
   wire signed [9:0] m90_10;
   assign m90_10 =10'b0;

   // m90_11 = W*in
   wire signed [9:0] m90_11;
   assign m90_11 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_12 = W*in
   wire signed [9:0] m90_12;
   assign m90_12 =10'b0;

   // m90_13 = W*in
   wire signed [9:0] m90_13;
   assign m90_13 =10'b0;

   // m90_14 = W*in
   wire signed [9:0] m90_14;
   assign m90_14 =10'b0;

   // m90_15 = W*in
   wire signed [9:0] m90_15;
   assign m90_15 =10'b0;

   // m90_16 = W*in
   wire signed [9:0] m90_16;
   assign m90_16 =10'b0;

   // m90_17 = W*in
   wire signed [9:0] m90_17;
   assign m90_17 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_18 = W*in
   wire signed [9:0] m90_18;
   assign m90_18 =10'b0;

   // m90_19 = W*in
   wire signed [9:0] m90_19;
   assign m90_19 =10'b0;

   // m90_20 = W*in
   wire signed [9:0] m90_20;
   assign m90_20 =10'b0;

   // m90_21 = W*in
   wire signed [9:0] m90_21;
   assign m90_21 =10'b0;

   // m90_22 = W*in
   wire signed [9:0] m90_22;
   assign m90_22 =10'b0;

   // m90_23 = W*in
   wire signed [9:0] m90_23;
   assign m90_23 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_24 = W*in
   wire signed [9:0] m90_24;
   assign m90_24 =10'b0;

   // m90_25 = W*in
   wire signed [9:0] m90_25;
   assign m90_25 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_26 = W*in
   wire signed [9:0] m90_26;
   assign m90_26 =10'b0;

   // m90_27 = W*in
   wire signed [9:0] m90_27;
   assign m90_27 =10'b0;

   // m90_28 = W*in
   wire signed [9:0] m90_28;
   assign m90_28 =10'b0;

   // m90_29 = W*in
   wire signed [9:0] m90_29;
   assign m90_29 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_30 = W*in
   wire signed [9:0] m90_30;
   assign m90_30 =10'b0;

   // m90_31 = W*in
   wire signed [9:0] m90_31;
   assign m90_31 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_32 = W*in
   wire signed [9:0] m90_32;
   assign m90_32 =10'b0;

   // m90_33 = W*in
   wire signed [9:0] m90_33;
   assign m90_33 =10'b0;

   // m90_34 = W*in
   wire signed [9:0] m90_34;
   assign m90_34 =10'b0;

   // m90_35 = W*in
   wire signed [9:0] m90_35;
   assign m90_35 =10'b0;

   // m90_36 = W*in
   wire signed [9:0] m90_36;
   assign m90_36 =10'b0;

   // m90_37 = W*in
   wire signed [9:0] m90_37;
   assign m90_37 =10'b0;

   // m90_38 = W*in
   wire signed [9:0] m90_38;
   assign m90_38 =10'b0;

   // m90_39 = W*in
   wire signed [9:0] m90_39;
   assign m90_39 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_40 = W*in
   wire signed [9:0] m90_40;
   assign m90_40 =10'b0;

   // m90_41 = W*in
   wire signed [9:0] m90_41;
   assign m90_41 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_42 = W*in
   wire signed [9:0] m90_42;
   assign m90_42 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_43 = W*in
   wire signed [9:0] m90_43;
   assign m90_43 =10'b0;

   // m90_44 = W*in
   wire signed [9:0] m90_44;
   assign m90_44 =10'b0;

   // m90_45 = W*in
   wire signed [9:0] m90_45;
   assign m90_45 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_46 = W*in
   wire signed [9:0] m90_46;
   assign m90_46 =10'b0;

   // m90_47 = W*in
   wire signed [9:0] m90_47;
   assign m90_47 =10'b0;

   // m90_48 = W*in
   wire signed [9:0] m90_48;
   assign m90_48 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_49 = W*in
   wire signed [9:0] m90_49;
   assign m90_49 ={ {2{in90[5]}} , in90 , {2{1'b0}} };

   // m90_50 = W*in
   wire signed [9:0] m90_50;
   assign m90_50 =10'b0;

   // m90_51 = W*in
   wire signed [9:0] m90_51;
   assign m90_51 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_52 = W*in
   wire signed [9:0] m90_52;
   assign m90_52 =10'b0;

   // m90_53 = W*in
   wire signed [9:0] m90_53;
   assign m90_53 =10'b0;

   // m90_54 = W*in
   wire signed [9:0] m90_54;
   assign m90_54 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_55 = W*in
   wire signed [9:0] m90_55;
   assign m90_55 ={ {2{in90[5]}} , in90 , {2{1'b0}} };

   // m90_56 = W*in
   wire signed [9:0] m90_56;
   assign m90_56 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_57 = W*in
   wire signed [9:0] m90_57;
   assign m90_57 =10'b0;

   // m90_58 = W*in
   wire signed [9:0] m90_58;
   assign m90_58 =10'b0;

   // m90_59 = W*in
   wire signed [9:0] m90_59;
   assign m90_59 =10'b0;

   // m90_60 = W*in
   wire signed [9:0] m90_60;
   assign m90_60 =10'b0;

   // m90_61 = W*in
   wire signed [9:0] m90_61;
   assign m90_61 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_62 = W*in
   wire signed [9:0] m90_62;
   assign m90_62 =10'b0;

   // m90_63 = W*in
   wire signed [9:0] m90_63;
   assign m90_63 ={ {3{neg90[5]}} , neg90 , {1{1'b0}} };

   // m90_64 = W*in
   wire signed [9:0] m90_64;
   assign m90_64 ={ {2{in90[5]}} , in90 , {2{1'b0}} };

   // m90_65 = W*in
   wire signed [9:0] m90_65;
   assign m90_65 =10'b0;

   // m90_66 = W*in
   wire signed [9:0] m90_66;
   assign m90_66 =10'b0;

   // m90_67 = W*in
   wire signed [9:0] m90_67;
   assign m90_67 ={ {2{in90[5]}} , in90 , {2{1'b0}} };

   // m90_68 = W*in
   wire signed [9:0] m90_68;
   assign m90_68 =10'b0;

   // m90_69 = W*in
   wire signed [9:0] m90_69;
   assign m90_69 =10'b0;

   // m90_70 = W*in
   wire signed [9:0] m90_70;
   assign m90_70 ={ {3{in90[5]}} , in90 , {1{1'b0}} };

   // m90_71 = W*in
   wire signed [9:0] m90_71;
   assign m90_71 =10'b0;

   // m90_72 = W*in
   wire signed [9:0] m90_72;
   assign m90_72 =10'b0;

   // m90_73 = W*in
   wire signed [9:0] m90_73;
   assign m90_73 =10'b0;

   // m90_74 = W*in
   wire signed [9:0] m90_74;
   assign m90_74 =10'b0;

   // m90_75 = W*in
   wire signed [9:0] m90_75;
   assign m90_75 ={ {2{in90[5]}} , in90 , {2{1'b0}} };

   // m90_76 = W*in
   wire signed [9:0] m90_76;
   assign m90_76 =10'b0;

   // m90_77 = W*in
   wire signed [9:0] m90_77;
   assign m90_77 =10'b0;

   // m90_78 = W*in
   wire signed [9:0] m90_78;
   assign m90_78 =10'b0;

   // m90_79 = W*in
   wire signed [9:0] m90_79;
   assign m90_79 =10'b0;

   // m90_80 = W*in
   wire signed [9:0] m90_80;
   assign m90_80 =10'b0;

   // m90_81 = W*in
   wire signed [9:0] m90_81;
   assign m90_81 =10'b0;

   // m91_1 = W*in
   wire signed [9:0] m91_1;
   assign m91_1 =10'b0;

   // m91_2 = W*in
   wire signed [9:0] m91_2;
   assign m91_2 =10'b0;

   // m91_3 = W*in
   wire signed [9:0] m91_3;
   assign m91_3 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_4 = W*in
   wire signed [9:0] m91_4;
   assign m91_4 =10'b0;

   // m91_5 = W*in
   wire signed [9:0] m91_5;
   assign m91_5 =10'b0;

   // m91_6 = W*in
   wire signed [9:0] m91_6;
   assign m91_6 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_7 = W*in
   wire signed [9:0] m91_7;
   assign m91_7 =10'b0;

   // m91_8 = W*in
   wire signed [9:0] m91_8;
   assign m91_8 =10'b0;

   // m91_9 = W*in
   wire signed [9:0] m91_9;
   assign m91_9 =10'b0;

   // m91_10 = W*in
   wire signed [9:0] m91_10;
   assign m91_10 =10'b0;

   // m91_11 = W*in
   wire signed [9:0] m91_11;
   assign m91_11 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_12 = W*in
   wire signed [9:0] m91_12;
   assign m91_12 =10'b0;

   // m91_13 = W*in
   wire signed [9:0] m91_13;
   assign m91_13 =10'b0;

   // m91_14 = W*in
   wire signed [9:0] m91_14;
   assign m91_14 =10'b0;

   // m91_15 = W*in
   wire signed [9:0] m91_15;
   assign m91_15 =10'b0;

   // m91_16 = W*in
   wire signed [9:0] m91_16;
   assign m91_16 =10'b0;

   // m91_17 = W*in
   wire signed [9:0] m91_17;
   assign m91_17 =10'b0;

   // m91_18 = W*in
   wire signed [9:0] m91_18;
   assign m91_18 =10'b0;

   // m91_19 = W*in
   wire signed [9:0] m91_19;
   assign m91_19 =10'b0;

   // m91_20 = W*in
   wire signed [9:0] m91_20;
   assign m91_20 =10'b0;

   // m91_21 = W*in
   wire signed [9:0] m91_21;
   assign m91_21 =10'b0;

   // m91_22 = W*in
   wire signed [9:0] m91_22;
   assign m91_22 =10'b0;

   // m91_23 = W*in
   wire signed [9:0] m91_23;
   assign m91_23 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_24 = W*in
   wire signed [9:0] m91_24;
   assign m91_24 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_25 = W*in
   wire signed [9:0] m91_25;
   assign m91_25 =10'b0;

   // m91_26 = W*in
   wire signed [9:0] m91_26;
   assign m91_26 =10'b0;

   // m91_27 = W*in
   wire signed [9:0] m91_27;
   assign m91_27 =10'b0;

   // m91_28 = W*in
   wire signed [9:0] m91_28;
   assign m91_28 =10'b0;

   // m91_29 = W*in
   wire signed [9:0] m91_29;
   assign m91_29 =10'b0;

   // m91_30 = W*in
   wire signed [9:0] m91_30;
   assign m91_30 =10'b0;

   // m91_31 = W*in
   wire signed [9:0] m91_31;
   assign m91_31 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_32 = W*in
   wire signed [9:0] m91_32;
   assign m91_32 =10'b0;

   // m91_33 = W*in
   wire signed [9:0] m91_33;
   assign m91_33 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_34 = W*in
   wire signed [9:0] m91_34;
   assign m91_34 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_35 = W*in
   wire signed [9:0] m91_35;
   assign m91_35 =10'b0;

   // m91_36 = W*in
   wire signed [9:0] m91_36;
   assign m91_36 =10'b0;

   // m91_37 = W*in
   wire signed [9:0] m91_37;
   assign m91_37 =10'b0;

   // m91_38 = W*in
   wire signed [9:0] m91_38;
   assign m91_38 =10'b0;

   // m91_39 = W*in
   wire signed [9:0] m91_39;
   assign m91_39 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_40 = W*in
   wire signed [9:0] m91_40;
   assign m91_40 =10'b0;

   // m91_41 = W*in
   wire signed [9:0] m91_41;
   assign m91_41 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_42 = W*in
   wire signed [9:0] m91_42;
   assign m91_42 =10'b0;

   // m91_43 = W*in
   wire signed [9:0] m91_43;
   assign m91_43 =10'b0;

   // m91_44 = W*in
   wire signed [9:0] m91_44;
   assign m91_44 =10'b0;

   // m91_45 = W*in
   wire signed [9:0] m91_45;
   assign m91_45 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_46 = W*in
   wire signed [9:0] m91_46;
   assign m91_46 =10'b0;

   // m91_47 = W*in
   wire signed [9:0] m91_47;
   assign m91_47 =10'b0;

   // m91_48 = W*in
   wire signed [9:0] m91_48;
   assign m91_48 =10'b0;

   // m91_49 = W*in
   wire signed [9:0] m91_49;
   assign m91_49 =10'b0;

   // m91_50 = W*in
   wire signed [9:0] m91_50;
   assign m91_50 =10'b0;

   // m91_51 = W*in
   wire signed [9:0] m91_51;
   assign m91_51 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_52 = W*in
   wire signed [9:0] m91_52;
   assign m91_52 =10'b0;

   // m91_53 = W*in
   wire signed [9:0] m91_53;
   assign m91_53 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_54 = W*in
   wire signed [9:0] m91_54;
   assign m91_54 =10'b0;

   // m91_55 = W*in
   wire signed [9:0] m91_55;
   assign m91_55 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_56 = W*in
   wire signed [9:0] m91_56;
   assign m91_56 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_57 = W*in
   wire signed [9:0] m91_57;
   assign m91_57 =10'b0;

   // m91_58 = W*in
   wire signed [9:0] m91_58;
   assign m91_58 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_59 = W*in
   wire signed [9:0] m91_59;
   assign m91_59 =10'b0;

   // m91_60 = W*in
   wire signed [9:0] m91_60;
   assign m91_60 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_61 = W*in
   wire signed [9:0] m91_61;
   assign m91_61 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_62 = W*in
   wire signed [9:0] m91_62;
   assign m91_62 =10'b0;

   // m91_63 = W*in
   wire signed [9:0] m91_63;
   assign m91_63 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_64 = W*in
   wire signed [9:0] m91_64;
   assign m91_64 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_65 = W*in
   wire signed [9:0] m91_65;
   assign m91_65 =10'b0;

   // m91_66 = W*in
   wire signed [9:0] m91_66;
   assign m91_66 =10'b0;

   // m91_67 = W*in
   wire signed [9:0] m91_67;
   assign m91_67 =10'b0;

   // m91_68 = W*in
   wire signed [9:0] m91_68;
   assign m91_68 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_69 = W*in
   wire signed [9:0] m91_69;
   assign m91_69 ={ {2{in91[5]}} , in91 , {2{1'b0}} };

   // m91_70 = W*in
   wire signed [9:0] m91_70;
   assign m91_70 =10'b0;

   // m91_71 = W*in
   wire signed [9:0] m91_71;
   assign m91_71 =10'b0;

   // m91_72 = W*in
   wire signed [9:0] m91_72;
   assign m91_72 =10'b0;

   // m91_73 = W*in
   wire signed [9:0] m91_73;
   assign m91_73 =10'b0;

   // m91_74 = W*in
   wire signed [9:0] m91_74;
   assign m91_74 =10'b0;

   // m91_75 = W*in
   wire signed [9:0] m91_75;
   assign m91_75 =10'b0;

   // m91_76 = W*in
   wire signed [9:0] m91_76;
   assign m91_76 =10'b0;

   // m91_77 = W*in
   wire signed [9:0] m91_77;
   assign m91_77 ={ {3{in91[5]}} , in91 , {1{1'b0}} };

   // m91_78 = W*in
   wire signed [9:0] m91_78;
   assign m91_78 ={ {3{neg91[5]}} , neg91 , {1{1'b0}} };

   // m91_79 = W*in
   wire signed [9:0] m91_79;
   assign m91_79 =10'b0;

   // m91_80 = W*in
   wire signed [9:0] m91_80;
   assign m91_80 =10'b0;

   // m91_81 = W*in
   wire signed [9:0] m91_81;
   assign m91_81 =10'b0;

   // m92_1 = W*in
   wire signed [9:0] m92_1;
   assign m92_1 =10'b0;

   // m92_2 = W*in
   wire signed [9:0] m92_2;
   assign m92_2 =10'b0;

   // m92_3 = W*in
   wire signed [9:0] m92_3;
   assign m92_3 =10'b0;

   // m92_4 = W*in
   wire signed [9:0] m92_4;
   assign m92_4 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_5 = W*in
   wire signed [9:0] m92_5;
   assign m92_5 =10'b0;

   // m92_6 = W*in
   wire signed [9:0] m92_6;
   assign m92_6 =10'b0;

   // m92_7 = W*in
   wire signed [9:0] m92_7;
   assign m92_7 =10'b0;

   // m92_8 = W*in
   wire signed [9:0] m92_8;
   assign m92_8 =10'b0;

   // m92_9 = W*in
   wire signed [9:0] m92_9;
   assign m92_9 =10'b0;

   // m92_10 = W*in
   wire signed [9:0] m92_10;
   assign m92_10 =10'b0;

   // m92_11 = W*in
   wire signed [9:0] m92_11;
   assign m92_11 =10'b0;

   // m92_12 = W*in
   wire signed [9:0] m92_12;
   assign m92_12 =10'b0;

   // m92_13 = W*in
   wire signed [9:0] m92_13;
   assign m92_13 =10'b0;

   // m92_14 = W*in
   wire signed [9:0] m92_14;
   assign m92_14 ={ {3{neg92[5]}} , neg92 , {1{1'b0}} };

   // m92_15 = W*in
   wire signed [9:0] m92_15;
   assign m92_15 =10'b0;

   // m92_16 = W*in
   wire signed [9:0] m92_16;
   assign m92_16 =10'b0;

   // m92_17 = W*in
   wire signed [9:0] m92_17;
   assign m92_17 =10'b0;

   // m92_18 = W*in
   wire signed [9:0] m92_18;
   assign m92_18 =10'b0;

   // m92_19 = W*in
   wire signed [9:0] m92_19;
   assign m92_19 =10'b0;

   // m92_20 = W*in
   wire signed [9:0] m92_20;
   assign m92_20 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_21 = W*in
   wire signed [9:0] m92_21;
   assign m92_21 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_22 = W*in
   wire signed [9:0] m92_22;
   assign m92_22 =10'b0;

   // m92_23 = W*in
   wire signed [9:0] m92_23;
   assign m92_23 =10'b0;

   // m92_24 = W*in
   wire signed [9:0] m92_24;
   assign m92_24 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_25 = W*in
   wire signed [9:0] m92_25;
   assign m92_25 =10'b0;

   // m92_26 = W*in
   wire signed [9:0] m92_26;
   assign m92_26 =10'b0;

   // m92_27 = W*in
   wire signed [9:0] m92_27;
   assign m92_27 =10'b0;

   // m92_28 = W*in
   wire signed [9:0] m92_28;
   assign m92_28 =10'b0;

   // m92_29 = W*in
   wire signed [9:0] m92_29;
   assign m92_29 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_30 = W*in
   wire signed [9:0] m92_30;
   assign m92_30 =10'b0;

   // m92_31 = W*in
   wire signed [9:0] m92_31;
   assign m92_31 ={ {3{neg92[5]}} , neg92 , {1{1'b0}} };

   // m92_32 = W*in
   wire signed [9:0] m92_32;
   assign m92_32 =10'b0;

   // m92_33 = W*in
   wire signed [9:0] m92_33;
   assign m92_33 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_34 = W*in
   wire signed [9:0] m92_34;
   assign m92_34 =10'b0;

   // m92_35 = W*in
   wire signed [9:0] m92_35;
   assign m92_35 ={ {3{neg92[5]}} , neg92 , {1{1'b0}} };

   // m92_36 = W*in
   wire signed [9:0] m92_36;
   assign m92_36 =10'b0;

   // m92_37 = W*in
   wire signed [9:0] m92_37;
   assign m92_37 =10'b0;

   // m92_38 = W*in
   wire signed [9:0] m92_38;
   assign m92_38 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_39 = W*in
   wire signed [9:0] m92_39;
   assign m92_39 =10'b0;

   // m92_40 = W*in
   wire signed [9:0] m92_40;
   assign m92_40 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_41 = W*in
   wire signed [9:0] m92_41;
   assign m92_41 =10'b0;

   // m92_42 = W*in
   wire signed [9:0] m92_42;
   assign m92_42 =10'b0;

   // m92_43 = W*in
   wire signed [9:0] m92_43;
   assign m92_43 ={ {3{neg92[5]}} , neg92 , {1{1'b0}} };

   // m92_44 = W*in
   wire signed [9:0] m92_44;
   assign m92_44 =10'b0;

   // m92_45 = W*in
   wire signed [9:0] m92_45;
   assign m92_45 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_46 = W*in
   wire signed [9:0] m92_46;
   assign m92_46 =10'b0;

   // m92_47 = W*in
   wire signed [9:0] m92_47;
   assign m92_47 =10'b0;

   // m92_48 = W*in
   wire signed [9:0] m92_48;
   assign m92_48 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_49 = W*in
   wire signed [9:0] m92_49;
   assign m92_49 =10'b0;

   // m92_50 = W*in
   wire signed [9:0] m92_50;
   assign m92_50 =10'b0;

   // m92_51 = W*in
   wire signed [9:0] m92_51;
   assign m92_51 =10'b0;

   // m92_52 = W*in
   wire signed [9:0] m92_52;
   assign m92_52 =10'b0;

   // m92_53 = W*in
   wire signed [9:0] m92_53;
   assign m92_53 =10'b0;

   // m92_54 = W*in
   wire signed [9:0] m92_54;
   assign m92_54 =10'b0;

   // m92_55 = W*in
   wire signed [9:0] m92_55;
   assign m92_55 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_56 = W*in
   wire signed [9:0] m92_56;
   assign m92_56 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_57 = W*in
   wire signed [9:0] m92_57;
   assign m92_57 =10'b0;

   // m92_58 = W*in
   wire signed [9:0] m92_58;
   assign m92_58 =10'b0;

   // m92_59 = W*in
   wire signed [9:0] m92_59;
   assign m92_59 =10'b0;

   // m92_60 = W*in
   wire signed [9:0] m92_60;
   assign m92_60 =10'b0;

   // m92_61 = W*in
   wire signed [9:0] m92_61;
   assign m92_61 ={ {3{neg92[5]}} , neg92 , {1{1'b0}} };

   // m92_62 = W*in
   wire signed [9:0] m92_62;
   assign m92_62 =10'b0;

   // m92_63 = W*in
   wire signed [9:0] m92_63;
   assign m92_63 =10'b0;

   // m92_64 = W*in
   wire signed [9:0] m92_64;
   assign m92_64 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_65 = W*in
   wire signed [9:0] m92_65;
   assign m92_65 =10'b0;

   // m92_66 = W*in
   wire signed [9:0] m92_66;
   assign m92_66 =10'b0;

   // m92_67 = W*in
   wire signed [9:0] m92_67;
   assign m92_67 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_68 = W*in
   wire signed [9:0] m92_68;
   assign m92_68 ={ {3{in92[5]}} , in92 , {1{1'b0}} };

   // m92_69 = W*in
   wire signed [9:0] m92_69;
   assign m92_69 =10'b0;

   // m92_70 = W*in
   wire signed [9:0] m92_70;
   assign m92_70 =10'b0;

   // m92_71 = W*in
   wire signed [9:0] m92_71;
   assign m92_71 =10'b0;

   // m92_72 = W*in
   wire signed [9:0] m92_72;
   assign m92_72 =10'b0;

   // m92_73 = W*in
   wire signed [9:0] m92_73;
   assign m92_73 =10'b0;

   // m92_74 = W*in
   wire signed [9:0] m92_74;
   assign m92_74 ={ {2{in92[5]}} , in92 , {2{1'b0}} };

   // m92_75 = W*in
   wire signed [9:0] m92_75;
   assign m92_75 ={ {2{in92[5]}} , in92 , {2{1'b0}} };

   // m92_76 = W*in
   wire signed [9:0] m92_76;
   assign m92_76 =10'b0;

   // m92_77 = W*in
   wire signed [9:0] m92_77;
   assign m92_77 =10'b0;

   // m92_78 = W*in
   wire signed [9:0] m92_78;
   assign m92_78 =10'b0;

   // m92_79 = W*in
   wire signed [9:0] m92_79;
   assign m92_79 =10'b0;

   // m92_80 = W*in
   wire signed [9:0] m92_80;
   assign m92_80 =10'b0;

   // m92_81 = W*in
   wire signed [9:0] m92_81;
   assign m92_81 =10'b0;

   // m93_1 = W*in
   wire signed [9:0] m93_1;
   assign m93_1 =10'b0;

   // m93_2 = W*in
   wire signed [9:0] m93_2;
   assign m93_2 =10'b0;

   // m93_3 = W*in
   wire signed [9:0] m93_3;
   assign m93_3 =10'b0;

   // m93_4 = W*in
   wire signed [9:0] m93_4;
   assign m93_4 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_5 = W*in
   wire signed [9:0] m93_5;
   assign m93_5 =10'b0;

   // m93_6 = W*in
   wire signed [9:0] m93_6;
   assign m93_6 =10'b0;

   // m93_7 = W*in
   wire signed [9:0] m93_7;
   assign m93_7 =10'b0;

   // m93_8 = W*in
   wire signed [9:0] m93_8;
   assign m93_8 =10'b0;

   // m93_9 = W*in
   wire signed [9:0] m93_9;
   assign m93_9 =10'b0;

   // m93_10 = W*in
   wire signed [9:0] m93_10;
   assign m93_10 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_11 = W*in
   wire signed [9:0] m93_11;
   assign m93_11 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_12 = W*in
   wire signed [9:0] m93_12;
   assign m93_12 =10'b0;

   // m93_13 = W*in
   wire signed [9:0] m93_13;
   assign m93_13 =10'b0;

   // m93_14 = W*in
   wire signed [9:0] m93_14;
   assign m93_14 =10'b0;

   // m93_15 = W*in
   wire signed [9:0] m93_15;
   assign m93_15 =10'b0;

   // m93_16 = W*in
   wire signed [9:0] m93_16;
   assign m93_16 =10'b0;

   // m93_17 = W*in
   wire signed [9:0] m93_17;
   assign m93_17 =10'b0;

   // m93_18 = W*in
   wire signed [9:0] m93_18;
   assign m93_18 =10'b0;

   // m93_19 = W*in
   wire signed [9:0] m93_19;
   assign m93_19 =10'b0;

   // m93_20 = W*in
   wire signed [9:0] m93_20;
   assign m93_20 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_21 = W*in
   wire signed [9:0] m93_21;
   assign m93_21 =10'b0;

   // m93_22 = W*in
   wire signed [9:0] m93_22;
   assign m93_22 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_23 = W*in
   wire signed [9:0] m93_23;
   assign m93_23 =10'b0;

   // m93_24 = W*in
   wire signed [9:0] m93_24;
   assign m93_24 =10'b0;

   // m93_25 = W*in
   wire signed [9:0] m93_25;
   assign m93_25 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_26 = W*in
   wire signed [9:0] m93_26;
   assign m93_26 =10'b0;

   // m93_27 = W*in
   wire signed [9:0] m93_27;
   assign m93_27 =10'b0;

   // m93_28 = W*in
   wire signed [9:0] m93_28;
   assign m93_28 =10'b0;

   // m93_29 = W*in
   wire signed [9:0] m93_29;
   assign m93_29 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_30 = W*in
   wire signed [9:0] m93_30;
   assign m93_30 =10'b0;

   // m93_31 = W*in
   wire signed [9:0] m93_31;
   assign m93_31 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_32 = W*in
   wire signed [9:0] m93_32;
   assign m93_32 =10'b0;

   // m93_33 = W*in
   wire signed [9:0] m93_33;
   assign m93_33 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_34 = W*in
   wire signed [9:0] m93_34;
   assign m93_34 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_35 = W*in
   wire signed [9:0] m93_35;
   assign m93_35 =10'b0;

   // m93_36 = W*in
   wire signed [9:0] m93_36;
   assign m93_36 =10'b0;

   // m93_37 = W*in
   wire signed [9:0] m93_37;
   assign m93_37 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_38 = W*in
   wire signed [9:0] m93_38;
   assign m93_38 =10'b0;

   // m93_39 = W*in
   wire signed [9:0] m93_39;
   assign m93_39 =10'b0;

   // m93_40 = W*in
   wire signed [9:0] m93_40;
   assign m93_40 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_41 = W*in
   wire signed [9:0] m93_41;
   assign m93_41 =10'b0;

   // m93_42 = W*in
   wire signed [9:0] m93_42;
   assign m93_42 =10'b0;

   // m93_43 = W*in
   wire signed [9:0] m93_43;
   assign m93_43 =10'b0;

   // m93_44 = W*in
   wire signed [9:0] m93_44;
   assign m93_44 =10'b0;

   // m93_45 = W*in
   wire signed [9:0] m93_45;
   assign m93_45 =10'b0;

   // m93_46 = W*in
   wire signed [9:0] m93_46;
   assign m93_46 =10'b0;

   // m93_47 = W*in
   wire signed [9:0] m93_47;
   assign m93_47 =10'b0;

   // m93_48 = W*in
   wire signed [9:0] m93_48;
   assign m93_48 =10'b0;

   // m93_49 = W*in
   wire signed [9:0] m93_49;
   assign m93_49 =10'b0;

   // m93_50 = W*in
   wire signed [9:0] m93_50;
   assign m93_50 =10'b0;

   // m93_51 = W*in
   wire signed [9:0] m93_51;
   assign m93_51 =10'b0;

   // m93_52 = W*in
   wire signed [9:0] m93_52;
   assign m93_52 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_53 = W*in
   wire signed [9:0] m93_53;
   assign m93_53 =10'b0;

   // m93_54 = W*in
   wire signed [9:0] m93_54;
   assign m93_54 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_55 = W*in
   wire signed [9:0] m93_55;
   assign m93_55 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_56 = W*in
   wire signed [9:0] m93_56;
   assign m93_56 =10'b0;

   // m93_57 = W*in
   wire signed [9:0] m93_57;
   assign m93_57 =10'b0;

   // m93_58 = W*in
   wire signed [9:0] m93_58;
   assign m93_58 =10'b0;

   // m93_59 = W*in
   wire signed [9:0] m93_59;
   assign m93_59 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_60 = W*in
   wire signed [9:0] m93_60;
   assign m93_60 =10'b0;

   // m93_61 = W*in
   wire signed [9:0] m93_61;
   assign m93_61 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_62 = W*in
   wire signed [9:0] m93_62;
   assign m93_62 =10'b0;

   // m93_63 = W*in
   wire signed [9:0] m93_63;
   assign m93_63 =10'b0;

   // m93_64 = W*in
   wire signed [9:0] m93_64;
   assign m93_64 =10'b0;

   // m93_65 = W*in
   wire signed [9:0] m93_65;
   assign m93_65 =10'b0;

   // m93_66 = W*in
   wire signed [9:0] m93_66;
   assign m93_66 =10'b0;

   // m93_67 = W*in
   wire signed [9:0] m93_67;
   assign m93_67 =10'b0;

   // m93_68 = W*in
   wire signed [9:0] m93_68;
   assign m93_68 =10'b0;

   // m93_69 = W*in
   wire signed [9:0] m93_69;
   assign m93_69 =10'b0;

   // m93_70 = W*in
   wire signed [9:0] m93_70;
   assign m93_70 =10'b0;

   // m93_71 = W*in
   wire signed [9:0] m93_71;
   assign m93_71 =10'b0;

   // m93_72 = W*in
   wire signed [9:0] m93_72;
   assign m93_72 =10'b0;

   // m93_73 = W*in
   wire signed [9:0] m93_73;
   assign m93_73 =10'b0;

   // m93_74 = W*in
   wire signed [9:0] m93_74;
   assign m93_74 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_75 = W*in
   wire signed [9:0] m93_75;
   assign m93_75 =10'b0;

   // m93_76 = W*in
   wire signed [9:0] m93_76;
   assign m93_76 ={ {2{in93[5]}} , in93 , {2{1'b0}} };

   // m93_77 = W*in
   wire signed [9:0] m93_77;
   assign m93_77 ={ {3{in93[5]}} , in93 , {1{1'b0}} };

   // m93_78 = W*in
   wire signed [9:0] m93_78;
   assign m93_78 =10'b0;

   // m93_79 = W*in
   wire signed [9:0] m93_79;
   assign m93_79 ={ {3{neg93[5]}} , neg93 , {1{1'b0}} };

   // m93_80 = W*in
   wire signed [9:0] m93_80;
   assign m93_80 =10'b0;

   // m93_81 = W*in
   wire signed [9:0] m93_81;
   assign m93_81 =10'b0;

   // m94_1 = W*in
   wire signed [9:0] m94_1;
   assign m94_1 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_2 = W*in
   wire signed [9:0] m94_2;
   assign m94_2 =10'b0;

   // m94_3 = W*in
   wire signed [9:0] m94_3;
   assign m94_3 ={ {3{in94[5]}} , in94 , {1{1'b0}} };

   // m94_4 = W*in
   wire signed [9:0] m94_4;
   assign m94_4 =10'b0;

   // m94_5 = W*in
   wire signed [9:0] m94_5;
   assign m94_5 =10'b0;

   // m94_6 = W*in
   wire signed [9:0] m94_6;
   assign m94_6 =10'b0;

   // m94_7 = W*in
   wire signed [9:0] m94_7;
   assign m94_7 =10'b0;

   // m94_8 = W*in
   wire signed [9:0] m94_8;
   assign m94_8 =10'b0;

   // m94_9 = W*in
   wire signed [9:0] m94_9;
   assign m94_9 ={ {3{in94[5]}} , in94 , {1{1'b0}} };

   // m94_10 = W*in
   wire signed [9:0] m94_10;
   assign m94_10 =10'b0;

   // m94_11 = W*in
   wire signed [9:0] m94_11;
   assign m94_11 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_12 = W*in
   wire signed [9:0] m94_12;
   assign m94_12 =10'b0;

   // m94_13 = W*in
   wire signed [9:0] m94_13;
   assign m94_13 =10'b0;

   // m94_14 = W*in
   wire signed [9:0] m94_14;
   assign m94_14 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_15 = W*in
   wire signed [9:0] m94_15;
   assign m94_15 =10'b0;

   // m94_16 = W*in
   wire signed [9:0] m94_16;
   assign m94_16 =10'b0;

   // m94_17 = W*in
   wire signed [9:0] m94_17;
   assign m94_17 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_18 = W*in
   wire signed [9:0] m94_18;
   assign m94_18 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_19 = W*in
   wire signed [9:0] m94_19;
   assign m94_19 ={ {3{in94[5]}} , in94 , {1{1'b0}} };

   // m94_20 = W*in
   wire signed [9:0] m94_20;
   assign m94_20 =10'b0;

   // m94_21 = W*in
   wire signed [9:0] m94_21;
   assign m94_21 =10'b0;

   // m94_22 = W*in
   wire signed [9:0] m94_22;
   assign m94_22 ={ {3{in94[5]}} , in94 , {1{1'b0}} };

   // m94_23 = W*in
   wire signed [9:0] m94_23;
   assign m94_23 =10'b0;

   // m94_24 = W*in
   wire signed [9:0] m94_24;
   assign m94_24 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_25 = W*in
   wire signed [9:0] m94_25;
   assign m94_25 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_26 = W*in
   wire signed [9:0] m94_26;
   assign m94_26 =10'b0;

   // m94_27 = W*in
   wire signed [9:0] m94_27;
   assign m94_27 =10'b0;

   // m94_28 = W*in
   wire signed [9:0] m94_28;
   assign m94_28 =10'b0;

   // m94_29 = W*in
   wire signed [9:0] m94_29;
   assign m94_29 =10'b0;

   // m94_30 = W*in
   wire signed [9:0] m94_30;
   assign m94_30 =10'b0;

   // m94_31 = W*in
   wire signed [9:0] m94_31;
   assign m94_31 ={ {3{in94[5]}} , in94 , {1{1'b0}} };

   // m94_32 = W*in
   wire signed [9:0] m94_32;
   assign m94_32 =10'b0;

   // m94_33 = W*in
   wire signed [9:0] m94_33;
   assign m94_33 =10'b0;

   // m94_34 = W*in
   wire signed [9:0] m94_34;
   assign m94_34 =10'b0;

   // m94_35 = W*in
   wire signed [9:0] m94_35;
   assign m94_35 =10'b0;

   // m94_36 = W*in
   wire signed [9:0] m94_36;
   assign m94_36 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_37 = W*in
   wire signed [9:0] m94_37;
   assign m94_37 =10'b0;

   // m94_38 = W*in
   wire signed [9:0] m94_38;
   assign m94_38 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_39 = W*in
   wire signed [9:0] m94_39;
   assign m94_39 =10'b0;

   // m94_40 = W*in
   wire signed [9:0] m94_40;
   assign m94_40 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_41 = W*in
   wire signed [9:0] m94_41;
   assign m94_41 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_42 = W*in
   wire signed [9:0] m94_42;
   assign m94_42 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_43 = W*in
   wire signed [9:0] m94_43;
   assign m94_43 =10'b0;

   // m94_44 = W*in
   wire signed [9:0] m94_44;
   assign m94_44 =10'b0;

   // m94_45 = W*in
   wire signed [9:0] m94_45;
   assign m94_45 =10'b0;

   // m94_46 = W*in
   wire signed [9:0] m94_46;
   assign m94_46 =10'b0;

   // m94_47 = W*in
   wire signed [9:0] m94_47;
   assign m94_47 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_48 = W*in
   wire signed [9:0] m94_48;
   assign m94_48 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_49 = W*in
   wire signed [9:0] m94_49;
   assign m94_49 =10'b0;

   // m94_50 = W*in
   wire signed [9:0] m94_50;
   assign m94_50 ={ {2{in94[5]}} , in94 , {2{1'b0}} };

   // m94_51 = W*in
   wire signed [9:0] m94_51;
   assign m94_51 =10'b0;

   // m94_52 = W*in
   wire signed [9:0] m94_52;
   assign m94_52 =10'b0;

   // m94_53 = W*in
   wire signed [9:0] m94_53;
   assign m94_53 =10'b0;

   // m94_54 = W*in
   wire signed [9:0] m94_54;
   assign m94_54 =10'b0;

   // m94_55 = W*in
   wire signed [9:0] m94_55;
   assign m94_55 =10'b0;

   // m94_56 = W*in
   wire signed [9:0] m94_56;
   assign m94_56 =10'b0;

   // m94_57 = W*in
   wire signed [9:0] m94_57;
   assign m94_57 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_58 = W*in
   wire signed [9:0] m94_58;
   assign m94_58 =10'b0;

   // m94_59 = W*in
   wire signed [9:0] m94_59;
   assign m94_59 =10'b0;

   // m94_60 = W*in
   wire signed [9:0] m94_60;
   assign m94_60 =10'b0;

   // m94_61 = W*in
   wire signed [9:0] m94_61;
   assign m94_61 ={ {3{in94[5]}} , in94 , {1{1'b0}} };

   // m94_62 = W*in
   wire signed [9:0] m94_62;
   assign m94_62 =10'b0;

   // m94_63 = W*in
   wire signed [9:0] m94_63;
   assign m94_63 =10'b0;

   // m94_64 = W*in
   wire signed [9:0] m94_64;
   assign m94_64 =10'b0;

   // m94_65 = W*in
   wire signed [9:0] m94_65;
   assign m94_65 =10'b0;

   // m94_66 = W*in
   wire signed [9:0] m94_66;
   assign m94_66 =10'b0;

   // m94_67 = W*in
   wire signed [9:0] m94_67;
   assign m94_67 =10'b0;

   // m94_68 = W*in
   wire signed [9:0] m94_68;
   assign m94_68 =10'b0;

   // m94_69 = W*in
   wire signed [9:0] m94_69;
   assign m94_69 ={ {3{neg94[5]}} , neg94 , {1{1'b0}} };

   // m94_70 = W*in
   wire signed [9:0] m94_70;
   assign m94_70 =10'b0;

   // m94_71 = W*in
   wire signed [9:0] m94_71;
   assign m94_71 =10'b0;

   // m94_72 = W*in
   wire signed [9:0] m94_72;
   assign m94_72 =10'b0;

   // m94_73 = W*in
   wire signed [9:0] m94_73;
   assign m94_73 =10'b0;

   // m94_74 = W*in
   wire signed [9:0] m94_74;
   assign m94_74 =10'b0;

   // m94_75 = W*in
   wire signed [9:0] m94_75;
   assign m94_75 =10'b0;

   // m94_76 = W*in
   wire signed [9:0] m94_76;
   assign m94_76 =10'b0;

   // m94_77 = W*in
   wire signed [9:0] m94_77;
   assign m94_77 =10'b0;

   // m94_78 = W*in
   wire signed [9:0] m94_78;
   assign m94_78 =10'b0;

   // m94_79 = W*in
   wire signed [9:0] m94_79;
   assign m94_79 =10'b0;

   // m94_80 = W*in
   wire signed [9:0] m94_80;
   assign m94_80 =10'b0;

   // m94_81 = W*in
   wire signed [9:0] m94_81;
   assign m94_81 =10'b0;

   // m95_1 = W*in
   wire signed [9:0] m95_1;
   assign m95_1 =10'b0;

   // m95_2 = W*in
   wire signed [9:0] m95_2;
   assign m95_2 =10'b0;

   // m95_3 = W*in
   wire signed [9:0] m95_3;
   assign m95_3 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_4 = W*in
   wire signed [9:0] m95_4;
   assign m95_4 =10'b0;

   // m95_5 = W*in
   wire signed [9:0] m95_5;
   assign m95_5 =10'b0;

   // m95_6 = W*in
   wire signed [9:0] m95_6;
   assign m95_6 =10'b0;

   // m95_7 = W*in
   wire signed [9:0] m95_7;
   assign m95_7 =10'b0;

   // m95_8 = W*in
   wire signed [9:0] m95_8;
   assign m95_8 =10'b0;

   // m95_9 = W*in
   wire signed [9:0] m95_9;
   assign m95_9 =10'b0;

   // m95_10 = W*in
   wire signed [9:0] m95_10;
   assign m95_10 =10'b0;

   // m95_11 = W*in
   wire signed [9:0] m95_11;
   assign m95_11 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_12 = W*in
   wire signed [9:0] m95_12;
   assign m95_12 =10'b0;

   // m95_13 = W*in
   wire signed [9:0] m95_13;
   assign m95_13 =10'b0;

   // m95_14 = W*in
   wire signed [9:0] m95_14;
   assign m95_14 =10'b0;

   // m95_15 = W*in
   wire signed [9:0] m95_15;
   assign m95_15 ={ {2{in95[5]}} , in95 , {2{1'b0}} };

   // m95_16 = W*in
   wire signed [9:0] m95_16;
   assign m95_16 =10'b0;

   // m95_17 = W*in
   wire signed [9:0] m95_17;
   assign m95_17 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_18 = W*in
   wire signed [9:0] m95_18;
   assign m95_18 =10'b0;

   // m95_19 = W*in
   wire signed [9:0] m95_19;
   assign m95_19 =10'b0;

   // m95_20 = W*in
   wire signed [9:0] m95_20;
   assign m95_20 =10'b0;

   // m95_21 = W*in
   wire signed [9:0] m95_21;
   assign m95_21 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_22 = W*in
   wire signed [9:0] m95_22;
   assign m95_22 =10'b0;

   // m95_23 = W*in
   wire signed [9:0] m95_23;
   assign m95_23 =10'b0;

   // m95_24 = W*in
   wire signed [9:0] m95_24;
   assign m95_24 =10'b0;

   // m95_25 = W*in
   wire signed [9:0] m95_25;
   assign m95_25 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_26 = W*in
   wire signed [9:0] m95_26;
   assign m95_26 =10'b0;

   // m95_27 = W*in
   wire signed [9:0] m95_27;
   assign m95_27 =10'b0;

   // m95_28 = W*in
   wire signed [9:0] m95_28;
   assign m95_28 =10'b0;

   // m95_29 = W*in
   wire signed [9:0] m95_29;
   assign m95_29 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_30 = W*in
   wire signed [9:0] m95_30;
   assign m95_30 =10'b0;

   // m95_31 = W*in
   wire signed [9:0] m95_31;
   assign m95_31 =10'b0;

   // m95_32 = W*in
   wire signed [9:0] m95_32;
   assign m95_32 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_33 = W*in
   wire signed [9:0] m95_33;
   assign m95_33 =10'b0;

   // m95_34 = W*in
   wire signed [9:0] m95_34;
   assign m95_34 =10'b0;

   // m95_35 = W*in
   wire signed [9:0] m95_35;
   assign m95_35 =10'b0;

   // m95_36 = W*in
   wire signed [9:0] m95_36;
   assign m95_36 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_37 = W*in
   wire signed [9:0] m95_37;
   assign m95_37 =10'b0;

   // m95_38 = W*in
   wire signed [9:0] m95_38;
   assign m95_38 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_39 = W*in
   wire signed [9:0] m95_39;
   assign m95_39 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_40 = W*in
   wire signed [9:0] m95_40;
   assign m95_40 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_41 = W*in
   wire signed [9:0] m95_41;
   assign m95_41 =10'b0;

   // m95_42 = W*in
   wire signed [9:0] m95_42;
   assign m95_42 =10'b0;

   // m95_43 = W*in
   wire signed [9:0] m95_43;
   assign m95_43 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_44 = W*in
   wire signed [9:0] m95_44;
   assign m95_44 =10'b0;

   // m95_45 = W*in
   wire signed [9:0] m95_45;
   assign m95_45 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_46 = W*in
   wire signed [9:0] m95_46;
   assign m95_46 =10'b0;

   // m95_47 = W*in
   wire signed [9:0] m95_47;
   assign m95_47 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_48 = W*in
   wire signed [9:0] m95_48;
   assign m95_48 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_49 = W*in
   wire signed [9:0] m95_49;
   assign m95_49 =10'b0;

   // m95_50 = W*in
   wire signed [9:0] m95_50;
   assign m95_50 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_51 = W*in
   wire signed [9:0] m95_51;
   assign m95_51 =10'b0;

   // m95_52 = W*in
   wire signed [9:0] m95_52;
   assign m95_52 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_53 = W*in
   wire signed [9:0] m95_53;
   assign m95_53 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_54 = W*in
   wire signed [9:0] m95_54;
   assign m95_54 ={ {2{in95[5]}} , in95 , {2{1'b0}} };

   // m95_55 = W*in
   wire signed [9:0] m95_55;
   assign m95_55 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_56 = W*in
   wire signed [9:0] m95_56;
   assign m95_56 =10'b0;

   // m95_57 = W*in
   wire signed [9:0] m95_57;
   assign m95_57 ={ {2{in95[5]}} , in95 , {2{1'b0}} };

   // m95_58 = W*in
   wire signed [9:0] m95_58;
   assign m95_58 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_59 = W*in
   wire signed [9:0] m95_59;
   assign m95_59 =10'b0;

   // m95_60 = W*in
   wire signed [9:0] m95_60;
   assign m95_60 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_61 = W*in
   wire signed [9:0] m95_61;
   assign m95_61 =10'b0;

   // m95_62 = W*in
   wire signed [9:0] m95_62;
   assign m95_62 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_63 = W*in
   wire signed [9:0] m95_63;
   assign m95_63 =10'b0;

   // m95_64 = W*in
   wire signed [9:0] m95_64;
   assign m95_64 =10'b0;

   // m95_65 = W*in
   wire signed [9:0] m95_65;
   assign m95_65 =10'b0;

   // m95_66 = W*in
   wire signed [9:0] m95_66;
   assign m95_66 =10'b0;

   // m95_67 = W*in
   wire signed [9:0] m95_67;
   assign m95_67 =10'b0;

   // m95_68 = W*in
   wire signed [9:0] m95_68;
   assign m95_68 =10'b0;

   // m95_69 = W*in
   wire signed [9:0] m95_69;
   assign m95_69 ={ {3{in95[5]}} , in95 , {1{1'b0}} };

   // m95_70 = W*in
   wire signed [9:0] m95_70;
   assign m95_70 =10'b0;

   // m95_71 = W*in
   wire signed [9:0] m95_71;
   assign m95_71 =10'b0;

   // m95_72 = W*in
   wire signed [9:0] m95_72;
   assign m95_72 =10'b0;

   // m95_73 = W*in
   wire signed [9:0] m95_73;
   assign m95_73 =10'b0;

   // m95_74 = W*in
   wire signed [9:0] m95_74;
   assign m95_74 =10'b0;

   // m95_75 = W*in
   wire signed [9:0] m95_75;
   assign m95_75 =10'b0;

   // m95_76 = W*in
   wire signed [9:0] m95_76;
   assign m95_76 =10'b0;

   // m95_77 = W*in
   wire signed [9:0] m95_77;
   assign m95_77 =10'b0;

   // m95_78 = W*in
   wire signed [9:0] m95_78;
   assign m95_78 ={ {3{neg95[5]}} , neg95 , {1{1'b0}} };

   // m95_79 = W*in
   wire signed [9:0] m95_79;
   assign m95_79 =10'b0;

   // m95_80 = W*in
   wire signed [9:0] m95_80;
   assign m95_80 =10'b0;

   // m95_81 = W*in
   wire signed [9:0] m95_81;
   assign m95_81 =10'b0;

   // m96_1 = W*in
   wire signed [9:0] m96_1;
   assign m96_1 =10'b0;

   // m96_2 = W*in
   wire signed [9:0] m96_2;
   assign m96_2 =10'b0;

   // m96_3 = W*in
   wire signed [9:0] m96_3;
   assign m96_3 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_4 = W*in
   wire signed [9:0] m96_4;
   assign m96_4 =10'b0;

   // m96_5 = W*in
   wire signed [9:0] m96_5;
   assign m96_5 =10'b0;

   // m96_6 = W*in
   wire signed [9:0] m96_6;
   assign m96_6 =10'b0;

   // m96_7 = W*in
   wire signed [9:0] m96_7;
   assign m96_7 =10'b0;

   // m96_8 = W*in
   wire signed [9:0] m96_8;
   assign m96_8 =10'b0;

   // m96_9 = W*in
   wire signed [9:0] m96_9;
   assign m96_9 =10'b0;

   // m96_10 = W*in
   wire signed [9:0] m96_10;
   assign m96_10 =10'b0;

   // m96_11 = W*in
   wire signed [9:0] m96_11;
   assign m96_11 =10'b0;

   // m96_12 = W*in
   wire signed [9:0] m96_12;
   assign m96_12 =10'b0;

   // m96_13 = W*in
   wire signed [9:0] m96_13;
   assign m96_13 =10'b0;

   // m96_14 = W*in
   wire signed [9:0] m96_14;
   assign m96_14 =10'b0;

   // m96_15 = W*in
   wire signed [9:0] m96_15;
   assign m96_15 =10'b0;

   // m96_16 = W*in
   wire signed [9:0] m96_16;
   assign m96_16 =10'b0;

   // m96_17 = W*in
   wire signed [9:0] m96_17;
   assign m96_17 ={ {3{neg96[5]}} , neg96 , {1{1'b0}} };

   // m96_18 = W*in
   wire signed [9:0] m96_18;
   assign m96_18 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_19 = W*in
   wire signed [9:0] m96_19;
   assign m96_19 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_20 = W*in
   wire signed [9:0] m96_20;
   assign m96_20 =10'b0;

   // m96_21 = W*in
   wire signed [9:0] m96_21;
   assign m96_21 =10'b0;

   // m96_22 = W*in
   wire signed [9:0] m96_22;
   assign m96_22 =10'b0;

   // m96_23 = W*in
   wire signed [9:0] m96_23;
   assign m96_23 =10'b0;

   // m96_24 = W*in
   wire signed [9:0] m96_24;
   assign m96_24 =10'b0;

   // m96_25 = W*in
   wire signed [9:0] m96_25;
   assign m96_25 =10'b0;

   // m96_26 = W*in
   wire signed [9:0] m96_26;
   assign m96_26 =10'b0;

   // m96_27 = W*in
   wire signed [9:0] m96_27;
   assign m96_27 =10'b0;

   // m96_28 = W*in
   wire signed [9:0] m96_28;
   assign m96_28 =10'b0;

   // m96_29 = W*in
   wire signed [9:0] m96_29;
   assign m96_29 =10'b0;

   // m96_30 = W*in
   wire signed [9:0] m96_30;
   assign m96_30 =10'b0;

   // m96_31 = W*in
   wire signed [9:0] m96_31;
   assign m96_31 =10'b0;

   // m96_32 = W*in
   wire signed [9:0] m96_32;
   assign m96_32 =10'b0;

   // m96_33 = W*in
   wire signed [9:0] m96_33;
   assign m96_33 =10'b0;

   // m96_34 = W*in
   wire signed [9:0] m96_34;
   assign m96_34 =10'b0;

   // m96_35 = W*in
   wire signed [9:0] m96_35;
   assign m96_35 =10'b0;

   // m96_36 = W*in
   wire signed [9:0] m96_36;
   assign m96_36 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_37 = W*in
   wire signed [9:0] m96_37;
   assign m96_37 =10'b0;

   // m96_38 = W*in
   wire signed [9:0] m96_38;
   assign m96_38 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_39 = W*in
   wire signed [9:0] m96_39;
   assign m96_39 =10'b0;

   // m96_40 = W*in
   wire signed [9:0] m96_40;
   assign m96_40 =10'b0;

   // m96_41 = W*in
   wire signed [9:0] m96_41;
   assign m96_41 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_42 = W*in
   wire signed [9:0] m96_42;
   assign m96_42 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_43 = W*in
   wire signed [9:0] m96_43;
   assign m96_43 =10'b0;

   // m96_44 = W*in
   wire signed [9:0] m96_44;
   assign m96_44 =10'b0;

   // m96_45 = W*in
   wire signed [9:0] m96_45;
   assign m96_45 =10'b0;

   // m96_46 = W*in
   wire signed [9:0] m96_46;
   assign m96_46 =10'b0;

   // m96_47 = W*in
   wire signed [9:0] m96_47;
   assign m96_47 =10'b0;

   // m96_48 = W*in
   wire signed [9:0] m96_48;
   assign m96_48 ={ {3{neg96[5]}} , neg96 , {1{1'b0}} };

   // m96_49 = W*in
   wire signed [9:0] m96_49;
   assign m96_49 ={ {3{neg96[5]}} , neg96 , {1{1'b0}} };

   // m96_50 = W*in
   wire signed [9:0] m96_50;
   assign m96_50 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_51 = W*in
   wire signed [9:0] m96_51;
   assign m96_51 =10'b0;

   // m96_52 = W*in
   wire signed [9:0] m96_52;
   assign m96_52 =10'b0;

   // m96_53 = W*in
   wire signed [9:0] m96_53;
   assign m96_53 =10'b0;

   // m96_54 = W*in
   wire signed [9:0] m96_54;
   assign m96_54 =10'b0;

   // m96_55 = W*in
   wire signed [9:0] m96_55;
   assign m96_55 =10'b0;

   // m96_56 = W*in
   wire signed [9:0] m96_56;
   assign m96_56 =10'b0;

   // m96_57 = W*in
   wire signed [9:0] m96_57;
   assign m96_57 =10'b0;

   // m96_58 = W*in
   wire signed [9:0] m96_58;
   assign m96_58 =10'b0;

   // m96_59 = W*in
   wire signed [9:0] m96_59;
   assign m96_59 =10'b0;

   // m96_60 = W*in
   wire signed [9:0] m96_60;
   assign m96_60 =10'b0;

   // m96_61 = W*in
   wire signed [9:0] m96_61;
   assign m96_61 =10'b0;

   // m96_62 = W*in
   wire signed [9:0] m96_62;
   assign m96_62 =10'b0;

   // m96_63 = W*in
   wire signed [9:0] m96_63;
   assign m96_63 =10'b0;

   // m96_64 = W*in
   wire signed [9:0] m96_64;
   assign m96_64 =10'b0;

   // m96_65 = W*in
   wire signed [9:0] m96_65;
   assign m96_65 =10'b0;

   // m96_66 = W*in
   wire signed [9:0] m96_66;
   assign m96_66 =10'b0;

   // m96_67 = W*in
   wire signed [9:0] m96_67;
   assign m96_67 =10'b0;

   // m96_68 = W*in
   wire signed [9:0] m96_68;
   assign m96_68 =10'b0;

   // m96_69 = W*in
   wire signed [9:0] m96_69;
   assign m96_69 =10'b0;

   // m96_70 = W*in
   wire signed [9:0] m96_70;
   assign m96_70 =10'b0;

   // m96_71 = W*in
   wire signed [9:0] m96_71;
   assign m96_71 =10'b0;

   // m96_72 = W*in
   wire signed [9:0] m96_72;
   assign m96_72 =10'b0;

   // m96_73 = W*in
   wire signed [9:0] m96_73;
   assign m96_73 =10'b0;

   // m96_74 = W*in
   wire signed [9:0] m96_74;
   assign m96_74 =10'b0;

   // m96_75 = W*in
   wire signed [9:0] m96_75;
   assign m96_75 =10'b0;

   // m96_76 = W*in
   wire signed [9:0] m96_76;
   assign m96_76 =10'b0;

   // m96_77 = W*in
   wire signed [9:0] m96_77;
   assign m96_77 =10'b0;

   // m96_78 = W*in
   wire signed [9:0] m96_78;
   assign m96_78 ={ {3{in96[5]}} , in96 , {1{1'b0}} };

   // m96_79 = W*in
   wire signed [9:0] m96_79;
   assign m96_79 =10'b0;

   // m96_80 = W*in
   wire signed [9:0] m96_80;
   assign m96_80 =10'b0;

   // m96_81 = W*in
   wire signed [9:0] m96_81;
   assign m96_81 =10'b0;

   // m97_1 = W*in
   wire signed [9:0] m97_1;
   assign m97_1 =10'b0;

   // m97_2 = W*in
   wire signed [9:0] m97_2;
   assign m97_2 =10'b0;

   // m97_3 = W*in
   wire signed [9:0] m97_3;
   assign m97_3 =10'b0;

   // m97_4 = W*in
   wire signed [9:0] m97_4;
   assign m97_4 =10'b0;

   // m97_5 = W*in
   wire signed [9:0] m97_5;
   assign m97_5 =10'b0;

   // m97_6 = W*in
   wire signed [9:0] m97_6;
   assign m97_6 ={ {2{in97[5]}} , in97 , {2{1'b0}} };

   // m97_7 = W*in
   wire signed [9:0] m97_7;
   assign m97_7 =10'b0;

   // m97_8 = W*in
   wire signed [9:0] m97_8;
   assign m97_8 ={ {2{in97[5]}} , in97 , {2{1'b0}} };

   // m97_9 = W*in
   wire signed [9:0] m97_9;
   assign m97_9 =10'b0;

   // m97_10 = W*in
   wire signed [9:0] m97_10;
   assign m97_10 =10'b0;

   // m97_11 = W*in
   wire signed [9:0] m97_11;
   assign m97_11 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_12 = W*in
   wire signed [9:0] m97_12;
   assign m97_12 =10'b0;

   // m97_13 = W*in
   wire signed [9:0] m97_13;
   assign m97_13 =10'b0;

   // m97_14 = W*in
   wire signed [9:0] m97_14;
   assign m97_14 =10'b0;

   // m97_15 = W*in
   wire signed [9:0] m97_15;
   assign m97_15 =10'b0;

   // m97_16 = W*in
   wire signed [9:0] m97_16;
   assign m97_16 =10'b0;

   // m97_17 = W*in
   wire signed [9:0] m97_17;
   assign m97_17 =10'b0;

   // m97_18 = W*in
   wire signed [9:0] m97_18;
   assign m97_18 =10'b0;

   // m97_19 = W*in
   wire signed [9:0] m97_19;
   assign m97_19 =10'b0;

   // m97_20 = W*in
   wire signed [9:0] m97_20;
   assign m97_20 =10'b0;

   // m97_21 = W*in
   wire signed [9:0] m97_21;
   assign m97_21 =10'b0;

   // m97_22 = W*in
   wire signed [9:0] m97_22;
   assign m97_22 =10'b0;

   // m97_23 = W*in
   wire signed [9:0] m97_23;
   assign m97_23 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_24 = W*in
   wire signed [9:0] m97_24;
   assign m97_24 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_25 = W*in
   wire signed [9:0] m97_25;
   assign m97_25 =10'b0;

   // m97_26 = W*in
   wire signed [9:0] m97_26;
   assign m97_26 =10'b0;

   // m97_27 = W*in
   wire signed [9:0] m97_27;
   assign m97_27 =10'b0;

   // m97_28 = W*in
   wire signed [9:0] m97_28;
   assign m97_28 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_29 = W*in
   wire signed [9:0] m97_29;
   assign m97_29 =10'b0;

   // m97_30 = W*in
   wire signed [9:0] m97_30;
   assign m97_30 =10'b0;

   // m97_31 = W*in
   wire signed [9:0] m97_31;
   assign m97_31 =10'b0;

   // m97_32 = W*in
   wire signed [9:0] m97_32;
   assign m97_32 =10'b0;

   // m97_33 = W*in
   wire signed [9:0] m97_33;
   assign m97_33 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_34 = W*in
   wire signed [9:0] m97_34;
   assign m97_34 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_35 = W*in
   wire signed [9:0] m97_35;
   assign m97_35 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_36 = W*in
   wire signed [9:0] m97_36;
   assign m97_36 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_37 = W*in
   wire signed [9:0] m97_37;
   assign m97_37 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_38 = W*in
   wire signed [9:0] m97_38;
   assign m97_38 =10'b0;

   // m97_39 = W*in
   wire signed [9:0] m97_39;
   assign m97_39 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_40 = W*in
   wire signed [9:0] m97_40;
   assign m97_40 =10'b0;

   // m97_41 = W*in
   wire signed [9:0] m97_41;
   assign m97_41 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_42 = W*in
   wire signed [9:0] m97_42;
   assign m97_42 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_43 = W*in
   wire signed [9:0] m97_43;
   assign m97_43 =10'b0;

   // m97_44 = W*in
   wire signed [9:0] m97_44;
   assign m97_44 =10'b0;

   // m97_45 = W*in
   wire signed [9:0] m97_45;
   assign m97_45 =10'b0;

   // m97_46 = W*in
   wire signed [9:0] m97_46;
   assign m97_46 =10'b0;

   // m97_47 = W*in
   wire signed [9:0] m97_47;
   assign m97_47 =10'b0;

   // m97_48 = W*in
   wire signed [9:0] m97_48;
   assign m97_48 =10'b0;

   // m97_49 = W*in
   wire signed [9:0] m97_49;
   assign m97_49 =10'b0;

   // m97_50 = W*in
   wire signed [9:0] m97_50;
   assign m97_50 =10'b0;

   // m97_51 = W*in
   wire signed [9:0] m97_51;
   assign m97_51 ={ {2{in97[5]}} , in97 , {2{1'b0}} };

   // m97_52 = W*in
   wire signed [9:0] m97_52;
   assign m97_52 =10'b0;

   // m97_53 = W*in
   wire signed [9:0] m97_53;
   assign m97_53 =10'b0;

   // m97_54 = W*in
   wire signed [9:0] m97_54;
   assign m97_54 =10'b0;

   // m97_55 = W*in
   wire signed [9:0] m97_55;
   assign m97_55 =10'b0;

   // m97_56 = W*in
   wire signed [9:0] m97_56;
   assign m97_56 ={ {2{in97[5]}} , in97 , {2{1'b0}} };

   // m97_57 = W*in
   wire signed [9:0] m97_57;
   assign m97_57 =10'b0;

   // m97_58 = W*in
   wire signed [9:0] m97_58;
   assign m97_58 ={ {2{in97[5]}} , in97 , {2{1'b0}} };

   // m97_59 = W*in
   wire signed [9:0] m97_59;
   assign m97_59 =10'b0;

   // m97_60 = W*in
   wire signed [9:0] m97_60;
   assign m97_60 ={ {2{in97[5]}} , in97 , {2{1'b0}} };

   // m97_61 = W*in
   wire signed [9:0] m97_61;
   assign m97_61 =10'b0;

   // m97_62 = W*in
   wire signed [9:0] m97_62;
   assign m97_62 =10'b0;

   // m97_63 = W*in
   wire signed [9:0] m97_63;
   assign m97_63 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_64 = W*in
   wire signed [9:0] m97_64;
   assign m97_64 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_65 = W*in
   wire signed [9:0] m97_65;
   assign m97_65 =10'b0;

   // m97_66 = W*in
   wire signed [9:0] m97_66;
   assign m97_66 =10'b0;

   // m97_67 = W*in
   wire signed [9:0] m97_67;
   assign m97_67 =10'b0;

   // m97_68 = W*in
   wire signed [9:0] m97_68;
   assign m97_68 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_69 = W*in
   wire signed [9:0] m97_69;
   assign m97_69 =10'b0;

   // m97_70 = W*in
   wire signed [9:0] m97_70;
   assign m97_70 =10'b0;

   // m97_71 = W*in
   wire signed [9:0] m97_71;
   assign m97_71 =10'b0;

   // m97_72 = W*in
   wire signed [9:0] m97_72;
   assign m97_72 =10'b0;

   // m97_73 = W*in
   wire signed [9:0] m97_73;
   assign m97_73 =10'b0;

   // m97_74 = W*in
   wire signed [9:0] m97_74;
   assign m97_74 =10'b0;

   // m97_75 = W*in
   wire signed [9:0] m97_75;
   assign m97_75 =10'b0;

   // m97_76 = W*in
   wire signed [9:0] m97_76;
   assign m97_76 =10'b0;

   // m97_77 = W*in
   wire signed [9:0] m97_77;
   assign m97_77 =10'b0;

   // m97_78 = W*in
   wire signed [9:0] m97_78;
   assign m97_78 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_79 = W*in
   wire signed [9:0] m97_79;
   assign m97_79 =10'b0;

   // m97_80 = W*in
   wire signed [9:0] m97_80;
   assign m97_80 =10'b0;

   // m97_81 = W*in
   wire signed [9:0] m97_81;
   assign m97_81 =10'b0;

   // m98_1 = W*in
   wire signed [9:0] m98_1;
   assign m98_1 =10'b0;

   // m98_2 = W*in
   wire signed [9:0] m98_2;
   assign m98_2 =10'b0;

   // m98_3 = W*in
   wire signed [9:0] m98_3;
   assign m98_3 =10'b0;

   // m98_4 = W*in
   wire signed [9:0] m98_4;
   assign m98_4 =10'b0;

   // m98_5 = W*in
   wire signed [9:0] m98_5;
   assign m98_5 =10'b0;

   // m98_6 = W*in
   wire signed [9:0] m98_6;
   assign m98_6 =10'b0;

   // m98_7 = W*in
   wire signed [9:0] m98_7;
   assign m98_7 =10'b0;

   // m98_8 = W*in
   wire signed [9:0] m98_8;
   assign m98_8 =10'b0;

   // m98_9 = W*in
   wire signed [9:0] m98_9;
   assign m98_9 =10'b0;

   // m98_10 = W*in
   wire signed [9:0] m98_10;
   assign m98_10 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_11 = W*in
   wire signed [9:0] m98_11;
   assign m98_11 =10'b0;

   // m98_12 = W*in
   wire signed [9:0] m98_12;
   assign m98_12 =10'b0;

   // m98_13 = W*in
   wire signed [9:0] m98_13;
   assign m98_13 =10'b0;

   // m98_14 = W*in
   wire signed [9:0] m98_14;
   assign m98_14 =10'b0;

   // m98_15 = W*in
   wire signed [9:0] m98_15;
   assign m98_15 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_16 = W*in
   wire signed [9:0] m98_16;
   assign m98_16 =10'b0;

   // m98_17 = W*in
   wire signed [9:0] m98_17;
   assign m98_17 =10'b0;

   // m98_18 = W*in
   wire signed [9:0] m98_18;
   assign m98_18 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_19 = W*in
   wire signed [9:0] m98_19;
   assign m98_19 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_20 = W*in
   wire signed [9:0] m98_20;
   assign m98_20 =10'b0;

   // m98_21 = W*in
   wire signed [9:0] m98_21;
   assign m98_21 =10'b0;

   // m98_22 = W*in
   wire signed [9:0] m98_22;
   assign m98_22 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_23 = W*in
   wire signed [9:0] m98_23;
   assign m98_23 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_24 = W*in
   wire signed [9:0] m98_24;
   assign m98_24 =10'b0;

   // m98_25 = W*in
   wire signed [9:0] m98_25;
   assign m98_25 =10'b0;

   // m98_26 = W*in
   wire signed [9:0] m98_26;
   assign m98_26 =10'b0;

   // m98_27 = W*in
   wire signed [9:0] m98_27;
   assign m98_27 =10'b0;

   // m98_28 = W*in
   wire signed [9:0] m98_28;
   assign m98_28 =10'b0;

   // m98_29 = W*in
   wire signed [9:0] m98_29;
   assign m98_29 =10'b0;

   // m98_30 = W*in
   wire signed [9:0] m98_30;
   assign m98_30 =10'b0;

   // m98_31 = W*in
   wire signed [9:0] m98_31;
   assign m98_31 =10'b0;

   // m98_32 = W*in
   wire signed [9:0] m98_32;
   assign m98_32 =10'b0;

   // m98_33 = W*in
   wire signed [9:0] m98_33;
   assign m98_33 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_34 = W*in
   wire signed [9:0] m98_34;
   assign m98_34 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_35 = W*in
   wire signed [9:0] m98_35;
   assign m98_35 =10'b0;

   // m98_36 = W*in
   wire signed [9:0] m98_36;
   assign m98_36 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_37 = W*in
   wire signed [9:0] m98_37;
   assign m98_37 =10'b0;

   // m98_38 = W*in
   wire signed [9:0] m98_38;
   assign m98_38 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_39 = W*in
   wire signed [9:0] m98_39;
   assign m98_39 =10'b0;

   // m98_40 = W*in
   wire signed [9:0] m98_40;
   assign m98_40 ={ {2{in98[5]}} , in98 , {2{1'b0}} };

   // m98_41 = W*in
   wire signed [9:0] m98_41;
   assign m98_41 =10'b0;

   // m98_42 = W*in
   wire signed [9:0] m98_42;
   assign m98_42 =10'b0;

   // m98_43 = W*in
   wire signed [9:0] m98_43;
   assign m98_43 =10'b0;

   // m98_44 = W*in
   wire signed [9:0] m98_44;
   assign m98_44 =10'b0;

   // m98_45 = W*in
   wire signed [9:0] m98_45;
   assign m98_45 =10'b0;

   // m98_46 = W*in
   wire signed [9:0] m98_46;
   assign m98_46 =10'b0;

   // m98_47 = W*in
   wire signed [9:0] m98_47;
   assign m98_47 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_48 = W*in
   wire signed [9:0] m98_48;
   assign m98_48 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_49 = W*in
   wire signed [9:0] m98_49;
   assign m98_49 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_50 = W*in
   wire signed [9:0] m98_50;
   assign m98_50 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_51 = W*in
   wire signed [9:0] m98_51;
   assign m98_51 =10'b0;

   // m98_52 = W*in
   wire signed [9:0] m98_52;
   assign m98_52 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_53 = W*in
   wire signed [9:0] m98_53;
   assign m98_53 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_54 = W*in
   wire signed [9:0] m98_54;
   assign m98_54 =10'b0;

   // m98_55 = W*in
   wire signed [9:0] m98_55;
   assign m98_55 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_56 = W*in
   wire signed [9:0] m98_56;
   assign m98_56 =10'b0;

   // m98_57 = W*in
   wire signed [9:0] m98_57;
   assign m98_57 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_58 = W*in
   wire signed [9:0] m98_58;
   assign m98_58 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_59 = W*in
   wire signed [9:0] m98_59;
   assign m98_59 =10'b0;

   // m98_60 = W*in
   wire signed [9:0] m98_60;
   assign m98_60 ={ {3{in98[5]}} , in98 , {1{1'b0}} };

   // m98_61 = W*in
   wire signed [9:0] m98_61;
   assign m98_61 =10'b0;

   // m98_62 = W*in
   wire signed [9:0] m98_62;
   assign m98_62 =10'b0;

   // m98_63 = W*in
   wire signed [9:0] m98_63;
   assign m98_63 =10'b0;

   // m98_64 = W*in
   wire signed [9:0] m98_64;
   assign m98_64 =10'b0;

   // m98_65 = W*in
   wire signed [9:0] m98_65;
   assign m98_65 =10'b0;

   // m98_66 = W*in
   wire signed [9:0] m98_66;
   assign m98_66 =10'b0;

   // m98_67 = W*in
   wire signed [9:0] m98_67;
   assign m98_67 =10'b0;

   // m98_68 = W*in
   wire signed [9:0] m98_68;
   assign m98_68 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_69 = W*in
   wire signed [9:0] m98_69;
   assign m98_69 =10'b0;

   // m98_70 = W*in
   wire signed [9:0] m98_70;
   assign m98_70 ={ {2{in98[5]}} , in98 , {2{1'b0}} };

   // m98_71 = W*in
   wire signed [9:0] m98_71;
   assign m98_71 =10'b0;

   // m98_72 = W*in
   wire signed [9:0] m98_72;
   assign m98_72 ={ {2{in98[5]}} , in98 , {2{1'b0}} };

   // m98_73 = W*in
   wire signed [9:0] m98_73;
   assign m98_73 =10'b0;

   // m98_74 = W*in
   wire signed [9:0] m98_74;
   assign m98_74 =10'b0;

   // m98_75 = W*in
   wire signed [9:0] m98_75;
   assign m98_75 =10'b0;

   // m98_76 = W*in
   wire signed [9:0] m98_76;
   assign m98_76 =10'b0;

   // m98_77 = W*in
   wire signed [9:0] m98_77;
   assign m98_77 ={ {3{neg98[5]}} , neg98 , {1{1'b0}} };

   // m98_78 = W*in
   wire signed [9:0] m98_78;
   assign m98_78 =10'b0;

   // m98_79 = W*in
   wire signed [9:0] m98_79;
   assign m98_79 =10'b0;

   // m98_80 = W*in
   wire signed [9:0] m98_80;
   assign m98_80 =10'b0;

   // m98_81 = W*in
   wire signed [9:0] m98_81;
   assign m98_81 =10'b0;

   // m99_1 = W*in
   wire signed [9:0] m99_1;
   assign m99_1 =10'b0;

   // m99_2 = W*in
   wire signed [9:0] m99_2;
   assign m99_2 =10'b0;

   // m99_3 = W*in
   wire signed [9:0] m99_3;
   assign m99_3 =10'b0;

   // m99_4 = W*in
   wire signed [9:0] m99_4;
   assign m99_4 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_5 = W*in
   wire signed [9:0] m99_5;
   assign m99_5 =10'b0;

   // m99_6 = W*in
   wire signed [9:0] m99_6;
   assign m99_6 =10'b0;

   // m99_7 = W*in
   wire signed [9:0] m99_7;
   assign m99_7 =10'b0;

   // m99_8 = W*in
   wire signed [9:0] m99_8;
   assign m99_8 =10'b0;

   // m99_9 = W*in
   wire signed [9:0] m99_9;
   assign m99_9 =10'b0;

   // m99_10 = W*in
   wire signed [9:0] m99_10;
   assign m99_10 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_11 = W*in
   wire signed [9:0] m99_11;
   assign m99_11 =10'b0;

   // m99_12 = W*in
   wire signed [9:0] m99_12;
   assign m99_12 =10'b0;

   // m99_13 = W*in
   wire signed [9:0] m99_13;
   assign m99_13 =10'b0;

   // m99_14 = W*in
   wire signed [9:0] m99_14;
   assign m99_14 =10'b0;

   // m99_15 = W*in
   wire signed [9:0] m99_15;
   assign m99_15 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_16 = W*in
   wire signed [9:0] m99_16;
   assign m99_16 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_17 = W*in
   wire signed [9:0] m99_17;
   assign m99_17 =10'b0;

   // m99_18 = W*in
   wire signed [9:0] m99_18;
   assign m99_18 =10'b0;

   // m99_19 = W*in
   wire signed [9:0] m99_19;
   assign m99_19 =10'b0;

   // m99_20 = W*in
   wire signed [9:0] m99_20;
   assign m99_20 =10'b0;

   // m99_21 = W*in
   wire signed [9:0] m99_21;
   assign m99_21 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_22 = W*in
   wire signed [9:0] m99_22;
   assign m99_22 =10'b0;

   // m99_23 = W*in
   wire signed [9:0] m99_23;
   assign m99_23 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_24 = W*in
   wire signed [9:0] m99_24;
   assign m99_24 =10'b0;

   // m99_25 = W*in
   wire signed [9:0] m99_25;
   assign m99_25 =10'b0;

   // m99_26 = W*in
   wire signed [9:0] m99_26;
   assign m99_26 =10'b0;

   // m99_27 = W*in
   wire signed [9:0] m99_27;
   assign m99_27 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_28 = W*in
   wire signed [9:0] m99_28;
   assign m99_28 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_29 = W*in
   wire signed [9:0] m99_29;
   assign m99_29 =10'b0;

   // m99_30 = W*in
   wire signed [9:0] m99_30;
   assign m99_30 =10'b0;

   // m99_31 = W*in
   wire signed [9:0] m99_31;
   assign m99_31 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_32 = W*in
   wire signed [9:0] m99_32;
   assign m99_32 =10'b0;

   // m99_33 = W*in
   wire signed [9:0] m99_33;
   assign m99_33 =10'b0;

   // m99_34 = W*in
   wire signed [9:0] m99_34;
   assign m99_34 ={ {2{in99[5]}} , in99 , {2{1'b0}} };

   // m99_35 = W*in
   wire signed [9:0] m99_35;
   assign m99_35 =10'b0;

   // m99_36 = W*in
   wire signed [9:0] m99_36;
   assign m99_36 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_37 = W*in
   wire signed [9:0] m99_37;
   assign m99_37 =10'b0;

   // m99_38 = W*in
   wire signed [9:0] m99_38;
   assign m99_38 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_39 = W*in
   wire signed [9:0] m99_39;
   assign m99_39 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_40 = W*in
   wire signed [9:0] m99_40;
   assign m99_40 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_41 = W*in
   wire signed [9:0] m99_41;
   assign m99_41 =10'b0;

   // m99_42 = W*in
   wire signed [9:0] m99_42;
   assign m99_42 =10'b0;

   // m99_43 = W*in
   wire signed [9:0] m99_43;
   assign m99_43 =10'b0;

   // m99_44 = W*in
   wire signed [9:0] m99_44;
   assign m99_44 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_45 = W*in
   wire signed [9:0] m99_45;
   assign m99_45 =10'b0;

   // m99_46 = W*in
   wire signed [9:0] m99_46;
   assign m99_46 =10'b0;

   // m99_47 = W*in
   wire signed [9:0] m99_47;
   assign m99_47 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_48 = W*in
   wire signed [9:0] m99_48;
   assign m99_48 =10'b0;

   // m99_49 = W*in
   wire signed [9:0] m99_49;
   assign m99_49 =10'b0;

   // m99_50 = W*in
   wire signed [9:0] m99_50;
   assign m99_50 =10'b0;

   // m99_51 = W*in
   wire signed [9:0] m99_51;
   assign m99_51 =10'b0;

   // m99_52 = W*in
   wire signed [9:0] m99_52;
   assign m99_52 =10'b0;

   // m99_53 = W*in
   wire signed [9:0] m99_53;
   assign m99_53 =10'b0;

   // m99_54 = W*in
   wire signed [9:0] m99_54;
   assign m99_54 =10'b0;

   // m99_55 = W*in
   wire signed [9:0] m99_55;
   assign m99_55 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_56 = W*in
   wire signed [9:0] m99_56;
   assign m99_56 =10'b0;

   // m99_57 = W*in
   wire signed [9:0] m99_57;
   assign m99_57 =10'b0;

   // m99_58 = W*in
   wire signed [9:0] m99_58;
   assign m99_58 =10'b0;

   // m99_59 = W*in
   wire signed [9:0] m99_59;
   assign m99_59 =10'b0;

   // m99_60 = W*in
   wire signed [9:0] m99_60;
   assign m99_60 =10'b0;

   // m99_61 = W*in
   wire signed [9:0] m99_61;
   assign m99_61 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_62 = W*in
   wire signed [9:0] m99_62;
   assign m99_62 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_63 = W*in
   wire signed [9:0] m99_63;
   assign m99_63 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_64 = W*in
   wire signed [9:0] m99_64;
   assign m99_64 =10'b0;

   // m99_65 = W*in
   wire signed [9:0] m99_65;
   assign m99_65 =10'b0;

   // m99_66 = W*in
   wire signed [9:0] m99_66;
   assign m99_66 =10'b0;

   // m99_67 = W*in
   wire signed [9:0] m99_67;
   assign m99_67 =10'b0;

   // m99_68 = W*in
   wire signed [9:0] m99_68;
   assign m99_68 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_69 = W*in
   wire signed [9:0] m99_69;
   assign m99_69 ={ {3{neg99[5]}} , neg99 , {1{1'b0}} };

   // m99_70 = W*in
   wire signed [9:0] m99_70;
   assign m99_70 =10'b0;

   // m99_71 = W*in
   wire signed [9:0] m99_71;
   assign m99_71 =10'b0;

   // m99_72 = W*in
   wire signed [9:0] m99_72;
   assign m99_72 =10'b0;

   // m99_73 = W*in
   wire signed [9:0] m99_73;
   assign m99_73 =10'b0;

   // m99_74 = W*in
   wire signed [9:0] m99_74;
   assign m99_74 =10'b0;

   // m99_75 = W*in
   wire signed [9:0] m99_75;
   assign m99_75 =10'b0;

   // m99_76 = W*in
   wire signed [9:0] m99_76;
   assign m99_76 ={ {2{in99[5]}} , in99 , {2{1'b0}} };

   // m99_77 = W*in
   wire signed [9:0] m99_77;
   assign m99_77 ={ {3{in99[5]}} , in99 , {1{1'b0}} };

   // m99_78 = W*in
   wire signed [9:0] m99_78;
   assign m99_78 =10'b0;

   // m99_79 = W*in
   wire signed [9:0] m99_79;
   assign m99_79 =10'b0;

   // m99_80 = W*in
   wire signed [9:0] m99_80;
   assign m99_80 =10'b0;

   // m99_81 = W*in
   wire signed [9:0] m99_81;
   assign m99_81 =10'b0;

   // m100_1 = W*in
   wire signed [9:0] m100_1;
   assign m100_1 ={ {2{in100[5]}} , in100 , {2{1'b0}} };

   // m100_2 = W*in
   wire signed [9:0] m100_2;
   assign m100_2 =10'b0;

   // m100_3 = W*in
   wire signed [9:0] m100_3;
   assign m100_3 =10'b0;

   // m100_4 = W*in
   wire signed [9:0] m100_4;
   assign m100_4 =10'b0;

   // m100_5 = W*in
   wire signed [9:0] m100_5;
   assign m100_5 =10'b0;

   // m100_6 = W*in
   wire signed [9:0] m100_6;
   assign m100_6 =10'b0;

   // m100_7 = W*in
   wire signed [9:0] m100_7;
   assign m100_7 =10'b0;

   // m100_8 = W*in
   wire signed [9:0] m100_8;
   assign m100_8 =10'b0;

   // m100_9 = W*in
   wire signed [9:0] m100_9;
   assign m100_9 =10'b0;

   // m100_10 = W*in
   wire signed [9:0] m100_10;
   assign m100_10 =10'b0;

   // m100_11 = W*in
   wire signed [9:0] m100_11;
   assign m100_11 ={ {2{in100[5]}} , in100 , {2{1'b0}} };

   // m100_12 = W*in
   wire signed [9:0] m100_12;
   assign m100_12 =10'b0;

   // m100_13 = W*in
   wire signed [9:0] m100_13;
   assign m100_13 =10'b0;

   // m100_14 = W*in
   wire signed [9:0] m100_14;
   assign m100_14 =10'b0;

   // m100_15 = W*in
   wire signed [9:0] m100_15;
   assign m100_15 =10'b0;

   // m100_16 = W*in
   wire signed [9:0] m100_16;
   assign m100_16 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_17 = W*in
   wire signed [9:0] m100_17;
   assign m100_17 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_18 = W*in
   wire signed [9:0] m100_18;
   assign m100_18 ={ {2{in100[5]}} , in100 , {2{1'b0}} };

   // m100_19 = W*in
   wire signed [9:0] m100_19;
   assign m100_19 ={ {2{in100[5]}} , in100 , {2{1'b0}} };

   // m100_20 = W*in
   wire signed [9:0] m100_20;
   assign m100_20 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_21 = W*in
   wire signed [9:0] m100_21;
   assign m100_21 ={ {2{in100[5]}} , in100 , {2{1'b0}} };

   // m100_22 = W*in
   wire signed [9:0] m100_22;
   assign m100_22 =10'b0;

   // m100_23 = W*in
   wire signed [9:0] m100_23;
   assign m100_23 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_24 = W*in
   wire signed [9:0] m100_24;
   assign m100_24 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_25 = W*in
   wire signed [9:0] m100_25;
   assign m100_25 =10'b0;

   // m100_26 = W*in
   wire signed [9:0] m100_26;
   assign m100_26 =10'b0;

   // m100_27 = W*in
   wire signed [9:0] m100_27;
   assign m100_27 =10'b0;

   // m100_28 = W*in
   wire signed [9:0] m100_28;
   assign m100_28 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_29 = W*in
   wire signed [9:0] m100_29;
   assign m100_29 =10'b0;

   // m100_30 = W*in
   wire signed [9:0] m100_30;
   assign m100_30 =10'b0;

   // m100_31 = W*in
   wire signed [9:0] m100_31;
   assign m100_31 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_32 = W*in
   wire signed [9:0] m100_32;
   assign m100_32 =10'b0;

   // m100_33 = W*in
   wire signed [9:0] m100_33;
   assign m100_33 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_34 = W*in
   wire signed [9:0] m100_34;
   assign m100_34 =10'b0;

   // m100_35 = W*in
   wire signed [9:0] m100_35;
   assign m100_35 =10'b0;

   // m100_36 = W*in
   wire signed [9:0] m100_36;
   assign m100_36 =10'b0;

   // m100_37 = W*in
   wire signed [9:0] m100_37;
   assign m100_37 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_38 = W*in
   wire signed [9:0] m100_38;
   assign m100_38 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_39 = W*in
   wire signed [9:0] m100_39;
   assign m100_39 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_40 = W*in
   wire signed [9:0] m100_40;
   assign m100_40 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_41 = W*in
   wire signed [9:0] m100_41;
   assign m100_41 ={ {2{in100[5]}} , in100 , {2{1'b0}} };

   // m100_42 = W*in
   wire signed [9:0] m100_42;
   assign m100_42 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_43 = W*in
   wire signed [9:0] m100_43;
   assign m100_43 =10'b0;

   // m100_44 = W*in
   wire signed [9:0] m100_44;
   assign m100_44 =10'b0;

   // m100_45 = W*in
   wire signed [9:0] m100_45;
   assign m100_45 =10'b0;

   // m100_46 = W*in
   wire signed [9:0] m100_46;
   assign m100_46 =10'b0;

   // m100_47 = W*in
   wire signed [9:0] m100_47;
   assign m100_47 =10'b0;

   // m100_48 = W*in
   wire signed [9:0] m100_48;
   assign m100_48 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_49 = W*in
   wire signed [9:0] m100_49;
   assign m100_49 =10'b0;

   // m100_50 = W*in
   wire signed [9:0] m100_50;
   assign m100_50 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_51 = W*in
   wire signed [9:0] m100_51;
   assign m100_51 =10'b0;

   // m100_52 = W*in
   wire signed [9:0] m100_52;
   assign m100_52 =10'b0;

   // m100_53 = W*in
   wire signed [9:0] m100_53;
   assign m100_53 =10'b0;

   // m100_54 = W*in
   wire signed [9:0] m100_54;
   assign m100_54 =10'b0;

   // m100_55 = W*in
   wire signed [9:0] m100_55;
   assign m100_55 =10'b0;

   // m100_56 = W*in
   wire signed [9:0] m100_56;
   assign m100_56 =10'b0;

   // m100_57 = W*in
   wire signed [9:0] m100_57;
   assign m100_57 =10'b0;

   // m100_58 = W*in
   wire signed [9:0] m100_58;
   assign m100_58 =10'b0;

   // m100_59 = W*in
   wire signed [9:0] m100_59;
   assign m100_59 =10'b0;

   // m100_60 = W*in
   wire signed [9:0] m100_60;
   assign m100_60 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_61 = W*in
   wire signed [9:0] m100_61;
   assign m100_61 =10'b0;

   // m100_62 = W*in
   wire signed [9:0] m100_62;
   assign m100_62 ={ {3{in100[5]}} , in100 , {1{1'b0}} };

   // m100_63 = W*in
   wire signed [9:0] m100_63;
   assign m100_63 =10'b0;

   // m100_64 = W*in
   wire signed [9:0] m100_64;
   assign m100_64 =10'b0;

   // m100_65 = W*in
   wire signed [9:0] m100_65;
   assign m100_65 =10'b0;

   // m100_66 = W*in
   wire signed [9:0] m100_66;
   assign m100_66 =10'b0;

   // m100_67 = W*in
   wire signed [9:0] m100_67;
   assign m100_67 =10'b0;

   // m100_68 = W*in
   wire signed [9:0] m100_68;
   assign m100_68 ={ {3{neg100[5]}} , neg100 , {1{1'b0}} };

   // m100_69 = W*in
   wire signed [9:0] m100_69;
   assign m100_69 =10'b0;

   // m100_70 = W*in
   wire signed [9:0] m100_70;
   assign m100_70 =10'b0;

   // m100_71 = W*in
   wire signed [9:0] m100_71;
   assign m100_71 =10'b0;

   // m100_72 = W*in
   wire signed [9:0] m100_72;
   assign m100_72 =10'b0;

   // m100_73 = W*in
   wire signed [9:0] m100_73;
   assign m100_73 =10'b0;

   // m100_74 = W*in
   wire signed [9:0] m100_74;
   assign m100_74 =10'b0;

   // m100_75 = W*in
   wire signed [9:0] m100_75;
   assign m100_75 =10'b0;

   // m100_76 = W*in
   wire signed [9:0] m100_76;
   assign m100_76 =10'b0;

   // m100_77 = W*in
   wire signed [9:0] m100_77;
   assign m100_77 =10'b0;

   // m100_78 = W*in
   wire signed [9:0] m100_78;
   assign m100_78 =10'b0;

   // m100_79 = W*in
   wire signed [9:0] m100_79;
   assign m100_79 =10'b0;

   // m100_80 = W*in
   wire signed [9:0] m100_80;
   assign m100_80 =10'b0;

   // m100_81 = W*in
   wire signed [9:0] m100_81;
   assign m100_81 =10'b0;

   // m101_1 = W*in
   wire signed [9:0] m101_1;
   assign m101_1 =10'b0;

   // m101_2 = W*in
   wire signed [9:0] m101_2;
   assign m101_2 =10'b0;

   // m101_3 = W*in
   wire signed [9:0] m101_3;
   assign m101_3 =10'b0;

   // m101_4 = W*in
   wire signed [9:0] m101_4;
   assign m101_4 =10'b0;

   // m101_5 = W*in
   wire signed [9:0] m101_5;
   assign m101_5 =10'b0;

   // m101_6 = W*in
   wire signed [9:0] m101_6;
   assign m101_6 =10'b0;

   // m101_7 = W*in
   wire signed [9:0] m101_7;
   assign m101_7 =10'b0;

   // m101_8 = W*in
   wire signed [9:0] m101_8;
   assign m101_8 =10'b0;

   // m101_9 = W*in
   wire signed [9:0] m101_9;
   assign m101_9 =10'b0;

   // m101_10 = W*in
   wire signed [9:0] m101_10;
   assign m101_10 =10'b0;

   // m101_11 = W*in
   wire signed [9:0] m101_11;
   assign m101_11 =10'b0;

   // m101_12 = W*in
   wire signed [9:0] m101_12;
   assign m101_12 =10'b0;

   // m101_13 = W*in
   wire signed [9:0] m101_13;
   assign m101_13 =10'b0;

   // m101_14 = W*in
   wire signed [9:0] m101_14;
   assign m101_14 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_15 = W*in
   wire signed [9:0] m101_15;
   assign m101_15 =10'b0;

   // m101_16 = W*in
   wire signed [9:0] m101_16;
   assign m101_16 =10'b0;

   // m101_17 = W*in
   wire signed [9:0] m101_17;
   assign m101_17 =10'b0;

   // m101_18 = W*in
   wire signed [9:0] m101_18;
   assign m101_18 =10'b0;

   // m101_19 = W*in
   wire signed [9:0] m101_19;
   assign m101_19 =10'b0;

   // m101_20 = W*in
   wire signed [9:0] m101_20;
   assign m101_20 =10'b0;

   // m101_21 = W*in
   wire signed [9:0] m101_21;
   assign m101_21 =10'b0;

   // m101_22 = W*in
   wire signed [9:0] m101_22;
   assign m101_22 ={ {3{neg101[5]}} , neg101 , {1{1'b0}} };

   // m101_23 = W*in
   wire signed [9:0] m101_23;
   assign m101_23 =10'b0;

   // m101_24 = W*in
   wire signed [9:0] m101_24;
   assign m101_24 =10'b0;

   // m101_25 = W*in
   wire signed [9:0] m101_25;
   assign m101_25 =10'b0;

   // m101_26 = W*in
   wire signed [9:0] m101_26;
   assign m101_26 =10'b0;

   // m101_27 = W*in
   wire signed [9:0] m101_27;
   assign m101_27 =10'b0;

   // m101_28 = W*in
   wire signed [9:0] m101_28;
   assign m101_28 =10'b0;

   // m101_29 = W*in
   wire signed [9:0] m101_29;
   assign m101_29 =10'b0;

   // m101_30 = W*in
   wire signed [9:0] m101_30;
   assign m101_30 =10'b0;

   // m101_31 = W*in
   wire signed [9:0] m101_31;
   assign m101_31 =10'b0;

   // m101_32 = W*in
   wire signed [9:0] m101_32;
   assign m101_32 =10'b0;

   // m101_33 = W*in
   wire signed [9:0] m101_33;
   assign m101_33 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_34 = W*in
   wire signed [9:0] m101_34;
   assign m101_34 =10'b0;

   // m101_35 = W*in
   wire signed [9:0] m101_35;
   assign m101_35 =10'b0;

   // m101_36 = W*in
   wire signed [9:0] m101_36;
   assign m101_36 =10'b0;

   // m101_37 = W*in
   wire signed [9:0] m101_37;
   assign m101_37 =10'b0;

   // m101_38 = W*in
   wire signed [9:0] m101_38;
   assign m101_38 =10'b0;

   // m101_39 = W*in
   wire signed [9:0] m101_39;
   assign m101_39 =10'b0;

   // m101_40 = W*in
   wire signed [9:0] m101_40;
   assign m101_40 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_41 = W*in
   wire signed [9:0] m101_41;
   assign m101_41 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_42 = W*in
   wire signed [9:0] m101_42;
   assign m101_42 =10'b0;

   // m101_43 = W*in
   wire signed [9:0] m101_43;
   assign m101_43 =10'b0;

   // m101_44 = W*in
   wire signed [9:0] m101_44;
   assign m101_44 =10'b0;

   // m101_45 = W*in
   wire signed [9:0] m101_45;
   assign m101_45 =10'b0;

   // m101_46 = W*in
   wire signed [9:0] m101_46;
   assign m101_46 =10'b0;

   // m101_47 = W*in
   wire signed [9:0] m101_47;
   assign m101_47 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_48 = W*in
   wire signed [9:0] m101_48;
   assign m101_48 =10'b0;

   // m101_49 = W*in
   wire signed [9:0] m101_49;
   assign m101_49 ={ {3{neg101[5]}} , neg101 , {1{1'b0}} };

   // m101_50 = W*in
   wire signed [9:0] m101_50;
   assign m101_50 =10'b0;

   // m101_51 = W*in
   wire signed [9:0] m101_51;
   assign m101_51 =10'b0;

   // m101_52 = W*in
   wire signed [9:0] m101_52;
   assign m101_52 =10'b0;

   // m101_53 = W*in
   wire signed [9:0] m101_53;
   assign m101_53 =10'b0;

   // m101_54 = W*in
   wire signed [9:0] m101_54;
   assign m101_54 =10'b0;

   // m101_55 = W*in
   wire signed [9:0] m101_55;
   assign m101_55 =10'b0;

   // m101_56 = W*in
   wire signed [9:0] m101_56;
   assign m101_56 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_57 = W*in
   wire signed [9:0] m101_57;
   assign m101_57 =10'b0;

   // m101_58 = W*in
   wire signed [9:0] m101_58;
   assign m101_58 =10'b0;

   // m101_59 = W*in
   wire signed [9:0] m101_59;
   assign m101_59 =10'b0;

   // m101_60 = W*in
   wire signed [9:0] m101_60;
   assign m101_60 =10'b0;

   // m101_61 = W*in
   wire signed [9:0] m101_61;
   assign m101_61 =10'b0;

   // m101_62 = W*in
   wire signed [9:0] m101_62;
   assign m101_62 ={ {3{in101[5]}} , in101 , {1{1'b0}} };

   // m101_63 = W*in
   wire signed [9:0] m101_63;
   assign m101_63 =10'b0;

   // m101_64 = W*in
   wire signed [9:0] m101_64;
   assign m101_64 =10'b0;

   // m101_65 = W*in
   wire signed [9:0] m101_65;
   assign m101_65 =10'b0;

   // m101_66 = W*in
   wire signed [9:0] m101_66;
   assign m101_66 =10'b0;

   // m101_67 = W*in
   wire signed [9:0] m101_67;
   assign m101_67 =10'b0;

   // m101_68 = W*in
   wire signed [9:0] m101_68;
   assign m101_68 =10'b0;

   // m101_69 = W*in
   wire signed [9:0] m101_69;
   assign m101_69 =10'b0;

   // m101_70 = W*in
   wire signed [9:0] m101_70;
   assign m101_70 =10'b0;

   // m101_71 = W*in
   wire signed [9:0] m101_71;
   assign m101_71 =10'b0;

   // m101_72 = W*in
   wire signed [9:0] m101_72;
   assign m101_72 =10'b0;

   // m101_73 = W*in
   wire signed [9:0] m101_73;
   assign m101_73 =10'b0;

   // m101_74 = W*in
   wire signed [9:0] m101_74;
   assign m101_74 =10'b0;

   // m101_75 = W*in
   wire signed [9:0] m101_75;
   assign m101_75 =10'b0;

   // m101_76 = W*in
   wire signed [9:0] m101_76;
   assign m101_76 =10'b0;

   // m101_77 = W*in
   wire signed [9:0] m101_77;
   assign m101_77 =10'b0;

   // m101_78 = W*in
   wire signed [9:0] m101_78;
   assign m101_78 =10'b0;

   // m101_79 = W*in
   wire signed [9:0] m101_79;
   assign m101_79 =10'b0;

   // m101_80 = W*in
   wire signed [9:0] m101_80;
   assign m101_80 =10'b0;

   // m101_81 = W*in
   wire signed [9:0] m101_81;
   assign m101_81 =10'b0;

   // m102_1 = W*in
   wire signed [9:0] m102_1;
   assign m102_1 =10'b0;

   // m102_2 = W*in
   wire signed [9:0] m102_2;
   assign m102_2 =10'b0;

   // m102_3 = W*in
   wire signed [9:0] m102_3;
   assign m102_3 ={ {2{in102[5]}} , in102 , {2{1'b0}} };

   // m102_4 = W*in
   wire signed [9:0] m102_4;
   assign m102_4 =10'b0;

   // m102_5 = W*in
   wire signed [9:0] m102_5;
   assign m102_5 =10'b0;

   // m102_6 = W*in
   wire signed [9:0] m102_6;
   assign m102_6 =10'b0;

   // m102_7 = W*in
   wire signed [9:0] m102_7;
   assign m102_7 =10'b0;

   // m102_8 = W*in
   wire signed [9:0] m102_8;
   assign m102_8 =10'b0;

   // m102_9 = W*in
   wire signed [9:0] m102_9;
   assign m102_9 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_10 = W*in
   wire signed [9:0] m102_10;
   assign m102_10 =10'b0;

   // m102_11 = W*in
   wire signed [9:0] m102_11;
   assign m102_11 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_12 = W*in
   wire signed [9:0] m102_12;
   assign m102_12 =10'b0;

   // m102_13 = W*in
   wire signed [9:0] m102_13;
   assign m102_13 =10'b0;

   // m102_14 = W*in
   wire signed [9:0] m102_14;
   assign m102_14 =10'b0;

   // m102_15 = W*in
   wire signed [9:0] m102_15;
   assign m102_15 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_16 = W*in
   wire signed [9:0] m102_16;
   assign m102_16 =10'b0;

   // m102_17 = W*in
   wire signed [9:0] m102_17;
   assign m102_17 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_18 = W*in
   wire signed [9:0] m102_18;
   assign m102_18 =10'b0;

   // m102_19 = W*in
   wire signed [9:0] m102_19;
   assign m102_19 =10'b0;

   // m102_20 = W*in
   wire signed [9:0] m102_20;
   assign m102_20 =10'b0;

   // m102_21 = W*in
   wire signed [9:0] m102_21;
   assign m102_21 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_22 = W*in
   wire signed [9:0] m102_22;
   assign m102_22 =10'b0;

   // m102_23 = W*in
   wire signed [9:0] m102_23;
   assign m102_23 =10'b0;

   // m102_24 = W*in
   wire signed [9:0] m102_24;
   assign m102_24 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_25 = W*in
   wire signed [9:0] m102_25;
   assign m102_25 =10'b0;

   // m102_26 = W*in
   wire signed [9:0] m102_26;
   assign m102_26 =10'b0;

   // m102_27 = W*in
   wire signed [9:0] m102_27;
   assign m102_27 =10'b0;

   // m102_28 = W*in
   wire signed [9:0] m102_28;
   assign m102_28 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_29 = W*in
   wire signed [9:0] m102_29;
   assign m102_29 =10'b0;

   // m102_30 = W*in
   wire signed [9:0] m102_30;
   assign m102_30 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_31 = W*in
   wire signed [9:0] m102_31;
   assign m102_31 =10'b0;

   // m102_32 = W*in
   wire signed [9:0] m102_32;
   assign m102_32 =10'b0;

   // m102_33 = W*in
   wire signed [9:0] m102_33;
   assign m102_33 =10'b0;

   // m102_34 = W*in
   wire signed [9:0] m102_34;
   assign m102_34 =10'b0;

   // m102_35 = W*in
   wire signed [9:0] m102_35;
   assign m102_35 =10'b0;

   // m102_36 = W*in
   wire signed [9:0] m102_36;
   assign m102_36 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_37 = W*in
   wire signed [9:0] m102_37;
   assign m102_37 =10'b0;

   // m102_38 = W*in
   wire signed [9:0] m102_38;
   assign m102_38 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_39 = W*in
   wire signed [9:0] m102_39;
   assign m102_39 =10'b0;

   // m102_40 = W*in
   wire signed [9:0] m102_40;
   assign m102_40 =10'b0;

   // m102_41 = W*in
   wire signed [9:0] m102_41;
   assign m102_41 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_42 = W*in
   wire signed [9:0] m102_42;
   assign m102_42 =10'b0;

   // m102_43 = W*in
   wire signed [9:0] m102_43;
   assign m102_43 =10'b0;

   // m102_44 = W*in
   wire signed [9:0] m102_44;
   assign m102_44 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_45 = W*in
   wire signed [9:0] m102_45;
   assign m102_45 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_46 = W*in
   wire signed [9:0] m102_46;
   assign m102_46 =10'b0;

   // m102_47 = W*in
   wire signed [9:0] m102_47;
   assign m102_47 =10'b0;

   // m102_48 = W*in
   wire signed [9:0] m102_48;
   assign m102_48 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_49 = W*in
   wire signed [9:0] m102_49;
   assign m102_49 =10'b0;

   // m102_50 = W*in
   wire signed [9:0] m102_50;
   assign m102_50 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_51 = W*in
   wire signed [9:0] m102_51;
   assign m102_51 =10'b0;

   // m102_52 = W*in
   wire signed [9:0] m102_52;
   assign m102_52 =10'b0;

   // m102_53 = W*in
   wire signed [9:0] m102_53;
   assign m102_53 =10'b0;

   // m102_54 = W*in
   wire signed [9:0] m102_54;
   assign m102_54 =10'b0;

   // m102_55 = W*in
   wire signed [9:0] m102_55;
   assign m102_55 =10'b0;

   // m102_56 = W*in
   wire signed [9:0] m102_56;
   assign m102_56 =10'b0;

   // m102_57 = W*in
   wire signed [9:0] m102_57;
   assign m102_57 =10'b0;

   // m102_58 = W*in
   wire signed [9:0] m102_58;
   assign m102_58 =10'b0;

   // m102_59 = W*in
   wire signed [9:0] m102_59;
   assign m102_59 =10'b0;

   // m102_60 = W*in
   wire signed [9:0] m102_60;
   assign m102_60 =10'b0;

   // m102_61 = W*in
   wire signed [9:0] m102_61;
   assign m102_61 ={ {3{in102[5]}} , in102 , {1{1'b0}} };

   // m102_62 = W*in
   wire signed [9:0] m102_62;
   assign m102_62 ={ {2{in102[5]}} , in102 , {2{1'b0}} };

   // m102_63 = W*in
   wire signed [9:0] m102_63;
   assign m102_63 =10'b0;

   // m102_64 = W*in
   wire signed [9:0] m102_64;
   assign m102_64 =10'b0;

   // m102_65 = W*in
   wire signed [9:0] m102_65;
   assign m102_65 =10'b0;

   // m102_66 = W*in
   wire signed [9:0] m102_66;
   assign m102_66 =10'b0;

   // m102_67 = W*in
   wire signed [9:0] m102_67;
   assign m102_67 =10'b0;

   // m102_68 = W*in
   wire signed [9:0] m102_68;
   assign m102_68 =10'b0;

   // m102_69 = W*in
   wire signed [9:0] m102_69;
   assign m102_69 =10'b0;

   // m102_70 = W*in
   wire signed [9:0] m102_70;
   assign m102_70 ={ {3{neg102[5]}} , neg102 , {1{1'b0}} };

   // m102_71 = W*in
   wire signed [9:0] m102_71;
   assign m102_71 =10'b0;

   // m102_72 = W*in
   wire signed [9:0] m102_72;
   assign m102_72 =10'b0;

   // m102_73 = W*in
   wire signed [9:0] m102_73;
   assign m102_73 =10'b0;

   // m102_74 = W*in
   wire signed [9:0] m102_74;
   assign m102_74 =10'b0;

   // m102_75 = W*in
   wire signed [9:0] m102_75;
   assign m102_75 =10'b0;

   // m102_76 = W*in
   wire signed [9:0] m102_76;
   assign m102_76 =10'b0;

   // m102_77 = W*in
   wire signed [9:0] m102_77;
   assign m102_77 =10'b0;

   // m102_78 = W*in
   wire signed [9:0] m102_78;
   assign m102_78 =10'b0;

   // m102_79 = W*in
   wire signed [9:0] m102_79;
   assign m102_79 =10'b0;

   // m102_80 = W*in
   wire signed [9:0] m102_80;
   assign m102_80 =10'b0;

   // m102_81 = W*in
   wire signed [9:0] m102_81;
   assign m102_81 =10'b0;

   // m103_1 = W*in
   wire signed [9:0] m103_1;
   assign m103_1 =10'b0;

   // m103_2 = W*in
   wire signed [9:0] m103_2;
   assign m103_2 =10'b0;

   // m103_3 = W*in
   wire signed [9:0] m103_3;
   assign m103_3 =10'b0;

   // m103_4 = W*in
   wire signed [9:0] m103_4;
   assign m103_4 =10'b0;

   // m103_5 = W*in
   wire signed [9:0] m103_5;
   assign m103_5 =10'b0;

   // m103_6 = W*in
   wire signed [9:0] m103_6;
   assign m103_6 =10'b0;

   // m103_7 = W*in
   wire signed [9:0] m103_7;
   assign m103_7 =10'b0;

   // m103_8 = W*in
   wire signed [9:0] m103_8;
   assign m103_8 =10'b0;

   // m103_9 = W*in
   wire signed [9:0] m103_9;
   assign m103_9 =10'b0;

   // m103_10 = W*in
   wire signed [9:0] m103_10;
   assign m103_10 =10'b0;

   // m103_11 = W*in
   wire signed [9:0] m103_11;
   assign m103_11 =10'b0;

   // m103_12 = W*in
   wire signed [9:0] m103_12;
   assign m103_12 =10'b0;

   // m103_13 = W*in
   wire signed [9:0] m103_13;
   assign m103_13 =10'b0;

   // m103_14 = W*in
   wire signed [9:0] m103_14;
   assign m103_14 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_15 = W*in
   wire signed [9:0] m103_15;
   assign m103_15 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_16 = W*in
   wire signed [9:0] m103_16;
   assign m103_16 =10'b0;

   // m103_17 = W*in
   wire signed [9:0] m103_17;
   assign m103_17 =10'b0;

   // m103_18 = W*in
   wire signed [9:0] m103_18;
   assign m103_18 =10'b0;

   // m103_19 = W*in
   wire signed [9:0] m103_19;
   assign m103_19 =10'b0;

   // m103_20 = W*in
   wire signed [9:0] m103_20;
   assign m103_20 =10'b0;

   // m103_21 = W*in
   wire signed [9:0] m103_21;
   assign m103_21 =10'b0;

   // m103_22 = W*in
   wire signed [9:0] m103_22;
   assign m103_22 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_23 = W*in
   wire signed [9:0] m103_23;
   assign m103_23 =10'b0;

   // m103_24 = W*in
   wire signed [9:0] m103_24;
   assign m103_24 =10'b0;

   // m103_25 = W*in
   wire signed [9:0] m103_25;
   assign m103_25 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_26 = W*in
   wire signed [9:0] m103_26;
   assign m103_26 =10'b0;

   // m103_27 = W*in
   wire signed [9:0] m103_27;
   assign m103_27 =10'b0;

   // m103_28 = W*in
   wire signed [9:0] m103_28;
   assign m103_28 =10'b0;

   // m103_29 = W*in
   wire signed [9:0] m103_29;
   assign m103_29 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_30 = W*in
   wire signed [9:0] m103_30;
   assign m103_30 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_31 = W*in
   wire signed [9:0] m103_31;
   assign m103_31 =10'b0;

   // m103_32 = W*in
   wire signed [9:0] m103_32;
   assign m103_32 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_33 = W*in
   wire signed [9:0] m103_33;
   assign m103_33 =10'b0;

   // m103_34 = W*in
   wire signed [9:0] m103_34;
   assign m103_34 =10'b0;

   // m103_35 = W*in
   wire signed [9:0] m103_35;
   assign m103_35 =10'b0;

   // m103_36 = W*in
   wire signed [9:0] m103_36;
   assign m103_36 =10'b0;

   // m103_37 = W*in
   wire signed [9:0] m103_37;
   assign m103_37 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_38 = W*in
   wire signed [9:0] m103_38;
   assign m103_38 =10'b0;

   // m103_39 = W*in
   wire signed [9:0] m103_39;
   assign m103_39 =10'b0;

   // m103_40 = W*in
   wire signed [9:0] m103_40;
   assign m103_40 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_41 = W*in
   wire signed [9:0] m103_41;
   assign m103_41 =10'b0;

   // m103_42 = W*in
   wire signed [9:0] m103_42;
   assign m103_42 =10'b0;

   // m103_43 = W*in
   wire signed [9:0] m103_43;
   assign m103_43 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_44 = W*in
   wire signed [9:0] m103_44;
   assign m103_44 =10'b0;

   // m103_45 = W*in
   wire signed [9:0] m103_45;
   assign m103_45 =10'b0;

   // m103_46 = W*in
   wire signed [9:0] m103_46;
   assign m103_46 =10'b0;

   // m103_47 = W*in
   wire signed [9:0] m103_47;
   assign m103_47 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_48 = W*in
   wire signed [9:0] m103_48;
   assign m103_48 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_49 = W*in
   wire signed [9:0] m103_49;
   assign m103_49 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_50 = W*in
   wire signed [9:0] m103_50;
   assign m103_50 =10'b0;

   // m103_51 = W*in
   wire signed [9:0] m103_51;
   assign m103_51 =10'b0;

   // m103_52 = W*in
   wire signed [9:0] m103_52;
   assign m103_52 =10'b0;

   // m103_53 = W*in
   wire signed [9:0] m103_53;
   assign m103_53 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_54 = W*in
   wire signed [9:0] m103_54;
   assign m103_54 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_55 = W*in
   wire signed [9:0] m103_55;
   assign m103_55 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_56 = W*in
   wire signed [9:0] m103_56;
   assign m103_56 =10'b0;

   // m103_57 = W*in
   wire signed [9:0] m103_57;
   assign m103_57 =10'b0;

   // m103_58 = W*in
   wire signed [9:0] m103_58;
   assign m103_58 =10'b0;

   // m103_59 = W*in
   wire signed [9:0] m103_59;
   assign m103_59 =10'b0;

   // m103_60 = W*in
   wire signed [9:0] m103_60;
   assign m103_60 =10'b0;

   // m103_61 = W*in
   wire signed [9:0] m103_61;
   assign m103_61 =10'b0;

   // m103_62 = W*in
   wire signed [9:0] m103_62;
   assign m103_62 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_63 = W*in
   wire signed [9:0] m103_63;
   assign m103_63 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_64 = W*in
   wire signed [9:0] m103_64;
   assign m103_64 =10'b0;

   // m103_65 = W*in
   wire signed [9:0] m103_65;
   assign m103_65 =10'b0;

   // m103_66 = W*in
   wire signed [9:0] m103_66;
   assign m103_66 =10'b0;

   // m103_67 = W*in
   wire signed [9:0] m103_67;
   assign m103_67 =10'b0;

   // m103_68 = W*in
   wire signed [9:0] m103_68;
   assign m103_68 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_69 = W*in
   wire signed [9:0] m103_69;
   assign m103_69 =10'b0;

   // m103_70 = W*in
   wire signed [9:0] m103_70;
   assign m103_70 =10'b0;

   // m103_71 = W*in
   wire signed [9:0] m103_71;
   assign m103_71 =10'b0;

   // m103_72 = W*in
   wire signed [9:0] m103_72;
   assign m103_72 =10'b0;

   // m103_73 = W*in
   wire signed [9:0] m103_73;
   assign m103_73 =10'b0;

   // m103_74 = W*in
   wire signed [9:0] m103_74;
   assign m103_74 =10'b0;

   // m103_75 = W*in
   wire signed [9:0] m103_75;
   assign m103_75 =10'b0;

   // m103_76 = W*in
   wire signed [9:0] m103_76;
   assign m103_76 =10'b0;

   // m103_77 = W*in
   wire signed [9:0] m103_77;
   assign m103_77 ={ {3{neg103[5]}} , neg103 , {1{1'b0}} };

   // m103_78 = W*in
   wire signed [9:0] m103_78;
   assign m103_78 =10'b0;

   // m103_79 = W*in
   wire signed [9:0] m103_79;
   assign m103_79 ={ {3{in103[5]}} , in103 , {1{1'b0}} };

   // m103_80 = W*in
   wire signed [9:0] m103_80;
   assign m103_80 =10'b0;

   // m103_81 = W*in
   wire signed [9:0] m103_81;
   assign m103_81 =10'b0;

   // m104_1 = W*in
   wire signed [9:0] m104_1;
   assign m104_1 =10'b0;

   // m104_2 = W*in
   wire signed [9:0] m104_2;
   assign m104_2 =10'b0;

   // m104_3 = W*in
   wire signed [9:0] m104_3;
   assign m104_3 =10'b0;

   // m104_4 = W*in
   wire signed [9:0] m104_4;
   assign m104_4 =10'b0;

   // m104_5 = W*in
   wire signed [9:0] m104_5;
   assign m104_5 =10'b0;

   // m104_6 = W*in
   wire signed [9:0] m104_6;
   assign m104_6 =10'b0;

   // m104_7 = W*in
   wire signed [9:0] m104_7;
   assign m104_7 =10'b0;

   // m104_8 = W*in
   wire signed [9:0] m104_8;
   assign m104_8 =10'b0;

   // m104_9 = W*in
   wire signed [9:0] m104_9;
   assign m104_9 =10'b0;

   // m104_10 = W*in
   wire signed [9:0] m104_10;
   assign m104_10 =10'b0;

   // m104_11 = W*in
   wire signed [9:0] m104_11;
   assign m104_11 =10'b0;

   // m104_12 = W*in
   wire signed [9:0] m104_12;
   assign m104_12 =10'b0;

   // m104_13 = W*in
   wire signed [9:0] m104_13;
   assign m104_13 =10'b0;

   // m104_14 = W*in
   wire signed [9:0] m104_14;
   assign m104_14 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_15 = W*in
   wire signed [9:0] m104_15;
   assign m104_15 =10'b0;

   // m104_16 = W*in
   wire signed [9:0] m104_16;
   assign m104_16 =10'b0;

   // m104_17 = W*in
   wire signed [9:0] m104_17;
   assign m104_17 =10'b0;

   // m104_18 = W*in
   wire signed [9:0] m104_18;
   assign m104_18 =10'b0;

   // m104_19 = W*in
   wire signed [9:0] m104_19;
   assign m104_19 =10'b0;

   // m104_20 = W*in
   wire signed [9:0] m104_20;
   assign m104_20 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_21 = W*in
   wire signed [9:0] m104_21;
   assign m104_21 =10'b0;

   // m104_22 = W*in
   wire signed [9:0] m104_22;
   assign m104_22 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_23 = W*in
   wire signed [9:0] m104_23;
   assign m104_23 =10'b0;

   // m104_24 = W*in
   wire signed [9:0] m104_24;
   assign m104_24 =10'b0;

   // m104_25 = W*in
   wire signed [9:0] m104_25;
   assign m104_25 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_26 = W*in
   wire signed [9:0] m104_26;
   assign m104_26 =10'b0;

   // m104_27 = W*in
   wire signed [9:0] m104_27;
   assign m104_27 =10'b0;

   // m104_28 = W*in
   wire signed [9:0] m104_28;
   assign m104_28 =10'b0;

   // m104_29 = W*in
   wire signed [9:0] m104_29;
   assign m104_29 =10'b0;

   // m104_30 = W*in
   wire signed [9:0] m104_30;
   assign m104_30 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_31 = W*in
   wire signed [9:0] m104_31;
   assign m104_31 =10'b0;

   // m104_32 = W*in
   wire signed [9:0] m104_32;
   assign m104_32 =10'b0;

   // m104_33 = W*in
   wire signed [9:0] m104_33;
   assign m104_33 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_34 = W*in
   wire signed [9:0] m104_34;
   assign m104_34 =10'b0;

   // m104_35 = W*in
   wire signed [9:0] m104_35;
   assign m104_35 =10'b0;

   // m104_36 = W*in
   wire signed [9:0] m104_36;
   assign m104_36 =10'b0;

   // m104_37 = W*in
   wire signed [9:0] m104_37;
   assign m104_37 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_38 = W*in
   wire signed [9:0] m104_38;
   assign m104_38 =10'b0;

   // m104_39 = W*in
   wire signed [9:0] m104_39;
   assign m104_39 =10'b0;

   // m104_40 = W*in
   wire signed [9:0] m104_40;
   assign m104_40 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_41 = W*in
   wire signed [9:0] m104_41;
   assign m104_41 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_42 = W*in
   wire signed [9:0] m104_42;
   assign m104_42 =10'b0;

   // m104_43 = W*in
   wire signed [9:0] m104_43;
   assign m104_43 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_44 = W*in
   wire signed [9:0] m104_44;
   assign m104_44 =10'b0;

   // m104_45 = W*in
   wire signed [9:0] m104_45;
   assign m104_45 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_46 = W*in
   wire signed [9:0] m104_46;
   assign m104_46 =10'b0;

   // m104_47 = W*in
   wire signed [9:0] m104_47;
   assign m104_47 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_48 = W*in
   wire signed [9:0] m104_48;
   assign m104_48 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_49 = W*in
   wire signed [9:0] m104_49;
   assign m104_49 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_50 = W*in
   wire signed [9:0] m104_50;
   assign m104_50 =10'b0;

   // m104_51 = W*in
   wire signed [9:0] m104_51;
   assign m104_51 =10'b0;

   // m104_52 = W*in
   wire signed [9:0] m104_52;
   assign m104_52 =10'b0;

   // m104_53 = W*in
   wire signed [9:0] m104_53;
   assign m104_53 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_54 = W*in
   wire signed [9:0] m104_54;
   assign m104_54 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_55 = W*in
   wire signed [9:0] m104_55;
   assign m104_55 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_56 = W*in
   wire signed [9:0] m104_56;
   assign m104_56 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_57 = W*in
   wire signed [9:0] m104_57;
   assign m104_57 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_58 = W*in
   wire signed [9:0] m104_58;
   assign m104_58 =10'b0;

   // m104_59 = W*in
   wire signed [9:0] m104_59;
   assign m104_59 =10'b0;

   // m104_60 = W*in
   wire signed [9:0] m104_60;
   assign m104_60 =10'b0;

   // m104_61 = W*in
   wire signed [9:0] m104_61;
   assign m104_61 =10'b0;

   // m104_62 = W*in
   wire signed [9:0] m104_62;
   assign m104_62 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_63 = W*in
   wire signed [9:0] m104_63;
   assign m104_63 =10'b0;

   // m104_64 = W*in
   wire signed [9:0] m104_64;
   assign m104_64 =10'b0;

   // m104_65 = W*in
   wire signed [9:0] m104_65;
   assign m104_65 =10'b0;

   // m104_66 = W*in
   wire signed [9:0] m104_66;
   assign m104_66 =10'b0;

   // m104_67 = W*in
   wire signed [9:0] m104_67;
   assign m104_67 =10'b0;

   // m104_68 = W*in
   wire signed [9:0] m104_68;
   assign m104_68 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_69 = W*in
   wire signed [9:0] m104_69;
   assign m104_69 =10'b0;

   // m104_70 = W*in
   wire signed [9:0] m104_70;
   assign m104_70 =10'b0;

   // m104_71 = W*in
   wire signed [9:0] m104_71;
   assign m104_71 =10'b0;

   // m104_72 = W*in
   wire signed [9:0] m104_72;
   assign m104_72 =10'b0;

   // m104_73 = W*in
   wire signed [9:0] m104_73;
   assign m104_73 =10'b0;

   // m104_74 = W*in
   wire signed [9:0] m104_74;
   assign m104_74 =10'b0;

   // m104_75 = W*in
   wire signed [9:0] m104_75;
   assign m104_75 =10'b0;

   // m104_76 = W*in
   wire signed [9:0] m104_76;
   assign m104_76 =10'b0;

   // m104_77 = W*in
   wire signed [9:0] m104_77;
   assign m104_77 ={ {3{neg104[5]}} , neg104 , {1{1'b0}} };

   // m104_78 = W*in
   wire signed [9:0] m104_78;
   assign m104_78 =10'b0;

   // m104_79 = W*in
   wire signed [9:0] m104_79;
   assign m104_79 ={ {3{in104[5]}} , in104 , {1{1'b0}} };

   // m104_80 = W*in
   wire signed [9:0] m104_80;
   assign m104_80 =10'b0;

   // m104_81 = W*in
   wire signed [9:0] m104_81;
   assign m104_81 ={ {2{in104[5]}} , in104 , {2{1'b0}} };

   // m105_1 = W*in
   wire signed [9:0] m105_1;
   assign m105_1 =10'b0;

   // m105_2 = W*in
   wire signed [9:0] m105_2;
   assign m105_2 =10'b0;

   // m105_3 = W*in
   wire signed [9:0] m105_3;
   assign m105_3 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_4 = W*in
   wire signed [9:0] m105_4;
   assign m105_4 =10'b0;

   // m105_5 = W*in
   wire signed [9:0] m105_5;
   assign m105_5 =10'b0;

   // m105_6 = W*in
   wire signed [9:0] m105_6;
   assign m105_6 =10'b0;

   // m105_7 = W*in
   wire signed [9:0] m105_7;
   assign m105_7 =10'b0;

   // m105_8 = W*in
   wire signed [9:0] m105_8;
   assign m105_8 =10'b0;

   // m105_9 = W*in
   wire signed [9:0] m105_9;
   assign m105_9 =10'b0;

   // m105_10 = W*in
   wire signed [9:0] m105_10;
   assign m105_10 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_11 = W*in
   wire signed [9:0] m105_11;
   assign m105_11 =10'b0;

   // m105_12 = W*in
   wire signed [9:0] m105_12;
   assign m105_12 =10'b0;

   // m105_13 = W*in
   wire signed [9:0] m105_13;
   assign m105_13 =10'b0;

   // m105_14 = W*in
   wire signed [9:0] m105_14;
   assign m105_14 =10'b0;

   // m105_15 = W*in
   wire signed [9:0] m105_15;
   assign m105_15 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_16 = W*in
   wire signed [9:0] m105_16;
   assign m105_16 =10'b0;

   // m105_17 = W*in
   wire signed [9:0] m105_17;
   assign m105_17 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_18 = W*in
   wire signed [9:0] m105_18;
   assign m105_18 =10'b0;

   // m105_19 = W*in
   wire signed [9:0] m105_19;
   assign m105_19 =10'b0;

   // m105_20 = W*in
   wire signed [9:0] m105_20;
   assign m105_20 =10'b0;

   // m105_21 = W*in
   wire signed [9:0] m105_21;
   assign m105_21 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_22 = W*in
   wire signed [9:0] m105_22;
   assign m105_22 =10'b0;

   // m105_23 = W*in
   wire signed [9:0] m105_23;
   assign m105_23 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_24 = W*in
   wire signed [9:0] m105_24;
   assign m105_24 =10'b0;

   // m105_25 = W*in
   wire signed [9:0] m105_25;
   assign m105_25 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_26 = W*in
   wire signed [9:0] m105_26;
   assign m105_26 =10'b0;

   // m105_27 = W*in
   wire signed [9:0] m105_27;
   assign m105_27 =10'b0;

   // m105_28 = W*in
   wire signed [9:0] m105_28;
   assign m105_28 =10'b0;

   // m105_29 = W*in
   wire signed [9:0] m105_29;
   assign m105_29 =10'b0;

   // m105_30 = W*in
   wire signed [9:0] m105_30;
   assign m105_30 =10'b0;

   // m105_31 = W*in
   wire signed [9:0] m105_31;
   assign m105_31 =10'b0;

   // m105_32 = W*in
   wire signed [9:0] m105_32;
   assign m105_32 =10'b0;

   // m105_33 = W*in
   wire signed [9:0] m105_33;
   assign m105_33 =10'b0;

   // m105_34 = W*in
   wire signed [9:0] m105_34;
   assign m105_34 =10'b0;

   // m105_35 = W*in
   wire signed [9:0] m105_35;
   assign m105_35 =10'b0;

   // m105_36 = W*in
   wire signed [9:0] m105_36;
   assign m105_36 =10'b0;

   // m105_37 = W*in
   wire signed [9:0] m105_37;
   assign m105_37 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_38 = W*in
   wire signed [9:0] m105_38;
   assign m105_38 =10'b0;

   // m105_39 = W*in
   wire signed [9:0] m105_39;
   assign m105_39 =10'b0;

   // m105_40 = W*in
   wire signed [9:0] m105_40;
   assign m105_40 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_41 = W*in
   wire signed [9:0] m105_41;
   assign m105_41 =10'b0;

   // m105_42 = W*in
   wire signed [9:0] m105_42;
   assign m105_42 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_43 = W*in
   wire signed [9:0] m105_43;
   assign m105_43 =10'b0;

   // m105_44 = W*in
   wire signed [9:0] m105_44;
   assign m105_44 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_45 = W*in
   wire signed [9:0] m105_45;
   assign m105_45 =10'b0;

   // m105_46 = W*in
   wire signed [9:0] m105_46;
   assign m105_46 =10'b0;

   // m105_47 = W*in
   wire signed [9:0] m105_47;
   assign m105_47 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_48 = W*in
   wire signed [9:0] m105_48;
   assign m105_48 =10'b0;

   // m105_49 = W*in
   wire signed [9:0] m105_49;
   assign m105_49 =10'b0;

   // m105_50 = W*in
   wire signed [9:0] m105_50;
   assign m105_50 =10'b0;

   // m105_51 = W*in
   wire signed [9:0] m105_51;
   assign m105_51 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_52 = W*in
   wire signed [9:0] m105_52;
   assign m105_52 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_53 = W*in
   wire signed [9:0] m105_53;
   assign m105_53 =10'b0;

   // m105_54 = W*in
   wire signed [9:0] m105_54;
   assign m105_54 =10'b0;

   // m105_55 = W*in
   wire signed [9:0] m105_55;
   assign m105_55 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_56 = W*in
   wire signed [9:0] m105_56;
   assign m105_56 =10'b0;

   // m105_57 = W*in
   wire signed [9:0] m105_57;
   assign m105_57 =10'b0;

   // m105_58 = W*in
   wire signed [9:0] m105_58;
   assign m105_58 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_59 = W*in
   wire signed [9:0] m105_59;
   assign m105_59 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_60 = W*in
   wire signed [9:0] m105_60;
   assign m105_60 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_61 = W*in
   wire signed [9:0] m105_61;
   assign m105_61 =10'b0;

   // m105_62 = W*in
   wire signed [9:0] m105_62;
   assign m105_62 =10'b0;

   // m105_63 = W*in
   wire signed [9:0] m105_63;
   assign m105_63 =10'b0;

   // m105_64 = W*in
   wire signed [9:0] m105_64;
   assign m105_64 =10'b0;

   // m105_65 = W*in
   wire signed [9:0] m105_65;
   assign m105_65 =10'b0;

   // m105_66 = W*in
   wire signed [9:0] m105_66;
   assign m105_66 =10'b0;

   // m105_67 = W*in
   wire signed [9:0] m105_67;
   assign m105_67 =10'b0;

   // m105_68 = W*in
   wire signed [9:0] m105_68;
   assign m105_68 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_69 = W*in
   wire signed [9:0] m105_69;
   assign m105_69 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_70 = W*in
   wire signed [9:0] m105_70;
   assign m105_70 =10'b0;

   // m105_71 = W*in
   wire signed [9:0] m105_71;
   assign m105_71 =10'b0;

   // m105_72 = W*in
   wire signed [9:0] m105_72;
   assign m105_72 =10'b0;

   // m105_73 = W*in
   wire signed [9:0] m105_73;
   assign m105_73 =10'b0;

   // m105_74 = W*in
   wire signed [9:0] m105_74;
   assign m105_74 =10'b0;

   // m105_75 = W*in
   wire signed [9:0] m105_75;
   assign m105_75 =10'b0;

   // m105_76 = W*in
   wire signed [9:0] m105_76;
   assign m105_76 =10'b0;

   // m105_77 = W*in
   wire signed [9:0] m105_77;
   assign m105_77 ={ {3{neg105[5]}} , neg105 , {1{1'b0}} };

   // m105_78 = W*in
   wire signed [9:0] m105_78;
   assign m105_78 =10'b0;

   // m105_79 = W*in
   wire signed [9:0] m105_79;
   assign m105_79 ={ {3{in105[5]}} , in105 , {1{1'b0}} };

   // m105_80 = W*in
   wire signed [9:0] m105_80;
   assign m105_80 =10'b0;

   // m105_81 = W*in
   wire signed [9:0] m105_81;
   assign m105_81 =10'b0;

   // m106_1 = W*in
   wire signed [9:0] m106_1;
   assign m106_1 =10'b0;

   // m106_2 = W*in
   wire signed [9:0] m106_2;
   assign m106_2 =10'b0;

   // m106_3 = W*in
   wire signed [9:0] m106_3;
   assign m106_3 ={ {2{in106[5]}} , in106 , {2{1'b0}} };

   // m106_4 = W*in
   wire signed [9:0] m106_4;
   assign m106_4 =10'b0;

   // m106_5 = W*in
   wire signed [9:0] m106_5;
   assign m106_5 =10'b0;

   // m106_6 = W*in
   wire signed [9:0] m106_6;
   assign m106_6 =10'b0;

   // m106_7 = W*in
   wire signed [9:0] m106_7;
   assign m106_7 =10'b0;

   // m106_8 = W*in
   wire signed [9:0] m106_8;
   assign m106_8 =10'b0;

   // m106_9 = W*in
   wire signed [9:0] m106_9;
   assign m106_9 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_10 = W*in
   wire signed [9:0] m106_10;
   assign m106_10 =10'b0;

   // m106_11 = W*in
   wire signed [9:0] m106_11;
   assign m106_11 =10'b0;

   // m106_12 = W*in
   wire signed [9:0] m106_12;
   assign m106_12 =10'b0;

   // m106_13 = W*in
   wire signed [9:0] m106_13;
   assign m106_13 =10'b0;

   // m106_14 = W*in
   wire signed [9:0] m106_14;
   assign m106_14 =10'b0;

   // m106_15 = W*in
   wire signed [9:0] m106_15;
   assign m106_15 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_16 = W*in
   wire signed [9:0] m106_16;
   assign m106_16 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_17 = W*in
   wire signed [9:0] m106_17;
   assign m106_17 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_18 = W*in
   wire signed [9:0] m106_18;
   assign m106_18 =10'b0;

   // m106_19 = W*in
   wire signed [9:0] m106_19;
   assign m106_19 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_20 = W*in
   wire signed [9:0] m106_20;
   assign m106_20 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_21 = W*in
   wire signed [9:0] m106_21;
   assign m106_21 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_22 = W*in
   wire signed [9:0] m106_22;
   assign m106_22 =10'b0;

   // m106_23 = W*in
   wire signed [9:0] m106_23;
   assign m106_23 =10'b0;

   // m106_24 = W*in
   wire signed [9:0] m106_24;
   assign m106_24 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_25 = W*in
   wire signed [9:0] m106_25;
   assign m106_25 =10'b0;

   // m106_26 = W*in
   wire signed [9:0] m106_26;
   assign m106_26 =10'b0;

   // m106_27 = W*in
   wire signed [9:0] m106_27;
   assign m106_27 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_28 = W*in
   wire signed [9:0] m106_28;
   assign m106_28 =10'b0;

   // m106_29 = W*in
   wire signed [9:0] m106_29;
   assign m106_29 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_30 = W*in
   wire signed [9:0] m106_30;
   assign m106_30 ={ {2{in106[5]}} , in106 , {2{1'b0}} };

   // m106_31 = W*in
   wire signed [9:0] m106_31;
   assign m106_31 =10'b0;

   // m106_32 = W*in
   wire signed [9:0] m106_32;
   assign m106_32 =10'b0;

   // m106_33 = W*in
   wire signed [9:0] m106_33;
   assign m106_33 =10'b0;

   // m106_34 = W*in
   wire signed [9:0] m106_34;
   assign m106_34 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_35 = W*in
   wire signed [9:0] m106_35;
   assign m106_35 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_36 = W*in
   wire signed [9:0] m106_36;
   assign m106_36 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_37 = W*in
   wire signed [9:0] m106_37;
   assign m106_37 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_38 = W*in
   wire signed [9:0] m106_38;
   assign m106_38 =10'b0;

   // m106_39 = W*in
   wire signed [9:0] m106_39;
   assign m106_39 =10'b0;

   // m106_40 = W*in
   wire signed [9:0] m106_40;
   assign m106_40 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_41 = W*in
   wire signed [9:0] m106_41;
   assign m106_41 =10'b0;

   // m106_42 = W*in
   wire signed [9:0] m106_42;
   assign m106_42 =10'b0;

   // m106_43 = W*in
   wire signed [9:0] m106_43;
   assign m106_43 =10'b0;

   // m106_44 = W*in
   wire signed [9:0] m106_44;
   assign m106_44 =10'b0;

   // m106_45 = W*in
   wire signed [9:0] m106_45;
   assign m106_45 =10'b0;

   // m106_46 = W*in
   wire signed [9:0] m106_46;
   assign m106_46 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_47 = W*in
   wire signed [9:0] m106_47;
   assign m106_47 =10'b0;

   // m106_48 = W*in
   wire signed [9:0] m106_48;
   assign m106_48 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_49 = W*in
   wire signed [9:0] m106_49;
   assign m106_49 =10'b0;

   // m106_50 = W*in
   wire signed [9:0] m106_50;
   assign m106_50 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_51 = W*in
   wire signed [9:0] m106_51;
   assign m106_51 =10'b0;

   // m106_52 = W*in
   wire signed [9:0] m106_52;
   assign m106_52 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_53 = W*in
   wire signed [9:0] m106_53;
   assign m106_53 =10'b0;

   // m106_54 = W*in
   wire signed [9:0] m106_54;
   assign m106_54 =10'b0;

   // m106_55 = W*in
   wire signed [9:0] m106_55;
   assign m106_55 =10'b0;

   // m106_56 = W*in
   wire signed [9:0] m106_56;
   assign m106_56 =10'b0;

   // m106_57 = W*in
   wire signed [9:0] m106_57;
   assign m106_57 =10'b0;

   // m106_58 = W*in
   wire signed [9:0] m106_58;
   assign m106_58 =10'b0;

   // m106_59 = W*in
   wire signed [9:0] m106_59;
   assign m106_59 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_60 = W*in
   wire signed [9:0] m106_60;
   assign m106_60 =10'b0;

   // m106_61 = W*in
   wire signed [9:0] m106_61;
   assign m106_61 =10'b0;

   // m106_62 = W*in
   wire signed [9:0] m106_62;
   assign m106_62 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_63 = W*in
   wire signed [9:0] m106_63;
   assign m106_63 =10'b0;

   // m106_64 = W*in
   wire signed [9:0] m106_64;
   assign m106_64 =10'b0;

   // m106_65 = W*in
   wire signed [9:0] m106_65;
   assign m106_65 =10'b0;

   // m106_66 = W*in
   wire signed [9:0] m106_66;
   assign m106_66 =10'b0;

   // m106_67 = W*in
   wire signed [9:0] m106_67;
   assign m106_67 =10'b0;

   // m106_68 = W*in
   wire signed [9:0] m106_68;
   assign m106_68 =10'b0;

   // m106_69 = W*in
   wire signed [9:0] m106_69;
   assign m106_69 =10'b0;

   // m106_70 = W*in
   wire signed [9:0] m106_70;
   assign m106_70 =10'b0;

   // m106_71 = W*in
   wire signed [9:0] m106_71;
   assign m106_71 =10'b0;

   // m106_72 = W*in
   wire signed [9:0] m106_72;
   assign m106_72 =10'b0;

   // m106_73 = W*in
   wire signed [9:0] m106_73;
   assign m106_73 =10'b0;

   // m106_74 = W*in
   wire signed [9:0] m106_74;
   assign m106_74 =10'b0;

   // m106_75 = W*in
   wire signed [9:0] m106_75;
   assign m106_75 =10'b0;

   // m106_76 = W*in
   wire signed [9:0] m106_76;
   assign m106_76 =10'b0;

   // m106_77 = W*in
   wire signed [9:0] m106_77;
   assign m106_77 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_78 = W*in
   wire signed [9:0] m106_78;
   assign m106_78 =10'b0;

   // m106_79 = W*in
   wire signed [9:0] m106_79;
   assign m106_79 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_80 = W*in
   wire signed [9:0] m106_80;
   assign m106_80 =10'b0;

   // m106_81 = W*in
   wire signed [9:0] m106_81;
   assign m106_81 ={ {2{in106[5]}} , in106 , {2{1'b0}} };

   // m107_1 = W*in
   wire signed [9:0] m107_1;
   assign m107_1 =10'b0;

   // m107_2 = W*in
   wire signed [9:0] m107_2;
   assign m107_2 =10'b0;

   // m107_3 = W*in
   wire signed [9:0] m107_3;
   assign m107_3 =10'b0;

   // m107_4 = W*in
   wire signed [9:0] m107_4;
   assign m107_4 =10'b0;

   // m107_5 = W*in
   wire signed [9:0] m107_5;
   assign m107_5 =10'b0;

   // m107_6 = W*in
   wire signed [9:0] m107_6;
   assign m107_6 =10'b0;

   // m107_7 = W*in
   wire signed [9:0] m107_7;
   assign m107_7 =10'b0;

   // m107_8 = W*in
   wire signed [9:0] m107_8;
   assign m107_8 =10'b0;

   // m107_9 = W*in
   wire signed [9:0] m107_9;
   assign m107_9 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_10 = W*in
   wire signed [9:0] m107_10;
   assign m107_10 =10'b0;

   // m107_11 = W*in
   wire signed [9:0] m107_11;
   assign m107_11 =10'b0;

   // m107_12 = W*in
   wire signed [9:0] m107_12;
   assign m107_12 =10'b0;

   // m107_13 = W*in
   wire signed [9:0] m107_13;
   assign m107_13 =10'b0;

   // m107_14 = W*in
   wire signed [9:0] m107_14;
   assign m107_14 =10'b0;

   // m107_15 = W*in
   wire signed [9:0] m107_15;
   assign m107_15 ={ {2{in107[5]}} , in107 , {2{1'b0}} };

   // m107_16 = W*in
   wire signed [9:0] m107_16;
   assign m107_16 =10'b0;

   // m107_17 = W*in
   wire signed [9:0] m107_17;
   assign m107_17 =10'b0;

   // m107_18 = W*in
   wire signed [9:0] m107_18;
   assign m107_18 =10'b0;

   // m107_19 = W*in
   wire signed [9:0] m107_19;
   assign m107_19 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_20 = W*in
   wire signed [9:0] m107_20;
   assign m107_20 =10'b0;

   // m107_21 = W*in
   wire signed [9:0] m107_21;
   assign m107_21 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_22 = W*in
   wire signed [9:0] m107_22;
   assign m107_22 =10'b0;

   // m107_23 = W*in
   wire signed [9:0] m107_23;
   assign m107_23 =10'b0;

   // m107_24 = W*in
   wire signed [9:0] m107_24;
   assign m107_24 =10'b0;

   // m107_25 = W*in
   wire signed [9:0] m107_25;
   assign m107_25 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_26 = W*in
   wire signed [9:0] m107_26;
   assign m107_26 =10'b0;

   // m107_27 = W*in
   wire signed [9:0] m107_27;
   assign m107_27 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_28 = W*in
   wire signed [9:0] m107_28;
   assign m107_28 =10'b0;

   // m107_29 = W*in
   wire signed [9:0] m107_29;
   assign m107_29 =10'b0;

   // m107_30 = W*in
   wire signed [9:0] m107_30;
   assign m107_30 =10'b0;

   // m107_31 = W*in
   wire signed [9:0] m107_31;
   assign m107_31 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_32 = W*in
   wire signed [9:0] m107_32;
   assign m107_32 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_33 = W*in
   wire signed [9:0] m107_33;
   assign m107_33 =10'b0;

   // m107_34 = W*in
   wire signed [9:0] m107_34;
   assign m107_34 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_35 = W*in
   wire signed [9:0] m107_35;
   assign m107_35 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_36 = W*in
   wire signed [9:0] m107_36;
   assign m107_36 =10'b0;

   // m107_37 = W*in
   wire signed [9:0] m107_37;
   assign m107_37 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_38 = W*in
   wire signed [9:0] m107_38;
   assign m107_38 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_39 = W*in
   wire signed [9:0] m107_39;
   assign m107_39 =10'b0;

   // m107_40 = W*in
   wire signed [9:0] m107_40;
   assign m107_40 ={ {2{in107[5]}} , in107 , {2{1'b0}} };

   // m107_41 = W*in
   wire signed [9:0] m107_41;
   assign m107_41 =10'b0;

   // m107_42 = W*in
   wire signed [9:0] m107_42;
   assign m107_42 =10'b0;

   // m107_43 = W*in
   wire signed [9:0] m107_43;
   assign m107_43 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_44 = W*in
   wire signed [9:0] m107_44;
   assign m107_44 =10'b0;

   // m107_45 = W*in
   wire signed [9:0] m107_45;
   assign m107_45 =10'b0;

   // m107_46 = W*in
   wire signed [9:0] m107_46;
   assign m107_46 =10'b0;

   // m107_47 = W*in
   wire signed [9:0] m107_47;
   assign m107_47 ={ {2{in107[5]}} , in107 , {2{1'b0}} };

   // m107_48 = W*in
   wire signed [9:0] m107_48;
   assign m107_48 =10'b0;

   // m107_49 = W*in
   wire signed [9:0] m107_49;
   assign m107_49 =10'b0;

   // m107_50 = W*in
   wire signed [9:0] m107_50;
   assign m107_50 =10'b0;

   // m107_51 = W*in
   wire signed [9:0] m107_51;
   assign m107_51 =10'b0;

   // m107_52 = W*in
   wire signed [9:0] m107_52;
   assign m107_52 =10'b0;

   // m107_53 = W*in
   wire signed [9:0] m107_53;
   assign m107_53 =10'b0;

   // m107_54 = W*in
   wire signed [9:0] m107_54;
   assign m107_54 =10'b0;

   // m107_55 = W*in
   wire signed [9:0] m107_55;
   assign m107_55 ={ {2{in107[5]}} , in107 , {2{1'b0}} };

   // m107_56 = W*in
   wire signed [9:0] m107_56;
   assign m107_56 =10'b0;

   // m107_57 = W*in
   wire signed [9:0] m107_57;
   assign m107_57 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_58 = W*in
   wire signed [9:0] m107_58;
   assign m107_58 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_59 = W*in
   wire signed [9:0] m107_59;
   assign m107_59 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_60 = W*in
   wire signed [9:0] m107_60;
   assign m107_60 =10'b0;

   // m107_61 = W*in
   wire signed [9:0] m107_61;
   assign m107_61 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_62 = W*in
   wire signed [9:0] m107_62;
   assign m107_62 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_63 = W*in
   wire signed [9:0] m107_63;
   assign m107_63 =10'b0;

   // m107_64 = W*in
   wire signed [9:0] m107_64;
   assign m107_64 =10'b0;

   // m107_65 = W*in
   wire signed [9:0] m107_65;
   assign m107_65 =10'b0;

   // m107_66 = W*in
   wire signed [9:0] m107_66;
   assign m107_66 =10'b0;

   // m107_67 = W*in
   wire signed [9:0] m107_67;
   assign m107_67 =10'b0;

   // m107_68 = W*in
   wire signed [9:0] m107_68;
   assign m107_68 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_69 = W*in
   wire signed [9:0] m107_69;
   assign m107_69 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_70 = W*in
   wire signed [9:0] m107_70;
   assign m107_70 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_71 = W*in
   wire signed [9:0] m107_71;
   assign m107_71 =10'b0;

   // m107_72 = W*in
   wire signed [9:0] m107_72;
   assign m107_72 =10'b0;

   // m107_73 = W*in
   wire signed [9:0] m107_73;
   assign m107_73 =10'b0;

   // m107_74 = W*in
   wire signed [9:0] m107_74;
   assign m107_74 ={ {2{in107[5]}} , in107 , {2{1'b0}} };

   // m107_75 = W*in
   wire signed [9:0] m107_75;
   assign m107_75 =10'b0;

   // m107_76 = W*in
   wire signed [9:0] m107_76;
   assign m107_76 =10'b0;

   // m107_77 = W*in
   wire signed [9:0] m107_77;
   assign m107_77 ={ {3{neg107[5]}} , neg107 , {1{1'b0}} };

   // m107_78 = W*in
   wire signed [9:0] m107_78;
   assign m107_78 =10'b0;

   // m107_79 = W*in
   wire signed [9:0] m107_79;
   assign m107_79 =10'b0;

   // m107_80 = W*in
   wire signed [9:0] m107_80;
   assign m107_80 =10'b0;

   // m107_81 = W*in
   wire signed [9:0] m107_81;
   assign m107_81 =10'b0;

   // m108_1 = W*in
   wire signed [9:0] m108_1;
   assign m108_1 ={ {2{in108[5]}} , in108 , {2{1'b0}} };

   // m108_2 = W*in
   wire signed [9:0] m108_2;
   assign m108_2 =10'b0;

   // m108_3 = W*in
   wire signed [9:0] m108_3;
   assign m108_3 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_4 = W*in
   wire signed [9:0] m108_4;
   assign m108_4 =10'b0;

   // m108_5 = W*in
   wire signed [9:0] m108_5;
   assign m108_5 =10'b0;

   // m108_6 = W*in
   wire signed [9:0] m108_6;
   assign m108_6 ={ {2{neg108[5]}} , neg108 , {2{1'b0}} };

   // m108_7 = W*in
   wire signed [9:0] m108_7;
   assign m108_7 =10'b0;

   // m108_8 = W*in
   wire signed [9:0] m108_8;
   assign m108_8 =10'b0;

   // m108_9 = W*in
   wire signed [9:0] m108_9;
   assign m108_9 =10'b0;

   // m108_10 = W*in
   wire signed [9:0] m108_10;
   assign m108_10 =10'b0;

   // m108_11 = W*in
   wire signed [9:0] m108_11;
   assign m108_11 =10'b0;

   // m108_12 = W*in
   wire signed [9:0] m108_12;
   assign m108_12 =10'b0;

   // m108_13 = W*in
   wire signed [9:0] m108_13;
   assign m108_13 =10'b0;

   // m108_14 = W*in
   wire signed [9:0] m108_14;
   assign m108_14 =10'b0;

   // m108_15 = W*in
   wire signed [9:0] m108_15;
   assign m108_15 =10'b0;

   // m108_16 = W*in
   wire signed [9:0] m108_16;
   assign m108_16 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_17 = W*in
   wire signed [9:0] m108_17;
   assign m108_17 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_18 = W*in
   wire signed [9:0] m108_18;
   assign m108_18 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_19 = W*in
   wire signed [9:0] m108_19;
   assign m108_19 =10'b0;

   // m108_20 = W*in
   wire signed [9:0] m108_20;
   assign m108_20 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_21 = W*in
   wire signed [9:0] m108_21;
   assign m108_21 =10'b0;

   // m108_22 = W*in
   wire signed [9:0] m108_22;
   assign m108_22 =10'b0;

   // m108_23 = W*in
   wire signed [9:0] m108_23;
   assign m108_23 =10'b0;

   // m108_24 = W*in
   wire signed [9:0] m108_24;
   assign m108_24 =10'b0;

   // m108_25 = W*in
   wire signed [9:0] m108_25;
   assign m108_25 =10'b0;

   // m108_26 = W*in
   wire signed [9:0] m108_26;
   assign m108_26 =10'b0;

   // m108_27 = W*in
   wire signed [9:0] m108_27;
   assign m108_27 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_28 = W*in
   wire signed [9:0] m108_28;
   assign m108_28 =10'b0;

   // m108_29 = W*in
   wire signed [9:0] m108_29;
   assign m108_29 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_30 = W*in
   wire signed [9:0] m108_30;
   assign m108_30 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_31 = W*in
   wire signed [9:0] m108_31;
   assign m108_31 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_32 = W*in
   wire signed [9:0] m108_32;
   assign m108_32 =10'b0;

   // m108_33 = W*in
   wire signed [9:0] m108_33;
   assign m108_33 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_34 = W*in
   wire signed [9:0] m108_34;
   assign m108_34 =10'b0;

   // m108_35 = W*in
   wire signed [9:0] m108_35;
   assign m108_35 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_36 = W*in
   wire signed [9:0] m108_36;
   assign m108_36 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_37 = W*in
   wire signed [9:0] m108_37;
   assign m108_37 =10'b0;

   // m108_38 = W*in
   wire signed [9:0] m108_38;
   assign m108_38 =10'b0;

   // m108_39 = W*in
   wire signed [9:0] m108_39;
   assign m108_39 =10'b0;

   // m108_40 = W*in
   wire signed [9:0] m108_40;
   assign m108_40 =10'b0;

   // m108_41 = W*in
   wire signed [9:0] m108_41;
   assign m108_41 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_42 = W*in
   wire signed [9:0] m108_42;
   assign m108_42 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_43 = W*in
   wire signed [9:0] m108_43;
   assign m108_43 =10'b0;

   // m108_44 = W*in
   wire signed [9:0] m108_44;
   assign m108_44 =10'b0;

   // m108_45 = W*in
   wire signed [9:0] m108_45;
   assign m108_45 =10'b0;

   // m108_46 = W*in
   wire signed [9:0] m108_46;
   assign m108_46 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_47 = W*in
   wire signed [9:0] m108_47;
   assign m108_47 =10'b0;

   // m108_48 = W*in
   wire signed [9:0] m108_48;
   assign m108_48 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_49 = W*in
   wire signed [9:0] m108_49;
   assign m108_49 ={ {2{neg108[5]}} , neg108 , {2{1'b0}} };

   // m108_50 = W*in
   wire signed [9:0] m108_50;
   assign m108_50 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_51 = W*in
   wire signed [9:0] m108_51;
   assign m108_51 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_52 = W*in
   wire signed [9:0] m108_52;
   assign m108_52 =10'b0;

   // m108_53 = W*in
   wire signed [9:0] m108_53;
   assign m108_53 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_54 = W*in
   wire signed [9:0] m108_54;
   assign m108_54 =10'b0;

   // m108_55 = W*in
   wire signed [9:0] m108_55;
   assign m108_55 =10'b0;

   // m108_56 = W*in
   wire signed [9:0] m108_56;
   assign m108_56 ={ {2{neg108[5]}} , neg108 , {2{1'b0}} };

   // m108_57 = W*in
   wire signed [9:0] m108_57;
   assign m108_57 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_58 = W*in
   wire signed [9:0] m108_58;
   assign m108_58 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_59 = W*in
   wire signed [9:0] m108_59;
   assign m108_59 =10'b0;

   // m108_60 = W*in
   wire signed [9:0] m108_60;
   assign m108_60 =10'b0;

   // m108_61 = W*in
   wire signed [9:0] m108_61;
   assign m108_61 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_62 = W*in
   wire signed [9:0] m108_62;
   assign m108_62 =10'b0;

   // m108_63 = W*in
   wire signed [9:0] m108_63;
   assign m108_63 =10'b0;

   // m108_64 = W*in
   wire signed [9:0] m108_64;
   assign m108_64 =10'b0;

   // m108_65 = W*in
   wire signed [9:0] m108_65;
   assign m108_65 =10'b0;

   // m108_66 = W*in
   wire signed [9:0] m108_66;
   assign m108_66 =10'b0;

   // m108_67 = W*in
   wire signed [9:0] m108_67;
   assign m108_67 =10'b0;

   // m108_68 = W*in
   wire signed [9:0] m108_68;
   assign m108_68 ={ {3{neg108[5]}} , neg108 , {1{1'b0}} };

   // m108_69 = W*in
   wire signed [9:0] m108_69;
   assign m108_69 =10'b0;

   // m108_70 = W*in
   wire signed [9:0] m108_70;
   assign m108_70 =10'b0;

   // m108_71 = W*in
   wire signed [9:0] m108_71;
   assign m108_71 =10'b0;

   // m108_72 = W*in
   wire signed [9:0] m108_72;
   assign m108_72 ={ {2{in108[5]}} , in108 , {2{1'b0}} };

   // m108_73 = W*in
   wire signed [9:0] m108_73;
   assign m108_73 =10'b0;

   // m108_74 = W*in
   wire signed [9:0] m108_74;
   assign m108_74 =10'b0;

   // m108_75 = W*in
   wire signed [9:0] m108_75;
   assign m108_75 =10'b0;

   // m108_76 = W*in
   wire signed [9:0] m108_76;
   assign m108_76 =10'b0;

   // m108_77 = W*in
   wire signed [9:0] m108_77;
   assign m108_77 =10'b0;

   // m108_78 = W*in
   wire signed [9:0] m108_78;
   assign m108_78 ={ {2{in108[5]}} , in108 , {2{1'b0}} };

   // m108_79 = W*in
   wire signed [9:0] m108_79;
   assign m108_79 ={ {3{in108[5]}} , in108 , {1{1'b0}} };

   // m108_80 = W*in
   wire signed [9:0] m108_80;
   assign m108_80 =10'b0;

   // m108_81 = W*in
   wire signed [9:0] m108_81;
   assign m108_81 =10'b0;

   // m109_1 = W*in
   wire signed [9:0] m109_1;
   assign m109_1 =10'b0;

   // m109_2 = W*in
   wire signed [9:0] m109_2;
   assign m109_2 =10'b0;

   // m109_3 = W*in
   wire signed [9:0] m109_3;
   assign m109_3 ={ {2{in109[5]}} , in109 , {2{1'b0}} };

   // m109_4 = W*in
   wire signed [9:0] m109_4;
   assign m109_4 =10'b0;

   // m109_5 = W*in
   wire signed [9:0] m109_5;
   assign m109_5 =10'b0;

   // m109_6 = W*in
   wire signed [9:0] m109_6;
   assign m109_6 ={ {2{neg109[5]}} , neg109 , {2{1'b0}} };

   // m109_7 = W*in
   wire signed [9:0] m109_7;
   assign m109_7 =10'b0;

   // m109_8 = W*in
   wire signed [9:0] m109_8;
   assign m109_8 =10'b0;

   // m109_9 = W*in
   wire signed [9:0] m109_9;
   assign m109_9 =10'b0;

   // m109_10 = W*in
   wire signed [9:0] m109_10;
   assign m109_10 =10'b0;

   // m109_11 = W*in
   wire signed [9:0] m109_11;
   assign m109_11 =10'b0;

   // m109_12 = W*in
   wire signed [9:0] m109_12;
   assign m109_12 =10'b0;

   // m109_13 = W*in
   wire signed [9:0] m109_13;
   assign m109_13 =10'b0;

   // m109_14 = W*in
   wire signed [9:0] m109_14;
   assign m109_14 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_15 = W*in
   wire signed [9:0] m109_15;
   assign m109_15 =10'b0;

   // m109_16 = W*in
   wire signed [9:0] m109_16;
   assign m109_16 =10'b0;

   // m109_17 = W*in
   wire signed [9:0] m109_17;
   assign m109_17 ={ {3{neg109[5]}} , neg109 , {1{1'b0}} };

   // m109_18 = W*in
   wire signed [9:0] m109_18;
   assign m109_18 =10'b0;

   // m109_19 = W*in
   wire signed [9:0] m109_19;
   assign m109_19 =10'b0;

   // m109_20 = W*in
   wire signed [9:0] m109_20;
   assign m109_20 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_21 = W*in
   wire signed [9:0] m109_21;
   assign m109_21 =10'b0;

   // m109_22 = W*in
   wire signed [9:0] m109_22;
   assign m109_22 =10'b0;

   // m109_23 = W*in
   wire signed [9:0] m109_23;
   assign m109_23 =10'b0;

   // m109_24 = W*in
   wire signed [9:0] m109_24;
   assign m109_24 =10'b0;

   // m109_25 = W*in
   wire signed [9:0] m109_25;
   assign m109_25 =10'b0;

   // m109_26 = W*in
   wire signed [9:0] m109_26;
   assign m109_26 =10'b0;

   // m109_27 = W*in
   wire signed [9:0] m109_27;
   assign m109_27 =10'b0;

   // m109_28 = W*in
   wire signed [9:0] m109_28;
   assign m109_28 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_29 = W*in
   wire signed [9:0] m109_29;
   assign m109_29 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_30 = W*in
   wire signed [9:0] m109_30;
   assign m109_30 =10'b0;

   // m109_31 = W*in
   wire signed [9:0] m109_31;
   assign m109_31 =10'b0;

   // m109_32 = W*in
   wire signed [9:0] m109_32;
   assign m109_32 =10'b0;

   // m109_33 = W*in
   wire signed [9:0] m109_33;
   assign m109_33 ={ {3{neg109[5]}} , neg109 , {1{1'b0}} };

   // m109_34 = W*in
   wire signed [9:0] m109_34;
   assign m109_34 =10'b0;

   // m109_35 = W*in
   wire signed [9:0] m109_35;
   assign m109_35 ={ {2{in109[5]}} , in109 , {2{1'b0}} };

   // m109_36 = W*in
   wire signed [9:0] m109_36;
   assign m109_36 =10'b0;

   // m109_37 = W*in
   wire signed [9:0] m109_37;
   assign m109_37 =10'b0;

   // m109_38 = W*in
   wire signed [9:0] m109_38;
   assign m109_38 =10'b0;

   // m109_39 = W*in
   wire signed [9:0] m109_39;
   assign m109_39 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_40 = W*in
   wire signed [9:0] m109_40;
   assign m109_40 =10'b0;

   // m109_41 = W*in
   wire signed [9:0] m109_41;
   assign m109_41 =10'b0;

   // m109_42 = W*in
   wire signed [9:0] m109_42;
   assign m109_42 =10'b0;

   // m109_43 = W*in
   wire signed [9:0] m109_43;
   assign m109_43 =10'b0;

   // m109_44 = W*in
   wire signed [9:0] m109_44;
   assign m109_44 =10'b0;

   // m109_45 = W*in
   wire signed [9:0] m109_45;
   assign m109_45 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_46 = W*in
   wire signed [9:0] m109_46;
   assign m109_46 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_47 = W*in
   wire signed [9:0] m109_47;
   assign m109_47 =10'b0;

   // m109_48 = W*in
   wire signed [9:0] m109_48;
   assign m109_48 =10'b0;

   // m109_49 = W*in
   wire signed [9:0] m109_49;
   assign m109_49 ={ {3{neg109[5]}} , neg109 , {1{1'b0}} };

   // m109_50 = W*in
   wire signed [9:0] m109_50;
   assign m109_50 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_51 = W*in
   wire signed [9:0] m109_51;
   assign m109_51 =10'b0;

   // m109_52 = W*in
   wire signed [9:0] m109_52;
   assign m109_52 =10'b0;

   // m109_53 = W*in
   wire signed [9:0] m109_53;
   assign m109_53 ={ {2{neg109[5]}} , neg109 , {2{1'b0}} };

   // m109_54 = W*in
   wire signed [9:0] m109_54;
   assign m109_54 =10'b0;

   // m109_55 = W*in
   wire signed [9:0] m109_55;
   assign m109_55 =10'b0;

   // m109_56 = W*in
   wire signed [9:0] m109_56;
   assign m109_56 ={ {2{neg109[5]}} , neg109 , {2{1'b0}} };

   // m109_57 = W*in
   wire signed [9:0] m109_57;
   assign m109_57 ={ {3{neg109[5]}} , neg109 , {1{1'b0}} };

   // m109_58 = W*in
   wire signed [9:0] m109_58;
   assign m109_58 ={ {3{neg109[5]}} , neg109 , {1{1'b0}} };

   // m109_59 = W*in
   wire signed [9:0] m109_59;
   assign m109_59 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_60 = W*in
   wire signed [9:0] m109_60;
   assign m109_60 =10'b0;

   // m109_61 = W*in
   wire signed [9:0] m109_61;
   assign m109_61 =10'b0;

   // m109_62 = W*in
   wire signed [9:0] m109_62;
   assign m109_62 =10'b0;

   // m109_63 = W*in
   wire signed [9:0] m109_63;
   assign m109_63 =10'b0;

   // m109_64 = W*in
   wire signed [9:0] m109_64;
   assign m109_64 =10'b0;

   // m109_65 = W*in
   wire signed [9:0] m109_65;
   assign m109_65 ={ {2{in109[5]}} , in109 , {2{1'b0}} };

   // m109_66 = W*in
   wire signed [9:0] m109_66;
   assign m109_66 =10'b0;

   // m109_67 = W*in
   wire signed [9:0] m109_67;
   assign m109_67 =10'b0;

   // m109_68 = W*in
   wire signed [9:0] m109_68;
   assign m109_68 ={ {2{neg109[5]}} , neg109 , {2{1'b0}} };

   // m109_69 = W*in
   wire signed [9:0] m109_69;
   assign m109_69 =10'b0;

   // m109_70 = W*in
   wire signed [9:0] m109_70;
   assign m109_70 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_71 = W*in
   wire signed [9:0] m109_71;
   assign m109_71 =10'b0;

   // m109_72 = W*in
   wire signed [9:0] m109_72;
   assign m109_72 ={ {2{in109[5]}} , in109 , {2{1'b0}} };

   // m109_73 = W*in
   wire signed [9:0] m109_73;
   assign m109_73 =10'b0;

   // m109_74 = W*in
   wire signed [9:0] m109_74;
   assign m109_74 =10'b0;

   // m109_75 = W*in
   wire signed [9:0] m109_75;
   assign m109_75 =10'b0;

   // m109_76 = W*in
   wire signed [9:0] m109_76;
   assign m109_76 =10'b0;

   // m109_77 = W*in
   wire signed [9:0] m109_77;
   assign m109_77 ={ {3{neg109[5]}} , neg109 , {1{1'b0}} };

   // m109_78 = W*in
   wire signed [9:0] m109_78;
   assign m109_78 ={ {2{in109[5]}} , in109 , {2{1'b0}} };

   // m109_79 = W*in
   wire signed [9:0] m109_79;
   assign m109_79 ={ {3{in109[5]}} , in109 , {1{1'b0}} };

   // m109_80 = W*in
   wire signed [9:0] m109_80;
   assign m109_80 =10'b0;

   // m109_81 = W*in
   wire signed [9:0] m109_81;
   assign m109_81 =10'b0;

   // m110_1 = W*in
   wire signed [9:0] m110_1;
   assign m110_1 =10'b0;

   // m110_2 = W*in
   wire signed [9:0] m110_2;
   assign m110_2 =10'b0;

   // m110_3 = W*in
   wire signed [9:0] m110_3;
   assign m110_3 ={ {3{neg110[5]}} , neg110 , {1{1'b0}} };

   // m110_4 = W*in
   wire signed [9:0] m110_4;
   assign m110_4 =10'b0;

   // m110_5 = W*in
   wire signed [9:0] m110_5;
   assign m110_5 =10'b0;

   // m110_6 = W*in
   wire signed [9:0] m110_6;
   assign m110_6 =10'b0;

   // m110_7 = W*in
   wire signed [9:0] m110_7;
   assign m110_7 =10'b0;

   // m110_8 = W*in
   wire signed [9:0] m110_8;
   assign m110_8 =10'b0;

   // m110_9 = W*in
   wire signed [9:0] m110_9;
   assign m110_9 =10'b0;

   // m110_10 = W*in
   wire signed [9:0] m110_10;
   assign m110_10 =10'b0;

   // m110_11 = W*in
   wire signed [9:0] m110_11;
   assign m110_11 =10'b0;

   // m110_12 = W*in
   wire signed [9:0] m110_12;
   assign m110_12 =10'b0;

   // m110_13 = W*in
   wire signed [9:0] m110_13;
   assign m110_13 =10'b0;

   // m110_14 = W*in
   wire signed [9:0] m110_14;
   assign m110_14 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_15 = W*in
   wire signed [9:0] m110_15;
   assign m110_15 =10'b0;

   // m110_16 = W*in
   wire signed [9:0] m110_16;
   assign m110_16 =10'b0;

   // m110_17 = W*in
   wire signed [9:0] m110_17;
   assign m110_17 =10'b0;

   // m110_18 = W*in
   wire signed [9:0] m110_18;
   assign m110_18 =10'b0;

   // m110_19 = W*in
   wire signed [9:0] m110_19;
   assign m110_19 =10'b0;

   // m110_20 = W*in
   wire signed [9:0] m110_20;
   assign m110_20 =10'b0;

   // m110_21 = W*in
   wire signed [9:0] m110_21;
   assign m110_21 =10'b0;

   // m110_22 = W*in
   wire signed [9:0] m110_22;
   assign m110_22 =10'b0;

   // m110_23 = W*in
   wire signed [9:0] m110_23;
   assign m110_23 =10'b0;

   // m110_24 = W*in
   wire signed [9:0] m110_24;
   assign m110_24 =10'b0;

   // m110_25 = W*in
   wire signed [9:0] m110_25;
   assign m110_25 =10'b0;

   // m110_26 = W*in
   wire signed [9:0] m110_26;
   assign m110_26 =10'b0;

   // m110_27 = W*in
   wire signed [9:0] m110_27;
   assign m110_27 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_28 = W*in
   wire signed [9:0] m110_28;
   assign m110_28 =10'b0;

   // m110_29 = W*in
   wire signed [9:0] m110_29;
   assign m110_29 =10'b0;

   // m110_30 = W*in
   wire signed [9:0] m110_30;
   assign m110_30 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_31 = W*in
   wire signed [9:0] m110_31;
   assign m110_31 ={ {2{in110[5]}} , in110 , {2{1'b0}} };

   // m110_32 = W*in
   wire signed [9:0] m110_32;
   assign m110_32 =10'b0;

   // m110_33 = W*in
   wire signed [9:0] m110_33;
   assign m110_33 =10'b0;

   // m110_34 = W*in
   wire signed [9:0] m110_34;
   assign m110_34 ={ {2{in110[5]}} , in110 , {2{1'b0}} };

   // m110_35 = W*in
   wire signed [9:0] m110_35;
   assign m110_35 =10'b0;

   // m110_36 = W*in
   wire signed [9:0] m110_36;
   assign m110_36 =10'b0;

   // m110_37 = W*in
   wire signed [9:0] m110_37;
   assign m110_37 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_38 = W*in
   wire signed [9:0] m110_38;
   assign m110_38 =10'b0;

   // m110_39 = W*in
   wire signed [9:0] m110_39;
   assign m110_39 =10'b0;

   // m110_40 = W*in
   wire signed [9:0] m110_40;
   assign m110_40 ={ {3{neg110[5]}} , neg110 , {1{1'b0}} };

   // m110_41 = W*in
   wire signed [9:0] m110_41;
   assign m110_41 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_42 = W*in
   wire signed [9:0] m110_42;
   assign m110_42 =10'b0;

   // m110_43 = W*in
   wire signed [9:0] m110_43;
   assign m110_43 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_44 = W*in
   wire signed [9:0] m110_44;
   assign m110_44 =10'b0;

   // m110_45 = W*in
   wire signed [9:0] m110_45;
   assign m110_45 =10'b0;

   // m110_46 = W*in
   wire signed [9:0] m110_46;
   assign m110_46 =10'b0;

   // m110_47 = W*in
   wire signed [9:0] m110_47;
   assign m110_47 =10'b0;

   // m110_48 = W*in
   wire signed [9:0] m110_48;
   assign m110_48 =10'b0;

   // m110_49 = W*in
   wire signed [9:0] m110_49;
   assign m110_49 =10'b0;

   // m110_50 = W*in
   wire signed [9:0] m110_50;
   assign m110_50 =10'b0;

   // m110_51 = W*in
   wire signed [9:0] m110_51;
   assign m110_51 ={ {2{in110[5]}} , in110 , {2{1'b0}} };

   // m110_52 = W*in
   wire signed [9:0] m110_52;
   assign m110_52 =10'b0;

   // m110_53 = W*in
   wire signed [9:0] m110_53;
   assign m110_53 =10'b0;

   // m110_54 = W*in
   wire signed [9:0] m110_54;
   assign m110_54 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_55 = W*in
   wire signed [9:0] m110_55;
   assign m110_55 ={ {3{neg110[5]}} , neg110 , {1{1'b0}} };

   // m110_56 = W*in
   wire signed [9:0] m110_56;
   assign m110_56 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_57 = W*in
   wire signed [9:0] m110_57;
   assign m110_57 =10'b0;

   // m110_58 = W*in
   wire signed [9:0] m110_58;
   assign m110_58 =10'b0;

   // m110_59 = W*in
   wire signed [9:0] m110_59;
   assign m110_59 =10'b0;

   // m110_60 = W*in
   wire signed [9:0] m110_60;
   assign m110_60 ={ {2{in110[5]}} , in110 , {2{1'b0}} };

   // m110_61 = W*in
   wire signed [9:0] m110_61;
   assign m110_61 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_62 = W*in
   wire signed [9:0] m110_62;
   assign m110_62 =10'b0;

   // m110_63 = W*in
   wire signed [9:0] m110_63;
   assign m110_63 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_64 = W*in
   wire signed [9:0] m110_64;
   assign m110_64 =10'b0;

   // m110_65 = W*in
   wire signed [9:0] m110_65;
   assign m110_65 =10'b0;

   // m110_66 = W*in
   wire signed [9:0] m110_66;
   assign m110_66 =10'b0;

   // m110_67 = W*in
   wire signed [9:0] m110_67;
   assign m110_67 =10'b0;

   // m110_68 = W*in
   wire signed [9:0] m110_68;
   assign m110_68 ={ {3{in110[5]}} , in110 , {1{1'b0}} };

   // m110_69 = W*in
   wire signed [9:0] m110_69;
   assign m110_69 =10'b0;

   // m110_70 = W*in
   wire signed [9:0] m110_70;
   assign m110_70 ={ {3{neg110[5]}} , neg110 , {1{1'b0}} };

   // m110_71 = W*in
   wire signed [9:0] m110_71;
   assign m110_71 =10'b0;

   // m110_72 = W*in
   wire signed [9:0] m110_72;
   assign m110_72 =10'b0;

   // m110_73 = W*in
   wire signed [9:0] m110_73;
   assign m110_73 =10'b0;

   // m110_74 = W*in
   wire signed [9:0] m110_74;
   assign m110_74 =10'b0;

   // m110_75 = W*in
   wire signed [9:0] m110_75;
   assign m110_75 =10'b0;

   // m110_76 = W*in
   wire signed [9:0] m110_76;
   assign m110_76 =10'b0;

   // m110_77 = W*in
   wire signed [9:0] m110_77;
   assign m110_77 =10'b0;

   // m110_78 = W*in
   wire signed [9:0] m110_78;
   assign m110_78 =10'b0;

   // m110_79 = W*in
   wire signed [9:0] m110_79;
   assign m110_79 =10'b0;

   // m110_80 = W*in
   wire signed [9:0] m110_80;
   assign m110_80 =10'b0;

   // m110_81 = W*in
   wire signed [9:0] m110_81;
   assign m110_81 =10'b0;

   // m111_1 = W*in
   wire signed [9:0] m111_1;
   assign m111_1 =10'b0;

   // m111_2 = W*in
   wire signed [9:0] m111_2;
   assign m111_2 =10'b0;

   // m111_3 = W*in
   wire signed [9:0] m111_3;
   assign m111_3 =10'b0;

   // m111_4 = W*in
   wire signed [9:0] m111_4;
   assign m111_4 =10'b0;

   // m111_5 = W*in
   wire signed [9:0] m111_5;
   assign m111_5 =10'b0;

   // m111_6 = W*in
   wire signed [9:0] m111_6;
   assign m111_6 =10'b0;

   // m111_7 = W*in
   wire signed [9:0] m111_7;
   assign m111_7 =10'b0;

   // m111_8 = W*in
   wire signed [9:0] m111_8;
   assign m111_8 =10'b0;

   // m111_9 = W*in
   wire signed [9:0] m111_9;
   assign m111_9 =10'b0;

   // m111_10 = W*in
   wire signed [9:0] m111_10;
   assign m111_10 =10'b0;

   // m111_11 = W*in
   wire signed [9:0] m111_11;
   assign m111_11 =10'b0;

   // m111_12 = W*in
   wire signed [9:0] m111_12;
   assign m111_12 =10'b0;

   // m111_13 = W*in
   wire signed [9:0] m111_13;
   assign m111_13 =10'b0;

   // m111_14 = W*in
   wire signed [9:0] m111_14;
   assign m111_14 =10'b0;

   // m111_15 = W*in
   wire signed [9:0] m111_15;
   assign m111_15 =10'b0;

   // m111_16 = W*in
   wire signed [9:0] m111_16;
   assign m111_16 =10'b0;

   // m111_17 = W*in
   wire signed [9:0] m111_17;
   assign m111_17 =10'b0;

   // m111_18 = W*in
   wire signed [9:0] m111_18;
   assign m111_18 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_19 = W*in
   wire signed [9:0] m111_19;
   assign m111_19 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_20 = W*in
   wire signed [9:0] m111_20;
   assign m111_20 =10'b0;

   // m111_21 = W*in
   wire signed [9:0] m111_21;
   assign m111_21 =10'b0;

   // m111_22 = W*in
   wire signed [9:0] m111_22;
   assign m111_22 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_23 = W*in
   wire signed [9:0] m111_23;
   assign m111_23 ={ {2{in111[5]}} , in111 , {2{1'b0}} };

   // m111_24 = W*in
   wire signed [9:0] m111_24;
   assign m111_24 =10'b0;

   // m111_25 = W*in
   wire signed [9:0] m111_25;
   assign m111_25 ={ {2{in111[5]}} , in111 , {2{1'b0}} };

   // m111_26 = W*in
   wire signed [9:0] m111_26;
   assign m111_26 =10'b0;

   // m111_27 = W*in
   wire signed [9:0] m111_27;
   assign m111_27 =10'b0;

   // m111_28 = W*in
   wire signed [9:0] m111_28;
   assign m111_28 =10'b0;

   // m111_29 = W*in
   wire signed [9:0] m111_29;
   assign m111_29 =10'b0;

   // m111_30 = W*in
   wire signed [9:0] m111_30;
   assign m111_30 ={ {3{in111[5]}} , in111 , {1{1'b0}} };

   // m111_31 = W*in
   wire signed [9:0] m111_31;
   assign m111_31 =10'b0;

   // m111_32 = W*in
   wire signed [9:0] m111_32;
   assign m111_32 =10'b0;

   // m111_33 = W*in
   wire signed [9:0] m111_33;
   assign m111_33 =10'b0;

   // m111_34 = W*in
   wire signed [9:0] m111_34;
   assign m111_34 =10'b0;

   // m111_35 = W*in
   wire signed [9:0] m111_35;
   assign m111_35 =10'b0;

   // m111_36 = W*in
   wire signed [9:0] m111_36;
   assign m111_36 ={ {3{in111[5]}} , in111 , {1{1'b0}} };

   // m111_37 = W*in
   wire signed [9:0] m111_37;
   assign m111_37 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_38 = W*in
   wire signed [9:0] m111_38;
   assign m111_38 =10'b0;

   // m111_39 = W*in
   wire signed [9:0] m111_39;
   assign m111_39 ={ {2{in111[5]}} , in111 , {2{1'b0}} };

   // m111_40 = W*in
   wire signed [9:0] m111_40;
   assign m111_40 =10'b0;

   // m111_41 = W*in
   wire signed [9:0] m111_41;
   assign m111_41 =10'b0;

   // m111_42 = W*in
   wire signed [9:0] m111_42;
   assign m111_42 =10'b0;

   // m111_43 = W*in
   wire signed [9:0] m111_43;
   assign m111_43 ={ {3{in111[5]}} , in111 , {1{1'b0}} };

   // m111_44 = W*in
   wire signed [9:0] m111_44;
   assign m111_44 =10'b0;

   // m111_45 = W*in
   wire signed [9:0] m111_45;
   assign m111_45 =10'b0;

   // m111_46 = W*in
   wire signed [9:0] m111_46;
   assign m111_46 =10'b0;

   // m111_47 = W*in
   wire signed [9:0] m111_47;
   assign m111_47 =10'b0;

   // m111_48 = W*in
   wire signed [9:0] m111_48;
   assign m111_48 =10'b0;

   // m111_49 = W*in
   wire signed [9:0] m111_49;
   assign m111_49 ={ {3{in111[5]}} , in111 , {1{1'b0}} };

   // m111_50 = W*in
   wire signed [9:0] m111_50;
   assign m111_50 ={ {3{in111[5]}} , in111 , {1{1'b0}} };

   // m111_51 = W*in
   wire signed [9:0] m111_51;
   assign m111_51 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_52 = W*in
   wire signed [9:0] m111_52;
   assign m111_52 =10'b0;

   // m111_53 = W*in
   wire signed [9:0] m111_53;
   assign m111_53 =10'b0;

   // m111_54 = W*in
   wire signed [9:0] m111_54;
   assign m111_54 =10'b0;

   // m111_55 = W*in
   wire signed [9:0] m111_55;
   assign m111_55 =10'b0;

   // m111_56 = W*in
   wire signed [9:0] m111_56;
   assign m111_56 =10'b0;

   // m111_57 = W*in
   wire signed [9:0] m111_57;
   assign m111_57 =10'b0;

   // m111_58 = W*in
   wire signed [9:0] m111_58;
   assign m111_58 =10'b0;

   // m111_59 = W*in
   wire signed [9:0] m111_59;
   assign m111_59 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_60 = W*in
   wire signed [9:0] m111_60;
   assign m111_60 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_61 = W*in
   wire signed [9:0] m111_61;
   assign m111_61 =10'b0;

   // m111_62 = W*in
   wire signed [9:0] m111_62;
   assign m111_62 ={ {3{in111[5]}} , in111 , {1{1'b0}} };

   // m111_63 = W*in
   wire signed [9:0] m111_63;
   assign m111_63 =10'b0;

   // m111_64 = W*in
   wire signed [9:0] m111_64;
   assign m111_64 =10'b0;

   // m111_65 = W*in
   wire signed [9:0] m111_65;
   assign m111_65 =10'b0;

   // m111_66 = W*in
   wire signed [9:0] m111_66;
   assign m111_66 =10'b0;

   // m111_67 = W*in
   wire signed [9:0] m111_67;
   assign m111_67 =10'b0;

   // m111_68 = W*in
   wire signed [9:0] m111_68;
   assign m111_68 =10'b0;

   // m111_69 = W*in
   wire signed [9:0] m111_69;
   assign m111_69 =10'b0;

   // m111_70 = W*in
   wire signed [9:0] m111_70;
   assign m111_70 ={ {3{neg111[5]}} , neg111 , {1{1'b0}} };

   // m111_71 = W*in
   wire signed [9:0] m111_71;
   assign m111_71 ={ {2{in111[5]}} , in111 , {2{1'b0}} };

   // m111_72 = W*in
   wire signed [9:0] m111_72;
   assign m111_72 =10'b0;

   // m111_73 = W*in
   wire signed [9:0] m111_73;
   assign m111_73 =10'b0;

   // m111_74 = W*in
   wire signed [9:0] m111_74;
   assign m111_74 =10'b0;

   // m111_75 = W*in
   wire signed [9:0] m111_75;
   assign m111_75 =10'b0;

   // m111_76 = W*in
   wire signed [9:0] m111_76;
   assign m111_76 =10'b0;

   // m111_77 = W*in
   wire signed [9:0] m111_77;
   assign m111_77 =10'b0;

   // m111_78 = W*in
   wire signed [9:0] m111_78;
   assign m111_78 =10'b0;

   // m111_79 = W*in
   wire signed [9:0] m111_79;
   assign m111_79 =10'b0;

   // m111_80 = W*in
   wire signed [9:0] m111_80;
   assign m111_80 =10'b0;

   // m111_81 = W*in
   wire signed [9:0] m111_81;
   assign m111_81 =10'b0;

   // m112_1 = W*in
   wire signed [9:0] m112_1;
   assign m112_1 =10'b0;

   // m112_2 = W*in
   wire signed [9:0] m112_2;
   assign m112_2 =10'b0;

   // m112_3 = W*in
   wire signed [9:0] m112_3;
   assign m112_3 =10'b0;

   // m112_4 = W*in
   wire signed [9:0] m112_4;
   assign m112_4 =10'b0;

   // m112_5 = W*in
   wire signed [9:0] m112_5;
   assign m112_5 =10'b0;

   // m112_6 = W*in
   wire signed [9:0] m112_6;
   assign m112_6 =10'b0;

   // m112_7 = W*in
   wire signed [9:0] m112_7;
   assign m112_7 =10'b0;

   // m112_8 = W*in
   wire signed [9:0] m112_8;
   assign m112_8 =10'b0;

   // m112_9 = W*in
   wire signed [9:0] m112_9;
   assign m112_9 =10'b0;

   // m112_10 = W*in
   wire signed [9:0] m112_10;
   assign m112_10 =10'b0;

   // m112_11 = W*in
   wire signed [9:0] m112_11;
   assign m112_11 ={ {2{in112[5]}} , in112 , {2{1'b0}} };

   // m112_12 = W*in
   wire signed [9:0] m112_12;
   assign m112_12 =10'b0;

   // m112_13 = W*in
   wire signed [9:0] m112_13;
   assign m112_13 =10'b0;

   // m112_14 = W*in
   wire signed [9:0] m112_14;
   assign m112_14 =10'b0;

   // m112_15 = W*in
   wire signed [9:0] m112_15;
   assign m112_15 =10'b0;

   // m112_16 = W*in
   wire signed [9:0] m112_16;
   assign m112_16 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_17 = W*in
   wire signed [9:0] m112_17;
   assign m112_17 =10'b0;

   // m112_18 = W*in
   wire signed [9:0] m112_18;
   assign m112_18 ={ {2{in112[5]}} , in112 , {2{1'b0}} };

   // m112_19 = W*in
   wire signed [9:0] m112_19;
   assign m112_19 ={ {2{in112[5]}} , in112 , {2{1'b0}} };

   // m112_20 = W*in
   wire signed [9:0] m112_20;
   assign m112_20 =10'b0;

   // m112_21 = W*in
   wire signed [9:0] m112_21;
   assign m112_21 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_22 = W*in
   wire signed [9:0] m112_22;
   assign m112_22 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_23 = W*in
   wire signed [9:0] m112_23;
   assign m112_23 ={ {3{neg112[5]}} , neg112 , {1{1'b0}} };

   // m112_24 = W*in
   wire signed [9:0] m112_24;
   assign m112_24 ={ {3{neg112[5]}} , neg112 , {1{1'b0}} };

   // m112_25 = W*in
   wire signed [9:0] m112_25;
   assign m112_25 =10'b0;

   // m112_26 = W*in
   wire signed [9:0] m112_26;
   assign m112_26 =10'b0;

   // m112_27 = W*in
   wire signed [9:0] m112_27;
   assign m112_27 =10'b0;

   // m112_28 = W*in
   wire signed [9:0] m112_28;
   assign m112_28 ={ {3{neg112[5]}} , neg112 , {1{1'b0}} };

   // m112_29 = W*in
   wire signed [9:0] m112_29;
   assign m112_29 =10'b0;

   // m112_30 = W*in
   wire signed [9:0] m112_30;
   assign m112_30 =10'b0;

   // m112_31 = W*in
   wire signed [9:0] m112_31;
   assign m112_31 =10'b0;

   // m112_32 = W*in
   wire signed [9:0] m112_32;
   assign m112_32 =10'b0;

   // m112_33 = W*in
   wire signed [9:0] m112_33;
   assign m112_33 =10'b0;

   // m112_34 = W*in
   wire signed [9:0] m112_34;
   assign m112_34 =10'b0;

   // m112_35 = W*in
   wire signed [9:0] m112_35;
   assign m112_35 =10'b0;

   // m112_36 = W*in
   wire signed [9:0] m112_36;
   assign m112_36 =10'b0;

   // m112_37 = W*in
   wire signed [9:0] m112_37;
   assign m112_37 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_38 = W*in
   wire signed [9:0] m112_38;
   assign m112_38 =10'b0;

   // m112_39 = W*in
   wire signed [9:0] m112_39;
   assign m112_39 ={ {3{neg112[5]}} , neg112 , {1{1'b0}} };

   // m112_40 = W*in
   wire signed [9:0] m112_40;
   assign m112_40 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_41 = W*in
   wire signed [9:0] m112_41;
   assign m112_41 ={ {2{in112[5]}} , in112 , {2{1'b0}} };

   // m112_42 = W*in
   wire signed [9:0] m112_42;
   assign m112_42 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_43 = W*in
   wire signed [9:0] m112_43;
   assign m112_43 =10'b0;

   // m112_44 = W*in
   wire signed [9:0] m112_44;
   assign m112_44 =10'b0;

   // m112_45 = W*in
   wire signed [9:0] m112_45;
   assign m112_45 ={ {3{neg112[5]}} , neg112 , {1{1'b0}} };

   // m112_46 = W*in
   wire signed [9:0] m112_46;
   assign m112_46 =10'b0;

   // m112_47 = W*in
   wire signed [9:0] m112_47;
   assign m112_47 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_48 = W*in
   wire signed [9:0] m112_48;
   assign m112_48 =10'b0;

   // m112_49 = W*in
   wire signed [9:0] m112_49;
   assign m112_49 =10'b0;

   // m112_50 = W*in
   wire signed [9:0] m112_50;
   assign m112_50 =10'b0;

   // m112_51 = W*in
   wire signed [9:0] m112_51;
   assign m112_51 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_52 = W*in
   wire signed [9:0] m112_52;
   assign m112_52 =10'b0;

   // m112_53 = W*in
   wire signed [9:0] m112_53;
   assign m112_53 =10'b0;

   // m112_54 = W*in
   wire signed [9:0] m112_54;
   assign m112_54 =10'b0;

   // m112_55 = W*in
   wire signed [9:0] m112_55;
   assign m112_55 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_56 = W*in
   wire signed [9:0] m112_56;
   assign m112_56 =10'b0;

   // m112_57 = W*in
   wire signed [9:0] m112_57;
   assign m112_57 =10'b0;

   // m112_58 = W*in
   wire signed [9:0] m112_58;
   assign m112_58 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_59 = W*in
   wire signed [9:0] m112_59;
   assign m112_59 =10'b0;

   // m112_60 = W*in
   wire signed [9:0] m112_60;
   assign m112_60 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_61 = W*in
   wire signed [9:0] m112_61;
   assign m112_61 =10'b0;

   // m112_62 = W*in
   wire signed [9:0] m112_62;
   assign m112_62 ={ {3{in112[5]}} , in112 , {1{1'b0}} };

   // m112_63 = W*in
   wire signed [9:0] m112_63;
   assign m112_63 =10'b0;

   // m112_64 = W*in
   wire signed [9:0] m112_64;
   assign m112_64 =10'b0;

   // m112_65 = W*in
   wire signed [9:0] m112_65;
   assign m112_65 =10'b0;

   // m112_66 = W*in
   wire signed [9:0] m112_66;
   assign m112_66 =10'b0;

   // m112_67 = W*in
   wire signed [9:0] m112_67;
   assign m112_67 =10'b0;

   // m112_68 = W*in
   wire signed [9:0] m112_68;
   assign m112_68 ={ {3{neg112[5]}} , neg112 , {1{1'b0}} };

   // m112_69 = W*in
   wire signed [9:0] m112_69;
   assign m112_69 =10'b0;

   // m112_70 = W*in
   wire signed [9:0] m112_70;
   assign m112_70 =10'b0;

   // m112_71 = W*in
   wire signed [9:0] m112_71;
   assign m112_71 =10'b0;

   // m112_72 = W*in
   wire signed [9:0] m112_72;
   assign m112_72 =10'b0;

   // m112_73 = W*in
   wire signed [9:0] m112_73;
   assign m112_73 =10'b0;

   // m112_74 = W*in
   wire signed [9:0] m112_74;
   assign m112_74 =10'b0;

   // m112_75 = W*in
   wire signed [9:0] m112_75;
   assign m112_75 =10'b0;

   // m112_76 = W*in
   wire signed [9:0] m112_76;
   assign m112_76 =10'b0;

   // m112_77 = W*in
   wire signed [9:0] m112_77;
   assign m112_77 =10'b0;

   // m112_78 = W*in
   wire signed [9:0] m112_78;
   assign m112_78 =10'b0;

   // m112_79 = W*in
   wire signed [9:0] m112_79;
   assign m112_79 =10'b0;

   // m112_80 = W*in
   wire signed [9:0] m112_80;
   assign m112_80 =10'b0;

   // m112_81 = W*in
   wire signed [9:0] m112_81;
   assign m112_81 =10'b0;

   // m113_1 = W*in
   wire signed [9:0] m113_1;
   assign m113_1 =10'b0;

   // m113_2 = W*in
   wire signed [9:0] m113_2;
   assign m113_2 =10'b0;

   // m113_3 = W*in
   wire signed [9:0] m113_3;
   assign m113_3 =10'b0;

   // m113_4 = W*in
   wire signed [9:0] m113_4;
   assign m113_4 =10'b0;

   // m113_5 = W*in
   wire signed [9:0] m113_5;
   assign m113_5 =10'b0;

   // m113_6 = W*in
   wire signed [9:0] m113_6;
   assign m113_6 =10'b0;

   // m113_7 = W*in
   wire signed [9:0] m113_7;
   assign m113_7 =10'b0;

   // m113_8 = W*in
   wire signed [9:0] m113_8;
   assign m113_8 =10'b0;

   // m113_9 = W*in
   wire signed [9:0] m113_9;
   assign m113_9 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_10 = W*in
   wire signed [9:0] m113_10;
   assign m113_10 =10'b0;

   // m113_11 = W*in
   wire signed [9:0] m113_11;
   assign m113_11 =10'b0;

   // m113_12 = W*in
   wire signed [9:0] m113_12;
   assign m113_12 =10'b0;

   // m113_13 = W*in
   wire signed [9:0] m113_13;
   assign m113_13 =10'b0;

   // m113_14 = W*in
   wire signed [9:0] m113_14;
   assign m113_14 =10'b0;

   // m113_15 = W*in
   wire signed [9:0] m113_15;
   assign m113_15 =10'b0;

   // m113_16 = W*in
   wire signed [9:0] m113_16;
   assign m113_16 =10'b0;

   // m113_17 = W*in
   wire signed [9:0] m113_17;
   assign m113_17 ={ {2{in113[5]}} , in113 , {2{1'b0}} };

   // m113_18 = W*in
   wire signed [9:0] m113_18;
   assign m113_18 =10'b0;

   // m113_19 = W*in
   wire signed [9:0] m113_19;
   assign m113_19 =10'b0;

   // m113_20 = W*in
   wire signed [9:0] m113_20;
   assign m113_20 =10'b0;

   // m113_21 = W*in
   wire signed [9:0] m113_21;
   assign m113_21 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_22 = W*in
   wire signed [9:0] m113_22;
   assign m113_22 =10'b0;

   // m113_23 = W*in
   wire signed [9:0] m113_23;
   assign m113_23 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_24 = W*in
   wire signed [9:0] m113_24;
   assign m113_24 =10'b0;

   // m113_25 = W*in
   wire signed [9:0] m113_25;
   assign m113_25 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_26 = W*in
   wire signed [9:0] m113_26;
   assign m113_26 =10'b0;

   // m113_27 = W*in
   wire signed [9:0] m113_27;
   assign m113_27 =10'b0;

   // m113_28 = W*in
   wire signed [9:0] m113_28;
   assign m113_28 =10'b0;

   // m113_29 = W*in
   wire signed [9:0] m113_29;
   assign m113_29 =10'b0;

   // m113_30 = W*in
   wire signed [9:0] m113_30;
   assign m113_30 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_31 = W*in
   wire signed [9:0] m113_31;
   assign m113_31 ={ {3{neg113[5]}} , neg113 , {1{1'b0}} };

   // m113_32 = W*in
   wire signed [9:0] m113_32;
   assign m113_32 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_33 = W*in
   wire signed [9:0] m113_33;
   assign m113_33 =10'b0;

   // m113_34 = W*in
   wire signed [9:0] m113_34;
   assign m113_34 =10'b0;

   // m113_35 = W*in
   wire signed [9:0] m113_35;
   assign m113_35 =10'b0;

   // m113_36 = W*in
   wire signed [9:0] m113_36;
   assign m113_36 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_37 = W*in
   wire signed [9:0] m113_37;
   assign m113_37 ={ {2{neg113[5]}} , neg113 , {2{1'b0}} };

   // m113_38 = W*in
   wire signed [9:0] m113_38;
   assign m113_38 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_39 = W*in
   wire signed [9:0] m113_39;
   assign m113_39 =10'b0;

   // m113_40 = W*in
   wire signed [9:0] m113_40;
   assign m113_40 =10'b0;

   // m113_41 = W*in
   wire signed [9:0] m113_41;
   assign m113_41 =10'b0;

   // m113_42 = W*in
   wire signed [9:0] m113_42;
   assign m113_42 ={ {2{in113[5]}} , in113 , {2{1'b0}} };

   // m113_43 = W*in
   wire signed [9:0] m113_43;
   assign m113_43 =10'b0;

   // m113_44 = W*in
   wire signed [9:0] m113_44;
   assign m113_44 =10'b0;

   // m113_45 = W*in
   wire signed [9:0] m113_45;
   assign m113_45 =10'b0;

   // m113_46 = W*in
   wire signed [9:0] m113_46;
   assign m113_46 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_47 = W*in
   wire signed [9:0] m113_47;
   assign m113_47 =10'b0;

   // m113_48 = W*in
   wire signed [9:0] m113_48;
   assign m113_48 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_49 = W*in
   wire signed [9:0] m113_49;
   assign m113_49 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_50 = W*in
   wire signed [9:0] m113_50;
   assign m113_50 =10'b0;

   // m113_51 = W*in
   wire signed [9:0] m113_51;
   assign m113_51 ={ {3{neg113[5]}} , neg113 , {1{1'b0}} };

   // m113_52 = W*in
   wire signed [9:0] m113_52;
   assign m113_52 =10'b0;

   // m113_53 = W*in
   wire signed [9:0] m113_53;
   assign m113_53 =10'b0;

   // m113_54 = W*in
   wire signed [9:0] m113_54;
   assign m113_54 =10'b0;

   // m113_55 = W*in
   wire signed [9:0] m113_55;
   assign m113_55 =10'b0;

   // m113_56 = W*in
   wire signed [9:0] m113_56;
   assign m113_56 =10'b0;

   // m113_57 = W*in
   wire signed [9:0] m113_57;
   assign m113_57 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_58 = W*in
   wire signed [9:0] m113_58;
   assign m113_58 ={ {3{neg113[5]}} , neg113 , {1{1'b0}} };

   // m113_59 = W*in
   wire signed [9:0] m113_59;
   assign m113_59 ={ {3{neg113[5]}} , neg113 , {1{1'b0}} };

   // m113_60 = W*in
   wire signed [9:0] m113_60;
   assign m113_60 ={ {3{neg113[5]}} , neg113 , {1{1'b0}} };

   // m113_61 = W*in
   wire signed [9:0] m113_61;
   assign m113_61 =10'b0;

   // m113_62 = W*in
   wire signed [9:0] m113_62;
   assign m113_62 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_63 = W*in
   wire signed [9:0] m113_63;
   assign m113_63 =10'b0;

   // m113_64 = W*in
   wire signed [9:0] m113_64;
   assign m113_64 =10'b0;

   // m113_65 = W*in
   wire signed [9:0] m113_65;
   assign m113_65 =10'b0;

   // m113_66 = W*in
   wire signed [9:0] m113_66;
   assign m113_66 ={ {2{in113[5]}} , in113 , {2{1'b0}} };

   // m113_67 = W*in
   wire signed [9:0] m113_67;
   assign m113_67 =10'b0;

   // m113_68 = W*in
   wire signed [9:0] m113_68;
   assign m113_68 ={ {3{in113[5]}} , in113 , {1{1'b0}} };

   // m113_69 = W*in
   wire signed [9:0] m113_69;
   assign m113_69 ={ {3{neg113[5]}} , neg113 , {1{1'b0}} };

   // m113_70 = W*in
   wire signed [9:0] m113_70;
   assign m113_70 =10'b0;

   // m113_71 = W*in
   wire signed [9:0] m113_71;
   assign m113_71 ={ {2{in113[5]}} , in113 , {2{1'b0}} };

   // m113_72 = W*in
   wire signed [9:0] m113_72;
   assign m113_72 =10'b0;

   // m113_73 = W*in
   wire signed [9:0] m113_73;
   assign m113_73 =10'b0;

   // m113_74 = W*in
   wire signed [9:0] m113_74;
   assign m113_74 =10'b0;

   // m113_75 = W*in
   wire signed [9:0] m113_75;
   assign m113_75 =10'b0;

   // m113_76 = W*in
   wire signed [9:0] m113_76;
   assign m113_76 =10'b0;

   // m113_77 = W*in
   wire signed [9:0] m113_77;
   assign m113_77 =10'b0;

   // m113_78 = W*in
   wire signed [9:0] m113_78;
   assign m113_78 =10'b0;

   // m113_79 = W*in
   wire signed [9:0] m113_79;
   assign m113_79 =10'b0;

   // m113_80 = W*in
   wire signed [9:0] m113_80;
   assign m113_80 =10'b0;

   // m113_81 = W*in
   wire signed [9:0] m113_81;
   assign m113_81 =10'b0;

   // m114_1 = W*in
   wire signed [9:0] m114_1;
   assign m114_1 =10'b0;

   // m114_2 = W*in
   wire signed [9:0] m114_2;
   assign m114_2 =10'b0;

   // m114_3 = W*in
   wire signed [9:0] m114_3;
   assign m114_3 =10'b0;

   // m114_4 = W*in
   wire signed [9:0] m114_4;
   assign m114_4 =10'b0;

   // m114_5 = W*in
   wire signed [9:0] m114_5;
   assign m114_5 =10'b0;

   // m114_6 = W*in
   wire signed [9:0] m114_6;
   assign m114_6 =10'b0;

   // m114_7 = W*in
   wire signed [9:0] m114_7;
   assign m114_7 =10'b0;

   // m114_8 = W*in
   wire signed [9:0] m114_8;
   assign m114_8 =10'b0;

   // m114_9 = W*in
   wire signed [9:0] m114_9;
   assign m114_9 =10'b0;

   // m114_10 = W*in
   wire signed [9:0] m114_10;
   assign m114_10 =10'b0;

   // m114_11 = W*in
   wire signed [9:0] m114_11;
   assign m114_11 =10'b0;

   // m114_12 = W*in
   wire signed [9:0] m114_12;
   assign m114_12 =10'b0;

   // m114_13 = W*in
   wire signed [9:0] m114_13;
   assign m114_13 =10'b0;

   // m114_14 = W*in
   wire signed [9:0] m114_14;
   assign m114_14 ={ {2{in114[5]}} , in114 , {2{1'b0}} };

   // m114_15 = W*in
   wire signed [9:0] m114_15;
   assign m114_15 ={ {3{neg114[5]}} , neg114 , {1{1'b0}} };

   // m114_16 = W*in
   wire signed [9:0] m114_16;
   assign m114_16 =10'b0;

   // m114_17 = W*in
   wire signed [9:0] m114_17;
   assign m114_17 =10'b0;

   // m114_18 = W*in
   wire signed [9:0] m114_18;
   assign m114_18 =10'b0;

   // m114_19 = W*in
   wire signed [9:0] m114_19;
   assign m114_19 =10'b0;

   // m114_20 = W*in
   wire signed [9:0] m114_20;
   assign m114_20 =10'b0;

   // m114_21 = W*in
   wire signed [9:0] m114_21;
   assign m114_21 =10'b0;

   // m114_22 = W*in
   wire signed [9:0] m114_22;
   assign m114_22 =10'b0;

   // m114_23 = W*in
   wire signed [9:0] m114_23;
   assign m114_23 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_24 = W*in
   wire signed [9:0] m114_24;
   assign m114_24 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_25 = W*in
   wire signed [9:0] m114_25;
   assign m114_25 =10'b0;

   // m114_26 = W*in
   wire signed [9:0] m114_26;
   assign m114_26 =10'b0;

   // m114_27 = W*in
   wire signed [9:0] m114_27;
   assign m114_27 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_28 = W*in
   wire signed [9:0] m114_28;
   assign m114_28 ={ {2{in114[5]}} , in114 , {2{1'b0}} };

   // m114_29 = W*in
   wire signed [9:0] m114_29;
   assign m114_29 =10'b0;

   // m114_30 = W*in
   wire signed [9:0] m114_30;
   assign m114_30 =10'b0;

   // m114_31 = W*in
   wire signed [9:0] m114_31;
   assign m114_31 =10'b0;

   // m114_32 = W*in
   wire signed [9:0] m114_32;
   assign m114_32 =10'b0;

   // m114_33 = W*in
   wire signed [9:0] m114_33;
   assign m114_33 ={ {3{neg114[5]}} , neg114 , {1{1'b0}} };

   // m114_34 = W*in
   wire signed [9:0] m114_34;
   assign m114_34 =10'b0;

   // m114_35 = W*in
   wire signed [9:0] m114_35;
   assign m114_35 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_36 = W*in
   wire signed [9:0] m114_36;
   assign m114_36 =10'b0;

   // m114_37 = W*in
   wire signed [9:0] m114_37;
   assign m114_37 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_38 = W*in
   wire signed [9:0] m114_38;
   assign m114_38 =10'b0;

   // m114_39 = W*in
   wire signed [9:0] m114_39;
   assign m114_39 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_40 = W*in
   wire signed [9:0] m114_40;
   assign m114_40 =10'b0;

   // m114_41 = W*in
   wire signed [9:0] m114_41;
   assign m114_41 ={ {3{neg114[5]}} , neg114 , {1{1'b0}} };

   // m114_42 = W*in
   wire signed [9:0] m114_42;
   assign m114_42 =10'b0;

   // m114_43 = W*in
   wire signed [9:0] m114_43;
   assign m114_43 =10'b0;

   // m114_44 = W*in
   wire signed [9:0] m114_44;
   assign m114_44 =10'b0;

   // m114_45 = W*in
   wire signed [9:0] m114_45;
   assign m114_45 =10'b0;

   // m114_46 = W*in
   wire signed [9:0] m114_46;
   assign m114_46 ={ {3{in114[5]}} , in114 , {1{1'b0}} };

   // m114_47 = W*in
   wire signed [9:0] m114_47;
   assign m114_47 =10'b0;

   // m114_48 = W*in
   wire signed [9:0] m114_48;
   assign m114_48 =10'b0;

   // m114_49 = W*in
   wire signed [9:0] m114_49;
   assign m114_49 =10'b0;

   // m114_50 = W*in
   wire signed [9:0] m114_50;
   assign m114_50 =10'b0;

   // m114_51 = W*in
   wire signed [9:0] m114_51;
   assign m114_51 =10'b0;

   // m114_52 = W*in
   wire signed [9:0] m114_52;
   assign m114_52 =10'b0;

   // m114_53 = W*in
   wire signed [9:0] m114_53;
   assign m114_53 =10'b0;

   // m114_54 = W*in
   wire signed [9:0] m114_54;
   assign m114_54 =10'b0;

   // m114_55 = W*in
   wire signed [9:0] m114_55;
   assign m114_55 =10'b0;

   // m114_56 = W*in
   wire signed [9:0] m114_56;
   assign m114_56 =10'b0;

   // m114_57 = W*in
   wire signed [9:0] m114_57;
   assign m114_57 =10'b0;

   // m114_58 = W*in
   wire signed [9:0] m114_58;
   assign m114_58 =10'b0;

   // m114_59 = W*in
   wire signed [9:0] m114_59;
   assign m114_59 =10'b0;

   // m114_60 = W*in
   wire signed [9:0] m114_60;
   assign m114_60 =10'b0;

   // m114_61 = W*in
   wire signed [9:0] m114_61;
   assign m114_61 =10'b0;

   // m114_62 = W*in
   wire signed [9:0] m114_62;
   assign m114_62 =10'b0;

   // m114_63 = W*in
   wire signed [9:0] m114_63;
   assign m114_63 =10'b0;

   // m114_64 = W*in
   wire signed [9:0] m114_64;
   assign m114_64 =10'b0;

   // m114_65 = W*in
   wire signed [9:0] m114_65;
   assign m114_65 =10'b0;

   // m114_66 = W*in
   wire signed [9:0] m114_66;
   assign m114_66 =10'b0;

   // m114_67 = W*in
   wire signed [9:0] m114_67;
   assign m114_67 =10'b0;

   // m114_68 = W*in
   wire signed [9:0] m114_68;
   assign m114_68 =10'b0;

   // m114_69 = W*in
   wire signed [9:0] m114_69;
   assign m114_69 =10'b0;

   // m114_70 = W*in
   wire signed [9:0] m114_70;
   assign m114_70 =10'b0;

   // m114_71 = W*in
   wire signed [9:0] m114_71;
   assign m114_71 =10'b0;

   // m114_72 = W*in
   wire signed [9:0] m114_72;
   assign m114_72 =10'b0;

   // m114_73 = W*in
   wire signed [9:0] m114_73;
   assign m114_73 =10'b0;

   // m114_74 = W*in
   wire signed [9:0] m114_74;
   assign m114_74 =10'b0;

   // m114_75 = W*in
   wire signed [9:0] m114_75;
   assign m114_75 =10'b0;

   // m114_76 = W*in
   wire signed [9:0] m114_76;
   assign m114_76 =10'b0;

   // m114_77 = W*in
   wire signed [9:0] m114_77;
   assign m114_77 =10'b0;

   // m114_78 = W*in
   wire signed [9:0] m114_78;
   assign m114_78 =10'b0;

   // m114_79 = W*in
   wire signed [9:0] m114_79;
   assign m114_79 =10'b0;

   // m114_80 = W*in
   wire signed [9:0] m114_80;
   assign m114_80 =10'b0;

   // m114_81 = W*in
   wire signed [9:0] m114_81;
   assign m114_81 =10'b0;

   // m115_1 = W*in
   wire signed [9:0] m115_1;
   assign m115_1 =10'b0;

   // m115_2 = W*in
   wire signed [9:0] m115_2;
   assign m115_2 =10'b0;

   // m115_3 = W*in
   wire signed [9:0] m115_3;
   assign m115_3 =10'b0;

   // m115_4 = W*in
   wire signed [9:0] m115_4;
   assign m115_4 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_5 = W*in
   wire signed [9:0] m115_5;
   assign m115_5 =10'b0;

   // m115_6 = W*in
   wire signed [9:0] m115_6;
   assign m115_6 =10'b0;

   // m115_7 = W*in
   wire signed [9:0] m115_7;
   assign m115_7 =10'b0;

   // m115_8 = W*in
   wire signed [9:0] m115_8;
   assign m115_8 =10'b0;

   // m115_9 = W*in
   wire signed [9:0] m115_9;
   assign m115_9 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_10 = W*in
   wire signed [9:0] m115_10;
   assign m115_10 =10'b0;

   // m115_11 = W*in
   wire signed [9:0] m115_11;
   assign m115_11 =10'b0;

   // m115_12 = W*in
   wire signed [9:0] m115_12;
   assign m115_12 =10'b0;

   // m115_13 = W*in
   wire signed [9:0] m115_13;
   assign m115_13 =10'b0;

   // m115_14 = W*in
   wire signed [9:0] m115_14;
   assign m115_14 =10'b0;

   // m115_15 = W*in
   wire signed [9:0] m115_15;
   assign m115_15 =10'b0;

   // m115_16 = W*in
   wire signed [9:0] m115_16;
   assign m115_16 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_17 = W*in
   wire signed [9:0] m115_17;
   assign m115_17 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_18 = W*in
   wire signed [9:0] m115_18;
   assign m115_18 =10'b0;

   // m115_19 = W*in
   wire signed [9:0] m115_19;
   assign m115_19 =10'b0;

   // m115_20 = W*in
   wire signed [9:0] m115_20;
   assign m115_20 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_21 = W*in
   wire signed [9:0] m115_21;
   assign m115_21 =10'b0;

   // m115_22 = W*in
   wire signed [9:0] m115_22;
   assign m115_22 =10'b0;

   // m115_23 = W*in
   wire signed [9:0] m115_23;
   assign m115_23 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_24 = W*in
   wire signed [9:0] m115_24;
   assign m115_24 =10'b0;

   // m115_25 = W*in
   wire signed [9:0] m115_25;
   assign m115_25 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_26 = W*in
   wire signed [9:0] m115_26;
   assign m115_26 =10'b0;

   // m115_27 = W*in
   wire signed [9:0] m115_27;
   assign m115_27 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_28 = W*in
   wire signed [9:0] m115_28;
   assign m115_28 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_29 = W*in
   wire signed [9:0] m115_29;
   assign m115_29 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_30 = W*in
   wire signed [9:0] m115_30;
   assign m115_30 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_31 = W*in
   wire signed [9:0] m115_31;
   assign m115_31 =10'b0;

   // m115_32 = W*in
   wire signed [9:0] m115_32;
   assign m115_32 ={ {2{in115[5]}} , in115 , {2{1'b0}} };

   // m115_33 = W*in
   wire signed [9:0] m115_33;
   assign m115_33 =10'b0;

   // m115_34 = W*in
   wire signed [9:0] m115_34;
   assign m115_34 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_35 = W*in
   wire signed [9:0] m115_35;
   assign m115_35 ={ {2{in115[5]}} , in115 , {2{1'b0}} };

   // m115_36 = W*in
   wire signed [9:0] m115_36;
   assign m115_36 =10'b0;

   // m115_37 = W*in
   wire signed [9:0] m115_37;
   assign m115_37 =10'b0;

   // m115_38 = W*in
   wire signed [9:0] m115_38;
   assign m115_38 =10'b0;

   // m115_39 = W*in
   wire signed [9:0] m115_39;
   assign m115_39 =10'b0;

   // m115_40 = W*in
   wire signed [9:0] m115_40;
   assign m115_40 =10'b0;

   // m115_41 = W*in
   wire signed [9:0] m115_41;
   assign m115_41 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_42 = W*in
   wire signed [9:0] m115_42;
   assign m115_42 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_43 = W*in
   wire signed [9:0] m115_43;
   assign m115_43 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_44 = W*in
   wire signed [9:0] m115_44;
   assign m115_44 =10'b0;

   // m115_45 = W*in
   wire signed [9:0] m115_45;
   assign m115_45 =10'b0;

   // m115_46 = W*in
   wire signed [9:0] m115_46;
   assign m115_46 ={ {2{in115[5]}} , in115 , {2{1'b0}} };

   // m115_47 = W*in
   wire signed [9:0] m115_47;
   assign m115_47 =10'b0;

   // m115_48 = W*in
   wire signed [9:0] m115_48;
   assign m115_48 =10'b0;

   // m115_49 = W*in
   wire signed [9:0] m115_49;
   assign m115_49 =10'b0;

   // m115_50 = W*in
   wire signed [9:0] m115_50;
   assign m115_50 =10'b0;

   // m115_51 = W*in
   wire signed [9:0] m115_51;
   assign m115_51 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_52 = W*in
   wire signed [9:0] m115_52;
   assign m115_52 =10'b0;

   // m115_53 = W*in
   wire signed [9:0] m115_53;
   assign m115_53 =10'b0;

   // m115_54 = W*in
   wire signed [9:0] m115_54;
   assign m115_54 =10'b0;

   // m115_55 = W*in
   wire signed [9:0] m115_55;
   assign m115_55 =10'b0;

   // m115_56 = W*in
   wire signed [9:0] m115_56;
   assign m115_56 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_57 = W*in
   wire signed [9:0] m115_57;
   assign m115_57 =10'b0;

   // m115_58 = W*in
   wire signed [9:0] m115_58;
   assign m115_58 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_59 = W*in
   wire signed [9:0] m115_59;
   assign m115_59 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_60 = W*in
   wire signed [9:0] m115_60;
   assign m115_60 =10'b0;

   // m115_61 = W*in
   wire signed [9:0] m115_61;
   assign m115_61 =10'b0;

   // m115_62 = W*in
   wire signed [9:0] m115_62;
   assign m115_62 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_63 = W*in
   wire signed [9:0] m115_63;
   assign m115_63 ={ {3{in115[5]}} , in115 , {1{1'b0}} };

   // m115_64 = W*in
   wire signed [9:0] m115_64;
   assign m115_64 =10'b0;

   // m115_65 = W*in
   wire signed [9:0] m115_65;
   assign m115_65 =10'b0;

   // m115_66 = W*in
   wire signed [9:0] m115_66;
   assign m115_66 =10'b0;

   // m115_67 = W*in
   wire signed [9:0] m115_67;
   assign m115_67 =10'b0;

   // m115_68 = W*in
   wire signed [9:0] m115_68;
   assign m115_68 =10'b0;

   // m115_69 = W*in
   wire signed [9:0] m115_69;
   assign m115_69 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_70 = W*in
   wire signed [9:0] m115_70;
   assign m115_70 =10'b0;

   // m115_71 = W*in
   wire signed [9:0] m115_71;
   assign m115_71 =10'b0;

   // m115_72 = W*in
   wire signed [9:0] m115_72;
   assign m115_72 =10'b0;

   // m115_73 = W*in
   wire signed [9:0] m115_73;
   assign m115_73 =10'b0;

   // m115_74 = W*in
   wire signed [9:0] m115_74;
   assign m115_74 =10'b0;

   // m115_75 = W*in
   wire signed [9:0] m115_75;
   assign m115_75 =10'b0;

   // m115_76 = W*in
   wire signed [9:0] m115_76;
   assign m115_76 =10'b0;

   // m115_77 = W*in
   wire signed [9:0] m115_77;
   assign m115_77 ={ {3{neg115[5]}} , neg115 , {1{1'b0}} };

   // m115_78 = W*in
   wire signed [9:0] m115_78;
   assign m115_78 =10'b0;

   // m115_79 = W*in
   wire signed [9:0] m115_79;
   assign m115_79 =10'b0;

   // m115_80 = W*in
   wire signed [9:0] m115_80;
   assign m115_80 =10'b0;

   // m115_81 = W*in
   wire signed [9:0] m115_81;
   assign m115_81 =10'b0;

   // m116_1 = W*in
   wire signed [9:0] m116_1;
   assign m116_1 =10'b0;

   // m116_2 = W*in
   wire signed [9:0] m116_2;
   assign m116_2 =10'b0;

   // m116_3 = W*in
   wire signed [9:0] m116_3;
   assign m116_3 ={ {2{in116[5]}} , in116 , {2{1'b0}} };

   // m116_4 = W*in
   wire signed [9:0] m116_4;
   assign m116_4 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_5 = W*in
   wire signed [9:0] m116_5;
   assign m116_5 =10'b0;

   // m116_6 = W*in
   wire signed [9:0] m116_6;
   assign m116_6 =10'b0;

   // m116_7 = W*in
   wire signed [9:0] m116_7;
   assign m116_7 =10'b0;

   // m116_8 = W*in
   wire signed [9:0] m116_8;
   assign m116_8 =10'b0;

   // m116_9 = W*in
   wire signed [9:0] m116_9;
   assign m116_9 ={ {2{in116[5]}} , in116 , {2{1'b0}} };

   // m116_10 = W*in
   wire signed [9:0] m116_10;
   assign m116_10 =10'b0;

   // m116_11 = W*in
   wire signed [9:0] m116_11;
   assign m116_11 =10'b0;

   // m116_12 = W*in
   wire signed [9:0] m116_12;
   assign m116_12 =10'b0;

   // m116_13 = W*in
   wire signed [9:0] m116_13;
   assign m116_13 =10'b0;

   // m116_14 = W*in
   wire signed [9:0] m116_14;
   assign m116_14 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_15 = W*in
   wire signed [9:0] m116_15;
   assign m116_15 =10'b0;

   // m116_16 = W*in
   wire signed [9:0] m116_16;
   assign m116_16 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_17 = W*in
   wire signed [9:0] m116_17;
   assign m116_17 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_18 = W*in
   wire signed [9:0] m116_18;
   assign m116_18 ={ {2{in116[5]}} , in116 , {2{1'b0}} };

   // m116_19 = W*in
   wire signed [9:0] m116_19;
   assign m116_19 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_20 = W*in
   wire signed [9:0] m116_20;
   assign m116_20 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_21 = W*in
   wire signed [9:0] m116_21;
   assign m116_21 =10'b0;

   // m116_22 = W*in
   wire signed [9:0] m116_22;
   assign m116_22 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_23 = W*in
   wire signed [9:0] m116_23;
   assign m116_23 =10'b0;

   // m116_24 = W*in
   wire signed [9:0] m116_24;
   assign m116_24 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_25 = W*in
   wire signed [9:0] m116_25;
   assign m116_25 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_26 = W*in
   wire signed [9:0] m116_26;
   assign m116_26 =10'b0;

   // m116_27 = W*in
   wire signed [9:0] m116_27;
   assign m116_27 =10'b0;

   // m116_28 = W*in
   wire signed [9:0] m116_28;
   assign m116_28 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_29 = W*in
   wire signed [9:0] m116_29;
   assign m116_29 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_30 = W*in
   wire signed [9:0] m116_30;
   assign m116_30 =10'b0;

   // m116_31 = W*in
   wire signed [9:0] m116_31;
   assign m116_31 =10'b0;

   // m116_32 = W*in
   wire signed [9:0] m116_32;
   assign m116_32 =10'b0;

   // m116_33 = W*in
   wire signed [9:0] m116_33;
   assign m116_33 =10'b0;

   // m116_34 = W*in
   wire signed [9:0] m116_34;
   assign m116_34 =10'b0;

   // m116_35 = W*in
   wire signed [9:0] m116_35;
   assign m116_35 =10'b0;

   // m116_36 = W*in
   wire signed [9:0] m116_36;
   assign m116_36 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_37 = W*in
   wire signed [9:0] m116_37;
   assign m116_37 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_38 = W*in
   wire signed [9:0] m116_38;
   assign m116_38 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_39 = W*in
   wire signed [9:0] m116_39;
   assign m116_39 =10'b0;

   // m116_40 = W*in
   wire signed [9:0] m116_40;
   assign m116_40 =10'b0;

   // m116_41 = W*in
   wire signed [9:0] m116_41;
   assign m116_41 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_42 = W*in
   wire signed [9:0] m116_42;
   assign m116_42 ={ {2{in116[5]}} , in116 , {2{1'b0}} };

   // m116_43 = W*in
   wire signed [9:0] m116_43;
   assign m116_43 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_44 = W*in
   wire signed [9:0] m116_44;
   assign m116_44 =10'b0;

   // m116_45 = W*in
   wire signed [9:0] m116_45;
   assign m116_45 =10'b0;

   // m116_46 = W*in
   wire signed [9:0] m116_46;
   assign m116_46 =10'b0;

   // m116_47 = W*in
   wire signed [9:0] m116_47;
   assign m116_47 =10'b0;

   // m116_48 = W*in
   wire signed [9:0] m116_48;
   assign m116_48 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_49 = W*in
   wire signed [9:0] m116_49;
   assign m116_49 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_50 = W*in
   wire signed [9:0] m116_50;
   assign m116_50 ={ {2{in116[5]}} , in116 , {2{1'b0}} };

   // m116_51 = W*in
   wire signed [9:0] m116_51;
   assign m116_51 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_52 = W*in
   wire signed [9:0] m116_52;
   assign m116_52 =10'b0;

   // m116_53 = W*in
   wire signed [9:0] m116_53;
   assign m116_53 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_54 = W*in
   wire signed [9:0] m116_54;
   assign m116_54 =10'b0;

   // m116_55 = W*in
   wire signed [9:0] m116_55;
   assign m116_55 =10'b0;

   // m116_56 = W*in
   wire signed [9:0] m116_56;
   assign m116_56 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_57 = W*in
   wire signed [9:0] m116_57;
   assign m116_57 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_58 = W*in
   wire signed [9:0] m116_58;
   assign m116_58 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_59 = W*in
   wire signed [9:0] m116_59;
   assign m116_59 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_60 = W*in
   wire signed [9:0] m116_60;
   assign m116_60 =10'b0;

   // m116_61 = W*in
   wire signed [9:0] m116_61;
   assign m116_61 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_62 = W*in
   wire signed [9:0] m116_62;
   assign m116_62 =10'b0;

   // m116_63 = W*in
   wire signed [9:0] m116_63;
   assign m116_63 =10'b0;

   // m116_64 = W*in
   wire signed [9:0] m116_64;
   assign m116_64 =10'b0;

   // m116_65 = W*in
   wire signed [9:0] m116_65;
   assign m116_65 =10'b0;

   // m116_66 = W*in
   wire signed [9:0] m116_66;
   assign m116_66 =10'b0;

   // m116_67 = W*in
   wire signed [9:0] m116_67;
   assign m116_67 =10'b0;

   // m116_68 = W*in
   wire signed [9:0] m116_68;
   assign m116_68 ={ {3{neg116[5]}} , neg116 , {1{1'b0}} };

   // m116_69 = W*in
   wire signed [9:0] m116_69;
   assign m116_69 =10'b0;

   // m116_70 = W*in
   wire signed [9:0] m116_70;
   assign m116_70 =10'b0;

   // m116_71 = W*in
   wire signed [9:0] m116_71;
   assign m116_71 =10'b0;

   // m116_72 = W*in
   wire signed [9:0] m116_72;
   assign m116_72 =10'b0;

   // m116_73 = W*in
   wire signed [9:0] m116_73;
   assign m116_73 =10'b0;

   // m116_74 = W*in
   wire signed [9:0] m116_74;
   assign m116_74 =10'b0;

   // m116_75 = W*in
   wire signed [9:0] m116_75;
   assign m116_75 =10'b0;

   // m116_76 = W*in
   wire signed [9:0] m116_76;
   assign m116_76 =10'b0;

   // m116_77 = W*in
   wire signed [9:0] m116_77;
   assign m116_77 =10'b0;

   // m116_78 = W*in
   wire signed [9:0] m116_78;
   assign m116_78 ={ {3{in116[5]}} , in116 , {1{1'b0}} };

   // m116_79 = W*in
   wire signed [9:0] m116_79;
   assign m116_79 =10'b0;

   // m116_80 = W*in
   wire signed [9:0] m116_80;
   assign m116_80 =10'b0;

   // m116_81 = W*in
   wire signed [9:0] m116_81;
   assign m116_81 =10'b0;

   // m117_1 = W*in
   wire signed [9:0] m117_1;
   assign m117_1 =10'b0;

   // m117_2 = W*in
   wire signed [9:0] m117_2;
   assign m117_2 =10'b0;

   // m117_3 = W*in
   wire signed [9:0] m117_3;
   assign m117_3 =10'b0;

   // m117_4 = W*in
   wire signed [9:0] m117_4;
   assign m117_4 =10'b0;

   // m117_5 = W*in
   wire signed [9:0] m117_5;
   assign m117_5 =10'b0;

   // m117_6 = W*in
   wire signed [9:0] m117_6;
   assign m117_6 =10'b0;

   // m117_7 = W*in
   wire signed [9:0] m117_7;
   assign m117_7 =10'b0;

   // m117_8 = W*in
   wire signed [9:0] m117_8;
   assign m117_8 =10'b0;

   // m117_9 = W*in
   wire signed [9:0] m117_9;
   assign m117_9 =10'b0;

   // m117_10 = W*in
   wire signed [9:0] m117_10;
   assign m117_10 =10'b0;

   // m117_11 = W*in
   wire signed [9:0] m117_11;
   assign m117_11 =10'b0;

   // m117_12 = W*in
   wire signed [9:0] m117_12;
   assign m117_12 =10'b0;

   // m117_13 = W*in
   wire signed [9:0] m117_13;
   assign m117_13 =10'b0;

   // m117_14 = W*in
   wire signed [9:0] m117_14;
   assign m117_14 ={ {3{in117[5]}} , in117 , {1{1'b0}} };

   // m117_15 = W*in
   wire signed [9:0] m117_15;
   assign m117_15 ={ {3{in117[5]}} , in117 , {1{1'b0}} };

   // m117_16 = W*in
   wire signed [9:0] m117_16;
   assign m117_16 ={ {3{in117[5]}} , in117 , {1{1'b0}} };

   // m117_17 = W*in
   wire signed [9:0] m117_17;
   assign m117_17 =10'b0;

   // m117_18 = W*in
   wire signed [9:0] m117_18;
   assign m117_18 =10'b0;

   // m117_19 = W*in
   wire signed [9:0] m117_19;
   assign m117_19 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_20 = W*in
   wire signed [9:0] m117_20;
   assign m117_20 =10'b0;

   // m117_21 = W*in
   wire signed [9:0] m117_21;
   assign m117_21 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_22 = W*in
   wire signed [9:0] m117_22;
   assign m117_22 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_23 = W*in
   wire signed [9:0] m117_23;
   assign m117_23 =10'b0;

   // m117_24 = W*in
   wire signed [9:0] m117_24;
   assign m117_24 =10'b0;

   // m117_25 = W*in
   wire signed [9:0] m117_25;
   assign m117_25 =10'b0;

   // m117_26 = W*in
   wire signed [9:0] m117_26;
   assign m117_26 =10'b0;

   // m117_27 = W*in
   wire signed [9:0] m117_27;
   assign m117_27 ={ {3{in117[5]}} , in117 , {1{1'b0}} };

   // m117_28 = W*in
   wire signed [9:0] m117_28;
   assign m117_28 =10'b0;

   // m117_29 = W*in
   wire signed [9:0] m117_29;
   assign m117_29 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_30 = W*in
   wire signed [9:0] m117_30;
   assign m117_30 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   // m117_31 = W*in
   wire signed [9:0] m117_31;
   assign m117_31 =10'b0;

   // m117_32 = W*in
   wire signed [9:0] m117_32;
   assign m117_32 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   // m117_33 = W*in
   wire signed [9:0] m117_33;
   assign m117_33 =10'b0;

   // m117_34 = W*in
   wire signed [9:0] m117_34;
   assign m117_34 =10'b0;

   // m117_35 = W*in
   wire signed [9:0] m117_35;
   assign m117_35 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   // m117_36 = W*in
   wire signed [9:0] m117_36;
   assign m117_36 =10'b0;

   // m117_37 = W*in
   wire signed [9:0] m117_37;
   assign m117_37 =10'b0;

   // m117_38 = W*in
   wire signed [9:0] m117_38;
   assign m117_38 =10'b0;

   // m117_39 = W*in
   wire signed [9:0] m117_39;
   assign m117_39 =10'b0;

   // m117_40 = W*in
   wire signed [9:0] m117_40;
   assign m117_40 =10'b0;

   // m117_41 = W*in
   wire signed [9:0] m117_41;
   assign m117_41 =10'b0;

   // m117_42 = W*in
   wire signed [9:0] m117_42;
   assign m117_42 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_43 = W*in
   wire signed [9:0] m117_43;
   assign m117_43 ={ {3{in117[5]}} , in117 , {1{1'b0}} };

   // m117_44 = W*in
   wire signed [9:0] m117_44;
   assign m117_44 =10'b0;

   // m117_45 = W*in
   wire signed [9:0] m117_45;
   assign m117_45 =10'b0;

   // m117_46 = W*in
   wire signed [9:0] m117_46;
   assign m117_46 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   // m117_47 = W*in
   wire signed [9:0] m117_47;
   assign m117_47 =10'b0;

   // m117_48 = W*in
   wire signed [9:0] m117_48;
   assign m117_48 =10'b0;

   // m117_49 = W*in
   wire signed [9:0] m117_49;
   assign m117_49 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_50 = W*in
   wire signed [9:0] m117_50;
   assign m117_50 =10'b0;

   // m117_51 = W*in
   wire signed [9:0] m117_51;
   assign m117_51 =10'b0;

   // m117_52 = W*in
   wire signed [9:0] m117_52;
   assign m117_52 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_53 = W*in
   wire signed [9:0] m117_53;
   assign m117_53 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_54 = W*in
   wire signed [9:0] m117_54;
   assign m117_54 =10'b0;

   // m117_55 = W*in
   wire signed [9:0] m117_55;
   assign m117_55 =10'b0;

   // m117_56 = W*in
   wire signed [9:0] m117_56;
   assign m117_56 =10'b0;

   // m117_57 = W*in
   wire signed [9:0] m117_57;
   assign m117_57 =10'b0;

   // m117_58 = W*in
   wire signed [9:0] m117_58;
   assign m117_58 =10'b0;

   // m117_59 = W*in
   wire signed [9:0] m117_59;
   assign m117_59 =10'b0;

   // m117_60 = W*in
   wire signed [9:0] m117_60;
   assign m117_60 =10'b0;

   // m117_61 = W*in
   wire signed [9:0] m117_61;
   assign m117_61 =10'b0;

   // m117_62 = W*in
   wire signed [9:0] m117_62;
   assign m117_62 ={ {3{in117[5]}} , in117 , {1{1'b0}} };

   // m117_63 = W*in
   wire signed [9:0] m117_63;
   assign m117_63 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   // m117_64 = W*in
   wire signed [9:0] m117_64;
   assign m117_64 =10'b0;

   // m117_65 = W*in
   wire signed [9:0] m117_65;
   assign m117_65 =10'b0;

   // m117_66 = W*in
   wire signed [9:0] m117_66;
   assign m117_66 =10'b0;

   // m117_67 = W*in
   wire signed [9:0] m117_67;
   assign m117_67 =10'b0;

   // m117_68 = W*in
   wire signed [9:0] m117_68;
   assign m117_68 =10'b0;

   // m117_69 = W*in
   wire signed [9:0] m117_69;
   assign m117_69 =10'b0;

   // m117_70 = W*in
   wire signed [9:0] m117_70;
   assign m117_70 =10'b0;

   // m117_71 = W*in
   wire signed [9:0] m117_71;
   assign m117_71 =10'b0;

   // m117_72 = W*in
   wire signed [9:0] m117_72;
   assign m117_72 =10'b0;

   // m117_73 = W*in
   wire signed [9:0] m117_73;
   assign m117_73 =10'b0;

   // m117_74 = W*in
   wire signed [9:0] m117_74;
   assign m117_74 =10'b0;

   // m117_75 = W*in
   wire signed [9:0] m117_75;
   assign m117_75 =10'b0;

   // m117_76 = W*in
   wire signed [9:0] m117_76;
   assign m117_76 =10'b0;

   // m117_77 = W*in
   wire signed [9:0] m117_77;
   assign m117_77 ={ {3{neg117[5]}} , neg117 , {1{1'b0}} };

   // m117_78 = W*in
   wire signed [9:0] m117_78;
   assign m117_78 =10'b0;

   // m117_79 = W*in
   wire signed [9:0] m117_79;
   assign m117_79 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   // m117_80 = W*in
   wire signed [9:0] m117_80;
   assign m117_80 =10'b0;

   // m117_81 = W*in
   wire signed [9:0] m117_81;
   assign m117_81 ={ {2{in117[5]}} , in117 , {2{1'b0}} };

   //Perceptron Adders
   always @(posedge clk) out1 <= m1_1+m2_1+m3_1+m4_1+m5_1+m6_1+m7_1+m8_1+m9_1+m10_1+m11_1+m12_1+m13_1+m14_1+m15_1+m16_1+m17_1+m18_1+m19_1+m20_1+m21_1+m22_1+m23_1+m24_1+m25_1+m26_1+m27_1+m28_1+m29_1+m30_1+m31_1+m32_1+m33_1+m34_1+m35_1+m36_1+m37_1+m38_1+m39_1+m40_1+m41_1+m42_1+m43_1+m44_1+m45_1+m46_1+m47_1+m48_1+m49_1+m50_1+m51_1+m52_1+m53_1+m54_1+m55_1+m56_1+m57_1+m58_1+m59_1+m60_1+m61_1+m62_1+m63_1+m64_1+m65_1+m66_1+m67_1+m68_1+m69_1+m70_1+m71_1+m72_1+m73_1+m74_1+m75_1+m76_1+m77_1+m78_1+m79_1+m80_1+m81_1+m82_1+m83_1+m84_1+m85_1+m86_1+m87_1+m88_1+m89_1+m90_1+m91_1+m92_1+m93_1+m94_1+m95_1+m96_1+m97_1+m98_1+m99_1+m100_1+m101_1+m102_1+m103_1+m104_1+m105_1+m106_1+m107_1+m108_1+m109_1+m110_1+m111_1+m112_1+m113_1+m114_1+m115_1+m116_1+m117_1+b1;
   always @(posedge clk) out2 <= m1_2+m2_2+m3_2+m4_2+m5_2+m6_2+m7_2+m8_2+m9_2+m10_2+m11_2+m12_2+m13_2+m14_2+m15_2+m16_2+m17_2+m18_2+m19_2+m20_2+m21_2+m22_2+m23_2+m24_2+m25_2+m26_2+m27_2+m28_2+m29_2+m30_2+m31_2+m32_2+m33_2+m34_2+m35_2+m36_2+m37_2+m38_2+m39_2+m40_2+m41_2+m42_2+m43_2+m44_2+m45_2+m46_2+m47_2+m48_2+m49_2+m50_2+m51_2+m52_2+m53_2+m54_2+m55_2+m56_2+m57_2+m58_2+m59_2+m60_2+m61_2+m62_2+m63_2+m64_2+m65_2+m66_2+m67_2+m68_2+m69_2+m70_2+m71_2+m72_2+m73_2+m74_2+m75_2+m76_2+m77_2+m78_2+m79_2+m80_2+m81_2+m82_2+m83_2+m84_2+m85_2+m86_2+m87_2+m88_2+m89_2+m90_2+m91_2+m92_2+m93_2+m94_2+m95_2+m96_2+m97_2+m98_2+m99_2+m100_2+m101_2+m102_2+m103_2+m104_2+m105_2+m106_2+m107_2+m108_2+m109_2+m110_2+m111_2+m112_2+m113_2+m114_2+m115_2+m116_2+m117_2+b2;
   always @(posedge clk) out3 <= m1_3+m2_3+m3_3+m4_3+m5_3+m6_3+m7_3+m8_3+m9_3+m10_3+m11_3+m12_3+m13_3+m14_3+m15_3+m16_3+m17_3+m18_3+m19_3+m20_3+m21_3+m22_3+m23_3+m24_3+m25_3+m26_3+m27_3+m28_3+m29_3+m30_3+m31_3+m32_3+m33_3+m34_3+m35_3+m36_3+m37_3+m38_3+m39_3+m40_3+m41_3+m42_3+m43_3+m44_3+m45_3+m46_3+m47_3+m48_3+m49_3+m50_3+m51_3+m52_3+m53_3+m54_3+m55_3+m56_3+m57_3+m58_3+m59_3+m60_3+m61_3+m62_3+m63_3+m64_3+m65_3+m66_3+m67_3+m68_3+m69_3+m70_3+m71_3+m72_3+m73_3+m74_3+m75_3+m76_3+m77_3+m78_3+m79_3+m80_3+m81_3+m82_3+m83_3+m84_3+m85_3+m86_3+m87_3+m88_3+m89_3+m90_3+m91_3+m92_3+m93_3+m94_3+m95_3+m96_3+m97_3+m98_3+m99_3+m100_3+m101_3+m102_3+m103_3+m104_3+m105_3+m106_3+m107_3+m108_3+m109_3+m110_3+m111_3+m112_3+m113_3+m114_3+m115_3+m116_3+m117_3+b3;
   always @(posedge clk) out4 <= m1_4+m2_4+m3_4+m4_4+m5_4+m6_4+m7_4+m8_4+m9_4+m10_4+m11_4+m12_4+m13_4+m14_4+m15_4+m16_4+m17_4+m18_4+m19_4+m20_4+m21_4+m22_4+m23_4+m24_4+m25_4+m26_4+m27_4+m28_4+m29_4+m30_4+m31_4+m32_4+m33_4+m34_4+m35_4+m36_4+m37_4+m38_4+m39_4+m40_4+m41_4+m42_4+m43_4+m44_4+m45_4+m46_4+m47_4+m48_4+m49_4+m50_4+m51_4+m52_4+m53_4+m54_4+m55_4+m56_4+m57_4+m58_4+m59_4+m60_4+m61_4+m62_4+m63_4+m64_4+m65_4+m66_4+m67_4+m68_4+m69_4+m70_4+m71_4+m72_4+m73_4+m74_4+m75_4+m76_4+m77_4+m78_4+m79_4+m80_4+m81_4+m82_4+m83_4+m84_4+m85_4+m86_4+m87_4+m88_4+m89_4+m90_4+m91_4+m92_4+m93_4+m94_4+m95_4+m96_4+m97_4+m98_4+m99_4+m100_4+m101_4+m102_4+m103_4+m104_4+m105_4+m106_4+m107_4+m108_4+m109_4+m110_4+m111_4+m112_4+m113_4+m114_4+m115_4+m116_4+m117_4+b4;
   always @(posedge clk) out5 <= m1_5+m2_5+m3_5+m4_5+m5_5+m6_5+m7_5+m8_5+m9_5+m10_5+m11_5+m12_5+m13_5+m14_5+m15_5+m16_5+m17_5+m18_5+m19_5+m20_5+m21_5+m22_5+m23_5+m24_5+m25_5+m26_5+m27_5+m28_5+m29_5+m30_5+m31_5+m32_5+m33_5+m34_5+m35_5+m36_5+m37_5+m38_5+m39_5+m40_5+m41_5+m42_5+m43_5+m44_5+m45_5+m46_5+m47_5+m48_5+m49_5+m50_5+m51_5+m52_5+m53_5+m54_5+m55_5+m56_5+m57_5+m58_5+m59_5+m60_5+m61_5+m62_5+m63_5+m64_5+m65_5+m66_5+m67_5+m68_5+m69_5+m70_5+m71_5+m72_5+m73_5+m74_5+m75_5+m76_5+m77_5+m78_5+m79_5+m80_5+m81_5+m82_5+m83_5+m84_5+m85_5+m86_5+m87_5+m88_5+m89_5+m90_5+m91_5+m92_5+m93_5+m94_5+m95_5+m96_5+m97_5+m98_5+m99_5+m100_5+m101_5+m102_5+m103_5+m104_5+m105_5+m106_5+m107_5+m108_5+m109_5+m110_5+m111_5+m112_5+m113_5+m114_5+m115_5+m116_5+m117_5+b5;
   always @(posedge clk) out6 <= m1_6+m2_6+m3_6+m4_6+m5_6+m6_6+m7_6+m8_6+m9_6+m10_6+m11_6+m12_6+m13_6+m14_6+m15_6+m16_6+m17_6+m18_6+m19_6+m20_6+m21_6+m22_6+m23_6+m24_6+m25_6+m26_6+m27_6+m28_6+m29_6+m30_6+m31_6+m32_6+m33_6+m34_6+m35_6+m36_6+m37_6+m38_6+m39_6+m40_6+m41_6+m42_6+m43_6+m44_6+m45_6+m46_6+m47_6+m48_6+m49_6+m50_6+m51_6+m52_6+m53_6+m54_6+m55_6+m56_6+m57_6+m58_6+m59_6+m60_6+m61_6+m62_6+m63_6+m64_6+m65_6+m66_6+m67_6+m68_6+m69_6+m70_6+m71_6+m72_6+m73_6+m74_6+m75_6+m76_6+m77_6+m78_6+m79_6+m80_6+m81_6+m82_6+m83_6+m84_6+m85_6+m86_6+m87_6+m88_6+m89_6+m90_6+m91_6+m92_6+m93_6+m94_6+m95_6+m96_6+m97_6+m98_6+m99_6+m100_6+m101_6+m102_6+m103_6+m104_6+m105_6+m106_6+m107_6+m108_6+m109_6+m110_6+m111_6+m112_6+m113_6+m114_6+m115_6+m116_6+m117_6+b6;
   always @(posedge clk) out7 <= m1_7+m2_7+m3_7+m4_7+m5_7+m6_7+m7_7+m8_7+m9_7+m10_7+m11_7+m12_7+m13_7+m14_7+m15_7+m16_7+m17_7+m18_7+m19_7+m20_7+m21_7+m22_7+m23_7+m24_7+m25_7+m26_7+m27_7+m28_7+m29_7+m30_7+m31_7+m32_7+m33_7+m34_7+m35_7+m36_7+m37_7+m38_7+m39_7+m40_7+m41_7+m42_7+m43_7+m44_7+m45_7+m46_7+m47_7+m48_7+m49_7+m50_7+m51_7+m52_7+m53_7+m54_7+m55_7+m56_7+m57_7+m58_7+m59_7+m60_7+m61_7+m62_7+m63_7+m64_7+m65_7+m66_7+m67_7+m68_7+m69_7+m70_7+m71_7+m72_7+m73_7+m74_7+m75_7+m76_7+m77_7+m78_7+m79_7+m80_7+m81_7+m82_7+m83_7+m84_7+m85_7+m86_7+m87_7+m88_7+m89_7+m90_7+m91_7+m92_7+m93_7+m94_7+m95_7+m96_7+m97_7+m98_7+m99_7+m100_7+m101_7+m102_7+m103_7+m104_7+m105_7+m106_7+m107_7+m108_7+m109_7+m110_7+m111_7+m112_7+m113_7+m114_7+m115_7+m116_7+m117_7+b7;
   always @(posedge clk) out8 <= m1_8+m2_8+m3_8+m4_8+m5_8+m6_8+m7_8+m8_8+m9_8+m10_8+m11_8+m12_8+m13_8+m14_8+m15_8+m16_8+m17_8+m18_8+m19_8+m20_8+m21_8+m22_8+m23_8+m24_8+m25_8+m26_8+m27_8+m28_8+m29_8+m30_8+m31_8+m32_8+m33_8+m34_8+m35_8+m36_8+m37_8+m38_8+m39_8+m40_8+m41_8+m42_8+m43_8+m44_8+m45_8+m46_8+m47_8+m48_8+m49_8+m50_8+m51_8+m52_8+m53_8+m54_8+m55_8+m56_8+m57_8+m58_8+m59_8+m60_8+m61_8+m62_8+m63_8+m64_8+m65_8+m66_8+m67_8+m68_8+m69_8+m70_8+m71_8+m72_8+m73_8+m74_8+m75_8+m76_8+m77_8+m78_8+m79_8+m80_8+m81_8+m82_8+m83_8+m84_8+m85_8+m86_8+m87_8+m88_8+m89_8+m90_8+m91_8+m92_8+m93_8+m94_8+m95_8+m96_8+m97_8+m98_8+m99_8+m100_8+m101_8+m102_8+m103_8+m104_8+m105_8+m106_8+m107_8+m108_8+m109_8+m110_8+m111_8+m112_8+m113_8+m114_8+m115_8+m116_8+m117_8+b8;
   always @(posedge clk) out9 <= m1_9+m2_9+m3_9+m4_9+m5_9+m6_9+m7_9+m8_9+m9_9+m10_9+m11_9+m12_9+m13_9+m14_9+m15_9+m16_9+m17_9+m18_9+m19_9+m20_9+m21_9+m22_9+m23_9+m24_9+m25_9+m26_9+m27_9+m28_9+m29_9+m30_9+m31_9+m32_9+m33_9+m34_9+m35_9+m36_9+m37_9+m38_9+m39_9+m40_9+m41_9+m42_9+m43_9+m44_9+m45_9+m46_9+m47_9+m48_9+m49_9+m50_9+m51_9+m52_9+m53_9+m54_9+m55_9+m56_9+m57_9+m58_9+m59_9+m60_9+m61_9+m62_9+m63_9+m64_9+m65_9+m66_9+m67_9+m68_9+m69_9+m70_9+m71_9+m72_9+m73_9+m74_9+m75_9+m76_9+m77_9+m78_9+m79_9+m80_9+m81_9+m82_9+m83_9+m84_9+m85_9+m86_9+m87_9+m88_9+m89_9+m90_9+m91_9+m92_9+m93_9+m94_9+m95_9+m96_9+m97_9+m98_9+m99_9+m100_9+m101_9+m102_9+m103_9+m104_9+m105_9+m106_9+m107_9+m108_9+m109_9+m110_9+m111_9+m112_9+m113_9+m114_9+m115_9+m116_9+m117_9+b9;
   always @(posedge clk) out10 <= m1_10+m2_10+m3_10+m4_10+m5_10+m6_10+m7_10+m8_10+m9_10+m10_10+m11_10+m12_10+m13_10+m14_10+m15_10+m16_10+m17_10+m18_10+m19_10+m20_10+m21_10+m22_10+m23_10+m24_10+m25_10+m26_10+m27_10+m28_10+m29_10+m30_10+m31_10+m32_10+m33_10+m34_10+m35_10+m36_10+m37_10+m38_10+m39_10+m40_10+m41_10+m42_10+m43_10+m44_10+m45_10+m46_10+m47_10+m48_10+m49_10+m50_10+m51_10+m52_10+m53_10+m54_10+m55_10+m56_10+m57_10+m58_10+m59_10+m60_10+m61_10+m62_10+m63_10+m64_10+m65_10+m66_10+m67_10+m68_10+m69_10+m70_10+m71_10+m72_10+m73_10+m74_10+m75_10+m76_10+m77_10+m78_10+m79_10+m80_10+m81_10+m82_10+m83_10+m84_10+m85_10+m86_10+m87_10+m88_10+m89_10+m90_10+m91_10+m92_10+m93_10+m94_10+m95_10+m96_10+m97_10+m98_10+m99_10+m100_10+m101_10+m102_10+m103_10+m104_10+m105_10+m106_10+m107_10+m108_10+m109_10+m110_10+m111_10+m112_10+m113_10+m114_10+m115_10+m116_10+m117_10+b10;
   always @(posedge clk) out11 <= m1_11+m2_11+m3_11+m4_11+m5_11+m6_11+m7_11+m8_11+m9_11+m10_11+m11_11+m12_11+m13_11+m14_11+m15_11+m16_11+m17_11+m18_11+m19_11+m20_11+m21_11+m22_11+m23_11+m24_11+m25_11+m26_11+m27_11+m28_11+m29_11+m30_11+m31_11+m32_11+m33_11+m34_11+m35_11+m36_11+m37_11+m38_11+m39_11+m40_11+m41_11+m42_11+m43_11+m44_11+m45_11+m46_11+m47_11+m48_11+m49_11+m50_11+m51_11+m52_11+m53_11+m54_11+m55_11+m56_11+m57_11+m58_11+m59_11+m60_11+m61_11+m62_11+m63_11+m64_11+m65_11+m66_11+m67_11+m68_11+m69_11+m70_11+m71_11+m72_11+m73_11+m74_11+m75_11+m76_11+m77_11+m78_11+m79_11+m80_11+m81_11+m82_11+m83_11+m84_11+m85_11+m86_11+m87_11+m88_11+m89_11+m90_11+m91_11+m92_11+m93_11+m94_11+m95_11+m96_11+m97_11+m98_11+m99_11+m100_11+m101_11+m102_11+m103_11+m104_11+m105_11+m106_11+m107_11+m108_11+m109_11+m110_11+m111_11+m112_11+m113_11+m114_11+m115_11+m116_11+m117_11+b11;
   always @(posedge clk) out12 <= m1_12+m2_12+m3_12+m4_12+m5_12+m6_12+m7_12+m8_12+m9_12+m10_12+m11_12+m12_12+m13_12+m14_12+m15_12+m16_12+m17_12+m18_12+m19_12+m20_12+m21_12+m22_12+m23_12+m24_12+m25_12+m26_12+m27_12+m28_12+m29_12+m30_12+m31_12+m32_12+m33_12+m34_12+m35_12+m36_12+m37_12+m38_12+m39_12+m40_12+m41_12+m42_12+m43_12+m44_12+m45_12+m46_12+m47_12+m48_12+m49_12+m50_12+m51_12+m52_12+m53_12+m54_12+m55_12+m56_12+m57_12+m58_12+m59_12+m60_12+m61_12+m62_12+m63_12+m64_12+m65_12+m66_12+m67_12+m68_12+m69_12+m70_12+m71_12+m72_12+m73_12+m74_12+m75_12+m76_12+m77_12+m78_12+m79_12+m80_12+m81_12+m82_12+m83_12+m84_12+m85_12+m86_12+m87_12+m88_12+m89_12+m90_12+m91_12+m92_12+m93_12+m94_12+m95_12+m96_12+m97_12+m98_12+m99_12+m100_12+m101_12+m102_12+m103_12+m104_12+m105_12+m106_12+m107_12+m108_12+m109_12+m110_12+m111_12+m112_12+m113_12+m114_12+m115_12+m116_12+m117_12+b12;
   always @(posedge clk) out13 <= m1_13+m2_13+m3_13+m4_13+m5_13+m6_13+m7_13+m8_13+m9_13+m10_13+m11_13+m12_13+m13_13+m14_13+m15_13+m16_13+m17_13+m18_13+m19_13+m20_13+m21_13+m22_13+m23_13+m24_13+m25_13+m26_13+m27_13+m28_13+m29_13+m30_13+m31_13+m32_13+m33_13+m34_13+m35_13+m36_13+m37_13+m38_13+m39_13+m40_13+m41_13+m42_13+m43_13+m44_13+m45_13+m46_13+m47_13+m48_13+m49_13+m50_13+m51_13+m52_13+m53_13+m54_13+m55_13+m56_13+m57_13+m58_13+m59_13+m60_13+m61_13+m62_13+m63_13+m64_13+m65_13+m66_13+m67_13+m68_13+m69_13+m70_13+m71_13+m72_13+m73_13+m74_13+m75_13+m76_13+m77_13+m78_13+m79_13+m80_13+m81_13+m82_13+m83_13+m84_13+m85_13+m86_13+m87_13+m88_13+m89_13+m90_13+m91_13+m92_13+m93_13+m94_13+m95_13+m96_13+m97_13+m98_13+m99_13+m100_13+m101_13+m102_13+m103_13+m104_13+m105_13+m106_13+m107_13+m108_13+m109_13+m110_13+m111_13+m112_13+m113_13+m114_13+m115_13+m116_13+m117_13+b13;
   always @(posedge clk) out14 <= m1_14+m2_14+m3_14+m4_14+m5_14+m6_14+m7_14+m8_14+m9_14+m10_14+m11_14+m12_14+m13_14+m14_14+m15_14+m16_14+m17_14+m18_14+m19_14+m20_14+m21_14+m22_14+m23_14+m24_14+m25_14+m26_14+m27_14+m28_14+m29_14+m30_14+m31_14+m32_14+m33_14+m34_14+m35_14+m36_14+m37_14+m38_14+m39_14+m40_14+m41_14+m42_14+m43_14+m44_14+m45_14+m46_14+m47_14+m48_14+m49_14+m50_14+m51_14+m52_14+m53_14+m54_14+m55_14+m56_14+m57_14+m58_14+m59_14+m60_14+m61_14+m62_14+m63_14+m64_14+m65_14+m66_14+m67_14+m68_14+m69_14+m70_14+m71_14+m72_14+m73_14+m74_14+m75_14+m76_14+m77_14+m78_14+m79_14+m80_14+m81_14+m82_14+m83_14+m84_14+m85_14+m86_14+m87_14+m88_14+m89_14+m90_14+m91_14+m92_14+m93_14+m94_14+m95_14+m96_14+m97_14+m98_14+m99_14+m100_14+m101_14+m102_14+m103_14+m104_14+m105_14+m106_14+m107_14+m108_14+m109_14+m110_14+m111_14+m112_14+m113_14+m114_14+m115_14+m116_14+m117_14+b14;
   always @(posedge clk) out15 <= m1_15+m2_15+m3_15+m4_15+m5_15+m6_15+m7_15+m8_15+m9_15+m10_15+m11_15+m12_15+m13_15+m14_15+m15_15+m16_15+m17_15+m18_15+m19_15+m20_15+m21_15+m22_15+m23_15+m24_15+m25_15+m26_15+m27_15+m28_15+m29_15+m30_15+m31_15+m32_15+m33_15+m34_15+m35_15+m36_15+m37_15+m38_15+m39_15+m40_15+m41_15+m42_15+m43_15+m44_15+m45_15+m46_15+m47_15+m48_15+m49_15+m50_15+m51_15+m52_15+m53_15+m54_15+m55_15+m56_15+m57_15+m58_15+m59_15+m60_15+m61_15+m62_15+m63_15+m64_15+m65_15+m66_15+m67_15+m68_15+m69_15+m70_15+m71_15+m72_15+m73_15+m74_15+m75_15+m76_15+m77_15+m78_15+m79_15+m80_15+m81_15+m82_15+m83_15+m84_15+m85_15+m86_15+m87_15+m88_15+m89_15+m90_15+m91_15+m92_15+m93_15+m94_15+m95_15+m96_15+m97_15+m98_15+m99_15+m100_15+m101_15+m102_15+m103_15+m104_15+m105_15+m106_15+m107_15+m108_15+m109_15+m110_15+m111_15+m112_15+m113_15+m114_15+m115_15+m116_15+m117_15+b15;
   always @(posedge clk) out16 <= m1_16+m2_16+m3_16+m4_16+m5_16+m6_16+m7_16+m8_16+m9_16+m10_16+m11_16+m12_16+m13_16+m14_16+m15_16+m16_16+m17_16+m18_16+m19_16+m20_16+m21_16+m22_16+m23_16+m24_16+m25_16+m26_16+m27_16+m28_16+m29_16+m30_16+m31_16+m32_16+m33_16+m34_16+m35_16+m36_16+m37_16+m38_16+m39_16+m40_16+m41_16+m42_16+m43_16+m44_16+m45_16+m46_16+m47_16+m48_16+m49_16+m50_16+m51_16+m52_16+m53_16+m54_16+m55_16+m56_16+m57_16+m58_16+m59_16+m60_16+m61_16+m62_16+m63_16+m64_16+m65_16+m66_16+m67_16+m68_16+m69_16+m70_16+m71_16+m72_16+m73_16+m74_16+m75_16+m76_16+m77_16+m78_16+m79_16+m80_16+m81_16+m82_16+m83_16+m84_16+m85_16+m86_16+m87_16+m88_16+m89_16+m90_16+m91_16+m92_16+m93_16+m94_16+m95_16+m96_16+m97_16+m98_16+m99_16+m100_16+m101_16+m102_16+m103_16+m104_16+m105_16+m106_16+m107_16+m108_16+m109_16+m110_16+m111_16+m112_16+m113_16+m114_16+m115_16+m116_16+m117_16+b16;
   always @(posedge clk) out17 <= m1_17+m2_17+m3_17+m4_17+m5_17+m6_17+m7_17+m8_17+m9_17+m10_17+m11_17+m12_17+m13_17+m14_17+m15_17+m16_17+m17_17+m18_17+m19_17+m20_17+m21_17+m22_17+m23_17+m24_17+m25_17+m26_17+m27_17+m28_17+m29_17+m30_17+m31_17+m32_17+m33_17+m34_17+m35_17+m36_17+m37_17+m38_17+m39_17+m40_17+m41_17+m42_17+m43_17+m44_17+m45_17+m46_17+m47_17+m48_17+m49_17+m50_17+m51_17+m52_17+m53_17+m54_17+m55_17+m56_17+m57_17+m58_17+m59_17+m60_17+m61_17+m62_17+m63_17+m64_17+m65_17+m66_17+m67_17+m68_17+m69_17+m70_17+m71_17+m72_17+m73_17+m74_17+m75_17+m76_17+m77_17+m78_17+m79_17+m80_17+m81_17+m82_17+m83_17+m84_17+m85_17+m86_17+m87_17+m88_17+m89_17+m90_17+m91_17+m92_17+m93_17+m94_17+m95_17+m96_17+m97_17+m98_17+m99_17+m100_17+m101_17+m102_17+m103_17+m104_17+m105_17+m106_17+m107_17+m108_17+m109_17+m110_17+m111_17+m112_17+m113_17+m114_17+m115_17+m116_17+m117_17+b17;
   always @(posedge clk) out18 <= m1_18+m2_18+m3_18+m4_18+m5_18+m6_18+m7_18+m8_18+m9_18+m10_18+m11_18+m12_18+m13_18+m14_18+m15_18+m16_18+m17_18+m18_18+m19_18+m20_18+m21_18+m22_18+m23_18+m24_18+m25_18+m26_18+m27_18+m28_18+m29_18+m30_18+m31_18+m32_18+m33_18+m34_18+m35_18+m36_18+m37_18+m38_18+m39_18+m40_18+m41_18+m42_18+m43_18+m44_18+m45_18+m46_18+m47_18+m48_18+m49_18+m50_18+m51_18+m52_18+m53_18+m54_18+m55_18+m56_18+m57_18+m58_18+m59_18+m60_18+m61_18+m62_18+m63_18+m64_18+m65_18+m66_18+m67_18+m68_18+m69_18+m70_18+m71_18+m72_18+m73_18+m74_18+m75_18+m76_18+m77_18+m78_18+m79_18+m80_18+m81_18+m82_18+m83_18+m84_18+m85_18+m86_18+m87_18+m88_18+m89_18+m90_18+m91_18+m92_18+m93_18+m94_18+m95_18+m96_18+m97_18+m98_18+m99_18+m100_18+m101_18+m102_18+m103_18+m104_18+m105_18+m106_18+m107_18+m108_18+m109_18+m110_18+m111_18+m112_18+m113_18+m114_18+m115_18+m116_18+m117_18+b18;
   always @(posedge clk) out19 <= m1_19+m2_19+m3_19+m4_19+m5_19+m6_19+m7_19+m8_19+m9_19+m10_19+m11_19+m12_19+m13_19+m14_19+m15_19+m16_19+m17_19+m18_19+m19_19+m20_19+m21_19+m22_19+m23_19+m24_19+m25_19+m26_19+m27_19+m28_19+m29_19+m30_19+m31_19+m32_19+m33_19+m34_19+m35_19+m36_19+m37_19+m38_19+m39_19+m40_19+m41_19+m42_19+m43_19+m44_19+m45_19+m46_19+m47_19+m48_19+m49_19+m50_19+m51_19+m52_19+m53_19+m54_19+m55_19+m56_19+m57_19+m58_19+m59_19+m60_19+m61_19+m62_19+m63_19+m64_19+m65_19+m66_19+m67_19+m68_19+m69_19+m70_19+m71_19+m72_19+m73_19+m74_19+m75_19+m76_19+m77_19+m78_19+m79_19+m80_19+m81_19+m82_19+m83_19+m84_19+m85_19+m86_19+m87_19+m88_19+m89_19+m90_19+m91_19+m92_19+m93_19+m94_19+m95_19+m96_19+m97_19+m98_19+m99_19+m100_19+m101_19+m102_19+m103_19+m104_19+m105_19+m106_19+m107_19+m108_19+m109_19+m110_19+m111_19+m112_19+m113_19+m114_19+m115_19+m116_19+m117_19+b19;
   always @(posedge clk) out20 <= m1_20+m2_20+m3_20+m4_20+m5_20+m6_20+m7_20+m8_20+m9_20+m10_20+m11_20+m12_20+m13_20+m14_20+m15_20+m16_20+m17_20+m18_20+m19_20+m20_20+m21_20+m22_20+m23_20+m24_20+m25_20+m26_20+m27_20+m28_20+m29_20+m30_20+m31_20+m32_20+m33_20+m34_20+m35_20+m36_20+m37_20+m38_20+m39_20+m40_20+m41_20+m42_20+m43_20+m44_20+m45_20+m46_20+m47_20+m48_20+m49_20+m50_20+m51_20+m52_20+m53_20+m54_20+m55_20+m56_20+m57_20+m58_20+m59_20+m60_20+m61_20+m62_20+m63_20+m64_20+m65_20+m66_20+m67_20+m68_20+m69_20+m70_20+m71_20+m72_20+m73_20+m74_20+m75_20+m76_20+m77_20+m78_20+m79_20+m80_20+m81_20+m82_20+m83_20+m84_20+m85_20+m86_20+m87_20+m88_20+m89_20+m90_20+m91_20+m92_20+m93_20+m94_20+m95_20+m96_20+m97_20+m98_20+m99_20+m100_20+m101_20+m102_20+m103_20+m104_20+m105_20+m106_20+m107_20+m108_20+m109_20+m110_20+m111_20+m112_20+m113_20+m114_20+m115_20+m116_20+m117_20+b20;
   always @(posedge clk) out21 <= m1_21+m2_21+m3_21+m4_21+m5_21+m6_21+m7_21+m8_21+m9_21+m10_21+m11_21+m12_21+m13_21+m14_21+m15_21+m16_21+m17_21+m18_21+m19_21+m20_21+m21_21+m22_21+m23_21+m24_21+m25_21+m26_21+m27_21+m28_21+m29_21+m30_21+m31_21+m32_21+m33_21+m34_21+m35_21+m36_21+m37_21+m38_21+m39_21+m40_21+m41_21+m42_21+m43_21+m44_21+m45_21+m46_21+m47_21+m48_21+m49_21+m50_21+m51_21+m52_21+m53_21+m54_21+m55_21+m56_21+m57_21+m58_21+m59_21+m60_21+m61_21+m62_21+m63_21+m64_21+m65_21+m66_21+m67_21+m68_21+m69_21+m70_21+m71_21+m72_21+m73_21+m74_21+m75_21+m76_21+m77_21+m78_21+m79_21+m80_21+m81_21+m82_21+m83_21+m84_21+m85_21+m86_21+m87_21+m88_21+m89_21+m90_21+m91_21+m92_21+m93_21+m94_21+m95_21+m96_21+m97_21+m98_21+m99_21+m100_21+m101_21+m102_21+m103_21+m104_21+m105_21+m106_21+m107_21+m108_21+m109_21+m110_21+m111_21+m112_21+m113_21+m114_21+m115_21+m116_21+m117_21+b21;
   always @(posedge clk) out22 <= m1_22+m2_22+m3_22+m4_22+m5_22+m6_22+m7_22+m8_22+m9_22+m10_22+m11_22+m12_22+m13_22+m14_22+m15_22+m16_22+m17_22+m18_22+m19_22+m20_22+m21_22+m22_22+m23_22+m24_22+m25_22+m26_22+m27_22+m28_22+m29_22+m30_22+m31_22+m32_22+m33_22+m34_22+m35_22+m36_22+m37_22+m38_22+m39_22+m40_22+m41_22+m42_22+m43_22+m44_22+m45_22+m46_22+m47_22+m48_22+m49_22+m50_22+m51_22+m52_22+m53_22+m54_22+m55_22+m56_22+m57_22+m58_22+m59_22+m60_22+m61_22+m62_22+m63_22+m64_22+m65_22+m66_22+m67_22+m68_22+m69_22+m70_22+m71_22+m72_22+m73_22+m74_22+m75_22+m76_22+m77_22+m78_22+m79_22+m80_22+m81_22+m82_22+m83_22+m84_22+m85_22+m86_22+m87_22+m88_22+m89_22+m90_22+m91_22+m92_22+m93_22+m94_22+m95_22+m96_22+m97_22+m98_22+m99_22+m100_22+m101_22+m102_22+m103_22+m104_22+m105_22+m106_22+m107_22+m108_22+m109_22+m110_22+m111_22+m112_22+m113_22+m114_22+m115_22+m116_22+m117_22+b22;
   always @(posedge clk) out23 <= m1_23+m2_23+m3_23+m4_23+m5_23+m6_23+m7_23+m8_23+m9_23+m10_23+m11_23+m12_23+m13_23+m14_23+m15_23+m16_23+m17_23+m18_23+m19_23+m20_23+m21_23+m22_23+m23_23+m24_23+m25_23+m26_23+m27_23+m28_23+m29_23+m30_23+m31_23+m32_23+m33_23+m34_23+m35_23+m36_23+m37_23+m38_23+m39_23+m40_23+m41_23+m42_23+m43_23+m44_23+m45_23+m46_23+m47_23+m48_23+m49_23+m50_23+m51_23+m52_23+m53_23+m54_23+m55_23+m56_23+m57_23+m58_23+m59_23+m60_23+m61_23+m62_23+m63_23+m64_23+m65_23+m66_23+m67_23+m68_23+m69_23+m70_23+m71_23+m72_23+m73_23+m74_23+m75_23+m76_23+m77_23+m78_23+m79_23+m80_23+m81_23+m82_23+m83_23+m84_23+m85_23+m86_23+m87_23+m88_23+m89_23+m90_23+m91_23+m92_23+m93_23+m94_23+m95_23+m96_23+m97_23+m98_23+m99_23+m100_23+m101_23+m102_23+m103_23+m104_23+m105_23+m106_23+m107_23+m108_23+m109_23+m110_23+m111_23+m112_23+m113_23+m114_23+m115_23+m116_23+m117_23+b23;
   always @(posedge clk) out24 <= m1_24+m2_24+m3_24+m4_24+m5_24+m6_24+m7_24+m8_24+m9_24+m10_24+m11_24+m12_24+m13_24+m14_24+m15_24+m16_24+m17_24+m18_24+m19_24+m20_24+m21_24+m22_24+m23_24+m24_24+m25_24+m26_24+m27_24+m28_24+m29_24+m30_24+m31_24+m32_24+m33_24+m34_24+m35_24+m36_24+m37_24+m38_24+m39_24+m40_24+m41_24+m42_24+m43_24+m44_24+m45_24+m46_24+m47_24+m48_24+m49_24+m50_24+m51_24+m52_24+m53_24+m54_24+m55_24+m56_24+m57_24+m58_24+m59_24+m60_24+m61_24+m62_24+m63_24+m64_24+m65_24+m66_24+m67_24+m68_24+m69_24+m70_24+m71_24+m72_24+m73_24+m74_24+m75_24+m76_24+m77_24+m78_24+m79_24+m80_24+m81_24+m82_24+m83_24+m84_24+m85_24+m86_24+m87_24+m88_24+m89_24+m90_24+m91_24+m92_24+m93_24+m94_24+m95_24+m96_24+m97_24+m98_24+m99_24+m100_24+m101_24+m102_24+m103_24+m104_24+m105_24+m106_24+m107_24+m108_24+m109_24+m110_24+m111_24+m112_24+m113_24+m114_24+m115_24+m116_24+m117_24+b24;
   always @(posedge clk) out25 <= m1_25+m2_25+m3_25+m4_25+m5_25+m6_25+m7_25+m8_25+m9_25+m10_25+m11_25+m12_25+m13_25+m14_25+m15_25+m16_25+m17_25+m18_25+m19_25+m20_25+m21_25+m22_25+m23_25+m24_25+m25_25+m26_25+m27_25+m28_25+m29_25+m30_25+m31_25+m32_25+m33_25+m34_25+m35_25+m36_25+m37_25+m38_25+m39_25+m40_25+m41_25+m42_25+m43_25+m44_25+m45_25+m46_25+m47_25+m48_25+m49_25+m50_25+m51_25+m52_25+m53_25+m54_25+m55_25+m56_25+m57_25+m58_25+m59_25+m60_25+m61_25+m62_25+m63_25+m64_25+m65_25+m66_25+m67_25+m68_25+m69_25+m70_25+m71_25+m72_25+m73_25+m74_25+m75_25+m76_25+m77_25+m78_25+m79_25+m80_25+m81_25+m82_25+m83_25+m84_25+m85_25+m86_25+m87_25+m88_25+m89_25+m90_25+m91_25+m92_25+m93_25+m94_25+m95_25+m96_25+m97_25+m98_25+m99_25+m100_25+m101_25+m102_25+m103_25+m104_25+m105_25+m106_25+m107_25+m108_25+m109_25+m110_25+m111_25+m112_25+m113_25+m114_25+m115_25+m116_25+m117_25+b25;
   always @(posedge clk) out26 <= m1_26+m2_26+m3_26+m4_26+m5_26+m6_26+m7_26+m8_26+m9_26+m10_26+m11_26+m12_26+m13_26+m14_26+m15_26+m16_26+m17_26+m18_26+m19_26+m20_26+m21_26+m22_26+m23_26+m24_26+m25_26+m26_26+m27_26+m28_26+m29_26+m30_26+m31_26+m32_26+m33_26+m34_26+m35_26+m36_26+m37_26+m38_26+m39_26+m40_26+m41_26+m42_26+m43_26+m44_26+m45_26+m46_26+m47_26+m48_26+m49_26+m50_26+m51_26+m52_26+m53_26+m54_26+m55_26+m56_26+m57_26+m58_26+m59_26+m60_26+m61_26+m62_26+m63_26+m64_26+m65_26+m66_26+m67_26+m68_26+m69_26+m70_26+m71_26+m72_26+m73_26+m74_26+m75_26+m76_26+m77_26+m78_26+m79_26+m80_26+m81_26+m82_26+m83_26+m84_26+m85_26+m86_26+m87_26+m88_26+m89_26+m90_26+m91_26+m92_26+m93_26+m94_26+m95_26+m96_26+m97_26+m98_26+m99_26+m100_26+m101_26+m102_26+m103_26+m104_26+m105_26+m106_26+m107_26+m108_26+m109_26+m110_26+m111_26+m112_26+m113_26+m114_26+m115_26+m116_26+m117_26+b26;
   always @(posedge clk) out27 <= m1_27+m2_27+m3_27+m4_27+m5_27+m6_27+m7_27+m8_27+m9_27+m10_27+m11_27+m12_27+m13_27+m14_27+m15_27+m16_27+m17_27+m18_27+m19_27+m20_27+m21_27+m22_27+m23_27+m24_27+m25_27+m26_27+m27_27+m28_27+m29_27+m30_27+m31_27+m32_27+m33_27+m34_27+m35_27+m36_27+m37_27+m38_27+m39_27+m40_27+m41_27+m42_27+m43_27+m44_27+m45_27+m46_27+m47_27+m48_27+m49_27+m50_27+m51_27+m52_27+m53_27+m54_27+m55_27+m56_27+m57_27+m58_27+m59_27+m60_27+m61_27+m62_27+m63_27+m64_27+m65_27+m66_27+m67_27+m68_27+m69_27+m70_27+m71_27+m72_27+m73_27+m74_27+m75_27+m76_27+m77_27+m78_27+m79_27+m80_27+m81_27+m82_27+m83_27+m84_27+m85_27+m86_27+m87_27+m88_27+m89_27+m90_27+m91_27+m92_27+m93_27+m94_27+m95_27+m96_27+m97_27+m98_27+m99_27+m100_27+m101_27+m102_27+m103_27+m104_27+m105_27+m106_27+m107_27+m108_27+m109_27+m110_27+m111_27+m112_27+m113_27+m114_27+m115_27+m116_27+m117_27+b27;
   always @(posedge clk) out28 <= m1_28+m2_28+m3_28+m4_28+m5_28+m6_28+m7_28+m8_28+m9_28+m10_28+m11_28+m12_28+m13_28+m14_28+m15_28+m16_28+m17_28+m18_28+m19_28+m20_28+m21_28+m22_28+m23_28+m24_28+m25_28+m26_28+m27_28+m28_28+m29_28+m30_28+m31_28+m32_28+m33_28+m34_28+m35_28+m36_28+m37_28+m38_28+m39_28+m40_28+m41_28+m42_28+m43_28+m44_28+m45_28+m46_28+m47_28+m48_28+m49_28+m50_28+m51_28+m52_28+m53_28+m54_28+m55_28+m56_28+m57_28+m58_28+m59_28+m60_28+m61_28+m62_28+m63_28+m64_28+m65_28+m66_28+m67_28+m68_28+m69_28+m70_28+m71_28+m72_28+m73_28+m74_28+m75_28+m76_28+m77_28+m78_28+m79_28+m80_28+m81_28+m82_28+m83_28+m84_28+m85_28+m86_28+m87_28+m88_28+m89_28+m90_28+m91_28+m92_28+m93_28+m94_28+m95_28+m96_28+m97_28+m98_28+m99_28+m100_28+m101_28+m102_28+m103_28+m104_28+m105_28+m106_28+m107_28+m108_28+m109_28+m110_28+m111_28+m112_28+m113_28+m114_28+m115_28+m116_28+m117_28+b28;
   always @(posedge clk) out29 <= m1_29+m2_29+m3_29+m4_29+m5_29+m6_29+m7_29+m8_29+m9_29+m10_29+m11_29+m12_29+m13_29+m14_29+m15_29+m16_29+m17_29+m18_29+m19_29+m20_29+m21_29+m22_29+m23_29+m24_29+m25_29+m26_29+m27_29+m28_29+m29_29+m30_29+m31_29+m32_29+m33_29+m34_29+m35_29+m36_29+m37_29+m38_29+m39_29+m40_29+m41_29+m42_29+m43_29+m44_29+m45_29+m46_29+m47_29+m48_29+m49_29+m50_29+m51_29+m52_29+m53_29+m54_29+m55_29+m56_29+m57_29+m58_29+m59_29+m60_29+m61_29+m62_29+m63_29+m64_29+m65_29+m66_29+m67_29+m68_29+m69_29+m70_29+m71_29+m72_29+m73_29+m74_29+m75_29+m76_29+m77_29+m78_29+m79_29+m80_29+m81_29+m82_29+m83_29+m84_29+m85_29+m86_29+m87_29+m88_29+m89_29+m90_29+m91_29+m92_29+m93_29+m94_29+m95_29+m96_29+m97_29+m98_29+m99_29+m100_29+m101_29+m102_29+m103_29+m104_29+m105_29+m106_29+m107_29+m108_29+m109_29+m110_29+m111_29+m112_29+m113_29+m114_29+m115_29+m116_29+m117_29+b29;
   always @(posedge clk) out30 <= m1_30+m2_30+m3_30+m4_30+m5_30+m6_30+m7_30+m8_30+m9_30+m10_30+m11_30+m12_30+m13_30+m14_30+m15_30+m16_30+m17_30+m18_30+m19_30+m20_30+m21_30+m22_30+m23_30+m24_30+m25_30+m26_30+m27_30+m28_30+m29_30+m30_30+m31_30+m32_30+m33_30+m34_30+m35_30+m36_30+m37_30+m38_30+m39_30+m40_30+m41_30+m42_30+m43_30+m44_30+m45_30+m46_30+m47_30+m48_30+m49_30+m50_30+m51_30+m52_30+m53_30+m54_30+m55_30+m56_30+m57_30+m58_30+m59_30+m60_30+m61_30+m62_30+m63_30+m64_30+m65_30+m66_30+m67_30+m68_30+m69_30+m70_30+m71_30+m72_30+m73_30+m74_30+m75_30+m76_30+m77_30+m78_30+m79_30+m80_30+m81_30+m82_30+m83_30+m84_30+m85_30+m86_30+m87_30+m88_30+m89_30+m90_30+m91_30+m92_30+m93_30+m94_30+m95_30+m96_30+m97_30+m98_30+m99_30+m100_30+m101_30+m102_30+m103_30+m104_30+m105_30+m106_30+m107_30+m108_30+m109_30+m110_30+m111_30+m112_30+m113_30+m114_30+m115_30+m116_30+m117_30+b30;
   always @(posedge clk) out31 <= m1_31+m2_31+m3_31+m4_31+m5_31+m6_31+m7_31+m8_31+m9_31+m10_31+m11_31+m12_31+m13_31+m14_31+m15_31+m16_31+m17_31+m18_31+m19_31+m20_31+m21_31+m22_31+m23_31+m24_31+m25_31+m26_31+m27_31+m28_31+m29_31+m30_31+m31_31+m32_31+m33_31+m34_31+m35_31+m36_31+m37_31+m38_31+m39_31+m40_31+m41_31+m42_31+m43_31+m44_31+m45_31+m46_31+m47_31+m48_31+m49_31+m50_31+m51_31+m52_31+m53_31+m54_31+m55_31+m56_31+m57_31+m58_31+m59_31+m60_31+m61_31+m62_31+m63_31+m64_31+m65_31+m66_31+m67_31+m68_31+m69_31+m70_31+m71_31+m72_31+m73_31+m74_31+m75_31+m76_31+m77_31+m78_31+m79_31+m80_31+m81_31+m82_31+m83_31+m84_31+m85_31+m86_31+m87_31+m88_31+m89_31+m90_31+m91_31+m92_31+m93_31+m94_31+m95_31+m96_31+m97_31+m98_31+m99_31+m100_31+m101_31+m102_31+m103_31+m104_31+m105_31+m106_31+m107_31+m108_31+m109_31+m110_31+m111_31+m112_31+m113_31+m114_31+m115_31+m116_31+m117_31+b31;
   always @(posedge clk) out32 <= m1_32+m2_32+m3_32+m4_32+m5_32+m6_32+m7_32+m8_32+m9_32+m10_32+m11_32+m12_32+m13_32+m14_32+m15_32+m16_32+m17_32+m18_32+m19_32+m20_32+m21_32+m22_32+m23_32+m24_32+m25_32+m26_32+m27_32+m28_32+m29_32+m30_32+m31_32+m32_32+m33_32+m34_32+m35_32+m36_32+m37_32+m38_32+m39_32+m40_32+m41_32+m42_32+m43_32+m44_32+m45_32+m46_32+m47_32+m48_32+m49_32+m50_32+m51_32+m52_32+m53_32+m54_32+m55_32+m56_32+m57_32+m58_32+m59_32+m60_32+m61_32+m62_32+m63_32+m64_32+m65_32+m66_32+m67_32+m68_32+m69_32+m70_32+m71_32+m72_32+m73_32+m74_32+m75_32+m76_32+m77_32+m78_32+m79_32+m80_32+m81_32+m82_32+m83_32+m84_32+m85_32+m86_32+m87_32+m88_32+m89_32+m90_32+m91_32+m92_32+m93_32+m94_32+m95_32+m96_32+m97_32+m98_32+m99_32+m100_32+m101_32+m102_32+m103_32+m104_32+m105_32+m106_32+m107_32+m108_32+m109_32+m110_32+m111_32+m112_32+m113_32+m114_32+m115_32+m116_32+m117_32+b32;
   always @(posedge clk) out33 <= m1_33+m2_33+m3_33+m4_33+m5_33+m6_33+m7_33+m8_33+m9_33+m10_33+m11_33+m12_33+m13_33+m14_33+m15_33+m16_33+m17_33+m18_33+m19_33+m20_33+m21_33+m22_33+m23_33+m24_33+m25_33+m26_33+m27_33+m28_33+m29_33+m30_33+m31_33+m32_33+m33_33+m34_33+m35_33+m36_33+m37_33+m38_33+m39_33+m40_33+m41_33+m42_33+m43_33+m44_33+m45_33+m46_33+m47_33+m48_33+m49_33+m50_33+m51_33+m52_33+m53_33+m54_33+m55_33+m56_33+m57_33+m58_33+m59_33+m60_33+m61_33+m62_33+m63_33+m64_33+m65_33+m66_33+m67_33+m68_33+m69_33+m70_33+m71_33+m72_33+m73_33+m74_33+m75_33+m76_33+m77_33+m78_33+m79_33+m80_33+m81_33+m82_33+m83_33+m84_33+m85_33+m86_33+m87_33+m88_33+m89_33+m90_33+m91_33+m92_33+m93_33+m94_33+m95_33+m96_33+m97_33+m98_33+m99_33+m100_33+m101_33+m102_33+m103_33+m104_33+m105_33+m106_33+m107_33+m108_33+m109_33+m110_33+m111_33+m112_33+m113_33+m114_33+m115_33+m116_33+m117_33+b33;
   always @(posedge clk) out34 <= m1_34+m2_34+m3_34+m4_34+m5_34+m6_34+m7_34+m8_34+m9_34+m10_34+m11_34+m12_34+m13_34+m14_34+m15_34+m16_34+m17_34+m18_34+m19_34+m20_34+m21_34+m22_34+m23_34+m24_34+m25_34+m26_34+m27_34+m28_34+m29_34+m30_34+m31_34+m32_34+m33_34+m34_34+m35_34+m36_34+m37_34+m38_34+m39_34+m40_34+m41_34+m42_34+m43_34+m44_34+m45_34+m46_34+m47_34+m48_34+m49_34+m50_34+m51_34+m52_34+m53_34+m54_34+m55_34+m56_34+m57_34+m58_34+m59_34+m60_34+m61_34+m62_34+m63_34+m64_34+m65_34+m66_34+m67_34+m68_34+m69_34+m70_34+m71_34+m72_34+m73_34+m74_34+m75_34+m76_34+m77_34+m78_34+m79_34+m80_34+m81_34+m82_34+m83_34+m84_34+m85_34+m86_34+m87_34+m88_34+m89_34+m90_34+m91_34+m92_34+m93_34+m94_34+m95_34+m96_34+m97_34+m98_34+m99_34+m100_34+m101_34+m102_34+m103_34+m104_34+m105_34+m106_34+m107_34+m108_34+m109_34+m110_34+m111_34+m112_34+m113_34+m114_34+m115_34+m116_34+m117_34+b34;
   always @(posedge clk) out35 <= m1_35+m2_35+m3_35+m4_35+m5_35+m6_35+m7_35+m8_35+m9_35+m10_35+m11_35+m12_35+m13_35+m14_35+m15_35+m16_35+m17_35+m18_35+m19_35+m20_35+m21_35+m22_35+m23_35+m24_35+m25_35+m26_35+m27_35+m28_35+m29_35+m30_35+m31_35+m32_35+m33_35+m34_35+m35_35+m36_35+m37_35+m38_35+m39_35+m40_35+m41_35+m42_35+m43_35+m44_35+m45_35+m46_35+m47_35+m48_35+m49_35+m50_35+m51_35+m52_35+m53_35+m54_35+m55_35+m56_35+m57_35+m58_35+m59_35+m60_35+m61_35+m62_35+m63_35+m64_35+m65_35+m66_35+m67_35+m68_35+m69_35+m70_35+m71_35+m72_35+m73_35+m74_35+m75_35+m76_35+m77_35+m78_35+m79_35+m80_35+m81_35+m82_35+m83_35+m84_35+m85_35+m86_35+m87_35+m88_35+m89_35+m90_35+m91_35+m92_35+m93_35+m94_35+m95_35+m96_35+m97_35+m98_35+m99_35+m100_35+m101_35+m102_35+m103_35+m104_35+m105_35+m106_35+m107_35+m108_35+m109_35+m110_35+m111_35+m112_35+m113_35+m114_35+m115_35+m116_35+m117_35+b35;
   always @(posedge clk) out36 <= m1_36+m2_36+m3_36+m4_36+m5_36+m6_36+m7_36+m8_36+m9_36+m10_36+m11_36+m12_36+m13_36+m14_36+m15_36+m16_36+m17_36+m18_36+m19_36+m20_36+m21_36+m22_36+m23_36+m24_36+m25_36+m26_36+m27_36+m28_36+m29_36+m30_36+m31_36+m32_36+m33_36+m34_36+m35_36+m36_36+m37_36+m38_36+m39_36+m40_36+m41_36+m42_36+m43_36+m44_36+m45_36+m46_36+m47_36+m48_36+m49_36+m50_36+m51_36+m52_36+m53_36+m54_36+m55_36+m56_36+m57_36+m58_36+m59_36+m60_36+m61_36+m62_36+m63_36+m64_36+m65_36+m66_36+m67_36+m68_36+m69_36+m70_36+m71_36+m72_36+m73_36+m74_36+m75_36+m76_36+m77_36+m78_36+m79_36+m80_36+m81_36+m82_36+m83_36+m84_36+m85_36+m86_36+m87_36+m88_36+m89_36+m90_36+m91_36+m92_36+m93_36+m94_36+m95_36+m96_36+m97_36+m98_36+m99_36+m100_36+m101_36+m102_36+m103_36+m104_36+m105_36+m106_36+m107_36+m108_36+m109_36+m110_36+m111_36+m112_36+m113_36+m114_36+m115_36+m116_36+m117_36+b36;
   always @(posedge clk) out37 <= m1_37+m2_37+m3_37+m4_37+m5_37+m6_37+m7_37+m8_37+m9_37+m10_37+m11_37+m12_37+m13_37+m14_37+m15_37+m16_37+m17_37+m18_37+m19_37+m20_37+m21_37+m22_37+m23_37+m24_37+m25_37+m26_37+m27_37+m28_37+m29_37+m30_37+m31_37+m32_37+m33_37+m34_37+m35_37+m36_37+m37_37+m38_37+m39_37+m40_37+m41_37+m42_37+m43_37+m44_37+m45_37+m46_37+m47_37+m48_37+m49_37+m50_37+m51_37+m52_37+m53_37+m54_37+m55_37+m56_37+m57_37+m58_37+m59_37+m60_37+m61_37+m62_37+m63_37+m64_37+m65_37+m66_37+m67_37+m68_37+m69_37+m70_37+m71_37+m72_37+m73_37+m74_37+m75_37+m76_37+m77_37+m78_37+m79_37+m80_37+m81_37+m82_37+m83_37+m84_37+m85_37+m86_37+m87_37+m88_37+m89_37+m90_37+m91_37+m92_37+m93_37+m94_37+m95_37+m96_37+m97_37+m98_37+m99_37+m100_37+m101_37+m102_37+m103_37+m104_37+m105_37+m106_37+m107_37+m108_37+m109_37+m110_37+m111_37+m112_37+m113_37+m114_37+m115_37+m116_37+m117_37+b37;
   always @(posedge clk) out38 <= m1_38+m2_38+m3_38+m4_38+m5_38+m6_38+m7_38+m8_38+m9_38+m10_38+m11_38+m12_38+m13_38+m14_38+m15_38+m16_38+m17_38+m18_38+m19_38+m20_38+m21_38+m22_38+m23_38+m24_38+m25_38+m26_38+m27_38+m28_38+m29_38+m30_38+m31_38+m32_38+m33_38+m34_38+m35_38+m36_38+m37_38+m38_38+m39_38+m40_38+m41_38+m42_38+m43_38+m44_38+m45_38+m46_38+m47_38+m48_38+m49_38+m50_38+m51_38+m52_38+m53_38+m54_38+m55_38+m56_38+m57_38+m58_38+m59_38+m60_38+m61_38+m62_38+m63_38+m64_38+m65_38+m66_38+m67_38+m68_38+m69_38+m70_38+m71_38+m72_38+m73_38+m74_38+m75_38+m76_38+m77_38+m78_38+m79_38+m80_38+m81_38+m82_38+m83_38+m84_38+m85_38+m86_38+m87_38+m88_38+m89_38+m90_38+m91_38+m92_38+m93_38+m94_38+m95_38+m96_38+m97_38+m98_38+m99_38+m100_38+m101_38+m102_38+m103_38+m104_38+m105_38+m106_38+m107_38+m108_38+m109_38+m110_38+m111_38+m112_38+m113_38+m114_38+m115_38+m116_38+m117_38+b38;
   always @(posedge clk) out39 <= m1_39+m2_39+m3_39+m4_39+m5_39+m6_39+m7_39+m8_39+m9_39+m10_39+m11_39+m12_39+m13_39+m14_39+m15_39+m16_39+m17_39+m18_39+m19_39+m20_39+m21_39+m22_39+m23_39+m24_39+m25_39+m26_39+m27_39+m28_39+m29_39+m30_39+m31_39+m32_39+m33_39+m34_39+m35_39+m36_39+m37_39+m38_39+m39_39+m40_39+m41_39+m42_39+m43_39+m44_39+m45_39+m46_39+m47_39+m48_39+m49_39+m50_39+m51_39+m52_39+m53_39+m54_39+m55_39+m56_39+m57_39+m58_39+m59_39+m60_39+m61_39+m62_39+m63_39+m64_39+m65_39+m66_39+m67_39+m68_39+m69_39+m70_39+m71_39+m72_39+m73_39+m74_39+m75_39+m76_39+m77_39+m78_39+m79_39+m80_39+m81_39+m82_39+m83_39+m84_39+m85_39+m86_39+m87_39+m88_39+m89_39+m90_39+m91_39+m92_39+m93_39+m94_39+m95_39+m96_39+m97_39+m98_39+m99_39+m100_39+m101_39+m102_39+m103_39+m104_39+m105_39+m106_39+m107_39+m108_39+m109_39+m110_39+m111_39+m112_39+m113_39+m114_39+m115_39+m116_39+m117_39+b39;
   always @(posedge clk) out40 <= m1_40+m2_40+m3_40+m4_40+m5_40+m6_40+m7_40+m8_40+m9_40+m10_40+m11_40+m12_40+m13_40+m14_40+m15_40+m16_40+m17_40+m18_40+m19_40+m20_40+m21_40+m22_40+m23_40+m24_40+m25_40+m26_40+m27_40+m28_40+m29_40+m30_40+m31_40+m32_40+m33_40+m34_40+m35_40+m36_40+m37_40+m38_40+m39_40+m40_40+m41_40+m42_40+m43_40+m44_40+m45_40+m46_40+m47_40+m48_40+m49_40+m50_40+m51_40+m52_40+m53_40+m54_40+m55_40+m56_40+m57_40+m58_40+m59_40+m60_40+m61_40+m62_40+m63_40+m64_40+m65_40+m66_40+m67_40+m68_40+m69_40+m70_40+m71_40+m72_40+m73_40+m74_40+m75_40+m76_40+m77_40+m78_40+m79_40+m80_40+m81_40+m82_40+m83_40+m84_40+m85_40+m86_40+m87_40+m88_40+m89_40+m90_40+m91_40+m92_40+m93_40+m94_40+m95_40+m96_40+m97_40+m98_40+m99_40+m100_40+m101_40+m102_40+m103_40+m104_40+m105_40+m106_40+m107_40+m108_40+m109_40+m110_40+m111_40+m112_40+m113_40+m114_40+m115_40+m116_40+m117_40+b40;
   always @(posedge clk) out41 <= m1_41+m2_41+m3_41+m4_41+m5_41+m6_41+m7_41+m8_41+m9_41+m10_41+m11_41+m12_41+m13_41+m14_41+m15_41+m16_41+m17_41+m18_41+m19_41+m20_41+m21_41+m22_41+m23_41+m24_41+m25_41+m26_41+m27_41+m28_41+m29_41+m30_41+m31_41+m32_41+m33_41+m34_41+m35_41+m36_41+m37_41+m38_41+m39_41+m40_41+m41_41+m42_41+m43_41+m44_41+m45_41+m46_41+m47_41+m48_41+m49_41+m50_41+m51_41+m52_41+m53_41+m54_41+m55_41+m56_41+m57_41+m58_41+m59_41+m60_41+m61_41+m62_41+m63_41+m64_41+m65_41+m66_41+m67_41+m68_41+m69_41+m70_41+m71_41+m72_41+m73_41+m74_41+m75_41+m76_41+m77_41+m78_41+m79_41+m80_41+m81_41+m82_41+m83_41+m84_41+m85_41+m86_41+m87_41+m88_41+m89_41+m90_41+m91_41+m92_41+m93_41+m94_41+m95_41+m96_41+m97_41+m98_41+m99_41+m100_41+m101_41+m102_41+m103_41+m104_41+m105_41+m106_41+m107_41+m108_41+m109_41+m110_41+m111_41+m112_41+m113_41+m114_41+m115_41+m116_41+m117_41+b41;
   always @(posedge clk) out42 <= m1_42+m2_42+m3_42+m4_42+m5_42+m6_42+m7_42+m8_42+m9_42+m10_42+m11_42+m12_42+m13_42+m14_42+m15_42+m16_42+m17_42+m18_42+m19_42+m20_42+m21_42+m22_42+m23_42+m24_42+m25_42+m26_42+m27_42+m28_42+m29_42+m30_42+m31_42+m32_42+m33_42+m34_42+m35_42+m36_42+m37_42+m38_42+m39_42+m40_42+m41_42+m42_42+m43_42+m44_42+m45_42+m46_42+m47_42+m48_42+m49_42+m50_42+m51_42+m52_42+m53_42+m54_42+m55_42+m56_42+m57_42+m58_42+m59_42+m60_42+m61_42+m62_42+m63_42+m64_42+m65_42+m66_42+m67_42+m68_42+m69_42+m70_42+m71_42+m72_42+m73_42+m74_42+m75_42+m76_42+m77_42+m78_42+m79_42+m80_42+m81_42+m82_42+m83_42+m84_42+m85_42+m86_42+m87_42+m88_42+m89_42+m90_42+m91_42+m92_42+m93_42+m94_42+m95_42+m96_42+m97_42+m98_42+m99_42+m100_42+m101_42+m102_42+m103_42+m104_42+m105_42+m106_42+m107_42+m108_42+m109_42+m110_42+m111_42+m112_42+m113_42+m114_42+m115_42+m116_42+m117_42+b42;
   always @(posedge clk) out43 <= m1_43+m2_43+m3_43+m4_43+m5_43+m6_43+m7_43+m8_43+m9_43+m10_43+m11_43+m12_43+m13_43+m14_43+m15_43+m16_43+m17_43+m18_43+m19_43+m20_43+m21_43+m22_43+m23_43+m24_43+m25_43+m26_43+m27_43+m28_43+m29_43+m30_43+m31_43+m32_43+m33_43+m34_43+m35_43+m36_43+m37_43+m38_43+m39_43+m40_43+m41_43+m42_43+m43_43+m44_43+m45_43+m46_43+m47_43+m48_43+m49_43+m50_43+m51_43+m52_43+m53_43+m54_43+m55_43+m56_43+m57_43+m58_43+m59_43+m60_43+m61_43+m62_43+m63_43+m64_43+m65_43+m66_43+m67_43+m68_43+m69_43+m70_43+m71_43+m72_43+m73_43+m74_43+m75_43+m76_43+m77_43+m78_43+m79_43+m80_43+m81_43+m82_43+m83_43+m84_43+m85_43+m86_43+m87_43+m88_43+m89_43+m90_43+m91_43+m92_43+m93_43+m94_43+m95_43+m96_43+m97_43+m98_43+m99_43+m100_43+m101_43+m102_43+m103_43+m104_43+m105_43+m106_43+m107_43+m108_43+m109_43+m110_43+m111_43+m112_43+m113_43+m114_43+m115_43+m116_43+m117_43+b43;
   always @(posedge clk) out44 <= m1_44+m2_44+m3_44+m4_44+m5_44+m6_44+m7_44+m8_44+m9_44+m10_44+m11_44+m12_44+m13_44+m14_44+m15_44+m16_44+m17_44+m18_44+m19_44+m20_44+m21_44+m22_44+m23_44+m24_44+m25_44+m26_44+m27_44+m28_44+m29_44+m30_44+m31_44+m32_44+m33_44+m34_44+m35_44+m36_44+m37_44+m38_44+m39_44+m40_44+m41_44+m42_44+m43_44+m44_44+m45_44+m46_44+m47_44+m48_44+m49_44+m50_44+m51_44+m52_44+m53_44+m54_44+m55_44+m56_44+m57_44+m58_44+m59_44+m60_44+m61_44+m62_44+m63_44+m64_44+m65_44+m66_44+m67_44+m68_44+m69_44+m70_44+m71_44+m72_44+m73_44+m74_44+m75_44+m76_44+m77_44+m78_44+m79_44+m80_44+m81_44+m82_44+m83_44+m84_44+m85_44+m86_44+m87_44+m88_44+m89_44+m90_44+m91_44+m92_44+m93_44+m94_44+m95_44+m96_44+m97_44+m98_44+m99_44+m100_44+m101_44+m102_44+m103_44+m104_44+m105_44+m106_44+m107_44+m108_44+m109_44+m110_44+m111_44+m112_44+m113_44+m114_44+m115_44+m116_44+m117_44+b44;
   always @(posedge clk) out45 <= m1_45+m2_45+m3_45+m4_45+m5_45+m6_45+m7_45+m8_45+m9_45+m10_45+m11_45+m12_45+m13_45+m14_45+m15_45+m16_45+m17_45+m18_45+m19_45+m20_45+m21_45+m22_45+m23_45+m24_45+m25_45+m26_45+m27_45+m28_45+m29_45+m30_45+m31_45+m32_45+m33_45+m34_45+m35_45+m36_45+m37_45+m38_45+m39_45+m40_45+m41_45+m42_45+m43_45+m44_45+m45_45+m46_45+m47_45+m48_45+m49_45+m50_45+m51_45+m52_45+m53_45+m54_45+m55_45+m56_45+m57_45+m58_45+m59_45+m60_45+m61_45+m62_45+m63_45+m64_45+m65_45+m66_45+m67_45+m68_45+m69_45+m70_45+m71_45+m72_45+m73_45+m74_45+m75_45+m76_45+m77_45+m78_45+m79_45+m80_45+m81_45+m82_45+m83_45+m84_45+m85_45+m86_45+m87_45+m88_45+m89_45+m90_45+m91_45+m92_45+m93_45+m94_45+m95_45+m96_45+m97_45+m98_45+m99_45+m100_45+m101_45+m102_45+m103_45+m104_45+m105_45+m106_45+m107_45+m108_45+m109_45+m110_45+m111_45+m112_45+m113_45+m114_45+m115_45+m116_45+m117_45+b45;
   always @(posedge clk) out46 <= m1_46+m2_46+m3_46+m4_46+m5_46+m6_46+m7_46+m8_46+m9_46+m10_46+m11_46+m12_46+m13_46+m14_46+m15_46+m16_46+m17_46+m18_46+m19_46+m20_46+m21_46+m22_46+m23_46+m24_46+m25_46+m26_46+m27_46+m28_46+m29_46+m30_46+m31_46+m32_46+m33_46+m34_46+m35_46+m36_46+m37_46+m38_46+m39_46+m40_46+m41_46+m42_46+m43_46+m44_46+m45_46+m46_46+m47_46+m48_46+m49_46+m50_46+m51_46+m52_46+m53_46+m54_46+m55_46+m56_46+m57_46+m58_46+m59_46+m60_46+m61_46+m62_46+m63_46+m64_46+m65_46+m66_46+m67_46+m68_46+m69_46+m70_46+m71_46+m72_46+m73_46+m74_46+m75_46+m76_46+m77_46+m78_46+m79_46+m80_46+m81_46+m82_46+m83_46+m84_46+m85_46+m86_46+m87_46+m88_46+m89_46+m90_46+m91_46+m92_46+m93_46+m94_46+m95_46+m96_46+m97_46+m98_46+m99_46+m100_46+m101_46+m102_46+m103_46+m104_46+m105_46+m106_46+m107_46+m108_46+m109_46+m110_46+m111_46+m112_46+m113_46+m114_46+m115_46+m116_46+m117_46+b46;
   always @(posedge clk) out47 <= m1_47+m2_47+m3_47+m4_47+m5_47+m6_47+m7_47+m8_47+m9_47+m10_47+m11_47+m12_47+m13_47+m14_47+m15_47+m16_47+m17_47+m18_47+m19_47+m20_47+m21_47+m22_47+m23_47+m24_47+m25_47+m26_47+m27_47+m28_47+m29_47+m30_47+m31_47+m32_47+m33_47+m34_47+m35_47+m36_47+m37_47+m38_47+m39_47+m40_47+m41_47+m42_47+m43_47+m44_47+m45_47+m46_47+m47_47+m48_47+m49_47+m50_47+m51_47+m52_47+m53_47+m54_47+m55_47+m56_47+m57_47+m58_47+m59_47+m60_47+m61_47+m62_47+m63_47+m64_47+m65_47+m66_47+m67_47+m68_47+m69_47+m70_47+m71_47+m72_47+m73_47+m74_47+m75_47+m76_47+m77_47+m78_47+m79_47+m80_47+m81_47+m82_47+m83_47+m84_47+m85_47+m86_47+m87_47+m88_47+m89_47+m90_47+m91_47+m92_47+m93_47+m94_47+m95_47+m96_47+m97_47+m98_47+m99_47+m100_47+m101_47+m102_47+m103_47+m104_47+m105_47+m106_47+m107_47+m108_47+m109_47+m110_47+m111_47+m112_47+m113_47+m114_47+m115_47+m116_47+m117_47+b47;
   always @(posedge clk) out48 <= m1_48+m2_48+m3_48+m4_48+m5_48+m6_48+m7_48+m8_48+m9_48+m10_48+m11_48+m12_48+m13_48+m14_48+m15_48+m16_48+m17_48+m18_48+m19_48+m20_48+m21_48+m22_48+m23_48+m24_48+m25_48+m26_48+m27_48+m28_48+m29_48+m30_48+m31_48+m32_48+m33_48+m34_48+m35_48+m36_48+m37_48+m38_48+m39_48+m40_48+m41_48+m42_48+m43_48+m44_48+m45_48+m46_48+m47_48+m48_48+m49_48+m50_48+m51_48+m52_48+m53_48+m54_48+m55_48+m56_48+m57_48+m58_48+m59_48+m60_48+m61_48+m62_48+m63_48+m64_48+m65_48+m66_48+m67_48+m68_48+m69_48+m70_48+m71_48+m72_48+m73_48+m74_48+m75_48+m76_48+m77_48+m78_48+m79_48+m80_48+m81_48+m82_48+m83_48+m84_48+m85_48+m86_48+m87_48+m88_48+m89_48+m90_48+m91_48+m92_48+m93_48+m94_48+m95_48+m96_48+m97_48+m98_48+m99_48+m100_48+m101_48+m102_48+m103_48+m104_48+m105_48+m106_48+m107_48+m108_48+m109_48+m110_48+m111_48+m112_48+m113_48+m114_48+m115_48+m116_48+m117_48+b48;
   always @(posedge clk) out49 <= m1_49+m2_49+m3_49+m4_49+m5_49+m6_49+m7_49+m8_49+m9_49+m10_49+m11_49+m12_49+m13_49+m14_49+m15_49+m16_49+m17_49+m18_49+m19_49+m20_49+m21_49+m22_49+m23_49+m24_49+m25_49+m26_49+m27_49+m28_49+m29_49+m30_49+m31_49+m32_49+m33_49+m34_49+m35_49+m36_49+m37_49+m38_49+m39_49+m40_49+m41_49+m42_49+m43_49+m44_49+m45_49+m46_49+m47_49+m48_49+m49_49+m50_49+m51_49+m52_49+m53_49+m54_49+m55_49+m56_49+m57_49+m58_49+m59_49+m60_49+m61_49+m62_49+m63_49+m64_49+m65_49+m66_49+m67_49+m68_49+m69_49+m70_49+m71_49+m72_49+m73_49+m74_49+m75_49+m76_49+m77_49+m78_49+m79_49+m80_49+m81_49+m82_49+m83_49+m84_49+m85_49+m86_49+m87_49+m88_49+m89_49+m90_49+m91_49+m92_49+m93_49+m94_49+m95_49+m96_49+m97_49+m98_49+m99_49+m100_49+m101_49+m102_49+m103_49+m104_49+m105_49+m106_49+m107_49+m108_49+m109_49+m110_49+m111_49+m112_49+m113_49+m114_49+m115_49+m116_49+m117_49+b49;
   always @(posedge clk) out50 <= m1_50+m2_50+m3_50+m4_50+m5_50+m6_50+m7_50+m8_50+m9_50+m10_50+m11_50+m12_50+m13_50+m14_50+m15_50+m16_50+m17_50+m18_50+m19_50+m20_50+m21_50+m22_50+m23_50+m24_50+m25_50+m26_50+m27_50+m28_50+m29_50+m30_50+m31_50+m32_50+m33_50+m34_50+m35_50+m36_50+m37_50+m38_50+m39_50+m40_50+m41_50+m42_50+m43_50+m44_50+m45_50+m46_50+m47_50+m48_50+m49_50+m50_50+m51_50+m52_50+m53_50+m54_50+m55_50+m56_50+m57_50+m58_50+m59_50+m60_50+m61_50+m62_50+m63_50+m64_50+m65_50+m66_50+m67_50+m68_50+m69_50+m70_50+m71_50+m72_50+m73_50+m74_50+m75_50+m76_50+m77_50+m78_50+m79_50+m80_50+m81_50+m82_50+m83_50+m84_50+m85_50+m86_50+m87_50+m88_50+m89_50+m90_50+m91_50+m92_50+m93_50+m94_50+m95_50+m96_50+m97_50+m98_50+m99_50+m100_50+m101_50+m102_50+m103_50+m104_50+m105_50+m106_50+m107_50+m108_50+m109_50+m110_50+m111_50+m112_50+m113_50+m114_50+m115_50+m116_50+m117_50+b50;
   always @(posedge clk) out51 <= m1_51+m2_51+m3_51+m4_51+m5_51+m6_51+m7_51+m8_51+m9_51+m10_51+m11_51+m12_51+m13_51+m14_51+m15_51+m16_51+m17_51+m18_51+m19_51+m20_51+m21_51+m22_51+m23_51+m24_51+m25_51+m26_51+m27_51+m28_51+m29_51+m30_51+m31_51+m32_51+m33_51+m34_51+m35_51+m36_51+m37_51+m38_51+m39_51+m40_51+m41_51+m42_51+m43_51+m44_51+m45_51+m46_51+m47_51+m48_51+m49_51+m50_51+m51_51+m52_51+m53_51+m54_51+m55_51+m56_51+m57_51+m58_51+m59_51+m60_51+m61_51+m62_51+m63_51+m64_51+m65_51+m66_51+m67_51+m68_51+m69_51+m70_51+m71_51+m72_51+m73_51+m74_51+m75_51+m76_51+m77_51+m78_51+m79_51+m80_51+m81_51+m82_51+m83_51+m84_51+m85_51+m86_51+m87_51+m88_51+m89_51+m90_51+m91_51+m92_51+m93_51+m94_51+m95_51+m96_51+m97_51+m98_51+m99_51+m100_51+m101_51+m102_51+m103_51+m104_51+m105_51+m106_51+m107_51+m108_51+m109_51+m110_51+m111_51+m112_51+m113_51+m114_51+m115_51+m116_51+m117_51+b51;
   always @(posedge clk) out52 <= m1_52+m2_52+m3_52+m4_52+m5_52+m6_52+m7_52+m8_52+m9_52+m10_52+m11_52+m12_52+m13_52+m14_52+m15_52+m16_52+m17_52+m18_52+m19_52+m20_52+m21_52+m22_52+m23_52+m24_52+m25_52+m26_52+m27_52+m28_52+m29_52+m30_52+m31_52+m32_52+m33_52+m34_52+m35_52+m36_52+m37_52+m38_52+m39_52+m40_52+m41_52+m42_52+m43_52+m44_52+m45_52+m46_52+m47_52+m48_52+m49_52+m50_52+m51_52+m52_52+m53_52+m54_52+m55_52+m56_52+m57_52+m58_52+m59_52+m60_52+m61_52+m62_52+m63_52+m64_52+m65_52+m66_52+m67_52+m68_52+m69_52+m70_52+m71_52+m72_52+m73_52+m74_52+m75_52+m76_52+m77_52+m78_52+m79_52+m80_52+m81_52+m82_52+m83_52+m84_52+m85_52+m86_52+m87_52+m88_52+m89_52+m90_52+m91_52+m92_52+m93_52+m94_52+m95_52+m96_52+m97_52+m98_52+m99_52+m100_52+m101_52+m102_52+m103_52+m104_52+m105_52+m106_52+m107_52+m108_52+m109_52+m110_52+m111_52+m112_52+m113_52+m114_52+m115_52+m116_52+m117_52+b52;
   always @(posedge clk) out53 <= m1_53+m2_53+m3_53+m4_53+m5_53+m6_53+m7_53+m8_53+m9_53+m10_53+m11_53+m12_53+m13_53+m14_53+m15_53+m16_53+m17_53+m18_53+m19_53+m20_53+m21_53+m22_53+m23_53+m24_53+m25_53+m26_53+m27_53+m28_53+m29_53+m30_53+m31_53+m32_53+m33_53+m34_53+m35_53+m36_53+m37_53+m38_53+m39_53+m40_53+m41_53+m42_53+m43_53+m44_53+m45_53+m46_53+m47_53+m48_53+m49_53+m50_53+m51_53+m52_53+m53_53+m54_53+m55_53+m56_53+m57_53+m58_53+m59_53+m60_53+m61_53+m62_53+m63_53+m64_53+m65_53+m66_53+m67_53+m68_53+m69_53+m70_53+m71_53+m72_53+m73_53+m74_53+m75_53+m76_53+m77_53+m78_53+m79_53+m80_53+m81_53+m82_53+m83_53+m84_53+m85_53+m86_53+m87_53+m88_53+m89_53+m90_53+m91_53+m92_53+m93_53+m94_53+m95_53+m96_53+m97_53+m98_53+m99_53+m100_53+m101_53+m102_53+m103_53+m104_53+m105_53+m106_53+m107_53+m108_53+m109_53+m110_53+m111_53+m112_53+m113_53+m114_53+m115_53+m116_53+m117_53+b53;
   always @(posedge clk) out54 <= m1_54+m2_54+m3_54+m4_54+m5_54+m6_54+m7_54+m8_54+m9_54+m10_54+m11_54+m12_54+m13_54+m14_54+m15_54+m16_54+m17_54+m18_54+m19_54+m20_54+m21_54+m22_54+m23_54+m24_54+m25_54+m26_54+m27_54+m28_54+m29_54+m30_54+m31_54+m32_54+m33_54+m34_54+m35_54+m36_54+m37_54+m38_54+m39_54+m40_54+m41_54+m42_54+m43_54+m44_54+m45_54+m46_54+m47_54+m48_54+m49_54+m50_54+m51_54+m52_54+m53_54+m54_54+m55_54+m56_54+m57_54+m58_54+m59_54+m60_54+m61_54+m62_54+m63_54+m64_54+m65_54+m66_54+m67_54+m68_54+m69_54+m70_54+m71_54+m72_54+m73_54+m74_54+m75_54+m76_54+m77_54+m78_54+m79_54+m80_54+m81_54+m82_54+m83_54+m84_54+m85_54+m86_54+m87_54+m88_54+m89_54+m90_54+m91_54+m92_54+m93_54+m94_54+m95_54+m96_54+m97_54+m98_54+m99_54+m100_54+m101_54+m102_54+m103_54+m104_54+m105_54+m106_54+m107_54+m108_54+m109_54+m110_54+m111_54+m112_54+m113_54+m114_54+m115_54+m116_54+m117_54+b54;
   always @(posedge clk) out55 <= m1_55+m2_55+m3_55+m4_55+m5_55+m6_55+m7_55+m8_55+m9_55+m10_55+m11_55+m12_55+m13_55+m14_55+m15_55+m16_55+m17_55+m18_55+m19_55+m20_55+m21_55+m22_55+m23_55+m24_55+m25_55+m26_55+m27_55+m28_55+m29_55+m30_55+m31_55+m32_55+m33_55+m34_55+m35_55+m36_55+m37_55+m38_55+m39_55+m40_55+m41_55+m42_55+m43_55+m44_55+m45_55+m46_55+m47_55+m48_55+m49_55+m50_55+m51_55+m52_55+m53_55+m54_55+m55_55+m56_55+m57_55+m58_55+m59_55+m60_55+m61_55+m62_55+m63_55+m64_55+m65_55+m66_55+m67_55+m68_55+m69_55+m70_55+m71_55+m72_55+m73_55+m74_55+m75_55+m76_55+m77_55+m78_55+m79_55+m80_55+m81_55+m82_55+m83_55+m84_55+m85_55+m86_55+m87_55+m88_55+m89_55+m90_55+m91_55+m92_55+m93_55+m94_55+m95_55+m96_55+m97_55+m98_55+m99_55+m100_55+m101_55+m102_55+m103_55+m104_55+m105_55+m106_55+m107_55+m108_55+m109_55+m110_55+m111_55+m112_55+m113_55+m114_55+m115_55+m116_55+m117_55+b55;
   always @(posedge clk) out56 <= m1_56+m2_56+m3_56+m4_56+m5_56+m6_56+m7_56+m8_56+m9_56+m10_56+m11_56+m12_56+m13_56+m14_56+m15_56+m16_56+m17_56+m18_56+m19_56+m20_56+m21_56+m22_56+m23_56+m24_56+m25_56+m26_56+m27_56+m28_56+m29_56+m30_56+m31_56+m32_56+m33_56+m34_56+m35_56+m36_56+m37_56+m38_56+m39_56+m40_56+m41_56+m42_56+m43_56+m44_56+m45_56+m46_56+m47_56+m48_56+m49_56+m50_56+m51_56+m52_56+m53_56+m54_56+m55_56+m56_56+m57_56+m58_56+m59_56+m60_56+m61_56+m62_56+m63_56+m64_56+m65_56+m66_56+m67_56+m68_56+m69_56+m70_56+m71_56+m72_56+m73_56+m74_56+m75_56+m76_56+m77_56+m78_56+m79_56+m80_56+m81_56+m82_56+m83_56+m84_56+m85_56+m86_56+m87_56+m88_56+m89_56+m90_56+m91_56+m92_56+m93_56+m94_56+m95_56+m96_56+m97_56+m98_56+m99_56+m100_56+m101_56+m102_56+m103_56+m104_56+m105_56+m106_56+m107_56+m108_56+m109_56+m110_56+m111_56+m112_56+m113_56+m114_56+m115_56+m116_56+m117_56+b56;
   always @(posedge clk) out57 <= m1_57+m2_57+m3_57+m4_57+m5_57+m6_57+m7_57+m8_57+m9_57+m10_57+m11_57+m12_57+m13_57+m14_57+m15_57+m16_57+m17_57+m18_57+m19_57+m20_57+m21_57+m22_57+m23_57+m24_57+m25_57+m26_57+m27_57+m28_57+m29_57+m30_57+m31_57+m32_57+m33_57+m34_57+m35_57+m36_57+m37_57+m38_57+m39_57+m40_57+m41_57+m42_57+m43_57+m44_57+m45_57+m46_57+m47_57+m48_57+m49_57+m50_57+m51_57+m52_57+m53_57+m54_57+m55_57+m56_57+m57_57+m58_57+m59_57+m60_57+m61_57+m62_57+m63_57+m64_57+m65_57+m66_57+m67_57+m68_57+m69_57+m70_57+m71_57+m72_57+m73_57+m74_57+m75_57+m76_57+m77_57+m78_57+m79_57+m80_57+m81_57+m82_57+m83_57+m84_57+m85_57+m86_57+m87_57+m88_57+m89_57+m90_57+m91_57+m92_57+m93_57+m94_57+m95_57+m96_57+m97_57+m98_57+m99_57+m100_57+m101_57+m102_57+m103_57+m104_57+m105_57+m106_57+m107_57+m108_57+m109_57+m110_57+m111_57+m112_57+m113_57+m114_57+m115_57+m116_57+m117_57+b57;
   always @(posedge clk) out58 <= m1_58+m2_58+m3_58+m4_58+m5_58+m6_58+m7_58+m8_58+m9_58+m10_58+m11_58+m12_58+m13_58+m14_58+m15_58+m16_58+m17_58+m18_58+m19_58+m20_58+m21_58+m22_58+m23_58+m24_58+m25_58+m26_58+m27_58+m28_58+m29_58+m30_58+m31_58+m32_58+m33_58+m34_58+m35_58+m36_58+m37_58+m38_58+m39_58+m40_58+m41_58+m42_58+m43_58+m44_58+m45_58+m46_58+m47_58+m48_58+m49_58+m50_58+m51_58+m52_58+m53_58+m54_58+m55_58+m56_58+m57_58+m58_58+m59_58+m60_58+m61_58+m62_58+m63_58+m64_58+m65_58+m66_58+m67_58+m68_58+m69_58+m70_58+m71_58+m72_58+m73_58+m74_58+m75_58+m76_58+m77_58+m78_58+m79_58+m80_58+m81_58+m82_58+m83_58+m84_58+m85_58+m86_58+m87_58+m88_58+m89_58+m90_58+m91_58+m92_58+m93_58+m94_58+m95_58+m96_58+m97_58+m98_58+m99_58+m100_58+m101_58+m102_58+m103_58+m104_58+m105_58+m106_58+m107_58+m108_58+m109_58+m110_58+m111_58+m112_58+m113_58+m114_58+m115_58+m116_58+m117_58+b58;
   always @(posedge clk) out59 <= m1_59+m2_59+m3_59+m4_59+m5_59+m6_59+m7_59+m8_59+m9_59+m10_59+m11_59+m12_59+m13_59+m14_59+m15_59+m16_59+m17_59+m18_59+m19_59+m20_59+m21_59+m22_59+m23_59+m24_59+m25_59+m26_59+m27_59+m28_59+m29_59+m30_59+m31_59+m32_59+m33_59+m34_59+m35_59+m36_59+m37_59+m38_59+m39_59+m40_59+m41_59+m42_59+m43_59+m44_59+m45_59+m46_59+m47_59+m48_59+m49_59+m50_59+m51_59+m52_59+m53_59+m54_59+m55_59+m56_59+m57_59+m58_59+m59_59+m60_59+m61_59+m62_59+m63_59+m64_59+m65_59+m66_59+m67_59+m68_59+m69_59+m70_59+m71_59+m72_59+m73_59+m74_59+m75_59+m76_59+m77_59+m78_59+m79_59+m80_59+m81_59+m82_59+m83_59+m84_59+m85_59+m86_59+m87_59+m88_59+m89_59+m90_59+m91_59+m92_59+m93_59+m94_59+m95_59+m96_59+m97_59+m98_59+m99_59+m100_59+m101_59+m102_59+m103_59+m104_59+m105_59+m106_59+m107_59+m108_59+m109_59+m110_59+m111_59+m112_59+m113_59+m114_59+m115_59+m116_59+m117_59+b59;
   always @(posedge clk) out60 <= m1_60+m2_60+m3_60+m4_60+m5_60+m6_60+m7_60+m8_60+m9_60+m10_60+m11_60+m12_60+m13_60+m14_60+m15_60+m16_60+m17_60+m18_60+m19_60+m20_60+m21_60+m22_60+m23_60+m24_60+m25_60+m26_60+m27_60+m28_60+m29_60+m30_60+m31_60+m32_60+m33_60+m34_60+m35_60+m36_60+m37_60+m38_60+m39_60+m40_60+m41_60+m42_60+m43_60+m44_60+m45_60+m46_60+m47_60+m48_60+m49_60+m50_60+m51_60+m52_60+m53_60+m54_60+m55_60+m56_60+m57_60+m58_60+m59_60+m60_60+m61_60+m62_60+m63_60+m64_60+m65_60+m66_60+m67_60+m68_60+m69_60+m70_60+m71_60+m72_60+m73_60+m74_60+m75_60+m76_60+m77_60+m78_60+m79_60+m80_60+m81_60+m82_60+m83_60+m84_60+m85_60+m86_60+m87_60+m88_60+m89_60+m90_60+m91_60+m92_60+m93_60+m94_60+m95_60+m96_60+m97_60+m98_60+m99_60+m100_60+m101_60+m102_60+m103_60+m104_60+m105_60+m106_60+m107_60+m108_60+m109_60+m110_60+m111_60+m112_60+m113_60+m114_60+m115_60+m116_60+m117_60+b60;
   always @(posedge clk) out61 <= m1_61+m2_61+m3_61+m4_61+m5_61+m6_61+m7_61+m8_61+m9_61+m10_61+m11_61+m12_61+m13_61+m14_61+m15_61+m16_61+m17_61+m18_61+m19_61+m20_61+m21_61+m22_61+m23_61+m24_61+m25_61+m26_61+m27_61+m28_61+m29_61+m30_61+m31_61+m32_61+m33_61+m34_61+m35_61+m36_61+m37_61+m38_61+m39_61+m40_61+m41_61+m42_61+m43_61+m44_61+m45_61+m46_61+m47_61+m48_61+m49_61+m50_61+m51_61+m52_61+m53_61+m54_61+m55_61+m56_61+m57_61+m58_61+m59_61+m60_61+m61_61+m62_61+m63_61+m64_61+m65_61+m66_61+m67_61+m68_61+m69_61+m70_61+m71_61+m72_61+m73_61+m74_61+m75_61+m76_61+m77_61+m78_61+m79_61+m80_61+m81_61+m82_61+m83_61+m84_61+m85_61+m86_61+m87_61+m88_61+m89_61+m90_61+m91_61+m92_61+m93_61+m94_61+m95_61+m96_61+m97_61+m98_61+m99_61+m100_61+m101_61+m102_61+m103_61+m104_61+m105_61+m106_61+m107_61+m108_61+m109_61+m110_61+m111_61+m112_61+m113_61+m114_61+m115_61+m116_61+m117_61+b61;
   always @(posedge clk) out62 <= m1_62+m2_62+m3_62+m4_62+m5_62+m6_62+m7_62+m8_62+m9_62+m10_62+m11_62+m12_62+m13_62+m14_62+m15_62+m16_62+m17_62+m18_62+m19_62+m20_62+m21_62+m22_62+m23_62+m24_62+m25_62+m26_62+m27_62+m28_62+m29_62+m30_62+m31_62+m32_62+m33_62+m34_62+m35_62+m36_62+m37_62+m38_62+m39_62+m40_62+m41_62+m42_62+m43_62+m44_62+m45_62+m46_62+m47_62+m48_62+m49_62+m50_62+m51_62+m52_62+m53_62+m54_62+m55_62+m56_62+m57_62+m58_62+m59_62+m60_62+m61_62+m62_62+m63_62+m64_62+m65_62+m66_62+m67_62+m68_62+m69_62+m70_62+m71_62+m72_62+m73_62+m74_62+m75_62+m76_62+m77_62+m78_62+m79_62+m80_62+m81_62+m82_62+m83_62+m84_62+m85_62+m86_62+m87_62+m88_62+m89_62+m90_62+m91_62+m92_62+m93_62+m94_62+m95_62+m96_62+m97_62+m98_62+m99_62+m100_62+m101_62+m102_62+m103_62+m104_62+m105_62+m106_62+m107_62+m108_62+m109_62+m110_62+m111_62+m112_62+m113_62+m114_62+m115_62+m116_62+m117_62+b62;
   always @(posedge clk) out63 <= m1_63+m2_63+m3_63+m4_63+m5_63+m6_63+m7_63+m8_63+m9_63+m10_63+m11_63+m12_63+m13_63+m14_63+m15_63+m16_63+m17_63+m18_63+m19_63+m20_63+m21_63+m22_63+m23_63+m24_63+m25_63+m26_63+m27_63+m28_63+m29_63+m30_63+m31_63+m32_63+m33_63+m34_63+m35_63+m36_63+m37_63+m38_63+m39_63+m40_63+m41_63+m42_63+m43_63+m44_63+m45_63+m46_63+m47_63+m48_63+m49_63+m50_63+m51_63+m52_63+m53_63+m54_63+m55_63+m56_63+m57_63+m58_63+m59_63+m60_63+m61_63+m62_63+m63_63+m64_63+m65_63+m66_63+m67_63+m68_63+m69_63+m70_63+m71_63+m72_63+m73_63+m74_63+m75_63+m76_63+m77_63+m78_63+m79_63+m80_63+m81_63+m82_63+m83_63+m84_63+m85_63+m86_63+m87_63+m88_63+m89_63+m90_63+m91_63+m92_63+m93_63+m94_63+m95_63+m96_63+m97_63+m98_63+m99_63+m100_63+m101_63+m102_63+m103_63+m104_63+m105_63+m106_63+m107_63+m108_63+m109_63+m110_63+m111_63+m112_63+m113_63+m114_63+m115_63+m116_63+m117_63+b63;
   always @(posedge clk) out64 <= m1_64+m2_64+m3_64+m4_64+m5_64+m6_64+m7_64+m8_64+m9_64+m10_64+m11_64+m12_64+m13_64+m14_64+m15_64+m16_64+m17_64+m18_64+m19_64+m20_64+m21_64+m22_64+m23_64+m24_64+m25_64+m26_64+m27_64+m28_64+m29_64+m30_64+m31_64+m32_64+m33_64+m34_64+m35_64+m36_64+m37_64+m38_64+m39_64+m40_64+m41_64+m42_64+m43_64+m44_64+m45_64+m46_64+m47_64+m48_64+m49_64+m50_64+m51_64+m52_64+m53_64+m54_64+m55_64+m56_64+m57_64+m58_64+m59_64+m60_64+m61_64+m62_64+m63_64+m64_64+m65_64+m66_64+m67_64+m68_64+m69_64+m70_64+m71_64+m72_64+m73_64+m74_64+m75_64+m76_64+m77_64+m78_64+m79_64+m80_64+m81_64+m82_64+m83_64+m84_64+m85_64+m86_64+m87_64+m88_64+m89_64+m90_64+m91_64+m92_64+m93_64+m94_64+m95_64+m96_64+m97_64+m98_64+m99_64+m100_64+m101_64+m102_64+m103_64+m104_64+m105_64+m106_64+m107_64+m108_64+m109_64+m110_64+m111_64+m112_64+m113_64+m114_64+m115_64+m116_64+m117_64+b64;
   always @(posedge clk) out65 <= m1_65+m2_65+m3_65+m4_65+m5_65+m6_65+m7_65+m8_65+m9_65+m10_65+m11_65+m12_65+m13_65+m14_65+m15_65+m16_65+m17_65+m18_65+m19_65+m20_65+m21_65+m22_65+m23_65+m24_65+m25_65+m26_65+m27_65+m28_65+m29_65+m30_65+m31_65+m32_65+m33_65+m34_65+m35_65+m36_65+m37_65+m38_65+m39_65+m40_65+m41_65+m42_65+m43_65+m44_65+m45_65+m46_65+m47_65+m48_65+m49_65+m50_65+m51_65+m52_65+m53_65+m54_65+m55_65+m56_65+m57_65+m58_65+m59_65+m60_65+m61_65+m62_65+m63_65+m64_65+m65_65+m66_65+m67_65+m68_65+m69_65+m70_65+m71_65+m72_65+m73_65+m74_65+m75_65+m76_65+m77_65+m78_65+m79_65+m80_65+m81_65+m82_65+m83_65+m84_65+m85_65+m86_65+m87_65+m88_65+m89_65+m90_65+m91_65+m92_65+m93_65+m94_65+m95_65+m96_65+m97_65+m98_65+m99_65+m100_65+m101_65+m102_65+m103_65+m104_65+m105_65+m106_65+m107_65+m108_65+m109_65+m110_65+m111_65+m112_65+m113_65+m114_65+m115_65+m116_65+m117_65+b65;
   always @(posedge clk) out66 <= m1_66+m2_66+m3_66+m4_66+m5_66+m6_66+m7_66+m8_66+m9_66+m10_66+m11_66+m12_66+m13_66+m14_66+m15_66+m16_66+m17_66+m18_66+m19_66+m20_66+m21_66+m22_66+m23_66+m24_66+m25_66+m26_66+m27_66+m28_66+m29_66+m30_66+m31_66+m32_66+m33_66+m34_66+m35_66+m36_66+m37_66+m38_66+m39_66+m40_66+m41_66+m42_66+m43_66+m44_66+m45_66+m46_66+m47_66+m48_66+m49_66+m50_66+m51_66+m52_66+m53_66+m54_66+m55_66+m56_66+m57_66+m58_66+m59_66+m60_66+m61_66+m62_66+m63_66+m64_66+m65_66+m66_66+m67_66+m68_66+m69_66+m70_66+m71_66+m72_66+m73_66+m74_66+m75_66+m76_66+m77_66+m78_66+m79_66+m80_66+m81_66+m82_66+m83_66+m84_66+m85_66+m86_66+m87_66+m88_66+m89_66+m90_66+m91_66+m92_66+m93_66+m94_66+m95_66+m96_66+m97_66+m98_66+m99_66+m100_66+m101_66+m102_66+m103_66+m104_66+m105_66+m106_66+m107_66+m108_66+m109_66+m110_66+m111_66+m112_66+m113_66+m114_66+m115_66+m116_66+m117_66+b66;
   always @(posedge clk) out67 <= m1_67+m2_67+m3_67+m4_67+m5_67+m6_67+m7_67+m8_67+m9_67+m10_67+m11_67+m12_67+m13_67+m14_67+m15_67+m16_67+m17_67+m18_67+m19_67+m20_67+m21_67+m22_67+m23_67+m24_67+m25_67+m26_67+m27_67+m28_67+m29_67+m30_67+m31_67+m32_67+m33_67+m34_67+m35_67+m36_67+m37_67+m38_67+m39_67+m40_67+m41_67+m42_67+m43_67+m44_67+m45_67+m46_67+m47_67+m48_67+m49_67+m50_67+m51_67+m52_67+m53_67+m54_67+m55_67+m56_67+m57_67+m58_67+m59_67+m60_67+m61_67+m62_67+m63_67+m64_67+m65_67+m66_67+m67_67+m68_67+m69_67+m70_67+m71_67+m72_67+m73_67+m74_67+m75_67+m76_67+m77_67+m78_67+m79_67+m80_67+m81_67+m82_67+m83_67+m84_67+m85_67+m86_67+m87_67+m88_67+m89_67+m90_67+m91_67+m92_67+m93_67+m94_67+m95_67+m96_67+m97_67+m98_67+m99_67+m100_67+m101_67+m102_67+m103_67+m104_67+m105_67+m106_67+m107_67+m108_67+m109_67+m110_67+m111_67+m112_67+m113_67+m114_67+m115_67+m116_67+m117_67+b67;
   always @(posedge clk) out68 <= m1_68+m2_68+m3_68+m4_68+m5_68+m6_68+m7_68+m8_68+m9_68+m10_68+m11_68+m12_68+m13_68+m14_68+m15_68+m16_68+m17_68+m18_68+m19_68+m20_68+m21_68+m22_68+m23_68+m24_68+m25_68+m26_68+m27_68+m28_68+m29_68+m30_68+m31_68+m32_68+m33_68+m34_68+m35_68+m36_68+m37_68+m38_68+m39_68+m40_68+m41_68+m42_68+m43_68+m44_68+m45_68+m46_68+m47_68+m48_68+m49_68+m50_68+m51_68+m52_68+m53_68+m54_68+m55_68+m56_68+m57_68+m58_68+m59_68+m60_68+m61_68+m62_68+m63_68+m64_68+m65_68+m66_68+m67_68+m68_68+m69_68+m70_68+m71_68+m72_68+m73_68+m74_68+m75_68+m76_68+m77_68+m78_68+m79_68+m80_68+m81_68+m82_68+m83_68+m84_68+m85_68+m86_68+m87_68+m88_68+m89_68+m90_68+m91_68+m92_68+m93_68+m94_68+m95_68+m96_68+m97_68+m98_68+m99_68+m100_68+m101_68+m102_68+m103_68+m104_68+m105_68+m106_68+m107_68+m108_68+m109_68+m110_68+m111_68+m112_68+m113_68+m114_68+m115_68+m116_68+m117_68+b68;
   always @(posedge clk) out69 <= m1_69+m2_69+m3_69+m4_69+m5_69+m6_69+m7_69+m8_69+m9_69+m10_69+m11_69+m12_69+m13_69+m14_69+m15_69+m16_69+m17_69+m18_69+m19_69+m20_69+m21_69+m22_69+m23_69+m24_69+m25_69+m26_69+m27_69+m28_69+m29_69+m30_69+m31_69+m32_69+m33_69+m34_69+m35_69+m36_69+m37_69+m38_69+m39_69+m40_69+m41_69+m42_69+m43_69+m44_69+m45_69+m46_69+m47_69+m48_69+m49_69+m50_69+m51_69+m52_69+m53_69+m54_69+m55_69+m56_69+m57_69+m58_69+m59_69+m60_69+m61_69+m62_69+m63_69+m64_69+m65_69+m66_69+m67_69+m68_69+m69_69+m70_69+m71_69+m72_69+m73_69+m74_69+m75_69+m76_69+m77_69+m78_69+m79_69+m80_69+m81_69+m82_69+m83_69+m84_69+m85_69+m86_69+m87_69+m88_69+m89_69+m90_69+m91_69+m92_69+m93_69+m94_69+m95_69+m96_69+m97_69+m98_69+m99_69+m100_69+m101_69+m102_69+m103_69+m104_69+m105_69+m106_69+m107_69+m108_69+m109_69+m110_69+m111_69+m112_69+m113_69+m114_69+m115_69+m116_69+m117_69+b69;
   always @(posedge clk) out70 <= m1_70+m2_70+m3_70+m4_70+m5_70+m6_70+m7_70+m8_70+m9_70+m10_70+m11_70+m12_70+m13_70+m14_70+m15_70+m16_70+m17_70+m18_70+m19_70+m20_70+m21_70+m22_70+m23_70+m24_70+m25_70+m26_70+m27_70+m28_70+m29_70+m30_70+m31_70+m32_70+m33_70+m34_70+m35_70+m36_70+m37_70+m38_70+m39_70+m40_70+m41_70+m42_70+m43_70+m44_70+m45_70+m46_70+m47_70+m48_70+m49_70+m50_70+m51_70+m52_70+m53_70+m54_70+m55_70+m56_70+m57_70+m58_70+m59_70+m60_70+m61_70+m62_70+m63_70+m64_70+m65_70+m66_70+m67_70+m68_70+m69_70+m70_70+m71_70+m72_70+m73_70+m74_70+m75_70+m76_70+m77_70+m78_70+m79_70+m80_70+m81_70+m82_70+m83_70+m84_70+m85_70+m86_70+m87_70+m88_70+m89_70+m90_70+m91_70+m92_70+m93_70+m94_70+m95_70+m96_70+m97_70+m98_70+m99_70+m100_70+m101_70+m102_70+m103_70+m104_70+m105_70+m106_70+m107_70+m108_70+m109_70+m110_70+m111_70+m112_70+m113_70+m114_70+m115_70+m116_70+m117_70+b70;
   always @(posedge clk) out71 <= m1_71+m2_71+m3_71+m4_71+m5_71+m6_71+m7_71+m8_71+m9_71+m10_71+m11_71+m12_71+m13_71+m14_71+m15_71+m16_71+m17_71+m18_71+m19_71+m20_71+m21_71+m22_71+m23_71+m24_71+m25_71+m26_71+m27_71+m28_71+m29_71+m30_71+m31_71+m32_71+m33_71+m34_71+m35_71+m36_71+m37_71+m38_71+m39_71+m40_71+m41_71+m42_71+m43_71+m44_71+m45_71+m46_71+m47_71+m48_71+m49_71+m50_71+m51_71+m52_71+m53_71+m54_71+m55_71+m56_71+m57_71+m58_71+m59_71+m60_71+m61_71+m62_71+m63_71+m64_71+m65_71+m66_71+m67_71+m68_71+m69_71+m70_71+m71_71+m72_71+m73_71+m74_71+m75_71+m76_71+m77_71+m78_71+m79_71+m80_71+m81_71+m82_71+m83_71+m84_71+m85_71+m86_71+m87_71+m88_71+m89_71+m90_71+m91_71+m92_71+m93_71+m94_71+m95_71+m96_71+m97_71+m98_71+m99_71+m100_71+m101_71+m102_71+m103_71+m104_71+m105_71+m106_71+m107_71+m108_71+m109_71+m110_71+m111_71+m112_71+m113_71+m114_71+m115_71+m116_71+m117_71+b71;
   always @(posedge clk) out72 <= m1_72+m2_72+m3_72+m4_72+m5_72+m6_72+m7_72+m8_72+m9_72+m10_72+m11_72+m12_72+m13_72+m14_72+m15_72+m16_72+m17_72+m18_72+m19_72+m20_72+m21_72+m22_72+m23_72+m24_72+m25_72+m26_72+m27_72+m28_72+m29_72+m30_72+m31_72+m32_72+m33_72+m34_72+m35_72+m36_72+m37_72+m38_72+m39_72+m40_72+m41_72+m42_72+m43_72+m44_72+m45_72+m46_72+m47_72+m48_72+m49_72+m50_72+m51_72+m52_72+m53_72+m54_72+m55_72+m56_72+m57_72+m58_72+m59_72+m60_72+m61_72+m62_72+m63_72+m64_72+m65_72+m66_72+m67_72+m68_72+m69_72+m70_72+m71_72+m72_72+m73_72+m74_72+m75_72+m76_72+m77_72+m78_72+m79_72+m80_72+m81_72+m82_72+m83_72+m84_72+m85_72+m86_72+m87_72+m88_72+m89_72+m90_72+m91_72+m92_72+m93_72+m94_72+m95_72+m96_72+m97_72+m98_72+m99_72+m100_72+m101_72+m102_72+m103_72+m104_72+m105_72+m106_72+m107_72+m108_72+m109_72+m110_72+m111_72+m112_72+m113_72+m114_72+m115_72+m116_72+m117_72+b72;
   always @(posedge clk) out73 <= m1_73+m2_73+m3_73+m4_73+m5_73+m6_73+m7_73+m8_73+m9_73+m10_73+m11_73+m12_73+m13_73+m14_73+m15_73+m16_73+m17_73+m18_73+m19_73+m20_73+m21_73+m22_73+m23_73+m24_73+m25_73+m26_73+m27_73+m28_73+m29_73+m30_73+m31_73+m32_73+m33_73+m34_73+m35_73+m36_73+m37_73+m38_73+m39_73+m40_73+m41_73+m42_73+m43_73+m44_73+m45_73+m46_73+m47_73+m48_73+m49_73+m50_73+m51_73+m52_73+m53_73+m54_73+m55_73+m56_73+m57_73+m58_73+m59_73+m60_73+m61_73+m62_73+m63_73+m64_73+m65_73+m66_73+m67_73+m68_73+m69_73+m70_73+m71_73+m72_73+m73_73+m74_73+m75_73+m76_73+m77_73+m78_73+m79_73+m80_73+m81_73+m82_73+m83_73+m84_73+m85_73+m86_73+m87_73+m88_73+m89_73+m90_73+m91_73+m92_73+m93_73+m94_73+m95_73+m96_73+m97_73+m98_73+m99_73+m100_73+m101_73+m102_73+m103_73+m104_73+m105_73+m106_73+m107_73+m108_73+m109_73+m110_73+m111_73+m112_73+m113_73+m114_73+m115_73+m116_73+m117_73+b73;
   always @(posedge clk) out74 <= m1_74+m2_74+m3_74+m4_74+m5_74+m6_74+m7_74+m8_74+m9_74+m10_74+m11_74+m12_74+m13_74+m14_74+m15_74+m16_74+m17_74+m18_74+m19_74+m20_74+m21_74+m22_74+m23_74+m24_74+m25_74+m26_74+m27_74+m28_74+m29_74+m30_74+m31_74+m32_74+m33_74+m34_74+m35_74+m36_74+m37_74+m38_74+m39_74+m40_74+m41_74+m42_74+m43_74+m44_74+m45_74+m46_74+m47_74+m48_74+m49_74+m50_74+m51_74+m52_74+m53_74+m54_74+m55_74+m56_74+m57_74+m58_74+m59_74+m60_74+m61_74+m62_74+m63_74+m64_74+m65_74+m66_74+m67_74+m68_74+m69_74+m70_74+m71_74+m72_74+m73_74+m74_74+m75_74+m76_74+m77_74+m78_74+m79_74+m80_74+m81_74+m82_74+m83_74+m84_74+m85_74+m86_74+m87_74+m88_74+m89_74+m90_74+m91_74+m92_74+m93_74+m94_74+m95_74+m96_74+m97_74+m98_74+m99_74+m100_74+m101_74+m102_74+m103_74+m104_74+m105_74+m106_74+m107_74+m108_74+m109_74+m110_74+m111_74+m112_74+m113_74+m114_74+m115_74+m116_74+m117_74+b74;
   always @(posedge clk) out75 <= m1_75+m2_75+m3_75+m4_75+m5_75+m6_75+m7_75+m8_75+m9_75+m10_75+m11_75+m12_75+m13_75+m14_75+m15_75+m16_75+m17_75+m18_75+m19_75+m20_75+m21_75+m22_75+m23_75+m24_75+m25_75+m26_75+m27_75+m28_75+m29_75+m30_75+m31_75+m32_75+m33_75+m34_75+m35_75+m36_75+m37_75+m38_75+m39_75+m40_75+m41_75+m42_75+m43_75+m44_75+m45_75+m46_75+m47_75+m48_75+m49_75+m50_75+m51_75+m52_75+m53_75+m54_75+m55_75+m56_75+m57_75+m58_75+m59_75+m60_75+m61_75+m62_75+m63_75+m64_75+m65_75+m66_75+m67_75+m68_75+m69_75+m70_75+m71_75+m72_75+m73_75+m74_75+m75_75+m76_75+m77_75+m78_75+m79_75+m80_75+m81_75+m82_75+m83_75+m84_75+m85_75+m86_75+m87_75+m88_75+m89_75+m90_75+m91_75+m92_75+m93_75+m94_75+m95_75+m96_75+m97_75+m98_75+m99_75+m100_75+m101_75+m102_75+m103_75+m104_75+m105_75+m106_75+m107_75+m108_75+m109_75+m110_75+m111_75+m112_75+m113_75+m114_75+m115_75+m116_75+m117_75+b75;
   always @(posedge clk) out76 <= m1_76+m2_76+m3_76+m4_76+m5_76+m6_76+m7_76+m8_76+m9_76+m10_76+m11_76+m12_76+m13_76+m14_76+m15_76+m16_76+m17_76+m18_76+m19_76+m20_76+m21_76+m22_76+m23_76+m24_76+m25_76+m26_76+m27_76+m28_76+m29_76+m30_76+m31_76+m32_76+m33_76+m34_76+m35_76+m36_76+m37_76+m38_76+m39_76+m40_76+m41_76+m42_76+m43_76+m44_76+m45_76+m46_76+m47_76+m48_76+m49_76+m50_76+m51_76+m52_76+m53_76+m54_76+m55_76+m56_76+m57_76+m58_76+m59_76+m60_76+m61_76+m62_76+m63_76+m64_76+m65_76+m66_76+m67_76+m68_76+m69_76+m70_76+m71_76+m72_76+m73_76+m74_76+m75_76+m76_76+m77_76+m78_76+m79_76+m80_76+m81_76+m82_76+m83_76+m84_76+m85_76+m86_76+m87_76+m88_76+m89_76+m90_76+m91_76+m92_76+m93_76+m94_76+m95_76+m96_76+m97_76+m98_76+m99_76+m100_76+m101_76+m102_76+m103_76+m104_76+m105_76+m106_76+m107_76+m108_76+m109_76+m110_76+m111_76+m112_76+m113_76+m114_76+m115_76+m116_76+m117_76+b76;
   always @(posedge clk) out77 <= m1_77+m2_77+m3_77+m4_77+m5_77+m6_77+m7_77+m8_77+m9_77+m10_77+m11_77+m12_77+m13_77+m14_77+m15_77+m16_77+m17_77+m18_77+m19_77+m20_77+m21_77+m22_77+m23_77+m24_77+m25_77+m26_77+m27_77+m28_77+m29_77+m30_77+m31_77+m32_77+m33_77+m34_77+m35_77+m36_77+m37_77+m38_77+m39_77+m40_77+m41_77+m42_77+m43_77+m44_77+m45_77+m46_77+m47_77+m48_77+m49_77+m50_77+m51_77+m52_77+m53_77+m54_77+m55_77+m56_77+m57_77+m58_77+m59_77+m60_77+m61_77+m62_77+m63_77+m64_77+m65_77+m66_77+m67_77+m68_77+m69_77+m70_77+m71_77+m72_77+m73_77+m74_77+m75_77+m76_77+m77_77+m78_77+m79_77+m80_77+m81_77+m82_77+m83_77+m84_77+m85_77+m86_77+m87_77+m88_77+m89_77+m90_77+m91_77+m92_77+m93_77+m94_77+m95_77+m96_77+m97_77+m98_77+m99_77+m100_77+m101_77+m102_77+m103_77+m104_77+m105_77+m106_77+m107_77+m108_77+m109_77+m110_77+m111_77+m112_77+m113_77+m114_77+m115_77+m116_77+m117_77+b77;
   always @(posedge clk) out78 <= m1_78+m2_78+m3_78+m4_78+m5_78+m6_78+m7_78+m8_78+m9_78+m10_78+m11_78+m12_78+m13_78+m14_78+m15_78+m16_78+m17_78+m18_78+m19_78+m20_78+m21_78+m22_78+m23_78+m24_78+m25_78+m26_78+m27_78+m28_78+m29_78+m30_78+m31_78+m32_78+m33_78+m34_78+m35_78+m36_78+m37_78+m38_78+m39_78+m40_78+m41_78+m42_78+m43_78+m44_78+m45_78+m46_78+m47_78+m48_78+m49_78+m50_78+m51_78+m52_78+m53_78+m54_78+m55_78+m56_78+m57_78+m58_78+m59_78+m60_78+m61_78+m62_78+m63_78+m64_78+m65_78+m66_78+m67_78+m68_78+m69_78+m70_78+m71_78+m72_78+m73_78+m74_78+m75_78+m76_78+m77_78+m78_78+m79_78+m80_78+m81_78+m82_78+m83_78+m84_78+m85_78+m86_78+m87_78+m88_78+m89_78+m90_78+m91_78+m92_78+m93_78+m94_78+m95_78+m96_78+m97_78+m98_78+m99_78+m100_78+m101_78+m102_78+m103_78+m104_78+m105_78+m106_78+m107_78+m108_78+m109_78+m110_78+m111_78+m112_78+m113_78+m114_78+m115_78+m116_78+m117_78+b78;
   always @(posedge clk) out79 <= m1_79+m2_79+m3_79+m4_79+m5_79+m6_79+m7_79+m8_79+m9_79+m10_79+m11_79+m12_79+m13_79+m14_79+m15_79+m16_79+m17_79+m18_79+m19_79+m20_79+m21_79+m22_79+m23_79+m24_79+m25_79+m26_79+m27_79+m28_79+m29_79+m30_79+m31_79+m32_79+m33_79+m34_79+m35_79+m36_79+m37_79+m38_79+m39_79+m40_79+m41_79+m42_79+m43_79+m44_79+m45_79+m46_79+m47_79+m48_79+m49_79+m50_79+m51_79+m52_79+m53_79+m54_79+m55_79+m56_79+m57_79+m58_79+m59_79+m60_79+m61_79+m62_79+m63_79+m64_79+m65_79+m66_79+m67_79+m68_79+m69_79+m70_79+m71_79+m72_79+m73_79+m74_79+m75_79+m76_79+m77_79+m78_79+m79_79+m80_79+m81_79+m82_79+m83_79+m84_79+m85_79+m86_79+m87_79+m88_79+m89_79+m90_79+m91_79+m92_79+m93_79+m94_79+m95_79+m96_79+m97_79+m98_79+m99_79+m100_79+m101_79+m102_79+m103_79+m104_79+m105_79+m106_79+m107_79+m108_79+m109_79+m110_79+m111_79+m112_79+m113_79+m114_79+m115_79+m116_79+m117_79+b79;
   always @(posedge clk) out80 <= m1_80+m2_80+m3_80+m4_80+m5_80+m6_80+m7_80+m8_80+m9_80+m10_80+m11_80+m12_80+m13_80+m14_80+m15_80+m16_80+m17_80+m18_80+m19_80+m20_80+m21_80+m22_80+m23_80+m24_80+m25_80+m26_80+m27_80+m28_80+m29_80+m30_80+m31_80+m32_80+m33_80+m34_80+m35_80+m36_80+m37_80+m38_80+m39_80+m40_80+m41_80+m42_80+m43_80+m44_80+m45_80+m46_80+m47_80+m48_80+m49_80+m50_80+m51_80+m52_80+m53_80+m54_80+m55_80+m56_80+m57_80+m58_80+m59_80+m60_80+m61_80+m62_80+m63_80+m64_80+m65_80+m66_80+m67_80+m68_80+m69_80+m70_80+m71_80+m72_80+m73_80+m74_80+m75_80+m76_80+m77_80+m78_80+m79_80+m80_80+m81_80+m82_80+m83_80+m84_80+m85_80+m86_80+m87_80+m88_80+m89_80+m90_80+m91_80+m92_80+m93_80+m94_80+m95_80+m96_80+m97_80+m98_80+m99_80+m100_80+m101_80+m102_80+m103_80+m104_80+m105_80+m106_80+m107_80+m108_80+m109_80+m110_80+m111_80+m112_80+m113_80+m114_80+m115_80+m116_80+m117_80+b80;
   always @(posedge clk) out81 <= m1_81+m2_81+m3_81+m4_81+m5_81+m6_81+m7_81+m8_81+m9_81+m10_81+m11_81+m12_81+m13_81+m14_81+m15_81+m16_81+m17_81+m18_81+m19_81+m20_81+m21_81+m22_81+m23_81+m24_81+m25_81+m26_81+m27_81+m28_81+m29_81+m30_81+m31_81+m32_81+m33_81+m34_81+m35_81+m36_81+m37_81+m38_81+m39_81+m40_81+m41_81+m42_81+m43_81+m44_81+m45_81+m46_81+m47_81+m48_81+m49_81+m50_81+m51_81+m52_81+m53_81+m54_81+m55_81+m56_81+m57_81+m58_81+m59_81+m60_81+m61_81+m62_81+m63_81+m64_81+m65_81+m66_81+m67_81+m68_81+m69_81+m70_81+m71_81+m72_81+m73_81+m74_81+m75_81+m76_81+m77_81+m78_81+m79_81+m80_81+m81_81+m82_81+m83_81+m84_81+m85_81+m86_81+m87_81+m88_81+m89_81+m90_81+m91_81+m92_81+m93_81+m94_81+m95_81+m96_81+m97_81+m98_81+m99_81+m100_81+m101_81+m102_81+m103_81+m104_81+m105_81+m106_81+m107_81+m108_81+m109_81+m110_81+m111_81+m112_81+m113_81+m114_81+m115_81+m116_81+m117_81+b81;
endmodule