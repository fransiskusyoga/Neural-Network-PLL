`include "actifunc.v"
module layer_12(in1,in2,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   input signed [8:0] in1,in2;
   output signed [16:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   wire signed [19:0] m1_1,m1_2,m1_3,m1_4,m1_5,m1_6,m1_7,m1_8;
   wire signed [19:0] m2_9,m2_10;
   wire signed [11:0] w1_1 = $signed(12'h0);
   wire signed [11:0] w1_2 = $signed(12'hE5C);
   wire signed [11:0] w1_3 = $signed(12'hC1B);
   wire signed [11:0] w1_4 = $signed(12'hF02);
   wire signed [11:0] w1_5 = $signed(12'hD9C);
   wire signed [11:0] w1_6 = $signed(12'hD97);
   wire signed [11:0] w1_7 = $signed(12'hFFF);
   wire signed [11:0] w1_8 = $signed(12'hD8B);
   wire signed [11:0] w2_9 = $signed(12'h25);
   wire signed [11:0] w2_10 = $signed(12'h37);
   wire signed [16:0] b1 = $signed(17'h56);
   wire signed [16:0] b2 = $signed(17'hD3);
   wire signed [16:0] b3 = $signed(17'h44);
   wire signed [16:0] b4 = $signed(17'h80);
   wire signed [16:0] b5 = $signed(17'h6D);
   wire signed [16:0] b6 = $signed(17'hC1);
   wire signed [16:0] b7 = $signed(17'h1FFDF);
   wire signed [16:0] b8 = $signed(17'hAC);
   wire signed [16:0] b9 = $signed(17'h1FFAC);
   wire signed [16:0] b10 = $signed(17'h1FF2E);
   assign m1_1 = in1*w1_1;
   assign m1_2 = in1*w1_2;
   assign m1_3 = in1*w1_3;
   assign m1_4 = in1*w1_4;
   assign m1_5 = in1*w1_5;
   assign m1_6 = in1*w1_6;
   assign m1_7 = in1*w1_7;
   assign m1_8 = in1*w1_8;
   assign m2_9 = in2*w2_9;
   assign m2_10 = in2*w2_10;
   assign out1 = { {1{m1_1[19]}} , m1_1[19:4] }+b1;
   assign out2 = { {1{m1_2[19]}} , m1_2[19:4] }+b2;
   assign out3 = { {1{m1_3[19]}} , m1_3[19:4] }+b3;
   assign out4 = { {1{m1_4[19]}} , m1_4[19:4] }+b4;
   assign out5 = { {1{m1_5[19]}} , m1_5[19:4] }+b5;
   assign out6 = { {1{m1_6[19]}} , m1_6[19:4] }+b6;
   assign out7 = { {1{m1_7[19]}} , m1_7[19:4] }+b7;
   assign out8 = { {1{m1_8[19]}} , m1_8[19:4] }+b8;
   assign out9 = { {1{m2_9[19]}} , m2_9[19:4] }+b9;
   assign out10 = { {1{m2_10[19]}} , m2_10[19:4] }+b10;
endmodule