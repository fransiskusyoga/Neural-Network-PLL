module test_tb();
   reg [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36;
   wire [7:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   test_top TopModule(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   initial begin
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h4; in15=6'h0; in16=6'h2; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h4; in29=6'h0; in30=6'h0; in31=6'h9; in32=6'h0; in33=6'h0; in34=6'h7; in35=6'hA; in36=6'h9;
      #50 in1=6'h3; in2=6'h0; in3=6'h2; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h1; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h9; in13=6'h0; in14=6'h9; in15=6'h0; in16=6'h3; in17=6'h0; in18=6'h5; in19=6'h0; in20=6'h9; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h1; in29=6'h0; in30=6'h0; in31=6'h8; in32=6'h6; in33=6'h0; in34=6'h2; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h9; in3=6'h0; in4=6'hC; in5=6'h7; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h5; in12=6'h1; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h1; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h4; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h2;
      #50 in1=6'h0; in2=6'h1; in3=6'h0; in4=6'h2; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h1; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h8; in29=6'h0; in30=6'h0; in31=6'h3; in32=6'h0; in33=6'h0; in34=6'h1; in35=6'h6; in36=6'h6;
      #50 in1=6'h0; in2=6'h8; in3=6'h0; in4=6'h6; in5=6'h3; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h6; in12=6'h4; in13=6'h0; in14=6'h0; in15=6'h2; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h1; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h2; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h9; in12=6'h0; in13=6'h6; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h6; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h4; in22=6'h0; in23=6'h0; in24=6'h3; in25=6'h4; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h5; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h9; in3=6'h0; in4=6'hA; in5=6'h5; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h6; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h2; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h3;
      #50 in1=6'h4; in2=6'h3; in3=6'h7; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h5; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h2; in13=6'h7; in14=6'h0; in15=6'h4; in16=6'h0; in17=6'h2; in18=6'h8; in19=6'h0; in20=6'h0; in21=6'h1; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h6; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h7; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h8; in17=6'h0; in18=6'h4; in19=6'h2; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'hB; in26=6'h0; in27=6'h1; in28=6'hA; in29=6'h3; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h7; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h5; in11=6'h8; in12=6'h0; in13=6'h6; in14=6'h0; in15=6'h1; in16=6'h0; in17=6'h8; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h6; in22=6'h0; in23=6'h0; in24=6'h5; in25=6'h2; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h3; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h6; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h8; in27=6'h1; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h2; in34=6'h7; in35=6'h0; in36=6'h4;
      #50 in1=6'h0; in2=6'h3; in3=6'h0; in4=6'h3; in5=6'h4; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h8; in12=6'h0; in13=6'h2; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h7; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h1; in35=6'h0; in36=6'hB;
      #50 in1=6'h3; in2=6'h1; in3=6'h0; in4=6'h4; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h5; in13=6'h0; in14=6'h6; in15=6'h0; in16=6'h1; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h8; in23=6'h0; in24=6'h4; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h1; in32=6'h0; in33=6'h0; in34=6'h1; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h3; in13=6'h0; in14=6'h4; in15=6'h1; in16=6'h1; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h3; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h1; in26=6'h0; in27=6'h3; in28=6'h2; in29=6'h0; in30=6'h1; in31=6'h4; in32=6'h4; in33=6'h0; in34=6'h2; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'hA; in22=6'h0; in23=6'h0; in24=6'h9; in25=6'h7; in26=6'h0; in27=6'h0; in28=6'h4; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h6; in36=6'h0;
      #50 in1=6'h7; in2=6'h2; in3=6'h0; in4=6'h3; in5=6'h4; in6=6'h6; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h5; in13=6'h0; in14=6'h5; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h4; in23=6'h0; in24=6'h0; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h1; in32=6'h0; in33=6'h0; in34=6'h3; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h3; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h4; in7=6'hA; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h6; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h3; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h5; in34=6'h5; in35=6'h0; in36=6'h4;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h1; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h5; in20=6'h6; in21=6'h0; in22=6'h0; in23=6'h2; in24=6'h0; in25=6'h2; in26=6'h2; in27=6'h9; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h3; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h3; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h2; in9=6'h3; in10=6'h0; in11=6'h0; in12=6'h4; in13=6'h0; in14=6'h7; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h3; in19=6'h3; in20=6'h4; in21=6'h0; in22=6'h0; in23=6'h6; in24=6'h0; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h5; in32=6'h4; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h5; in2=6'h0; in3=6'h1; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h5; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h9; in13=6'h0; in14=6'h6; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h6; in19=6'h0; in20=6'hA; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'hA; in32=6'h9; in33=6'h0; in34=6'h1; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h3; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h8; in17=6'h0; in18=6'h2; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h8; in26=6'h0; in27=6'h0; in28=6'hB; in29=6'h8; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h5; in2=6'h5; in3=6'h6; in4=6'h0; in5=6'h1; in6=6'h0; in7=6'h1; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h2; in13=6'h2; in14=6'h0; in15=6'h1; in16=6'h0; in17=6'h3; in18=6'h5; in19=6'h0; in20=6'h0; in21=6'h2; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h6; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h5; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h1; in16=6'h0; in17=6'h0; in18=6'h4; in19=6'h4; in20=6'h4; in21=6'h3; in22=6'h0; in23=6'h5; in24=6'h0; in25=6'h6; in26=6'h2; in27=6'h9; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h5; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h7; in10=6'h1; in11=6'h1; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h1; in16=6'hA; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h2; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h4; in26=6'h0; in27=6'h0; in28=6'h6; in29=6'hA; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h1; in2=6'h4; in3=6'h0; in4=6'h5; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h1; in15=6'h2; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h5; in23=6'h0; in24=6'h2; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h4; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h2; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h3; in9=6'h0; in10=6'h0; in11=6'hC; in12=6'h0; in13=6'h6; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h5; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h8;
      #50 in1=6'h6; in2=6'h0; in3=6'h2; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h9; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'hA; in13=6'h0; in14=6'h4; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h6; in19=6'h0; in20=6'hA; in21=6'h0; in22=6'h0; in23=6'h2; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'hB; in32=6'hB; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h5; in15=6'h0; in16=6'h1; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h5; in29=6'h0; in30=6'h0; in31=6'hA; in32=6'h0; in33=6'h0; in34=6'h8; in35=6'hA; in36=6'h7;
      #50 in1=6'h2; in2=6'h1; in3=6'h0; in4=6'h4; in5=6'h0; in6=6'h2; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h5; in13=6'h0; in14=6'h6; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h7; in23=6'h0; in24=6'h2; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h2; in32=6'h0; in33=6'h0; in34=6'h3; in35=6'h0; in36=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h2; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h1; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h7; in29=6'h0; in30=6'h0; in31=6'h7; in32=6'h0; in33=6'h0; in34=6'h4; in35=6'h9; in36=6'h7;
   end
endmodule