module lenet300_tb();
   reg [14:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598;
   wire [15:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   lenet300_top TopModule(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   initial begin
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7D9A; in74=15'h1DE; in75=15'h3F8; in76=15'h3F8; in77=15'h1D6; in78=15'h1DE; in79=15'h3F8; in80=15'h3F8; in81=15'h2E7; in82=15'h7EAB; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7E42; in97=15'h3C0; in98=15'h390; in99=15'h3D0; in100=15'h3F0; in101=15'h3F0; in102=15'h390; in103=15'h2BF; in104=15'h367; in105=15'h3F0; in106=15'h3C8; in107=15'h7E3A; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7CB1; in120=15'h2A7; in121=15'h3F0; in122=15'h175; in123=15'h390; in124=15'h357; in125=15'h4C; in126=15'h7D11; in127=15'h7C48; in128=15'h7CE9; in129=15'h22E; in130=15'h3F8; in131=15'h7F9C; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7F94; in145=15'h3F0; in146=15'h2DF; in147=15'h7EFB; in148=15'h1CE; in149=15'h7D31; in150=15'h7C00; in151=15'h7C00; in152=15'h7C00; in153=15'h7D9A; in154=15'h357; in155=15'h3F8; in156=15'h7E8B; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7E32; in168=15'h3B0; in169=15'h3F8; in170=15'h7F3B; in171=15'h7C00; in172=15'h7C00; in173=15'h7C00; in174=15'h7C00; in175=15'h7C00; in176=15'h7D31; in177=15'h2EF; in178=15'h3F8; in179=15'h7FFC; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h10D; in194=15'h3F0; in195=15'h1AE; in196=15'h7C30; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7E42; in202=15'h35F; in203=15'h3F0; in204=15'h1CE; in205=15'h7C48; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7D9A; in219=15'h36F; in220=15'h3C8; in221=15'h7DD2; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C18; in226=15'h7FEC; in227=15'h3F8; in228=15'h3F0; in229=15'h1BE; in230=15'h7C68; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h1C6; in244=15'h3F8; in245=15'h5C; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C89; in250=15'h64; in251=15'h3F0; in252=15'h3F8; in253=15'hBD; in254=15'h7C68; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h1CE; in271=15'h3F8; in272=15'h7E93; in273=15'h7C00; in274=15'h7C00; in275=15'h7C99; in276=15'h266; in277=15'h3F8; in278=15'h3F8; in279=15'h7E22; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h1C6; in295=15'h3F8; in296=15'h1F6; in297=15'h7DDA; in298=15'h7C89; in299=15'h266; in300=15'h3F0; in301=15'h236; in302=15'h7CB9; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7E1A; in319=15'h3B0; in320=15'h3F0; in321=15'h3D0; in322=15'h307; in323=15'h3F8; in324=15'h276; in325=15'h7C48; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7D61; in345=15'h14D; in346=15'h3F0; in347=15'h3F0; in348=15'h3F8; in349=15'h7F9C; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h14; in371=15'h3F8; in372=15'h3F8; in373=15'h3F8; in374=15'h16D; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7F94; in394=15'h3E0; in395=15'h3F0; in396=15'h367; in397=15'h3F8; in398=15'h276; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C58; in416=15'hED; in417=15'h36F; in418=15'h388; in419=15'h7F8C; in420=15'h7DFA; in421=15'h3F8; in422=15'h276; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h1B6; in440=15'h3F0; in441=15'h3F8; in442=15'h7D82; in443=15'h7C00; in444=15'h7C00; in445=15'h3F8; in446=15'h276; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h287; in464=15'h3F8; in465=15'h7EEB; in466=15'h7C00; in467=15'h7C00; in468=15'h7EAB; in469=15'h400; in470=15'h27E; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7E52; in489=15'h3F0; in490=15'h1A6; in491=15'h7F4B; in492=15'h2B7; in493=15'h3C0; in494=15'h3F8; in495=15'h276; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7CA9; in512=15'h3B8; in513=15'h3F8; in514=15'h3F0; in515=15'h3F0; in516=15'h3A8; in517=15'h26E; in518=15'h7D71; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'hBD; in536=15'h3F8; in537=15'h256; in538=15'h7FBC; in539=15'h7D61; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C58; in97=15'h7FD4; in98=15'h24; in99=15'h400; in100=15'h3F0; in101=15'h367; in102=15'h24; in103=15'h24; in104=15'h7D49; in105=15'h7C18; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C99; in119=15'h7FDC; in120=15'h36F; in121=15'h3E8; in122=15'h3E8; in123=15'h3F0; in124=15'h3E8; in125=15'h3E8; in126=15'h3E8; in127=15'h3E8; in128=15'h3E8; in129=15'h7FAC; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C48; in143=15'h24E; in144=15'h3E8; in145=15'h3E8; in146=15'h2DF; in147=15'hF5; in148=15'h7F03; in149=15'h7F03; in150=15'h7F03; in151=15'h7F03; in152=15'h1F6; in153=15'h3E8; in154=15'h13D; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7D09; in166=15'h1EE; in167=15'h3E8; in168=15'h367; in169=15'hED; in170=15'h7C40; in171=15'h7C00; in172=15'h7C00; in173=15'h7C00; in174=15'h7C00; in175=15'h7C00; in176=15'h7DEA; in177=15'h3E8; in178=15'h13D; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h3C; in192=15'h3E8; in193=15'h3E8; in194=15'h5C; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h9D; in203=15'h3E8; in204=15'h5C; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7CE1; in217=15'h34F; in218=15'h3E8; in219=15'h115; in220=15'h7C60; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7D31; in228=15'h35F; in229=15'h115; in230=15'h7C60; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7CC9; in242=15'h307; in243=15'h3E8; in244=15'h1AE; in245=15'h7DCA; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h4; in252=15'h2B7; in253=15'h1FE; in254=15'h7D41; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h14D; in270=15'h3E8; in271=15'h3E8; in272=15'h388; in273=15'h7F94; in274=15'h7DC2; in275=15'h7C00; in276=15'h7C28; in277=15'h7F6B; in278=15'h30F; in279=15'h7E5A; in280=15'h7C50; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7D39; in294=15'h14D; in295=15'h3E8; in296=15'h3E8; in297=15'h3E8; in298=15'h398; in299=15'h32F; in300=15'h33F; in301=15'h3E8; in302=15'h3D0; in303=15'h4; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C18; in319=15'h7F43; in320=15'h1C; in321=15'h18E; in322=15'h3E8; in323=15'h3E8; in324=15'h3F0; in325=15'h3E8; in326=15'h3E8; in327=15'h3D8; in328=15'h1BE; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7C38; in350=15'h85; in351=15'h3F0; in352=15'h3F0; in353=15'hC; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7CC1; in375=15'h3E8; in376=15'h3E8; in377=15'h307; in378=15'h7CF9; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C91; in398=15'h287; in399=15'h3E8; in400=15'h3E8; in401=15'hC; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7CA9; in421=15'h25E; in422=15'h3F0; in423=15'h3E8; in424=15'h9D; in425=15'h7CE1; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7CC1; in444=15'h246; in445=15'h3E8; in446=15'h3F0; in447=15'h276; in448=15'h7CD9; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7F23; in467=15'h2C7; in468=15'h3E8; in469=15'h3E8; in470=15'h28F; in471=15'h7CD1; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7F23; in491=15'h3A0; in492=15'h3E8; in493=15'h3E8; in494=15'hD5; in495=15'h7CB9; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C99; in512=15'h1BE; in513=15'h3A8; in514=15'h3E8; in515=15'h3E8; in516=15'h125; in517=15'h7CC1; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'hF5; in535=15'h3E8; in536=15'h3E8; in537=15'h2C7; in538=15'h7F13; in539=15'h7C18; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h14D; in556=15'h3E8; in557=15'h105; in558=15'h7CF1; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C60; in14=15'h22E; in15=15'h7DBA; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7D49; in33=15'h3F8; in34=15'h2D7; in35=15'h7CD9; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7F63; in54=15'h3F8; in55=15'h3F8; in56=15'hFD; in57=15'h7C28; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7D69; in76=15'h3E8; in77=15'h14D; in78=15'h3F8; in79=15'h7F7B; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7CE9; in100=15'h7E72; in101=15'h7C89; in102=15'h28F; in103=15'h26E; in104=15'h7C20; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h7C00; in124=15'h7C00; in125=15'h7C00; in126=15'h7FDC; in127=15'h3F8; in128=15'h7E32; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h7C00; in150=15'h7C00; in151=15'h7CB1; in152=15'h388; in153=15'h7FEC; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h7C00; in174=15'h7C00; in175=15'h7C00; in176=15'h34F; in177=15'h7FEC; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h2A7; in203=15'h7FEC; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h2F7; in229=15'h7FEC; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7E1A; in253=15'h3E0; in254=15'h7F94; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C30; in279=15'h125; in280=15'h30F; in281=15'h7CA9; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C08; in293=15'h7EA3; in294=15'h1C6; in295=15'hD5; in296=15'h7D31; in297=15'h7C08; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h7C00; in302=15'h7F9C; in303=15'h3F8; in304=15'h7F73; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7D21; in317=15'h3F8; in318=15'h3F8; in319=15'h3F8; in320=15'h3F8; in321=15'hDD; in322=15'h7C50; in323=15'h7C00; in324=15'h7C00; in325=15'h7CF1; in326=15'h22E; in327=15'h1AE; in328=15'h7C40; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7EE3; in342=15'h3F8; in343=15'h3B8; in344=15'h7C48; in345=15'hCD; in346=15'h3D8; in347=15'h246; in348=15'h7CE1; in349=15'h7DDA; in350=15'h307; in351=15'h28F; in352=15'h7D49; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7E62; in367=15'h3F8; in368=15'h186; in369=15'h7C00; in370=15'h7C00; in371=15'h7FEC; in372=15'h3C8; in373=15'h36F; in374=15'h3D8; in375=15'h1B6; in376=15'h7D29; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7D21; in391=15'h3F8; in392=15'h7FFC; in393=15'h7C00; in394=15'h7E12; in395=15'h14; in396=15'h388; in397=15'h3F8; in398=15'h398; in399=15'h7CA9; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C38; in415=15'h10D; in416=15'h3F0; in417=15'h276; in418=15'h3F8; in419=15'h3C8; in420=15'h1A6; in421=15'h2BF; in422=15'h3F8; in423=15'h7F8C; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C30; in440=15'h4; in441=15'hBD; in442=15'h7FFC; in443=15'h7D82; in444=15'h7C00; in445=15'h7C40; in446=15'h276; in447=15'h337; in448=15'h7D39; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7C00; in468=15'h7C00; in469=15'h7C00; in470=15'h7D01; in471=15'h16D; in472=15'h256; in473=15'h7C18; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C78; in69=15'h1AE; in70=15'h7F4B; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7D19; in78=15'h7DFA; in79=15'h7ED3; in80=15'hF5; in81=15'h34F; in82=15'h400; in83=15'h20E; in84=15'h7C81; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h6C; in93=15'h3F8; in94=15'h398; in95=15'h4; in96=15'h7FF4; in97=15'h7FF4; in98=15'h7FF4; in99=15'h25E; in100=15'h2EF; in101=15'h37F; in102=15'h3F8; in103=15'h3F8; in104=15'h3F8; in105=15'h3F8; in106=15'h3F8; in107=15'h3F8; in108=15'h7DF2; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h30F; in117=15'h3F8; in118=15'h3F8; in119=15'h3F8; in120=15'h3F8; in121=15'h3F8; in122=15'h3F8; in123=15'h3F8; in124=15'h3F8; in125=15'h3F8; in126=15'h3F8; in127=15'h3F8; in128=15'h3F8; in129=15'h3F8; in130=15'h3F8; in131=15'h3F8; in132=15'h7DF2; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7F84; in141=15'h3F0; in142=15'h287; in143=15'h7ED3; in144=15'h3F8; in145=15'h3F8; in146=15'h3F8; in147=15'h3F8; in148=15'h3F8; in149=15'h3F8; in150=15'h3F8; in151=15'h32F; in152=15'h226; in153=15'h7F6B; in154=15'h7F2B; in155=15'h7F2B; in156=15'h7C78; in157=15'h7C08; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h1DE; in165=15'h3F8; in166=15'h7FEC; in167=15'h7E7A; in168=15'h357; in169=15'h3F8; in170=15'h36F; in171=15'h32F; in172=15'h307; in173=15'h2C; in174=15'h7E8B; in175=15'h7CB1; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C50; in190=15'h297; in191=15'h357; in192=15'h7CC9; in193=15'h7C00; in194=15'h7C78; in195=15'h7E42; in196=15'h7CB1; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7D8A; in216=15'h3F8; in217=15'h5C; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h145; in241=15'h3F8; in242=15'h7F2B; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h2EF; in268=15'h3F8; in269=15'h27E; in270=15'h24; in271=15'h7E93; in272=15'h7E0A; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h2EF; in292=15'h3F8; in293=15'h3F8; in294=15'h3F8; in295=15'h3F8; in296=15'h3E0; in297=15'h34F; in298=15'h85; in299=15'h7ED3; in300=15'h7C48; in301=15'h7C00; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7D82; in315=15'h3B8; in316=15'h3F8; in317=15'h3F8; in318=15'h3F8; in319=15'h3F8; in320=15'h3F8; in321=15'h3F8; in322=15'h3F8; in323=15'h3F8; in324=15'h297; in325=15'h7D49; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h11D; in341=15'h307; in342=15'h3F8; in343=15'h307; in344=15'h3F8; in345=15'h3F8; in346=15'h3F8; in347=15'h3F8; in348=15'h3F8; in349=15'h3F8; in350=15'h32F; in351=15'h7E3A; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C18; in366=15'h7C60; in367=15'h7C99; in368=15'h7C60; in369=15'h7C99; in370=15'h7D39; in371=15'h7F9C; in372=15'h8D; in373=15'h35F; in374=15'h3F8; in375=15'h3F8; in376=15'h3D8; in377=15'h7F33; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7CF1; in398=15'h165; in399=15'h3D8; in400=15'h3F8; in401=15'h327; in402=15'h7D41; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7DA2; in418=15'h7DD2; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7C00; in423=15'h16D; in424=15'h3F8; in425=15'h3F8; in426=15'h1AE; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7CB1; in441=15'h3C0; in442=15'h3D0; in443=15'h7C; in444=15'h7CD9; in445=15'h7C00; in446=15'h7C00; in447=15'h7D51; in448=15'h388; in449=15'h3F8; in450=15'h2E7; in451=15'h7C68; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C30; in465=15'h236; in466=15'h3F8; in467=15'h3F8; in468=15'h35F; in469=15'h22E; in470=15'h22E; in471=15'h35F; in472=15'h3F8; in473=15'h3F8; in474=15'h30F; in475=15'h7C70; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7FCC; in491=15'h3F8; in492=15'h3F8; in493=15'h3F8; in494=15'h3F8; in495=15'h3F8; in496=15'h3F8; in497=15'h3F8; in498=15'h3F8; in499=15'hE5; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C50; in514=15'h9D; in515=15'h3F8; in516=15'h3F8; in517=15'h3F8; in518=15'h3F8; in519=15'h3F8; in520=15'h3F8; in521=15'h1BE; in522=15'h7C50; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C68; in538=15'h7F53; in539=15'hED; in540=15'h3C8; in541=15'h3F8; in542=15'h1E6; in543=15'h7E2A; in544=15'h7C68; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7EAB; in93=15'h1F6; in94=15'h7C18; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7C00; in100=15'h7C00; in101=15'h7C00; in102=15'h7C00; in103=15'hFD; in104=15'h3E0; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7D41; in116=15'h2FF; in117=15'h3F8; in118=15'h7D71; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h7C00; in124=15'h7C00; in125=15'h7C00; in126=15'h7C00; in127=15'h33F; in128=15'h3D8; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'hD5; in141=15'h3F8; in142=15'h3F8; in143=15'h7C48; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h7C00; in150=15'h7C00; in151=15'h7C00; in152=15'h33F; in153=15'h3D8; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h186; in165=15'h3F8; in166=15'h14D; in167=15'h7C08; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h7C00; in174=15'h7C00; in175=15'h7D61; in176=15'h3B0; in177=15'h3D8; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7D61; in190=15'h3E8; in191=15'h3E8; in192=15'h7E7A; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7E4A; in202=15'h3F8; in203=15'h390; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7FEC; in216=15'h3F8; in217=15'h22E; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7E4A; in228=15'h3F8; in229=15'hCD; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h1E6; in241=15'h3F8; in242=15'h34; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7E4A; in253=15'h3F8; in254=15'hCD; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h1E6; in268=15'h3F8; in269=15'h30F; in270=15'h7E9B; in271=15'h7CA1; in272=15'h7C91; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C00; in279=15'hC5; in280=15'h3F8; in281=15'hCD; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7EE3; in292=15'h3F0; in293=15'h3F8; in294=15'h3F8; in295=15'h3F8; in296=15'h3D0; in297=15'h196; in298=15'h196; in299=15'h16D; in300=15'h7E9B; in301=15'h7E9B; in302=15'h7EB3; in303=15'h32F; in304=15'h3F8; in305=15'h1C6; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h18E; in317=15'h3F8; in318=15'h3F8; in319=15'h3F8; in320=15'h3F8; in321=15'h3F8; in322=15'h3F8; in323=15'h3F8; in324=15'h3F8; in325=15'h3F8; in326=15'h3F8; in327=15'h3F8; in328=15'h3F8; in329=15'h3F0; in330=15'h7E2A; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C58; in342=15'h7EF3; in343=15'h7C; in344=15'h36F; in345=15'h388; in346=15'h3B0; in347=15'h3F8; in348=15'h3F8; in349=15'h3B0; in350=15'h3C8; in351=15'h3F8; in352=15'h3F8; in353=15'h377; in354=15'h7F4B; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7CD9; in372=15'h7E93; in373=15'h7E93; in374=15'h7CD1; in375=15'h7D69; in376=15'hCD; in377=15'h3F8; in378=15'h1DE; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7C40; in400=15'h266; in401=15'h398; in402=15'h7CD9; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7C00; in423=15'h7EA3; in424=15'h3F8; in425=15'h1B6; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7C00; in445=15'h7C00; in446=15'h7C00; in447=15'h13D; in448=15'h3F8; in449=15'h1B6; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7C00; in468=15'h7C00; in469=15'h7C00; in470=15'h7C60; in471=15'h37F; in472=15'h3D0; in473=15'h7D92; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'hC5; in496=15'h3F8; in497=15'h155; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h16D; in519=15'h3F8; in520=15'h7EBB; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C68; in541=15'h3B8; in542=15'h25E; in543=15'h7C30; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C50; in562=15'h307; in563=15'h7F9C; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7D49; in46=15'h7F84; in47=15'hE5; in48=15'hE5; in49=15'h7E52; in50=15'h7D49; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C28; in66=15'h9D; in67=15'h390; in68=15'h3F0; in69=15'h3F0; in70=15'h3F8; in71=15'h3F0; in72=15'h390; in73=15'h23E; in74=15'h7FB4; in75=15'h7C81; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'hE5; in90=15'h3C0; in91=15'h85; in92=15'h7E72; in93=15'h7E72; in94=15'h7E72; in95=15'h105; in96=15'h23E; in97=15'h3F0; in98=15'h3F0; in99=15'h367; in100=15'h7FEC; in101=15'h7C00; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h3F8; in114=15'h7EDB; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C30; in121=15'h7D11; in122=15'h1FE; in123=15'h3F8; in124=15'h3E0; in125=15'h175; in126=15'h7C18; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h3F8; in139=15'h7D39; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h64; in149=15'h3F0; in150=15'h3F0; in151=15'h1C; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7F1B; in163=15'h7C78; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h24; in174=15'h3F8; in175=15'h377; in176=15'h7DDA; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C18; in200=15'h74; in201=15'h3F0; in202=15'h246; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7E7A; in227=15'h3F0; in228=15'h3F0; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C38; in248=15'h7D41; in249=15'h7D41; in250=15'h7E6A; in251=15'h7D69; in252=15'h377; in253=15'h3F0; in254=15'h7C81; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7E22; in274=15'h22E; in275=15'h3F0; in276=15'h3F8; in277=15'h3F0; in278=15'h3F0; in279=15'h3F0; in280=15'h3F0; in281=15'h21E; in282=15'h7C78; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7DDA; in296=15'h37F; in297=15'h3F8; in298=15'h3F8; in299=15'h3F8; in300=15'h226; in301=15'h2F7; in302=15'h3F8; in303=15'h3F8; in304=15'h3F8; in305=15'h400; in306=15'h3F8; in307=15'h1D6; in308=15'h7DCA; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C40; in319=15'h37F; in320=15'h3F0; in321=15'h37F; in322=15'h74; in323=15'h7DEA; in324=15'h7C00; in325=15'h7C91; in326=15'h7F4B; in327=15'h3F0; in328=15'h3F0; in329=15'hF5; in330=15'h34F; in331=15'h3C0; in332=15'h3C0; in333=15'h5C; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h4; in344=15'h3F8; in345=15'h28F; in346=15'h7CC1; in347=15'h7C00; in348=15'h7C00; in349=15'h7C00; in350=15'h7C00; in351=15'h7F6B; in352=15'h3F0; in353=15'h2F7; in354=15'h7C00; in355=15'h7C00; in356=15'h7DB2; in357=15'h7E72; in358=15'h7E72; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7ED3; in368=15'h3C8; in369=15'h2F7; in370=15'h7CC9; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7FE4; in376=15'h3C0; in377=15'h3F0; in378=15'h64; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h175; in392=15'h3F0; in393=15'h21E; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7E9B; in399=15'h3A8; in400=15'h3F0; in401=15'h2F7; in402=15'h7C70; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h35F; in416=15'h3F8; in417=15'h7F1B; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7D71; in422=15'h2CF; in423=15'h3F8; in424=15'h35F; in425=15'h7DAA; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h1EE; in440=15'h3F0; in441=15'h74; in442=15'h7C00; in443=15'h7C00; in444=15'h7E3A; in445=15'h2F7; in446=15'h3F8; in447=15'h1FE; in448=15'h7DCA; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h44; in464=15'h3F0; in465=15'h2AF; in466=15'h7E7A; in467=15'h7F6B; in468=15'h3C0; in469=15'h3F0; in470=15'h8D; in471=15'h7C60; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7CD1; in489=15'h276; in490=15'h3F8; in491=15'h3F0; in492=15'h3F0; in493=15'h33F; in494=15'h54; in495=15'h7C40; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7CB9; in513=15'hDD; in514=15'h9D; in515=15'h7F03; in516=15'h7CD9; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7DD2; in51=15'h1D6; in52=15'h3F8; in53=15'h196; in54=15'h7F0B; in55=15'h7C48; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7F3B; in72=15'h3C0; in73=15'h3C0; in74=15'h367; in75=15'h3F0; in76=15'h3F8; in77=15'h4; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h3C; in95=15'h3F8; in96=15'h2C7; in97=15'h7EA3; in98=15'h7C60; in99=15'h7F9C; in100=15'h3F8; in101=15'h3C0; in102=15'h7DB2; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7CB1; in118=15'h317; in119=15'h3F8; in120=15'h7E9B; in121=15'h7C00; in122=15'h7C00; in123=15'h7C00; in124=15'h377; in125=15'h3F0; in126=15'h7E72; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7E6A; in143=15'h3F0; in144=15'h33F; in145=15'h7CC1; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'hE5; in150=15'h3F0; in151=15'hC5; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'hFD; in167=15'h3F8; in168=15'h7F1B; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h7DDA; in174=15'h3F8; in175=15'h17D; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h317; in193=15'h3F0; in194=15'h9D; in195=15'h7C18; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7DDA; in200=15'h3F0; in201=15'h29F; in202=15'h7C48; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7DCA; in219=15'h35F; in220=15'h26E; in221=15'h7CD9; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7DDA; in226=15'h3F0; in227=15'h3F0; in228=15'h7C99; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C78; in245=15'h7C40; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7FFC; in251=15'h3F0; in252=15'h388; in253=15'h7C81; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h3F8; in278=15'h3F0; in279=15'h175; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h400; in302=15'h3F8; in303=15'h7E72; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C00; in322=15'h7C00; in323=15'h7C00; in324=15'h7EDB; in325=15'h3F8; in326=15'h3A0; in327=15'h7D51; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C68; in349=15'h2AF; in350=15'h3F8; in351=15'h12D; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C99; in372=15'h7E32; in373=15'hD5; in374=15'h3F0; in375=15'h3F8; in376=15'h23E; in377=15'h7E2A; in378=15'h7C18; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7FCC; in395=15'h2F7; in396=15'h3F0; in397=15'h3F0; in398=15'h3F0; in399=15'h3F8; in400=15'h3F0; in401=15'h3F0; in402=15'h95; in403=15'h7DE2; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7F63; in417=15'h33F; in418=15'h400; in419=15'h3F8; in420=15'h3F8; in421=15'h3F8; in422=15'h3F8; in423=15'h226; in424=15'h2F7; in425=15'h3F8; in426=15'h3F8; in427=15'h3F8; in428=15'h19E; in429=15'h226; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h357; in441=15'h3F0; in442=15'h1D6; in443=15'h246; in444=15'h3F0; in445=15'h3D8; in446=15'h7FCC; in447=15'h7C00; in448=15'h7C91; in449=15'h7F5B; in450=15'h1E6; in451=15'h34F; in452=15'h357; in453=15'h2FF; in454=15'h7CF1; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7DBA; in464=15'h3C0; in465=15'h3F0; in466=15'h307; in467=15'h3F0; in468=15'h3F0; in469=15'h7FA4; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C30; in489=15'h35F; in490=15'h3F0; in491=15'h3F8; in492=15'h3F0; in493=15'h12D; in494=15'h7C10; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7E2A; in513=15'h337; in514=15'h33F; in515=15'h7F7B; in516=15'h7C91; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7D9A; in75=15'h7E6A; in76=15'h7E6A; in77=15'h7FDC; in78=15'h7E6A; in79=15'h1BE; in80=15'h1CE; in81=15'h7DE2; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C10; in96=15'h7EE3; in97=15'h2C7; in98=15'h3A8; in99=15'h3F8; in100=15'h3F8; in101=15'h3F8; in102=15'h3F8; in103=15'h3F8; in104=15'h3F8; in105=15'h216; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7E52; in120=15'h3F8; in121=15'h3F8; in122=15'h3F8; in123=15'h3F8; in124=15'h3F8; in125=15'h3F8; in126=15'h3F8; in127=15'h3F8; in128=15'h3F8; in129=15'h3F8; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h11D; in145=15'h3F8; in146=15'h3F8; in147=15'h3F8; in148=15'h3F8; in149=15'h1CE; in150=15'h3F8; in151=15'h3F8; in152=15'h3F8; in153=15'h3F8; in154=15'h3F8; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7E02; in169=15'h3A8; in170=15'h6C; in171=15'h7DFA; in172=15'h7CD9; in173=15'h7CE9; in174=15'h3F8; in175=15'h3F8; in176=15'h3F8; in177=15'h2EF; in178=15'h7D51; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7D41; in199=15'h7FB4; in200=15'h3F8; in201=15'h3F8; in202=15'h31F; in203=15'h7F3B; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'hC; in224=15'h3A0; in225=15'h3F8; in226=15'h3F8; in227=15'h2DF; in228=15'h7CE9; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C10; in245=15'h7D41; in246=15'h125; in247=15'h1DE; in248=15'h3C8; in249=15'h3F8; in250=15'h3F8; in251=15'h2BF; in252=15'h7CF9; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7EBB; in272=15'h3F8; in273=15'h3F8; in274=15'h3F8; in275=15'h3F8; in276=15'h3F8; in277=15'h3A0; in278=15'h7D79; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7FF4; in296=15'h3F8; in297=15'h3F8; in298=15'h3F8; in299=15'h3F8; in300=15'h3F8; in301=15'h3F8; in302=15'h2D7; in303=15'h7F7B; in304=15'h7C10; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C38; in313=15'h7C18; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7FF4; in320=15'h3F8; in321=15'h3F8; in322=15'h3F0; in323=15'h34F; in324=15'h3D8; in325=15'h3F8; in326=15'h3F8; in327=15'h3F8; in328=15'h19E; in329=15'h7EFB; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7D29; in337=15'h7E6A; in338=15'h7F53; in339=15'h7CC9; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7D59; in345=15'h7EBB; in346=15'h7EBB; in347=15'h7E7A; in348=15'h7C00; in349=15'h7E32; in350=15'h1F6; in351=15'h21E; in352=15'h3B0; in353=15'h3F8; in354=15'h1C6; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C78; in363=15'h115; in364=15'h317; in365=15'h165; in366=15'h7C58; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7C00; in376=15'h7CD1; in377=15'h1B6; in378=15'h3F8; in379=15'h390; in380=15'h7CF9; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7F33; in388=15'hE5; in389=15'h3F8; in390=15'h390; in391=15'h7FA4; in392=15'h7C38; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7C18; in400=15'h196; in401=15'h3F8; in402=15'h3F8; in403=15'h17D; in404=15'h7C10; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7E1A; in413=15'h297; in414=15'h3F8; in415=15'h3F8; in416=15'h206; in417=15'h7FCC; in418=15'h7E12; in419=15'h7E12; in420=15'h7FD4; in421=15'h175; in422=15'h175; in423=15'h1B6; in424=15'h400; in425=15'h3F8; in426=15'hF5; in427=15'h7CC1; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C70; in438=15'h34F; in439=15'h3F8; in440=15'h3F8; in441=15'h3F8; in442=15'h3F8; in443=15'h3F8; in444=15'h3F8; in445=15'h3F8; in446=15'h3F8; in447=15'h3F8; in448=15'h3F8; in449=15'h7E72; in450=15'h7C99; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C70; in463=15'h2F7; in464=15'h3C0; in465=15'h3F8; in466=15'h3F8; in467=15'h3F8; in468=15'h3F8; in469=15'h3F8; in470=15'h327; in471=15'h7F53; in472=15'h7C28; in473=15'h7C08; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7DD2; in490=15'h4; in491=15'h1C6; in492=15'h1C6; in493=15'h7E93; in494=15'h7E62; in495=15'h7C78; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7E9B; in51=15'h34; in52=15'h3F0; in53=15'h3F0; in54=15'h400; in55=15'h7FFC; in56=15'h7C68; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7F63; in72=15'h3C8; in73=15'h3E8; in74=15'h3E8; in75=15'h3E8; in76=15'h3F0; in77=15'h3E8; in78=15'hC5; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7F73; in95=15'h3B0; in96=15'h3E8; in97=15'h3E8; in98=15'h22E; in99=15'hF5; in100=15'h266; in101=15'h3E8; in102=15'hF5; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7E22; in118=15'h3A8; in119=15'h3E8; in120=15'h3E8; in121=15'h1DE; in122=15'h7C89; in123=15'h7C00; in124=15'h7E9B; in125=15'h3C8; in126=15'h7FAC; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7E8B; in143=15'h3E8; in144=15'h3E8; in145=15'h33F; in146=15'h7D61; in147=15'h7C00; in148=15'h7C00; in149=15'h7C00; in150=15'h7D92; in151=15'h7C30; in152=15'h7C00; in153=15'h7C91; in154=15'h4C; in155=15'h7DCA; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7CA9; in167=15'h1CE; in168=15'h3E8; in169=15'h3E8; in170=15'h226; in171=15'h7CB9; in172=15'h7C00; in173=15'h7C00; in174=15'h7C00; in175=15'h7C00; in176=15'h7C00; in177=15'h7DAA; in178=15'h377; in179=15'h390; in180=15'h7F3B; in181=15'h7CB9; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7DCA; in194=15'h390; in195=15'h3E8; in196=15'h3E8; in197=15'h7FFC; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7C78; in202=15'h7D49; in203=15'h95; in204=15'h33F; in205=15'h3E8; in206=15'h3E8; in207=15'h7F53; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7F0B; in221=15'h3A0; in222=15'h3E8; in223=15'h3C0; in224=15'h7ED3; in225=15'h7CD9; in226=15'h7CD9; in227=15'h1A6; in228=15'h3E8; in229=15'h3E8; in230=15'h3E8; in231=15'h3E8; in232=15'h35F; in233=15'h7EFB; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7F03; in247=15'h3E8; in248=15'h3E8; in249=15'h3E8; in250=15'h3F0; in251=15'h3E8; in252=15'h3E8; in253=15'h3E8; in254=15'h3E8; in255=15'h398; in256=15'h9D; in257=15'h7D39; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7CE9; in273=15'hC5; in274=15'h3E8; in275=15'h3E8; in276=15'h3E8; in277=15'h3F0; in278=15'h3E8; in279=15'h3E8; in280=15'h3E8; in281=15'h95; in282=15'h7CF9; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7F33; in295=15'hDD; in296=15'h3F0; in297=15'h3F0; in298=15'h3F0; in299=15'h3F0; in300=15'h3F0; in301=15'h400; in302=15'h5C; in303=15'h2C; in304=15'h7CA9; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7D41; in318=15'h32F; in319=15'h3E8; in320=15'h3E8; in321=15'h35F; in322=15'hE5; in323=15'h3E8; in324=15'h3E8; in325=15'h3F0; in326=15'h7C68; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7D41; in342=15'h2F7; in343=15'h3E8; in344=15'h3E8; in345=15'h1BE; in346=15'h7E02; in347=15'h7C18; in348=15'hED; in349=15'h3E8; in350=15'h3F0; in351=15'h24; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7F5B; in367=15'h3E8; in368=15'h3E8; in369=15'hCD; in370=15'h7C58; in371=15'h7C00; in372=15'h7C00; in373=15'h95; in374=15'h3E8; in375=15'h3F0; in376=15'h35F; in377=15'h7CB1; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7F5B; in391=15'h3E8; in392=15'h3E8; in393=15'h7DAA; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h95; in398=15'h3E8; in399=15'h3F0; in400=15'h307; in401=15'h7C99; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7F5B; in415=15'h3E8; in416=15'h3E8; in417=15'h7DAA; in418=15'h7C00; in419=15'h7C00; in420=15'h7C30; in421=15'h14D; in422=15'h3E8; in423=15'h3F0; in424=15'h7FB4; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7F5B; in439=15'h3E8; in440=15'h3E8; in441=15'h7E52; in442=15'h7C00; in443=15'h7C00; in444=15'h7CD9; in445=15'h3E8; in446=15'h3E8; in447=15'h3F0; in448=15'h7C68; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7F03; in463=15'h3D0; in464=15'h3E8; in465=15'h31F; in466=15'h105; in467=15'h105; in468=15'h14D; in469=15'h3E8; in470=15'h3E8; in471=15'h18E; in472=15'h7C28; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h85; in489=15'h3D8; in490=15'h3E8; in491=15'h3E8; in492=15'h3E8; in493=15'h3E8; in494=15'h3E8; in495=15'h3B0; in496=15'h7DC2; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7F2B; in513=15'hD5; in514=15'h3E8; in515=15'h3E8; in516=15'h3E8; in517=15'h3E8; in518=15'h7FBC; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7E02; in75=15'h256; in76=15'h3F0; in77=15'h3F0; in78=15'h3F0; in79=15'h3F0; in80=15'h4; in81=15'h7C48; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C89; in98=15'h20E; in99=15'h3F0; in100=15'h3E8; in101=15'h3E8; in102=15'h3E8; in103=15'h3E8; in104=15'h3F0; in105=15'h216; in106=15'h7E0A; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h186; in122=15'h3E8; in123=15'h3F0; in124=15'h3E8; in125=15'h3E8; in126=15'h3E8; in127=15'h1EE; in128=15'h3F0; in129=15'h3E8; in130=15'h1BE; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7CD1; in146=15'h307; in147=15'h3E8; in148=15'h3F0; in149=15'h3E8; in150=15'h3E8; in151=15'h186; in152=15'h7C20; in153=15'h7FAC; in154=15'h3E8; in155=15'h388; in156=15'h7D29; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7CB1; in169=15'h26E; in170=15'h3E8; in171=15'h3E8; in172=15'h3A0; in173=15'h7E02; in174=15'h7CB1; in175=15'h7C70; in176=15'h7C00; in177=15'h7C18; in178=15'h14D; in179=15'h3E8; in180=15'h206; in181=15'h7C58; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C18; in194=15'h155; in195=15'h3F0; in196=15'h3F0; in197=15'h3A0; in198=15'h7F53; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h115; in205=15'h3F0; in206=15'h3F0; in207=15'h7CB9; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7FB4; in220=15'h3E8; in221=15'h3E8; in222=15'h3E8; in223=15'h7FAC; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h10D; in231=15'h3E8; in232=15'h3E8; in233=15'h7CB1; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7E02; in244=15'h3F0; in245=15'h3E8; in246=15'h3E8; in247=15'hCD; in248=15'h7C30; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h10D; in256=15'h3E8; in257=15'h31F; in258=15'h7C81; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h337; in271=15'h3F0; in272=15'h3E8; in273=15'h31F; in274=15'h7CE9; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C48; in282=15'h216; in283=15'h3E8; in284=15'h7FBC; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h44; in294=15'h3D8; in295=15'h3F0; in296=15'h297; in297=15'h7C81; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h7C00; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h4; in306=15'h3E8; in307=15'h1EE; in308=15'h7C20; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7E8B; in317=15'h3F0; in318=15'h3F0; in319=15'h3E8; in320=15'h3C; in321=15'h7C00; in322=15'h7C00; in323=15'h7C00; in324=15'h7C00; in325=15'h7C00; in326=15'h7C00; in327=15'h7C00; in328=15'h7E02; in329=15'h400; in330=15'h3F0; in331=15'h16D; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7CF1; in341=15'h22E; in342=15'h3E8; in343=15'h3E8; in344=15'hED; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7C00; in350=15'h7C00; in351=15'h7C00; in352=15'h7E8B; in353=15'h25E; in354=15'h3F0; in355=15'h256; in356=15'h7CC9; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h10D; in366=15'h3E8; in367=15'h3E8; in368=15'h3E8; in369=15'h7EA3; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7C00; in376=15'h7D9A; in377=15'h2E7; in378=15'h3E8; in379=15'h26E; in380=15'h7CC9; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h10D; in390=15'h3E8; in391=15'h3E8; in392=15'h297; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7E8B; in400=15'h388; in401=15'h3E8; in402=15'h3E8; in403=15'h7CA9; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7CB1; in413=15'h3A8; in414=15'h3E8; in415=15'h3E8; in416=15'h7D01; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7FFC; in423=15'h3A8; in424=15'h3E8; in425=15'h3E8; in426=15'h7EFB; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7CC1; in437=15'h3F0; in438=15'h3F0; in439=15'h3F0; in440=15'h7CB9; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7F94; in445=15'h3A0; in446=15'h400; in447=15'h3F0; in448=15'h367; in449=15'h7EF3; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7D69; in461=15'h3E8; in462=15'h3E8; in463=15'h20E; in464=15'h7C40; in465=15'h7C00; in466=15'h7D9A; in467=15'h10D; in468=15'h367; in469=15'h3E8; in470=15'h3D0; in471=15'h1CE; in472=15'h7CC9; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7DBA; in486=15'h3E8; in487=15'h3E8; in488=15'h1CE; in489=15'h7E32; in490=15'h1CE; in491=15'h327; in492=15'h3E8; in493=15'h3E8; in494=15'h3E8; in495=15'h7F9C; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C78; in509=15'h2DF; in510=15'h3E8; in511=15'h3E8; in512=15'h3E8; in513=15'h3F0; in514=15'h3E8; in515=15'h3E8; in516=15'h186; in517=15'h7F63; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7D21; in533=15'h4C; in534=15'h347; in535=15'h3E8; in536=15'h3F0; in537=15'h196; in538=15'h7DB2; in539=15'h7C20; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7D09; in96=15'h186; in97=15'h307; in98=15'h13D; in99=15'h13D; in100=15'h8D; in101=15'h7C40; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7F33; in118=15'h22E; in119=15'h3D0; in120=15'h3F8; in121=15'h3F8; in122=15'h400; in123=15'h3F8; in124=15'h3F8; in125=15'h236; in126=15'h7D71; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7EEB; in142=15'h3E0; in143=15'h3F8; in144=15'h3F8; in145=15'h3F8; in146=15'h29F; in147=15'h20E; in148=15'h206; in149=15'h327; in150=15'h3F8; in151=15'h16D; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h1C; in166=15'h3F8; in167=15'h11D; in168=15'h7CD1; in169=15'h7CD1; in170=15'h7C40; in171=15'h7C00; in172=15'h7C00; in173=15'h7E3A; in174=15'h3F8; in175=15'h297; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7E7A; in192=15'hDD; in193=15'h7C40; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7DF2; in200=15'h3F8; in201=15'h30F; in202=15'h7C78; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7DF2; in226=15'h3F8; in227=15'h297; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7DF2; in251=15'h3F8; in252=15'h297; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h7DF2; in278=15'h3F8; in279=15'h297; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h4; in302=15'h3F8; in303=15'h186; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C00; in322=15'h7C00; in323=15'h7C00; in324=15'h7C00; in325=15'h36F; in326=15'h3F8; in327=15'h7FDC; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7F13; in350=15'h3F8; in351=15'h377; in352=15'h7CC1; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7CB1; in374=15'h2BF; in375=15'h3F8; in376=15'h18E; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7F2B; in398=15'h3F8; in399=15'h3F8; in400=15'h7DF2; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C99; in421=15'h2BF; in422=15'h3F8; in423=15'h236; in424=15'h7C18; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7F43; in445=15'h400; in446=15'h390; in447=15'h7F1B; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7CA1; in468=15'h388; in469=15'h3F8; in470=15'h1BE; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h44; in493=15'h3F8; in494=15'h3F8; in495=15'h7E5A; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C68; in515=15'h347; in516=15'h3F8; in517=15'h3D0; in518=15'h7C40; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h1C6; in539=15'h3F8; in540=15'h26E; in541=15'h7C20; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'hD5; in560=15'h3F8; in561=15'h3F8; in562=15'h7E2A; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7D19; in56=15'h35F; in57=15'h1B6; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C38; in77=15'h125; in78=15'h3F8; in79=15'h21E; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7C00; in100=15'h7CC9; in101=15'h3F8; in102=15'h3F8; in103=15'h7E32; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h7C81; in124=15'hC5; in125=15'h3F8; in126=15'h226; in127=15'h7C20; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7EEB; in149=15'h3F8; in150=15'h3F8; in151=15'h7FD4; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7CD1; in172=15'h2BF; in173=15'h3F8; in174=15'h3E8; in175=15'h7D71; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7FDC; in198=15'h3F8; in199=15'h3F8; in200=15'h175; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C30; in223=15'h216; in224=15'h3F8; in225=15'h3C0; in226=15'h7DCA; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7E6A; in248=15'h3F8; in249=15'h3F8; in250=15'h19E; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h357; in275=15'h3F8; in276=15'h3F8; in277=15'h7DBA; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7D01; in298=15'h390; in299=15'h3F8; in300=15'h1AE; in301=15'h7C20; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C; in322=15'h3F8; in323=15'h3F8; in324=15'h7F5B; in325=15'h7C00; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7D09; in346=15'h35F; in347=15'h3F8; in348=15'h2D7; in349=15'h7C99; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7D92; in371=15'h3F8; in372=15'h3F8; in373=15'h7F8C; in374=15'h7C00; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C10; in394=15'h125; in395=15'h3F8; in396=15'h3B8; in397=15'h7D59; in398=15'h7C00; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7EB3; in418=15'h3F8; in419=15'h3F8; in420=15'h297; in421=15'h7C00; in422=15'h7C00; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h125; in442=15'h3F8; in443=15'h3F8; in444=15'h7EB3; in445=15'h7C00; in446=15'h7C00; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7D71; in465=15'h3A0; in466=15'h3F8; in467=15'h3F8; in468=15'h7CA9; in469=15'h7C00; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7E93; in490=15'h3F8; in491=15'h3F8; in492=15'h20E; in493=15'h7C38; in494=15'h7C00; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7D79; in513=15'h3A0; in514=15'h357; in515=15'h7D92; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7CB9; in77=15'h2A7; in78=15'h2FF; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7CE1; in99=15'h7FBC; in100=15'h297; in101=15'h3F8; in102=15'h3F8; in103=15'h7F03; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7D01; in121=15'h7F84; in122=15'h2A7; in123=15'h3F8; in124=15'h3F8; in125=15'h3F8; in126=15'h3F8; in127=15'h7F13; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7D21; in144=15'h2AF; in145=15'h390; in146=15'h3F8; in147=15'h3F8; in148=15'h3F8; in149=15'h1AE; in150=15'h2E7; in151=15'h307; in152=15'h7C40; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7D21; in167=15'h2D7; in168=15'h3F8; in169=15'h3F8; in170=15'h3F8; in171=15'h1AE; in172=15'hC; in173=15'h7C40; in174=15'h155; in175=15'h3E0; in176=15'h337; in177=15'hC5; in178=15'h7D59; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7D21; in192=15'hB5; in193=15'h3F8; in194=15'h3F8; in195=15'h327; in196=15'h7DF2; in197=15'h7C40; in198=15'h7C00; in199=15'h7C00; in200=15'h7D51; in201=15'h2F7; in202=15'h3F8; in203=15'h3F8; in204=15'h7F7B; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7D21; in217=15'h2D7; in218=15'h3F8; in219=15'h3F8; in220=15'h1C6; in221=15'h7DB2; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7E72; in227=15'h390; in228=15'h3F8; in229=15'h3C8; in230=15'h7E52; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7D19; in241=15'h2DF; in242=15'h3F8; in243=15'h3F8; in244=15'h7C; in245=15'h7C40; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C89; in250=15'h155; in251=15'h388; in252=15'h3F8; in253=15'h3F8; in254=15'h7FFC; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7F84; in268=15'h3F8; in269=15'h3F8; in270=15'h27E; in271=15'h7C99; in272=15'h7DE2; in273=15'h7E4A; in274=15'h7E4A; in275=15'h155; in276=15'h2B7; in277=15'h3F8; in278=15'h3F8; in279=15'h3F8; in280=15'h226; in281=15'h7CA9; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7CD1; in292=15'h388; in293=15'h3F8; in294=15'h3F8; in295=15'h26E; in296=15'h3A8; in297=15'h3F8; in298=15'h400; in299=15'h3F8; in300=15'h3F8; in301=15'h3F8; in302=15'h3F8; in303=15'h32F; in304=15'h7CB9; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7F94; in317=15'h3D0; in318=15'h3F8; in319=15'h3F8; in320=15'h3F8; in321=15'h3F8; in322=15'h3F8; in323=15'h3F8; in324=15'h3F8; in325=15'h3F8; in326=15'h3F8; in327=15'h1FE; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7F9C; in343=15'h256; in344=15'h256; in345=15'h256; in346=15'h256; in347=15'h7F2B; in348=15'h287; in349=15'h3F8; in350=15'h3F8; in351=15'h3B8; in352=15'h7E42; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7D71; in373=15'h35F; in374=15'h3F8; in375=15'h400; in376=15'h7FEC; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7EBB; in397=15'h3F8; in398=15'h3F8; in399=15'h3C0; in400=15'h7E42; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7D79; in420=15'h357; in421=15'h3F8; in422=15'h3F8; in423=15'h287; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7EB3; in444=15'h400; in445=15'h3F8; in446=15'h3D0; in447=15'h7FC4; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h25E; in468=15'h400; in469=15'h3F8; in470=15'h256; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h25E; in493=15'h3F8; in494=15'h3F8; in495=15'h4C; in496=15'h7C58; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h25E; in516=15'h400; in517=15'h3F8; in518=15'h3F8; in519=15'h287; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h3C; in539=15'h400; in540=15'h3F8; in541=15'h31F; in542=15'h7F33; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7FDC; in76=15'h3F0; in77=15'h3F0; in78=15'h7EA3; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7E83; in99=15'h3F0; in100=15'h3E8; in101=15'h367; in102=15'h7CA9; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7F9C; in123=15'h3F0; in124=15'h3E8; in125=15'h2F7; in126=15'h7C00; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7F94; in147=15'h37F; in148=15'h3F0; in149=15'h3E8; in150=15'h7F23; in151=15'h7C00; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h14D; in171=15'h3E8; in172=15'h3F0; in173=15'h3E8; in174=15'h7CA9; in175=15'h7C00; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7CB1; in196=15'h3F0; in197=15'h3F0; in198=15'h400; in199=15'h145; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7CB1; in222=15'h3E8; in223=15'h3E8; in224=15'h3F0; in225=15'h145; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7E5A; in247=15'h3E8; in248=15'h3E8; in249=15'h3F0; in250=15'h7E3A; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7FFC; in274=15'h3E8; in275=15'h3E8; in276=15'h3F0; in277=15'h7DFA; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7FFC; in298=15'h3E8; in299=15'h3E8; in300=15'h3F0; in301=15'h7DFA; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h1EE; in322=15'h3F0; in323=15'h3F0; in324=15'h337; in325=15'h7CD9; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7E02; in346=15'h3C0; in347=15'h3E8; in348=15'h3E8; in349=15'h29F; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7EAB; in371=15'h3E8; in372=15'h3E8; in373=15'h3E8; in374=15'h7F9C; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7CE1; in395=15'h37F; in396=15'h3E8; in397=15'h3E8; in398=15'h7D19; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'hFD; in419=15'h3D0; in420=15'h3E8; in421=15'h3E8; in422=15'h7C00; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h1FE; in443=15'h3F0; in444=15'h3F0; in445=15'h3F0; in446=15'h7C00; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h1F6; in467=15'h3E8; in468=15'h3E8; in469=15'h2CF; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h1F6; in492=15'h3E8; in493=15'h3E8; in494=15'h9D; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7F1B; in515=15'h3C0; in516=15'h3E8; in517=15'h9D; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h85; in539=15'h317; in540=15'h7D51; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7C00; in100=15'h7C00; in101=15'h7C00; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C28; in120=15'h7DDA; in121=15'hAD; in122=15'h33F; in123=15'h400; in124=15'h3F8; in125=15'h3F8; in126=15'h377; in127=15'h7FBC; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7CE1; in144=15'h12D; in145=15'h3F0; in146=15'h3F0; in147=15'h3F0; in148=15'h3F8; in149=15'h3F0; in150=15'h3F0; in151=15'h3F0; in152=15'h3F0; in153=15'h7C40; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'hE5; in168=15'h3F0; in169=15'h3F0; in170=15'h3F0; in171=15'h3F0; in172=15'h3F8; in173=15'h2F7; in174=15'h3F0; in175=15'h3F0; in176=15'h3F0; in177=15'h7F13; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7DAA; in193=15'h3F8; in194=15'h3F0; in195=15'h3F0; in196=15'h24E; in197=15'h7E7A; in198=15'h7C99; in199=15'h7E9B; in200=15'h3F0; in201=15'h3F0; in202=15'h3F0; in203=15'h7D69; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7F13; in219=15'h3F8; in220=15'h3F0; in221=15'h7FB4; in222=15'h7C28; in223=15'h7D31; in224=15'h7FCC; in225=15'h2F7; in226=15'h3F0; in227=15'h3F0; in228=15'h3F0; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7F1B; in244=15'h400; in245=15'h3F8; in246=15'h3F8; in247=15'h3F8; in248=15'h3F8; in249=15'h400; in250=15'h3F8; in251=15'h3F8; in252=15'h3F8; in253=15'h33F; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C78; in271=15'h24E; in272=15'h3F0; in273=15'h3F0; in274=15'h3F0; in275=15'h3F0; in276=15'h3F8; in277=15'h3F0; in278=15'h3F0; in279=15'h3D8; in280=15'h7F53; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C91; in296=15'h7FDC; in297=15'h32F; in298=15'h3F0; in299=15'h3F0; in300=15'h3F8; in301=15'h3F0; in302=15'h3F0; in303=15'h2AF; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C68; in322=15'h7C99; in323=15'h7C99; in324=15'h196; in325=15'h3F0; in326=15'h3F0; in327=15'h10D; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h3F8; in350=15'h3F0; in351=15'h2F7; in352=15'h7D11; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7FCC; in374=15'h400; in375=15'h3F8; in376=15'h17D; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h21E; in398=15'h3F8; in399=15'h3F0; in400=15'h7EE3; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7DD2; in421=15'h35F; in422=15'h3F8; in423=15'h37F; in424=15'h7CC1; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h1EE; in445=15'h3F0; in446=15'h3F8; in447=15'h74; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7F1B; in468=15'h3C8; in469=15'h3F0; in470=15'h33F; in471=15'h7D71; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7D59; in492=15'h3F8; in493=15'h3F8; in494=15'h3F8; in495=15'h3C; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h115; in515=15'h3F0; in516=15'h3F0; in517=15'h27E; in518=15'h7C78; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7D49; in537=15'h390; in538=15'h3F0; in539=15'h3F0; in540=15'h7EC3; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7DDA; in558=15'h3F0; in559=15'h3F0; in560=15'h33F; in561=15'h7CD9; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C70; in580=15'hA5; in581=15'h3F0; in582=15'h7F2B; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7C00; in100=15'h7C00; in101=15'h7C00; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7FF4; in119=15'h266; in120=15'h3F0; in121=15'h3F0; in122=15'h3F0; in123=15'h398; in124=15'h6C; in125=15'h7CF9; in126=15'h7C00; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7DFA; in142=15'h14D; in143=15'h3A0; in144=15'h3F0; in145=15'h3E8; in146=15'h3E8; in147=15'h256; in148=15'h25E; in149=15'h3E8; in150=15'h7F53; in151=15'h7CD1; in152=15'hED; in153=15'h7C99; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7D31; in164=15'h9D; in165=15'h357; in166=15'h3E8; in167=15'h18E; in168=15'h7F53; in169=15'h7DC2; in170=15'h7DC2; in171=15'h7C30; in172=15'h7C38; in173=15'h7DC2; in174=15'h7C68; in175=15'h246; in176=15'h3F0; in177=15'h15D; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h2AF; in190=15'h3F0; in191=15'h3E8; in192=15'h125; in193=15'h7C78; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7E62; in201=15'h3D0; in202=15'h3F0; in203=15'h8D; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7D82; in215=15'h390; in216=15'h37F; in217=15'h7FEC; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7D01; in226=15'h32F; in227=15'h3F0; in228=15'h37F; in229=15'h7D31; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h105; in240=15'h3E8; in241=15'h7F8C; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C38; in250=15'hB5; in251=15'h3E8; in252=15'h3E8; in253=15'hB5; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7F73; in267=15'h3E8; in268=15'h7F8C; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'hD5; in277=15'h3E8; in278=15'h3E8; in279=15'h3E8; in280=15'h7F8C; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7EAB; in291=15'h3E8; in292=15'h11D; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7C00; in299=15'hBD; in300=15'h3F0; in301=15'h3E8; in302=15'h3E8; in303=15'h3E8; in304=15'h7F8C; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h2B7; in316=15'h400; in317=15'hCD; in318=15'h7C99; in319=15'h7CD1; in320=15'h7CE9; in321=15'h7F43; in322=15'h32F; in323=15'h3F0; in324=15'h317; in325=15'h85; in326=15'h3F0; in327=15'h3F0; in328=15'h7D9A; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7D31; in341=15'h327; in342=15'h3E8; in343=15'h307; in344=15'h3A0; in345=15'h3F0; in346=15'h3E8; in347=15'h3E8; in348=15'hBD; in349=15'h7D31; in350=15'h7DCA; in351=15'h3E8; in352=15'h3E8; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7F43; in367=15'h3E8; in368=15'h3E8; in369=15'h2B7; in370=15'h145; in371=15'h74; in372=15'h7DC2; in373=15'h7C30; in374=15'h7C00; in375=15'h7DCA; in376=15'h3E8; in377=15'h125; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C20; in391=15'h7CE1; in392=15'h7FA4; in393=15'h7CE1; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7F5B; in400=15'h3E8; in401=15'h5C; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7C00; in423=15'h155; in424=15'h3F0; in425=15'h64; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7C00; in445=15'h7C00; in446=15'h7C00; in447=15'h14D; in448=15'h3E8; in449=15'h5C; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7C00; in468=15'h7C00; in469=15'h7C00; in470=15'h7C00; in471=15'h14D; in472=15'h3E8; in473=15'h5C; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'h7C00; in496=15'h14D; in497=15'h3E8; in498=15'h5C; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7DCA; in520=15'h3F0; in521=15'h7CE1; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7DCA; in543=15'h3E8; in544=15'h7DAA; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7DCA; in564=15'h3E8; in565=15'h5C; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7D01; in586=15'h327; in587=15'h5C; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'hCD; in68=15'h276; in69=15'h7C30; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C40; in76=15'h7E0A; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h44; in92=15'h3F8; in93=15'h7C58; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7F94; in100=15'h25E; in101=15'h7E0A; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h155; in116=15'h3F8; in117=15'h7D21; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h7D29; in124=15'h3E0; in125=15'h1C; in126=15'h7C00; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h287; in141=15'h3F8; in142=15'hC; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h3D8; in150=15'h3C0; in151=15'h7E12; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7DDA; in164=15'h3B8; in165=15'h3F8; in166=15'h7D09; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h3D8; in174=15'h3F8; in175=15'h1CE; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h18E; in190=15'h3F8; in191=15'h3F8; in192=15'h7C58; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h3D8; in200=15'h3F8; in201=15'h27E; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h1F6; in216=15'h3F8; in217=15'h256; in218=15'h7C30; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C18; in225=15'h3D8; in226=15'h3F8; in227=15'h337; in228=15'h7D31; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7CF9; in240=15'h317; in241=15'h3F8; in242=15'hED; in243=15'h7C10; in244=15'h7C00; in245=15'h7C20; in246=15'h7CC1; in247=15'h7CC1; in248=15'h7E2A; in249=15'h206; in250=15'h3F8; in251=15'h3F8; in252=15'h3F8; in253=15'h21E; in254=15'h7C28; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7DB2; in267=15'h3F8; in268=15'h3F8; in269=15'h3F8; in270=15'h125; in271=15'h105; in272=15'h186; in273=15'h3F8; in274=15'h3F8; in275=15'h3F8; in276=15'h3F8; in277=15'h3F8; in278=15'h3F8; in279=15'h3F8; in280=15'h2AF; in281=15'h7CA1; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C89; in291=15'h28F; in292=15'h3F8; in293=15'h3F8; in294=15'h3F8; in295=15'h3F8; in296=15'h3F8; in297=15'h400; in298=15'h3F8; in299=15'h400; in300=15'h3F8; in301=15'h3F8; in302=15'h400; in303=15'h3F8; in304=15'h7F53; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7E72; in316=15'h266; in317=15'h3F8; in318=15'h3F8; in319=15'h3F8; in320=15'h3F8; in321=15'h3F8; in322=15'h3F8; in323=15'h3F8; in324=15'h3F8; in325=15'h3F8; in326=15'h3F8; in327=15'h347; in328=15'h7D31; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C78; in342=15'h7D49; in343=15'hD5; in344=15'hA5; in345=15'h1C; in346=15'h347; in347=15'hFD; in348=15'hFD; in349=15'h7F5B; in350=15'h3D8; in351=15'h3F8; in352=15'h3F8; in353=15'h7E3A; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C20; in371=15'h7C91; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7ECB; in376=15'h3F8; in377=15'h3F8; in378=15'h7E3A; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7C60; in400=15'h3F8; in401=15'h3F8; in402=15'h7E3A; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7C00; in423=15'h7C60; in424=15'h400; in425=15'h3F8; in426=15'h7EAB; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7C00; in445=15'h7C00; in446=15'h7C00; in447=15'h7C28; in448=15'h1CE; in449=15'h3F8; in450=15'h347; in451=15'h7D19; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7C00; in468=15'h7C00; in469=15'h7C00; in470=15'h7C00; in471=15'h7C00; in472=15'hA5; in473=15'h3F8; in474=15'h3F8; in475=15'h7DAA; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'h7C00; in496=15'h7C00; in497=15'hA5; in498=15'h3F8; in499=15'h3F8; in500=15'h7DAA; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'hA5; in521=15'h3F8; in522=15'h3F8; in523=15'h7DAA; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7D31; in544=15'h3F8; in545=15'h307; in546=15'h7CE1; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C70; in66=15'h7D59; in67=15'h7C; in68=15'h7F4B; in69=15'h5C; in70=15'h3F0; in71=15'h3F0; in72=15'hED; in73=15'h388; in74=15'h2E7; in75=15'h297; in76=15'h7C; in77=15'h7C; in78=15'h1B6; in79=15'h9D; in80=15'h7C68; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7EFB; in89=15'h1DE; in90=15'h3E8; in91=15'h3E8; in92=15'h3E8; in93=15'h3E8; in94=15'h3E8; in95=15'h3E8; in96=15'h3E8; in97=15'h3F0; in98=15'h3E8; in99=15'h3E8; in100=15'h3E8; in101=15'h3E8; in102=15'h3E8; in103=15'h3E8; in104=15'h1D6; in105=15'h7C91; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7DCA; in112=15'h276; in113=15'h3E8; in114=15'h3E8; in115=15'h3E8; in116=15'h3E8; in117=15'h3E8; in118=15'h3E8; in119=15'h3E8; in120=15'h3E8; in121=15'h388; in122=15'h19E; in123=15'h3E8; in124=15'h3E8; in125=15'h3E8; in126=15'h3E8; in127=15'h3E8; in128=15'h3E8; in129=15'hE5; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h2C; in137=15'h3E8; in138=15'h3E8; in139=15'h390; in140=15'h337; in141=15'h7C; in142=15'h7E22; in143=15'h7C50; in144=15'h7C50; in145=15'h7C50; in146=15'h7C48; in147=15'h7C18; in148=15'h7C50; in149=15'h7C60; in150=15'h186; in151=15'h3E8; in152=15'h3E8; in153=15'h3E8; in154=15'h17D; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7CD1; in161=15'h22E; in162=15'h7F5B; in163=15'h7D51; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7E12; in173=15'h16D; in174=15'h3E8; in175=15'h3E8; in176=15'h3E8; in177=15'h2FF; in178=15'h7DEA; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7CC1; in198=15'h24E; in199=15'h3E8; in200=15'h3E8; in201=15'h3E8; in202=15'h3C8; in203=15'h7EC3; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7CA9; in223=15'hDD; in224=15'h3E8; in225=15'h3E8; in226=15'h3E8; in227=15'h3C0; in228=15'h7EC3; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C70; in246=15'h7D69; in247=15'h297; in248=15'h3E8; in249=15'h3E8; in250=15'h3C8; in251=15'h1C6; in252=15'h7DC2; in253=15'h7C48; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7E72; in273=15'h3E8; in274=15'h3F0; in275=15'h3E8; in276=15'h3E8; in277=15'h337; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7D39; in296=15'h337; in297=15'h3E8; in298=15'h3F0; in299=15'h3E8; in300=15'h3E8; in301=15'h7D31; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7D69; in320=15'h3F0; in321=15'h3F0; in322=15'h400; in323=15'h3F0; in324=15'h3F0; in325=15'h226; in326=15'h7E02; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7D09; in345=15'h276; in346=15'h3E8; in347=15'h3F0; in348=15'h3E8; in349=15'h3E8; in350=15'h3E8; in351=15'h367; in352=15'h186; in353=15'h7D61; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C70; in371=15'h7D61; in372=15'h7F53; in373=15'h19E; in374=15'h3E8; in375=15'h3E8; in376=15'h3E8; in377=15'h3E8; in378=15'h31F; in379=15'h7E93; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C18; in398=15'h7DB2; in399=15'h196; in400=15'h3B0; in401=15'h3E8; in402=15'h3E8; in403=15'h3E0; in404=15'h7E4A; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7C00; in423=15'h7C00; in424=15'h7E32; in425=15'h32F; in426=15'h3E8; in427=15'h3E8; in428=15'h17D; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7D39; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7C00; in445=15'h7C00; in446=15'h7C00; in447=15'h7EAB; in448=15'h165; in449=15'h3E8; in450=15'h3E8; in451=15'h3E8; in452=15'h256; in453=15'h7C60; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C40; in463=15'h20E; in464=15'h196; in465=15'h7FD4; in466=15'h7FD4; in467=15'h2CF; in468=15'h155; in469=15'hB5; in470=15'h33F; in471=15'h3E0; in472=15'h3E8; in473=15'h3E8; in474=15'h3E8; in475=15'h3E8; in476=15'h18E; in477=15'h7C18; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'hDD; in488=15'h3A0; in489=15'h3E8; in490=15'h3E8; in491=15'h3E8; in492=15'h3E8; in493=15'h3F0; in494=15'h3E8; in495=15'h3E8; in496=15'h3E8; in497=15'h3E8; in498=15'h3E8; in499=15'h3E8; in500=15'h3B0; in501=15'h7DB2; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7CE9; in511=15'h7FAC; in512=15'h3E8; in513=15'h3E8; in514=15'h3E8; in515=15'h3E8; in516=15'h3F0; in517=15'h3E8; in518=15'h3E8; in519=15'h3E8; in520=15'h3E8; in521=15'h3E8; in522=15'h4; in523=15'h7DB2; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C60; in535=15'h2C; in536=15'h10D; in537=15'h266; in538=15'h3E8; in539=15'h26E; in540=15'h3E8; in541=15'h28F; in542=15'h74; in543=15'h74; in544=15'h7DC2; in545=15'h7C18; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C58; in97=15'h7D9A; in98=15'hC5; in99=15'hC5; in100=15'h7EE3; in101=15'h7CF9; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7D49; in120=15'h16D; in121=15'h3E8; in122=15'h3F0; in123=15'h3E8; in124=15'h3F0; in125=15'h347; in126=15'h7E93; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7F33; in145=15'h3F8; in146=15'h3F0; in147=15'h3F8; in148=15'h3F0; in149=15'h3F8; in150=15'h3F0; in151=15'h357; in152=15'h7D9A; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h1BE; in169=15'h3F0; in170=15'h3E8; in171=15'h3F0; in172=15'h3E8; in173=15'h3F0; in174=15'h3E8; in175=15'h3F0; in176=15'h347; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7E93; in195=15'h3F8; in196=15'h3F0; in197=15'h3F8; in198=15'h3F0; in199=15'h307; in200=15'h3A0; in201=15'h3F8; in202=15'h3F0; in203=15'h11D; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7E3A; in222=15'hBD; in223=15'hBD; in224=15'h7E32; in225=15'h7CA1; in226=15'h25E; in227=15'h3F0; in228=15'h3E8; in229=15'h25E; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C58; in251=15'h2AF; in252=15'h3F8; in253=15'h3F0; in254=15'h3F8; in255=15'h7D92; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7D49; in269=15'h7F33; in270=15'h74; in271=15'h25E; in272=15'h25E; in273=15'h1BE; in274=15'h7DEA; in275=15'h7C00; in276=15'h7C00; in277=15'h16D; in278=15'h3E8; in279=15'h3F0; in280=15'h3E8; in281=15'h3F0; in282=15'h7D92; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7CA9; in291=15'h16D; in292=15'h3F0; in293=15'h3F8; in294=15'h3F0; in295=15'h3F8; in296=15'h3F0; in297=15'h3F8; in298=15'h3F0; in299=15'h3F8; in300=15'h3F0; in301=15'h3F8; in302=15'h3F0; in303=15'h3F8; in304=15'h3F0; in305=15'h3F8; in306=15'h7D92; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7CA9; in314=15'h25E; in315=15'h3F0; in316=15'h3E8; in317=15'h3F0; in318=15'h3E8; in319=15'h3F0; in320=15'h3E8; in321=15'h3F0; in322=15'h3E8; in323=15'h3F0; in324=15'h3E8; in325=15'h3F0; in326=15'h3E8; in327=15'h3F0; in328=15'h3E8; in329=15'h34F; in330=15'h7CF1; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'hC5; in339=15'h3F0; in340=15'h3F8; in341=15'h3F0; in342=15'h3F8; in343=15'h3F0; in344=15'h3F8; in345=15'h3F0; in346=15'h3F8; in347=15'h3F0; in348=15'h3F8; in349=15'h3F0; in350=15'h3F8; in351=15'h3F0; in352=15'h3F8; in353=15'h3F0; in354=15'h2B7; in355=15'h7C50; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h34F; in364=15'h3E8; in365=15'h3F0; in366=15'h3E8; in367=15'h3F0; in368=15'h3E8; in369=15'h3F0; in370=15'h3E8; in371=15'h3F0; in372=15'h3E8; in373=15'h3F0; in374=15'h3E8; in375=15'h3F0; in376=15'h3E8; in377=15'h3F0; in378=15'h3E8; in379=15'h3F0; in380=15'h2A7; in381=15'h7E93; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h357; in388=15'h3F0; in389=15'h3F8; in390=15'h3F0; in391=15'h3F8; in392=15'h3F0; in393=15'h3F8; in394=15'h3F0; in395=15'h3F8; in396=15'h3F0; in397=15'h3F8; in398=15'h165; in399=15'h7F33; in400=15'h1BE; in401=15'h357; in402=15'h3F0; in403=15'h3F8; in404=15'h3F0; in405=15'h357; in406=15'h7D9A; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7F84; in412=15'h3E8; in413=15'h3F0; in414=15'h3E8; in415=15'h3F0; in416=15'h3E8; in417=15'h3F0; in418=15'h3E8; in419=15'h34F; in420=15'hBD; in421=15'h7D92; in422=15'h7C50; in423=15'h7C00; in424=15'h7C00; in425=15'h7CF1; in426=15'h1C; in427=15'h165; in428=15'h3E8; in429=15'h3F0; in430=15'h347; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7FDC; in437=15'h357; in438=15'h3F0; in439=15'h400; in440=15'h2AF; in441=15'h1BE; in442=15'h7DEA; in443=15'h7C00; in444=15'h7C00; in445=15'h7C00; in446=15'h7C00; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7E93; in453=15'h25E; in454=15'h7FD4; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7CF1; in462=15'h7D92; in463=15'h7D92; in464=15'h7C50; in465=15'h7C00; in466=15'h7C00; in467=15'h7C00; in468=15'h7C00; in469=15'h7C00; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C40; in54=15'h7F8C; in55=15'h3E8; in56=15'h3E8; in57=15'h3E8; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7F8C; in76=15'h3D8; in77=15'h3D8; in78=15'h3D8; in79=15'h3D8; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h3E8; in100=15'h3D8; in101=15'h3D8; in102=15'h3D8; in103=15'h3D8; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h3E8; in124=15'h3D8; in125=15'h3D8; in126=15'h3D8; in127=15'h3D8; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h18E; in148=15'h3E8; in149=15'h3D8; in150=15'h3D8; in151=15'h3D8; in152=15'h7E52; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7CE9; in171=15'h2DF; in172=15'h3F8; in173=15'h3E8; in174=15'h3E8; in175=15'h307; in176=15'h7D11; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7D59; in196=15'h226; in197=15'h3D8; in198=15'h3E8; in199=15'h3D8; in200=15'h287; in201=15'h7DBA; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7FFC; in222=15'h3D8; in223=15'h3D8; in224=15'h3E8; in225=15'h3D8; in226=15'h7FEC; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7FFC; in247=15'h3D8; in248=15'h3D8; in249=15'h3E8; in250=15'h3D8; in251=15'h7FEC; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7E3A; in273=15'h337; in274=15'h3D8; in275=15'h3D8; in276=15'h3E8; in277=15'h3D8; in278=15'h7FEC; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C40; in296=15'h7F8C; in297=15'h3E8; in298=15'h3E8; in299=15'h3E8; in300=15'h400; in301=15'h13D; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7F8C; in320=15'h3D8; in321=15'h3D8; in322=15'h3D8; in323=15'h3D8; in324=15'h377; in325=15'h7F7B; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h3E8; in345=15'h3D8; in346=15'h3D8; in347=15'h3D8; in348=15'h3D8; in349=15'h7F4B; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h3E8; in370=15'h3D8; in371=15'h3D8; in372=15'h3D8; in373=15'h3D8; in374=15'h7C00; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h3E8; in394=15'h3D8; in395=15'h3D8; in396=15'h3D8; in397=15'h3D8; in398=15'h7C00; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h3F8; in418=15'h3E8; in419=15'h3E8; in420=15'h3E8; in421=15'h3E8; in422=15'h7C00; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h3E8; in442=15'h3D8; in443=15'h3D8; in444=15'h3D8; in445=15'h3D8; in446=15'h7EB3; in447=15'h7EAB; in448=15'h7D51; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h3E8; in466=15'h3D8; in467=15'h3D8; in468=15'h3D8; in469=15'h3D8; in470=15'h3E8; in471=15'h287; in472=15'h7DF2; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h3E8; in491=15'h3D8; in492=15'h3D8; in493=15'h3D8; in494=15'h3D8; in495=15'h307; in496=15'h7DBA; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7E62; in514=15'h3D8; in515=15'h3D8; in516=15'h3D8; in517=15'h3D8; in518=15'h7D11; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7CD1; in51=15'h6C; in52=15'h1FE; in53=15'h32F; in54=15'h3F0; in55=15'h186; in56=15'h7DFA; in57=15'h7C50; in58=15'h7C20; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7DCA; in72=15'h20E; in73=15'h3F0; in74=15'h3E8; in75=15'h3E8; in76=15'h3E8; in77=15'h17D; in78=15'hB5; in79=15'h22E; in80=15'h4; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7DFA; in95=15'h1C; in96=15'h3A0; in97=15'h276; in98=15'h44; in99=15'h256; in100=15'h3E8; in101=15'h7F23; in102=15'h1C; in103=15'h1D6; in104=15'h3A0; in105=15'h7ECB; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7CD1; in118=15'h1DE; in119=15'h7C00; in120=15'h7CC9; in121=15'h7C68; in122=15'h7F5B; in123=15'h125; in124=15'h7D41; in125=15'h7C00; in126=15'h7C38; in127=15'h7C30; in128=15'h30F; in129=15'h317; in130=15'h7D31; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h11D; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7F43; in147=15'h3F0; in148=15'h7E2A; in149=15'h7C00; in150=15'h7C00; in151=15'h7C00; in152=15'h7C00; in153=15'h24E; in154=15'h400; in155=15'h22E; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7F8C; in167=15'h7C00; in168=15'h7C00; in169=15'h7D9A; in170=15'h3F0; in171=15'h3E8; in172=15'h26E; in173=15'h7C68; in174=15'h7C00; in175=15'h7C00; in176=15'h7C00; in177=15'h7CD1; in178=15'h3F0; in179=15'h226; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7CC9; in193=15'h7C00; in194=15'h7C00; in195=15'h30F; in196=15'h3F0; in197=15'h34F; in198=15'h7DF2; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7F8C; in204=15'h3F0; in205=15'h226; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h30F; in222=15'h25E; in223=15'h8D; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C68; in230=15'h7F3B; in231=15'h226; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7CB9; in246=15'h266; in247=15'h7F94; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7D49; in256=15'h22E; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7D31; in272=15'h7F3B; in273=15'h7C48; in274=15'h7D31; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h2C7; in283=15'h226; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h85; in296=15'h1AE; in297=15'h7C68; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h7C00; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7ECB; in306=15'h3F0; in307=15'h226; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h186; in319=15'h2D7; in320=15'h7D59; in321=15'h7C00; in322=15'h7C00; in323=15'h7C00; in324=15'h7C00; in325=15'h7C00; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h2AF; in330=15'h327; in331=15'h7CB1; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C50; in342=15'h32F; in343=15'h37F; in344=15'h7EC3; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7C00; in350=15'h7C00; in351=15'h7C00; in352=15'h7D01; in353=15'h196; in354=15'h3F0; in355=15'h317; in356=15'h7D31; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7EAB; in367=15'h3E8; in368=15'h246; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7C00; in376=15'h7D01; in377=15'h7FF4; in378=15'h327; in379=15'h31F; in380=15'h7D31; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7EAB; in391=15'h3E8; in392=15'h7F8C; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7C00; in400=15'h196; in401=15'h3E8; in402=15'h3E8; in403=15'h7DA2; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h34; in415=15'h3E8; in416=15'h2AF; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7ECB; in423=15'h2AF; in424=15'h3F0; in425=15'h3E8; in426=15'h2B7; in427=15'h7C78; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7D01; in438=15'h32F; in439=15'h3F0; in440=15'h7F94; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7F43; in445=15'h25E; in446=15'h3F0; in447=15'h3F0; in448=15'h186; in449=15'h7EC3; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7DCA; in462=15'h3E8; in463=15'h3E8; in464=15'h27E; in465=15'h14D; in466=15'h14D; in467=15'h7FBC; in468=15'h3F0; in469=15'h3E8; in470=15'h3E8; in471=15'hBD; in472=15'h7D31; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7D31; in487=15'h357; in488=15'h3E8; in489=15'h3F0; in490=15'h3E8; in491=15'h3E8; in492=15'h3E8; in493=15'h3F0; in494=15'h226; in495=15'h14; in496=15'h7C30; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7CB1; in511=15'h327; in512=15'h3F0; in513=15'h3E8; in514=15'h3E8; in515=15'hBD; in516=15'h7E72; in517=15'h7C48; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7CE9; in75=15'h390; in76=15'h7E62; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7D61; in99=15'h3F8; in100=15'h2C; in101=15'h7C00; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7E2A; in123=15'h3F8; in124=15'h2C; in125=15'h7C00; in126=15'h7C00; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h14; in148=15'h3F8; in149=15'h2C; in150=15'h7C00; in151=15'h7C00; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h14; in172=15'h3F8; in173=15'h7DAA; in174=15'h7C00; in175=15'h7C00; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h14; in198=15'h347; in199=15'h7CA1; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h14; in224=15'h2BF; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h14; in249=15'h5C; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h95; in276=15'hC; in277=15'h7C00; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7C00; in299=15'h2C7; in300=15'hC; in301=15'h7C00; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C00; in322=15'h7C00; in323=15'h2C7; in324=15'hC; in325=15'h7C00; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h2C7; in349=15'h7DDA; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'hED; in374=15'h7E9B; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h2C7; in398=15'hC; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7CA9; in421=15'h34F; in422=15'hC; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7D82; in445=15'h3F8; in446=15'hC; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h7C00; in468=15'h7F84; in469=15'h3F8; in470=15'hC; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h34; in494=15'h3F8; in495=15'hC; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7F43; in517=15'h3F8; in518=15'h7E2A; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7D82; in540=15'h297; in541=15'h7CE9; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h400; in52=15'h3F0; in53=15'hAD; in54=15'h7D79; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7D51; in73=15'h3F0; in74=15'h3E8; in75=15'h3E8; in76=15'h7F63; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7D79; in96=15'h2EF; in97=15'h3F0; in98=15'h3E8; in99=15'h3E8; in100=15'h4; in101=15'h7C00; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h1AE; in120=15'h3E8; in121=15'h3F0; in122=15'h3E8; in123=15'h3E8; in124=15'h3E8; in125=15'h7C00; in126=15'h7C00; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7FBC; in145=15'h3E8; in146=15'h3F0; in147=15'h3E8; in148=15'h3E8; in149=15'h3E8; in150=15'h7C00; in151=15'h7C00; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7CD1; in169=15'h2EF; in170=15'h3F0; in171=15'h3E8; in172=15'h3E8; in173=15'h3E8; in174=15'h7C00; in175=15'h7C00; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h85; in196=15'h3F0; in197=15'h3E8; in198=15'h3E8; in199=15'hA5; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h85; in222=15'h3F0; in223=15'h3E8; in224=15'h3E8; in225=15'h7F63; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7CA9; in246=15'h27E; in247=15'h400; in248=15'h3F0; in249=15'h3F0; in250=15'h1FE; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h85; in274=15'h3F0; in275=15'h3E8; in276=15'h3E8; in277=15'h347; in278=15'h7D51; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h85; in298=15'h3F0; in299=15'h3E8; in300=15'h3E8; in301=15'h3E8; in302=15'h2F7; in303=15'h7CC9; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7DF2; in322=15'h3F0; in323=15'h3E8; in324=15'h3E8; in325=15'h3E8; in326=15'h1FE; in327=15'h7C78; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h8D; in347=15'h400; in348=15'h3F0; in349=15'h3F0; in350=15'h3F0; in351=15'h8D; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7F43; in372=15'h3F0; in373=15'h3E8; in374=15'h3E8; in375=15'h3E8; in376=15'h186; in377=15'h7C50; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7CA9; in396=15'h3F0; in397=15'h3E8; in398=15'h3E8; in399=15'h3E8; in400=15'h36F; in401=15'h7CF1; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h85; in420=15'h3F0; in421=15'h3E8; in422=15'h3E8; in423=15'h3E8; in424=15'h85; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C81; in443=15'h1FE; in444=15'h400; in445=15'h3F0; in446=15'h3F0; in447=15'h3F0; in448=15'h206; in449=15'h7C78; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C28; in467=15'hFD; in468=15'h3F0; in469=15'h3E8; in470=15'h3E8; in471=15'h3E8; in472=15'h2F7; in473=15'h7CC9; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7D49; in493=15'h3F0; in494=15'h3E8; in495=15'h3E8; in496=15'h33F; in497=15'h7D49; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h3F0; in517=15'h3E8; in518=15'hA5; in519=15'h7D71; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h236; in57=15'h317; in58=15'h7EB3; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7CE9; in71=15'h7EB3; in72=15'h155; in73=15'h155; in74=15'h7F94; in75=15'h7CE9; in76=15'h7C00; in77=15'h7EB3; in78=15'h400; in79=15'h400; in80=15'h400; in81=15'h7EB3; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7EB3; in94=15'h317; in95=15'h400; in96=15'h400; in97=15'h317; in98=15'h400; in99=15'h236; in100=15'h7CE9; in101=15'h7EB3; in102=15'h400; in103=15'h155; in104=15'h400; in105=15'h400; in106=15'h7CE9; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h155; in117=15'h400; in118=15'h317; in119=15'h7F94; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h6C; in124=15'h6C; in125=15'h7DCA; in126=15'h7CE9; in127=15'h7C00; in128=15'h7F94; in129=15'h400; in130=15'h236; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h155; in141=15'h400; in142=15'h317; in143=15'h7EB3; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h7EB3; in150=15'h7EB3; in151=15'h7C00; in152=15'h7C00; in153=15'h7C00; in154=15'h236; in155=15'h400; in156=15'h7DCA; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h6C; in164=15'h400; in165=15'h400; in166=15'h7EB3; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h7C00; in174=15'h7DCA; in175=15'h7C00; in176=15'h7C00; in177=15'h7C00; in178=15'h155; in179=15'h400; in180=15'h7EB3; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7CE9; in189=15'h400; in190=15'h400; in191=15'h6C; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h155; in205=15'h400; in206=15'h6C; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7EB3; in215=15'h400; in216=15'h317; in217=15'h7CE9; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h155; in231=15'h400; in232=15'h155; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h155; in240=15'h400; in241=15'h6C; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h155; in256=15'h400; in257=15'h155; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7DCA; in266=15'h400; in267=15'h317; in268=15'h7CE9; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7CE9; in282=15'h400; in283=15'h400; in284=15'h7F94; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7EB3; in290=15'h400; in291=15'h155; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h7C00; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7F94; in306=15'h400; in307=15'h236; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7F94; in314=15'h400; in315=15'h6C; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C00; in322=15'h7C00; in323=15'h7C00; in324=15'h7C00; in325=15'h7C00; in326=15'h7C00; in327=15'h7C00; in328=15'h7CE9; in329=15'h317; in330=15'h400; in331=15'h155; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h155; in339=15'h400; in340=15'h7EB3; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7C00; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7F94; in354=15'h400; in355=15'h400; in356=15'h7EB3; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h6C; in364=15'h400; in365=15'h7EB3; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7C00; in376=15'h7C00; in377=15'h7EB3; in378=15'h400; in379=15'h400; in380=15'h6C; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h6C; in388=15'h400; in389=15'h7EB3; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7C00; in399=15'h7C00; in400=15'h155; in401=15'h400; in402=15'h400; in403=15'h317; in404=15'h7CE9; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7EB3; in412=15'h400; in413=15'h7F94; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C00; in422=15'h7CE9; in423=15'h155; in424=15'h400; in425=15'h400; in426=15'h317; in427=15'h7DCA; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7DCA; in436=15'h400; in437=15'h155; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7DCA; in445=15'h7F94; in446=15'h400; in447=15'h400; in448=15'h400; in449=15'h236; in450=15'h7DCA; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h6C; in461=15'h400; in462=15'h155; in463=15'h7EB3; in464=15'h7EB3; in465=15'h7EB3; in466=15'h6C; in467=15'h236; in468=15'h400; in469=15'h400; in470=15'h400; in471=15'h400; in472=15'h6C; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7CE9; in486=15'h317; in487=15'h400; in488=15'h400; in489=15'h400; in490=15'h400; in491=15'h400; in492=15'h400; in493=15'h400; in494=15'h400; in495=15'h155; in496=15'h7CE9; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7CE9; in510=15'h7F94; in511=15'h236; in512=15'h400; in513=15'h400; in514=15'h400; in515=15'h317; in516=15'h6C; in517=15'h7CE9; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7EDB; in100=15'h287; in101=15'h3F8; in102=15'h3F8; in103=15'hAD; in104=15'h7C60; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7D59; in122=15'h24E; in123=15'h3F8; in124=15'h3F0; in125=15'h3F0; in126=15'h37F; in127=15'h3F0; in128=15'h14; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7EBB; in146=15'h3B0; in147=15'h3F0; in148=15'h3F8; in149=15'h21E; in150=15'h7E8B; in151=15'h7D69; in152=15'h1B6; in153=15'h7E9B; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7CD1; in169=15'h3C0; in170=15'h3F0; in171=15'h3F0; in172=15'h1AE; in173=15'h7C50; in174=15'h1C; in175=15'h3F0; in176=15'h7F84; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C58; in194=15'h2AF; in195=15'h3F0; in196=15'h3F0; in197=15'hA5; in198=15'h7C38; in199=15'h7DAA; in200=15'h3D0; in201=15'h3F0; in202=15'h23E; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7DEA; in220=15'h3F0; in221=15'h3F0; in222=15'h1AE; in223=15'h7C60; in224=15'h7C60; in225=15'h17D; in226=15'h3F0; in227=15'h3F0; in228=15'h7FDC; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C81; in244=15'h216; in245=15'h3F0; in246=15'h3F0; in247=15'h7D29; in248=15'h7C00; in249=15'h1FE; in250=15'h3F0; in251=15'h3F0; in252=15'h23E; in253=15'h7C30; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7D82; in271=15'h3F0; in272=15'h3F0; in273=15'h74; in274=15'h7EFB; in275=15'h2E7; in276=15'h3F8; in277=15'h3F0; in278=15'h3E0; in279=15'h7E2A; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7D82; in295=15'h3F0; in296=15'h3F0; in297=15'h33F; in298=15'h3C0; in299=15'h3F0; in300=15'h3F8; in301=15'h3F0; in302=15'h11D; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7D82; in319=15'h3F0; in320=15'h3F0; in321=15'h3F0; in322=15'h3F0; in323=15'h3F0; in324=15'h3F8; in325=15'h3F0; in326=15'h7F9C; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7FE4; in345=15'h3F8; in346=15'h3F8; in347=15'h3F8; in348=15'h3F8; in349=15'h400; in350=15'hE5; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C18; in370=15'h7CE1; in371=15'h226; in372=15'h3F0; in373=15'h3F0; in374=15'h3A8; in375=15'h7E2A; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h307; in396=15'h3F0; in397=15'h3F0; in398=15'h7F9C; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7EAB; in419=15'h3D8; in420=15'h3F0; in421=15'h3F0; in422=15'h7D01; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C91; in442=15'h3C0; in443=15'h3F0; in444=15'h3F0; in445=15'h7F94; in446=15'h7C00; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7F03; in466=15'h3F0; in467=15'h3F0; in468=15'h3F0; in469=15'h7E0A; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C81; in490=15'h216; in491=15'h3F0; in492=15'h3F0; in493=15'h3F0; in494=15'h7E0A; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7D82; in513=15'h3F0; in514=15'h3F0; in515=15'h3F0; in516=15'h7E7A; in517=15'h7C18; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7EEB; in536=15'h3F0; in537=15'h3F0; in538=15'h216; in539=15'h7C30; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7E42; in557=15'h3F0; in558=15'h2EF; in559=15'h7CF1; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C00; in76=15'h7C00; in77=15'h7C00; in78=15'h7C00; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7C00; in100=15'h7C00; in101=15'h7C00; in102=15'h7C00; in103=15'h7C00; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h7C00; in124=15'h7C00; in125=15'h7C00; in126=15'h7C00; in127=15'h7C00; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C68; in147=15'h7D41; in148=15'h7D41; in149=15'h7D41; in150=15'h7D41; in151=15'h7D41; in152=15'h7D41; in153=15'h7D41; in154=15'h7D41; in155=15'h7EAB; in156=15'h44; in157=15'hBD; in158=15'h2DF; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7FA4; in171=15'h3F0; in172=15'h3F0; in173=15'h3F8; in174=15'h3F0; in175=15'h3F0; in176=15'h3F0; in177=15'h3F0; in178=15'h3F8; in179=15'h3F0; in180=15'h3F0; in181=15'h115; in182=15'h7F03; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7F03; in196=15'h307; in197=15'h3F8; in198=15'h33F; in199=15'h2D7; in200=15'h21E; in201=15'h21E; in202=15'h3D0; in203=15'h3F8; in204=15'h226; in205=15'hB5; in206=15'h7E22; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7E4A; in221=15'h347; in222=15'h3F0; in223=15'h175; in224=15'h7CC1; in225=15'h7C78; in226=15'h7C00; in227=15'h7C00; in228=15'h7D21; in229=15'h7D39; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C68; in244=15'h7FA4; in245=15'h307; in246=15'h3F0; in247=15'h3F0; in248=15'h7D8A; in249=15'h7CF9; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7E6A; in271=15'h3F0; in272=15'h3F8; in273=15'h3F0; in274=15'h3F0; in275=15'h35F; in276=15'h390; in277=15'h7F9C; in278=15'h7CA9; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'hC5; in295=15'h3F0; in296=15'h3F8; in297=15'h3F0; in298=15'h3F0; in299=15'h3F0; in300=15'h3F0; in301=15'h3F8; in302=15'h1AE; in303=15'h7CF1; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7E22; in319=15'h21E; in320=15'h16D; in321=15'h7EDB; in322=15'h7C00; in323=15'h7C00; in324=15'h7F1B; in325=15'h400; in326=15'h3B8; in327=15'h7F6B; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7C78; in350=15'h11D; in351=15'h3F0; in352=15'h390; in353=15'h7CC1; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7D8A; in366=15'h7E4A; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7FFC; in376=15'h3F0; in377=15'h3F0; in378=15'h7E7A; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h3B8; in390=15'h3A8; in391=15'h7F5B; in392=15'h7C91; in393=15'h7C00; in394=15'h7C00; in395=15'h7C20; in396=15'h7D41; in397=15'h85; in398=15'h357; in399=15'h3B8; in400=15'h3F0; in401=15'h21E; in402=15'h7C81; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h196; in414=15'h3F0; in415=15'h3F0; in416=15'h2EF; in417=15'h21E; in418=15'hF5; in419=15'h23E; in420=15'h3F0; in421=15'h3F0; in422=15'h3F0; in423=15'h3F8; in424=15'h36F; in425=15'h7C91; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7DEA; in438=15'h74; in439=15'h367; in440=15'h3F8; in441=15'h3F8; in442=15'h400; in443=15'h3F8; in444=15'h3F8; in445=15'h2F7; in446=15'hED; in447=15'h7E62; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7DCA; in464=15'h3C; in465=15'h3C; in466=15'h44; in467=15'h4; in468=15'h7D39; in469=15'h7C91; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C00; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C28; in71=15'h7FDC; in72=15'h2C; in73=15'h34; in74=15'h2C; in75=15'h2C; in76=15'hE5; in77=15'h226; in78=15'h3F8; in79=15'h3F8; in80=15'h25E; in81=15'h7C60; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7EC3; in95=15'h3E0; in96=15'h3F0; in97=15'h398; in98=15'h32F; in99=15'h32F; in100=15'h32F; in101=15'h32F; in102=15'h3C8; in103=15'h3F0; in104=15'hE5; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7EC3; in120=15'h7F03; in121=15'h7D71; in122=15'h7C00; in123=15'h7C00; in124=15'h7C00; in125=15'h7DC2; in126=15'h33F; in127=15'h3F0; in128=15'hE5; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h7D09; in150=15'h337; in151=15'h3F0; in152=15'h3F0; in153=15'h2C; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C30; in172=15'h7DEA; in173=15'hDD; in174=15'h3F0; in175=15'h367; in176=15'hC5; in177=15'h7C50; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7D39; in197=15'h7EDB; in198=15'h3F0; in199=15'h3F0; in200=15'h3F0; in201=15'h367; in202=15'h7D29; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7D29; in221=15'h7C; in222=15'h347; in223=15'h3F0; in224=15'h3F0; in225=15'h3F0; in226=15'h3F0; in227=15'h3F0; in228=15'h95; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'hDD; in246=15'h3F0; in247=15'h3F8; in248=15'h3F0; in249=15'h3F0; in250=15'h1E6; in251=15'h7E32; in252=15'h256; in253=15'h390; in254=15'h165; in255=15'h7C48; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7D01; in270=15'h7F73; in271=15'h2AF; in272=15'h3E0; in273=15'h3F0; in274=15'h22E; in275=15'h85; in276=15'h7E2A; in277=15'h7C40; in278=15'h7CD9; in279=15'h2DF; in280=15'h3F0; in281=15'h29F; in282=15'h7C70; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7E4A; in294=15'h3F0; in295=15'h3F0; in296=15'h24E; in297=15'h7E5A; in298=15'h7C30; in299=15'h7C00; in300=15'h7C00; in301=15'h7C00; in302=15'h7DEA; in303=15'h3F0; in304=15'h3F0; in305=15'hE5; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7E32; in318=15'h85; in319=15'h7E5A; in320=15'h7C00; in321=15'h7C00; in322=15'h7C00; in323=15'h7C00; in324=15'h7C00; in325=15'h7C00; in326=15'h7FC4; in327=15'h3F8; in328=15'h3F8; in329=15'h7D51; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C00; in346=15'h7C00; in347=15'h7C00; in348=15'h7C00; in349=15'h7C00; in350=15'h7C00; in351=15'h14; in352=15'h3F0; in353=15'h3B0; in354=15'h7EA3; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7C00; in371=15'h7C00; in372=15'h7C00; in373=15'h7C00; in374=15'h7C00; in375=15'h7F53; in376=15'h317; in377=15'h3F0; in378=15'h7EF3; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7C00; in395=15'h7C00; in396=15'h7C00; in397=15'h7C00; in398=15'h7D82; in399=15'h317; in400=15'h3F0; in401=15'h37F; in402=15'h7D39; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h7C00; in419=15'h7C00; in420=15'h7C00; in421=15'h7C91; in422=15'h317; in423=15'h3F0; in424=15'h307; in425=15'h7E12; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7C00; in442=15'h7C00; in443=15'h7C00; in444=15'h7D69; in445=15'h23E; in446=15'h3F0; in447=15'h3F0; in448=15'h165; in449=15'h7C70; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C48; in460=15'h7D09; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h7C00; in466=15'h7C00; in467=15'h5C; in468=15'h347; in469=15'h3F0; in470=15'h390; in471=15'h7EC3; in472=15'h7C70; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h4; in485=15'h2B7; in486=15'h7D09; in487=15'h7C00; in488=15'h7C00; in489=15'h7E83; in490=15'h7C; in491=15'h2D7; in492=15'h3E8; in493=15'h3F8; in494=15'h1D6; in495=15'h7CF9; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7EF3; in508=15'h3F0; in509=15'h377; in510=15'h337; in511=15'h337; in512=15'h3D0; in513=15'h3F0; in514=15'h3F0; in515=15'h3F0; in516=15'h7E93; in517=15'h7C50; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C10; in531=15'h7EBB; in532=15'hDD; in533=15'h3F0; in534=15'h3F0; in535=15'h3F0; in536=15'h3F0; in537=15'h7C; in538=15'h7C89; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7E93; in55=15'h400; in56=15'h7F53; in57=15'h7C00; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7C08; in76=15'h11D; in77=15'h3F0; in78=15'h85; in79=15'h7C00; in80=15'h7C00; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7C00; in99=15'h7CF9; in100=15'h3F0; in101=15'h3F0; in102=15'h32F; in103=15'h7C99; in104=15'h7C00; in105=15'h7C00; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7C00; in123=15'h7F8C; in124=15'h3F8; in125=15'h20E; in126=15'h7D11; in127=15'h7C20; in128=15'h7C00; in129=15'h7C00; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7E02; in148=15'h377; in149=15'h3F8; in150=15'h54; in151=15'h7C00; in152=15'h7C00; in153=15'h7C00; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h388; in172=15'h3F0; in173=15'h35F; in174=15'h7FDC; in175=15'h7C00; in176=15'h7C00; in177=15'h7C00; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h3D0; in198=15'h3F0; in199=15'h7EF3; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h85; in223=15'h3F0; in224=15'h3F0; in225=15'h7EF3; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7CF9; in247=15'h388; in248=15'h3F0; in249=15'h2A7; in250=15'h7CB1; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7DE2; in274=15'h3F0; in275=15'h3F0; in276=15'hC; in277=15'h7C00; in278=15'h7C00; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h5C; in298=15'h3F0; in299=15'h3F0; in300=15'h7EDB; in301=15'h7C00; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h256; in322=15'h3F8; in323=15'h3F0; in324=15'h7EBB; in325=15'h7C00; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7C30; in346=15'h388; in347=15'h3F0; in348=15'h29F; in349=15'h7C40; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7C00; in370=15'h7EAB; in371=15'h3F0; in372=15'h3F0; in373=15'h25E; in374=15'h7C00; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7C00; in393=15'h7C00; in394=15'h7EFB; in395=15'h3F8; in396=15'h3F8; in397=15'h3A0; in398=15'h7D39; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7C00; in416=15'h7C00; in417=15'h7C00; in418=15'h1C6; in419=15'h3F0; in420=15'h3F0; in421=15'h25E; in422=15'h7C00; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C00; in439=15'h7C00; in440=15'h7C00; in441=15'h7D51; in442=15'h3C8; in443=15'h3F8; in444=15'h3F8; in445=15'h266; in446=15'h7C00; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C00; in463=15'h7C00; in464=15'h7C00; in465=15'h14; in466=15'h3F8; in467=15'h3F0; in468=15'h3F8; in469=15'hC; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7E22; in491=15'h287; in492=15'h3E0; in493=15'h3F8; in494=15'h7D79; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7E1A; in516=15'h337; in517=15'h7C20; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7C00; in52=15'h7C00; in53=15'h7C00; in54=15'h7C00; in55=15'h7C00; in56=15'h7C28; in57=15'h7C58; in58=15'h7C30; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7C00; in71=15'h7C00; in72=15'h7C00; in73=15'h7C00; in74=15'h7C00; in75=15'h7E02; in76=15'h7E0A; in77=15'h7F4B; in78=15'h7FEC; in79=15'h3F0; in80=15'h246; in81=15'h7C99; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'h7C00; in93=15'h7C00; in94=15'h7C00; in95=15'h7C00; in96=15'h7C00; in97=15'h7C00; in98=15'h7EEB; in99=15'h3E0; in100=15'h3F0; in101=15'h3D0; in102=15'h327; in103=15'h34F; in104=15'h3E0; in105=15'hFD; in106=15'h7C48; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h7C00; in117=15'h7C00; in118=15'h7C00; in119=15'h7C00; in120=15'h7C00; in121=15'h7C00; in122=15'h7DEA; in123=15'h18E; in124=15'h18E; in125=15'h7DEA; in126=15'h7D01; in127=15'h7C00; in128=15'h21E; in129=15'h3F0; in130=15'h7D8A; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7C00; in142=15'h7C00; in143=15'h7C00; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h7C00; in150=15'h7C00; in151=15'h7C00; in152=15'h7C00; in153=15'h7D01; in154=15'h26E; in155=15'h7FC4; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h7C00; in174=15'h7C00; in175=15'h7C00; in176=15'h7C00; in177=15'h7C99; in178=15'h10D; in179=15'h7FC4; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h7C00; in200=15'h7C00; in201=15'h7C00; in202=15'h7C00; in203=15'h7F23; in204=15'h1AE; in205=15'h7E02; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7C00; in225=15'h7C00; in226=15'h7C00; in227=15'h7C00; in228=15'h7C00; in229=15'h7C50; in230=15'h9D; in231=15'h7CA1; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C00; in249=15'h7C00; in250=15'h7C00; in251=15'h7C00; in252=15'h7C00; in253=15'h7C00; in254=15'h2EF; in255=15'h7F9C; in256=15'h7C08; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7C00; in276=15'h7C00; in277=15'h7C00; in278=15'h7C00; in279=15'h7D41; in280=15'h7E42; in281=15'h1BE; in282=15'h7D61; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7C00; in299=15'h7C00; in300=15'h7C00; in301=15'h7C00; in302=15'h7D82; in303=15'h7ED3; in304=15'h4; in305=15'h7C58; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C00; in321=15'h7C00; in322=15'h7C18; in323=15'h7C78; in324=15'h7E5A; in325=15'h7FAC; in326=15'h13D; in327=15'h7D11; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7D8A; in345=15'h7E93; in346=15'h7F13; in347=15'h18E; in348=15'h3F0; in349=15'h3F0; in350=15'h3F0; in351=15'h3F0; in352=15'h8D; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C78; in367=15'h7EB3; in368=15'h24; in369=15'h3A8; in370=15'h3F0; in371=15'h2B7; in372=15'h3F0; in373=15'h3F0; in374=15'h3D0; in375=15'h327; in376=15'h1AE; in377=15'h7C81; in378=15'h7C00; in379=15'h7C00; in380=15'h7C00; in381=15'h7C00; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7F33; in390=15'h2A7; in391=15'h3F0; in392=15'h3F0; in393=15'h3F0; in394=15'h3F0; in395=15'h2E7; in396=15'h1CE; in397=15'h206; in398=15'h7F2B; in399=15'h7C00; in400=15'h7C00; in401=15'h7C00; in402=15'h7C00; in403=15'h7C00; in404=15'h7C00; in405=15'h7C00; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h3F8; in414=15'h3F0; in415=15'h3F0; in416=15'h3F0; in417=15'h3F0; in418=15'h367; in419=15'h95; in420=15'h7C50; in421=15'h7C28; in422=15'h7C00; in423=15'h7C00; in424=15'h7C00; in425=15'h7C00; in426=15'h7C00; in427=15'h7C00; in428=15'h7C00; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7D41; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7FF4; in438=15'h377; in439=15'h3F0; in440=15'h29F; in441=15'h14D; in442=15'h7D01; in443=15'h7C00; in444=15'h7C00; in445=15'h7C00; in446=15'h7C00; in447=15'h7C00; in448=15'h7C00; in449=15'h7C00; in450=15'h7C00; in451=15'h7C00; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7C40; in463=15'h7C48; in464=15'h7C28; in465=15'h7C20; in466=15'h7C00; in467=15'h7C00; in468=15'h7C00; in469=15'h7C00; in470=15'h7C00; in471=15'h7C00; in472=15'h7C00; in473=15'h7C00; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7C00; in488=15'h7C00; in489=15'h7C00; in490=15'h7C00; in491=15'h7C00; in492=15'h7C00; in493=15'h7C00; in494=15'h7C00; in495=15'h7C00; in496=15'h7C00; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7C00; in512=15'h7C00; in513=15'h7C00; in514=15'h7C00; in515=15'h7C00; in516=15'h7C00; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
      #50 in1=15'h7C00; in2=15'h7C00; in3=15'h7C00; in4=15'h7C00; in5=15'h7C00; in6=15'h7C00; in7=15'h7C00; in8=15'h7C00; in9=15'h7C00; in10=15'h7C00; in11=15'h7C00; in12=15'h7C00; in13=15'h7C00; in14=15'h7C00; in15=15'h7C00; in16=15'h7C00; in17=15'h7C00; in18=15'h7C00; in19=15'h7C00; in20=15'h7C00; in21=15'h7C00; in22=15'h7C00; in23=15'h7C00; in24=15'h7C00; in25=15'h7C00; in26=15'h7C00; in27=15'h7C00; in28=15'h7C00; in29=15'h7C00; in30=15'h7C00; in31=15'h7C00; in32=15'h7C00; in33=15'h7C00; in34=15'h7C00; in35=15'h7C00; in36=15'h7C00; in37=15'h7C00; in38=15'h7C00; in39=15'h7C00; in40=15'h7C00; in41=15'h7C00; in42=15'h7C00; in43=15'h7C00; in44=15'h7C00; in45=15'h7C00; in46=15'h7C00; in47=15'h7C00; in48=15'h7C00; in49=15'h7C00; in50=15'h7C00; in51=15'h7F23; in52=15'hED; in53=15'h3F8; in54=15'h327; in55=15'h7FEC; in56=15'h7FEC; in57=15'h7F6B; in58=15'h7C00; in59=15'h7C00; in60=15'h7C00; in61=15'h7C00; in62=15'h7C00; in63=15'h7C00; in64=15'h7C00; in65=15'h7C00; in66=15'h7C00; in67=15'h7C00; in68=15'h7C00; in69=15'h7C00; in70=15'h7F43; in71=15'h10D; in72=15'h3C8; in73=15'h3E8; in74=15'h3F0; in75=15'h3F0; in76=15'h3F0; in77=15'h3F0; in78=15'h3F0; in79=15'h3F0; in80=15'hDD; in81=15'h7C00; in82=15'h7C00; in83=15'h7C00; in84=15'h7C00; in85=15'h7C00; in86=15'h7C00; in87=15'h7C00; in88=15'h7C00; in89=15'h7C00; in90=15'h7C00; in91=15'h7C00; in92=15'hED; in93=15'h390; in94=15'h3E8; in95=15'h3F0; in96=15'h3F0; in97=15'h3F0; in98=15'h30F; in99=15'h30F; in100=15'h3F0; in101=15'h3F0; in102=15'h3F0; in103=15'h3F0; in104=15'h377; in105=15'h7D71; in106=15'h7C00; in107=15'h7C00; in108=15'h7C00; in109=15'h7C00; in110=15'h7C00; in111=15'h7C00; in112=15'h7C00; in113=15'h7C00; in114=15'h7C00; in115=15'h7C00; in116=15'h35F; in117=15'h3F0; in118=15'h115; in119=15'h7F53; in120=15'h7C99; in121=15'h7C99; in122=15'h7C70; in123=15'h7C70; in124=15'h7C99; in125=15'h7DEA; in126=15'h3F0; in127=15'h3F0; in128=15'h398; in129=15'h7DEA; in130=15'h7C00; in131=15'h7C00; in132=15'h7C00; in133=15'h7C00; in134=15'h7C00; in135=15'h7C00; in136=15'h7C00; in137=15'h7C00; in138=15'h7C00; in139=15'h7C00; in140=15'h7C00; in141=15'h7CC1; in142=15'h7CC9; in143=15'h7C20; in144=15'h7C00; in145=15'h7C00; in146=15'h7C00; in147=15'h7C00; in148=15'h7C00; in149=15'h7C00; in150=15'h7D71; in151=15'h3F0; in152=15'h3F0; in153=15'h31F; in154=15'h7C00; in155=15'h7C00; in156=15'h7C00; in157=15'h7C00; in158=15'h7C00; in159=15'h7C00; in160=15'h7C00; in161=15'h7C00; in162=15'h7C00; in163=15'h7C00; in164=15'h7C00; in165=15'h7C00; in166=15'h7C00; in167=15'h7C00; in168=15'h7C00; in169=15'h7C00; in170=15'h7C00; in171=15'h7C00; in172=15'h7C00; in173=15'h7C99; in174=15'h1E6; in175=15'h3F0; in176=15'h390; in177=15'h7E7A; in178=15'h7C00; in179=15'h7C00; in180=15'h7C00; in181=15'h7C00; in182=15'h7C00; in183=15'h7C00; in184=15'h7C00; in185=15'h7C00; in186=15'h7C00; in187=15'h7C00; in188=15'h7C00; in189=15'h7C00; in190=15'h7C00; in191=15'h7C00; in192=15'h7C00; in193=15'h7C00; in194=15'h7C00; in195=15'h7C00; in196=15'h7C00; in197=15'h7C00; in198=15'h7C00; in199=15'h11D; in200=15'h3F0; in201=15'h3F0; in202=15'h18E; in203=15'h7C00; in204=15'h7C00; in205=15'h7C00; in206=15'h7C00; in207=15'h7C00; in208=15'h7C00; in209=15'h7C00; in210=15'h7C00; in211=15'h7C00; in212=15'h7C00; in213=15'h7C00; in214=15'h7C00; in215=15'h7C00; in216=15'h7C00; in217=15'h7C00; in218=15'h7C00; in219=15'h7C00; in220=15'h7C00; in221=15'h7C00; in222=15'h7C00; in223=15'h7C00; in224=15'h7D8A; in225=15'h390; in226=15'h3F0; in227=15'h24E; in228=15'h7DFA; in229=15'h7C00; in230=15'h7C00; in231=15'h7C00; in232=15'h7C00; in233=15'h7C00; in234=15'h7C00; in235=15'h7C00; in236=15'h7C00; in237=15'h7C00; in238=15'h7C00; in239=15'h7C00; in240=15'h7C00; in241=15'h7C00; in242=15'h7C00; in243=15'h7C00; in244=15'h7C00; in245=15'h7C00; in246=15'h7C00; in247=15'h7C00; in248=15'h7C99; in249=15'h1AE; in250=15'h3F0; in251=15'h2CF; in252=15'h7C89; in253=15'h7C00; in254=15'h7C00; in255=15'h7C00; in256=15'h7C00; in257=15'h7C00; in258=15'h7C00; in259=15'h7C00; in260=15'h7C00; in261=15'h7C00; in262=15'h7C00; in263=15'h7C00; in264=15'h7C00; in265=15'h7C00; in266=15'h7C00; in267=15'h7C00; in268=15'h7C00; in269=15'h7C00; in270=15'h7C00; in271=15'h7C00; in272=15'h7C00; in273=15'h7C00; in274=15'h7C00; in275=15'h7F23; in276=15'h3F0; in277=15'h388; in278=15'h7EBB; in279=15'h7C00; in280=15'h7C00; in281=15'h7C00; in282=15'h7C00; in283=15'h7C00; in284=15'h7C00; in285=15'h7C00; in286=15'h7C00; in287=15'h7C00; in288=15'h7C00; in289=15'h7C00; in290=15'h7C00; in291=15'h7C00; in292=15'h7C00; in293=15'h7C00; in294=15'h7C00; in295=15'h7C00; in296=15'h7C00; in297=15'h7C00; in298=15'h7EAB; in299=15'h37F; in300=15'h3F0; in301=15'h7F43; in302=15'h7C00; in303=15'h7C00; in304=15'h7C00; in305=15'h7C00; in306=15'h7C00; in307=15'h7C00; in308=15'h7C00; in309=15'h7C00; in310=15'h7C00; in311=15'h7C00; in312=15'h7C00; in313=15'h7C00; in314=15'h7C00; in315=15'h7C00; in316=15'h7C00; in317=15'h7C00; in318=15'h7C00; in319=15'h7C00; in320=15'h7C91; in321=15'h7EEB; in322=15'h37F; in323=15'h3F0; in324=15'h1C6; in325=15'h7CA1; in326=15'h7C00; in327=15'h7C00; in328=15'h7C00; in329=15'h7C00; in330=15'h7C00; in331=15'h7C00; in332=15'h7C00; in333=15'h7C00; in334=15'h7C00; in335=15'h7C00; in336=15'h7C00; in337=15'h7C00; in338=15'h7C00; in339=15'h7C00; in340=15'h7C00; in341=15'h7C00; in342=15'h7C00; in343=15'h7C00; in344=15'h7C00; in345=15'h7F6B; in346=15'h3F0; in347=15'h3F0; in348=15'h287; in349=15'h7CA1; in350=15'h7C00; in351=15'h7C00; in352=15'h7C00; in353=15'h7C00; in354=15'h7C00; in355=15'h7C00; in356=15'h7C00; in357=15'h7C00; in358=15'h7C00; in359=15'h7C00; in360=15'h7C00; in361=15'h7C00; in362=15'h7C00; in363=15'h7C00; in364=15'h7C00; in365=15'h7C00; in366=15'h7C00; in367=15'h7C00; in368=15'h7C00; in369=15'h7E93; in370=15'h390; in371=15'h3F0; in372=15'h1CE; in373=15'h7DFA; in374=15'h7C00; in375=15'h7C00; in376=15'h7C00; in377=15'h7C00; in378=15'h7C00; in379=15'h7C28; in380=15'h7D41; in381=15'h7C89; in382=15'h7C00; in383=15'h7C00; in384=15'h7C00; in385=15'h7C00; in386=15'h7C00; in387=15'h7C00; in388=15'h7C00; in389=15'h7C00; in390=15'h7C00; in391=15'h7C00; in392=15'h7E8B; in393=15'h398; in394=15'h3F0; in395=15'h25E; in396=15'h7C99; in397=15'h7C00; in398=15'h7C00; in399=15'h7C00; in400=15'h7C30; in401=15'h7D09; in402=15'h7FAC; in403=15'h165; in404=15'h390; in405=15'h7D41; in406=15'h7C00; in407=15'h7C00; in408=15'h7C00; in409=15'h7C00; in410=15'h7C00; in411=15'h7C00; in412=15'h7C00; in413=15'h7C00; in414=15'h7C00; in415=15'h7E0A; in416=15'h3A8; in417=15'h3F0; in418=15'h24E; in419=15'h7E1A; in420=15'h7C40; in421=15'h7CD9; in422=15'h7DCA; in423=15'hE5; in424=15'h175; in425=15'h3F0; in426=15'h3F0; in427=15'h307; in428=15'h7ED3; in429=15'h7C00; in430=15'h7C00; in431=15'h7C00; in432=15'h7C00; in433=15'h7C00; in434=15'h7C00; in435=15'h7C00; in436=15'h7C00; in437=15'h7C00; in438=15'h7C48; in439=15'h1BE; in440=15'h3F0; in441=15'h3F0; in442=15'h17D; in443=15'h4; in444=15'h19E; in445=15'h3F0; in446=15'h3F0; in447=15'h3F0; in448=15'h3F0; in449=15'h3D8; in450=15'hAD; in451=15'h7D41; in452=15'h7C00; in453=15'h7C00; in454=15'h7C00; in455=15'h7C00; in456=15'h7C00; in457=15'h7C00; in458=15'h7C00; in459=15'h7C00; in460=15'h7C00; in461=15'h7C00; in462=15'h7F84; in463=15'h3F0; in464=15'h3F0; in465=15'h3F0; in466=15'h3F0; in467=15'h3F0; in468=15'h3F0; in469=15'h3F0; in470=15'h3F0; in471=15'h3A8; in472=15'h2CF; in473=15'h7EEB; in474=15'h7C00; in475=15'h7C00; in476=15'h7C00; in477=15'h7C00; in478=15'h7C00; in479=15'h7C00; in480=15'h7C00; in481=15'h7C00; in482=15'h7C00; in483=15'h7C00; in484=15'h7C00; in485=15'h7C00; in486=15'h7C00; in487=15'h7F6B; in488=15'h3F0; in489=15'h3F0; in490=15'h3F0; in491=15'h3F0; in492=15'h3F0; in493=15'h3C8; in494=15'h2AF; in495=15'h7FAC; in496=15'h7D09; in497=15'h7C00; in498=15'h7C00; in499=15'h7C00; in500=15'h7C00; in501=15'h7C00; in502=15'h7C00; in503=15'h7C00; in504=15'h7C00; in505=15'h7C00; in506=15'h7C00; in507=15'h7C00; in508=15'h7C00; in509=15'h7C00; in510=15'h7C00; in511=15'h7F9C; in512=15'h388; in513=15'h3F0; in514=15'h28F; in515=15'h7FDC; in516=15'h7CC9; in517=15'h7C00; in518=15'h7C00; in519=15'h7C00; in520=15'h7C00; in521=15'h7C00; in522=15'h7C00; in523=15'h7C00; in524=15'h7C00; in525=15'h7C00; in526=15'h7C00; in527=15'h7C00; in528=15'h7C00; in529=15'h7C00; in530=15'h7C00; in531=15'h7C00; in532=15'h7C00; in533=15'h7C00; in534=15'h7C00; in535=15'h7C00; in536=15'h7C00; in537=15'h7C00; in538=15'h7C00; in539=15'h7C00; in540=15'h7C00; in541=15'h7C00; in542=15'h7C00; in543=15'h7C00; in544=15'h7C00; in545=15'h7C00; in546=15'h7C00; in547=15'h7C00; in548=15'h7C00; in549=15'h7C00; in550=15'h7C00; in551=15'h7C00; in552=15'h7C00; in553=15'h7C00; in554=15'h7C00; in555=15'h7C00; in556=15'h7C00; in557=15'h7C00; in558=15'h7C00; in559=15'h7C00; in560=15'h7C00; in561=15'h7C00; in562=15'h7C00; in563=15'h7C00; in564=15'h7C00; in565=15'h7C00; in566=15'h7C00; in567=15'h7C00; in568=15'h7C00; in569=15'h7C00; in570=15'h7C00; in571=15'h7C00; in572=15'h7C00; in573=15'h7C00; in574=15'h7C00; in575=15'h7C00; in576=15'h7C00; in577=15'h7C00; in578=15'h7C00; in579=15'h7C00; in580=15'h7C00; in581=15'h7C00; in582=15'h7C00; in583=15'h7C00; in584=15'h7C00; in585=15'h7C00; in586=15'h7C00; in587=15'h7C00; in588=15'h7C00; in589=15'h7C00; in590=15'h7C00; in591=15'h7C00; in592=15'h7C00; in593=15'h7C00; in594=15'h7C00; in595=15'h7C00; in596=15'h7C00; in597=15'h7C00; in598=15'h7C00;
   end
endmodule