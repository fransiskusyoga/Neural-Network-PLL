module lenet5_layer_1(clk,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81,out82,out83,out84,out85,out86,out87,out88,out89,out90,out91,out92,out93,out94,out95,out96,out97,out98,out99,out100,out101,out102,out103,out104,out105,out106,out107,out108,out109,out110,out111,out112,out113,out114,out115,out116,out117);
   input clk;
   input signed [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381;
   output reg signed [9:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81,out82,out83,out84,out85,out86,out87,out88,out89,out90,out91,out92,out93,out94,out95,out96,out97,out98,out99,out100,out101,out102,out103,out104,out105,out106,out107,out108,out109,out110,out111,out112,out113,out114,out115,out116,out117;
   wire signed [5:0] neg1,neg2,neg3,neg4,neg5,neg6,neg7,neg8,neg9,neg10,neg11,neg12,neg13,neg14,neg15,neg16,neg17,neg18,neg19,neg20,neg21,neg22,neg23,neg24,neg25,neg26,neg27,neg28,neg29,neg30,neg31,neg32,neg33,neg34,neg35,neg36,neg37,neg38,neg39,neg40,neg41,neg42,neg43,neg44,neg45,neg46,neg47,neg48,neg49,neg50,neg51,neg52,neg53,neg54,neg55,neg56,neg57,neg58,neg59,neg60,neg61,neg62,neg63,neg64,neg65,neg66,neg67,neg68,neg69,neg70,neg71,neg72,neg73,neg74,neg75,neg76,neg77,neg78,neg79,neg80,neg81,neg82,neg83,neg84,neg85,neg86,neg87,neg88,neg89,neg90,neg91,neg92,neg93,neg94,neg95,neg96,neg97,neg98,neg99,neg100,neg101,neg102,neg103,neg104,neg105,neg106,neg107,neg108,neg109,neg110,neg111,neg112,neg113,neg114,neg115,neg116,neg117,neg118,neg119,neg120,neg121,neg122,neg123,neg124,neg125,neg126,neg127,neg128,neg129,neg130,neg131,neg132,neg133,neg134,neg135,neg136,neg137,neg138,neg139,neg140,neg141,neg142,neg143,neg144,neg145,neg146,neg147,neg148,neg149,neg150,neg151,neg152,neg153,neg154,neg155,neg156,neg157,neg158,neg159,neg160,neg161,neg162,neg163,neg164,neg165,neg166,neg167,neg168,neg169,neg170,neg171,neg172,neg173,neg174,neg175,neg176,neg177,neg178,neg179,neg180,neg181,neg182,neg183,neg184,neg185,neg186,neg187,neg188,neg189,neg190,neg191,neg192,neg193,neg194,neg195,neg196,neg197,neg198,neg199,neg200,neg201,neg202,neg203,neg204,neg205,neg206,neg207,neg208,neg209,neg210,neg211,neg212,neg213,neg214,neg215,neg216,neg217,neg218,neg219,neg220,neg221,neg222,neg223,neg224,neg225,neg226,neg227,neg228,neg229,neg230,neg231,neg232,neg233,neg234,neg235,neg236,neg237,neg238,neg239,neg240,neg241,neg242,neg243,neg244,neg245,neg246,neg247,neg248,neg249,neg250,neg251,neg252,neg253,neg254,neg255,neg256,neg257,neg258,neg259,neg260,neg261,neg262,neg263,neg264,neg265,neg266,neg267,neg268,neg269,neg270,neg271,neg272,neg273,neg274,neg275,neg276,neg277,neg278,neg279,neg280,neg281,neg282,neg283,neg284,neg285,neg286,neg287,neg288,neg289,neg290,neg291,neg292,neg293,neg294,neg295,neg296,neg297,neg298,neg299,neg300,neg301,neg302,neg303,neg304,neg305,neg306,neg307,neg308,neg309,neg310,neg311,neg312,neg313,neg314,neg315,neg316,neg317,neg318,neg319,neg320,neg321,neg322,neg323,neg324,neg325,neg326,neg327,neg328,neg329,neg330,neg331,neg332,neg333,neg334,neg335,neg336,neg337,neg338,neg339,neg340,neg341,neg342,neg343,neg344,neg345,neg346,neg347,neg348,neg349,neg350,neg351,neg352,neg353,neg354,neg355,neg356,neg357,neg358,neg359,neg360,neg361,neg362,neg363,neg364,neg365,neg366,neg367,neg368,neg369,neg370,neg371,neg372,neg373,neg374,neg375,neg376,neg377,neg378,neg379,neg380,neg381;

   //Bias value
   wire signed [9:0] b1 = $signed(10'h0);
   wire signed [9:0] b2 = $signed(10'h1);
   wire signed [9:0] b3 = $signed(10'h0);
   wire signed [9:0] b4 = $signed(10'h0);
   wire signed [9:0] b5 = $signed(10'h0);
   wire signed [9:0] b6 = $signed(10'h1);
   wire signed [9:0] b7 = $signed(10'h3FF);
   wire signed [9:0] b8 = $signed(10'h0);
   wire signed [9:0] b9 = $signed(10'h0);
   wire signed [9:0] b10 = $signed(10'h1);
   wire signed [9:0] b11 = $signed(10'h0);
   wire signed [9:0] b12 = $signed(10'h0);
   wire signed [9:0] b13 = $signed(10'h3FF);
   wire signed [9:0] b14 = $signed(10'h1);
   wire signed [9:0] b15 = $signed(10'h1);
   wire signed [9:0] b16 = $signed(10'h3FF);
   wire signed [9:0] b17 = $signed(10'h0);
   wire signed [9:0] b18 = $signed(10'h1);
   wire signed [9:0] b19 = $signed(10'h0);
   wire signed [9:0] b20 = $signed(10'h3FF);
   wire signed [9:0] b21 = $signed(10'h0);
   wire signed [9:0] b22 = $signed(10'h1);
   wire signed [9:0] b23 = $signed(10'h0);
   wire signed [9:0] b24 = $signed(10'h0);
   wire signed [9:0] b25 = $signed(10'h3FF);
   wire signed [9:0] b26 = $signed(10'h1);
   wire signed [9:0] b27 = $signed(10'h0);
   wire signed [9:0] b28 = $signed(10'h3FF);
   wire signed [9:0] b29 = $signed(10'h1);
   wire signed [9:0] b30 = $signed(10'h3FF);
   wire signed [9:0] b31 = $signed(10'h0);
   wire signed [9:0] b32 = $signed(10'h1);
   wire signed [9:0] b33 = $signed(10'h3FF);
   wire signed [9:0] b34 = $signed(10'h1);
   wire signed [9:0] b35 = $signed(10'h3FF);
   wire signed [9:0] b36 = $signed(10'h0);
   wire signed [9:0] b37 = $signed(10'h0);
   wire signed [9:0] b38 = $signed(10'h1);
   wire signed [9:0] b39 = $signed(10'h0);
   wire signed [9:0] b40 = $signed(10'h0);
   wire signed [9:0] b41 = $signed(10'h3FF);
   wire signed [9:0] b42 = $signed(10'h0);
   wire signed [9:0] b43 = $signed(10'h0);
   wire signed [9:0] b44 = $signed(10'h0);
   wire signed [9:0] b45 = $signed(10'h0);
   wire signed [9:0] b46 = $signed(10'h0);
   wire signed [9:0] b47 = $signed(10'h0);
   wire signed [9:0] b48 = $signed(10'h0);
   wire signed [9:0] b49 = $signed(10'h0);
   wire signed [9:0] b50 = $signed(10'h0);
   wire signed [9:0] b51 = $signed(10'h1);
   wire signed [9:0] b52 = $signed(10'h1);
   wire signed [9:0] b53 = $signed(10'h1);
   wire signed [9:0] b54 = $signed(10'h0);
   wire signed [9:0] b55 = $signed(10'h0);
   wire signed [9:0] b56 = $signed(10'h3FF);
   wire signed [9:0] b57 = $signed(10'h0);
   wire signed [9:0] b58 = $signed(10'h0);
   wire signed [9:0] b59 = $signed(10'h0);
   wire signed [9:0] b60 = $signed(10'h0);
   wire signed [9:0] b61 = $signed(10'h3FF);
   wire signed [9:0] b62 = $signed(10'h0);
   wire signed [9:0] b63 = $signed(10'h0);
   wire signed [9:0] b64 = $signed(10'h0);
   wire signed [9:0] b65 = $signed(10'h0);
   wire signed [9:0] b66 = $signed(10'h0);
   wire signed [9:0] b67 = $signed(10'h0);
   wire signed [9:0] b68 = $signed(10'h1);
   wire signed [9:0] b69 = $signed(10'h0);
   wire signed [9:0] b70 = $signed(10'h0);
   wire signed [9:0] b71 = $signed(10'h0);
   wire signed [9:0] b72 = $signed(10'h0);
   wire signed [9:0] b73 = $signed(10'h0);
   wire signed [9:0] b74 = $signed(10'h0);
   wire signed [9:0] b75 = $signed(10'h3FF);
   wire signed [9:0] b76 = $signed(10'h1);
   wire signed [9:0] b77 = $signed(10'h0);
   wire signed [9:0] b78 = $signed(10'h0);
   wire signed [9:0] b79 = $signed(10'h3FF);
   wire signed [9:0] b80 = $signed(10'h0);
   wire signed [9:0] b81 = $signed(10'h0);
   wire signed [9:0] b82 = $signed(10'h0);
   wire signed [9:0] b83 = $signed(10'h0);
   wire signed [9:0] b84 = $signed(10'h0);
   wire signed [9:0] b85 = $signed(10'h0);
   wire signed [9:0] b86 = $signed(10'h0);
   wire signed [9:0] b87 = $signed(10'h0);
   wire signed [9:0] b88 = $signed(10'h0);
   wire signed [9:0] b89 = $signed(10'h0);
   wire signed [9:0] b90 = $signed(10'h1);
   wire signed [9:0] b91 = $signed(10'h1);
   wire signed [9:0] b92 = $signed(10'h0);
   wire signed [9:0] b93 = $signed(10'h0);
   wire signed [9:0] b94 = $signed(10'h3FF);
   wire signed [9:0] b95 = $signed(10'h0);
   wire signed [9:0] b96 = $signed(10'h3FF);
   wire signed [9:0] b97 = $signed(10'h1);
   wire signed [9:0] b98 = $signed(10'h1);
   wire signed [9:0] b99 = $signed(10'h1);
   wire signed [9:0] b100 = $signed(10'h0);
   wire signed [9:0] b101 = $signed(10'h3FF);
   wire signed [9:0] b102 = $signed(10'h3FE);
   wire signed [9:0] b103 = $signed(10'h3FF);
   wire signed [9:0] b104 = $signed(10'h3FF);
   wire signed [9:0] b105 = $signed(10'h0);
   wire signed [9:0] b106 = $signed(10'h3FF);
   wire signed [9:0] b107 = $signed(10'h0);
   wire signed [9:0] b108 = $signed(10'h3FF);
   wire signed [9:0] b109 = $signed(10'h0);
   wire signed [9:0] b110 = $signed(10'h1);
   wire signed [9:0] b111 = $signed(10'h0);
   wire signed [9:0] b112 = $signed(10'h0);
   wire signed [9:0] b113 = $signed(10'h0);
   wire signed [9:0] b114 = $signed(10'h0);
   wire signed [9:0] b115 = $signed(10'h0);
   wire signed [9:0] b116 = $signed(10'h3FE);
   wire signed [9:0] b117 = $signed(10'h3FF);

   //Negation modules
   negate #(6) N1(in1,neg1);
   negate #(6) N2(in2,neg2);
   negate #(6) N3(in3,neg3);
   negate #(6) N4(in4,neg4);
   negate #(6) N5(in5,neg5);
   negate #(6) N6(in6,neg6);
   negate #(6) N7(in7,neg7);
   negate #(6) N8(in8,neg8);
   negate #(6) N9(in9,neg9);
   negate #(6) N10(in10,neg10);
   negate #(6) N11(in11,neg11);
   negate #(6) N12(in12,neg12);
   negate #(6) N13(in13,neg13);
   negate #(6) N14(in14,neg14);
   negate #(6) N15(in15,neg15);
   negate #(6) N16(in16,neg16);
   negate #(6) N17(in17,neg17);
   negate #(6) N18(in18,neg18);
   negate #(6) N19(in19,neg19);
   negate #(6) N20(in20,neg20);
   negate #(6) N21(in21,neg21);
   negate #(6) N22(in22,neg22);
   negate #(6) N23(in23,neg23);
   negate #(6) N24(in24,neg24);
   negate #(6) N25(in25,neg25);
   negate #(6) N26(in26,neg26);
   negate #(6) N27(in27,neg27);
   negate #(6) N28(in28,neg28);
   negate #(6) N29(in29,neg29);
   negate #(6) N30(in30,neg30);
   negate #(6) N31(in31,neg31);
   negate #(6) N32(in32,neg32);
   negate #(6) N33(in33,neg33);
   negate #(6) N34(in34,neg34);
   negate #(6) N35(in35,neg35);
   negate #(6) N36(in36,neg36);
   negate #(6) N37(in37,neg37);
   negate #(6) N38(in38,neg38);
   negate #(6) N39(in39,neg39);
   negate #(6) N40(in40,neg40);
   negate #(6) N41(in41,neg41);
   negate #(6) N42(in42,neg42);
   negate #(6) N43(in43,neg43);
   negate #(6) N44(in44,neg44);
   negate #(6) N45(in45,neg45);
   negate #(6) N46(in46,neg46);
   negate #(6) N47(in47,neg47);
   negate #(6) N48(in48,neg48);
   negate #(6) N49(in49,neg49);
   negate #(6) N50(in50,neg50);
   negate #(6) N51(in51,neg51);
   negate #(6) N52(in52,neg52);
   negate #(6) N53(in53,neg53);
   negate #(6) N54(in54,neg54);
   negate #(6) N55(in55,neg55);
   negate #(6) N56(in56,neg56);
   negate #(6) N57(in57,neg57);
   negate #(6) N58(in58,neg58);
   negate #(6) N59(in59,neg59);
   negate #(6) N60(in60,neg60);
   negate #(6) N61(in61,neg61);
   negate #(6) N62(in62,neg62);
   negate #(6) N63(in63,neg63);
   negate #(6) N64(in64,neg64);
   negate #(6) N65(in65,neg65);
   negate #(6) N66(in66,neg66);
   negate #(6) N67(in67,neg67);
   negate #(6) N68(in68,neg68);
   negate #(6) N69(in69,neg69);
   negate #(6) N70(in70,neg70);
   negate #(6) N71(in71,neg71);
   negate #(6) N72(in72,neg72);
   negate #(6) N73(in73,neg73);
   negate #(6) N74(in74,neg74);
   negate #(6) N75(in75,neg75);
   negate #(6) N76(in76,neg76);
   negate #(6) N77(in77,neg77);
   negate #(6) N78(in78,neg78);
   negate #(6) N79(in79,neg79);
   negate #(6) N80(in80,neg80);
   negate #(6) N81(in81,neg81);
   negate #(6) N82(in82,neg82);
   negate #(6) N83(in83,neg83);
   negate #(6) N84(in84,neg84);
   negate #(6) N85(in85,neg85);
   negate #(6) N86(in86,neg86);
   negate #(6) N87(in87,neg87);
   negate #(6) N88(in88,neg88);
   negate #(6) N89(in89,neg89);
   negate #(6) N90(in90,neg90);
   negate #(6) N91(in91,neg91);
   negate #(6) N92(in92,neg92);
   negate #(6) N93(in93,neg93);
   negate #(6) N94(in94,neg94);
   negate #(6) N95(in95,neg95);
   negate #(6) N96(in96,neg96);
   negate #(6) N97(in97,neg97);
   negate #(6) N98(in98,neg98);
   negate #(6) N99(in99,neg99);
   negate #(6) N100(in100,neg100);
   negate #(6) N101(in101,neg101);
   negate #(6) N102(in102,neg102);
   negate #(6) N103(in103,neg103);
   negate #(6) N104(in104,neg104);
   negate #(6) N105(in105,neg105);
   negate #(6) N106(in106,neg106);
   negate #(6) N107(in107,neg107);
   negate #(6) N108(in108,neg108);
   negate #(6) N109(in109,neg109);
   negate #(6) N110(in110,neg110);
   negate #(6) N111(in111,neg111);
   negate #(6) N112(in112,neg112);
   negate #(6) N113(in113,neg113);
   negate #(6) N114(in114,neg114);
   negate #(6) N115(in115,neg115);
   negate #(6) N116(in116,neg116);
   negate #(6) N117(in117,neg117);
   negate #(6) N118(in118,neg118);
   negate #(6) N119(in119,neg119);
   negate #(6) N120(in120,neg120);
   negate #(6) N121(in121,neg121);
   negate #(6) N122(in122,neg122);
   negate #(6) N123(in123,neg123);
   negate #(6) N124(in124,neg124);
   negate #(6) N125(in125,neg125);
   negate #(6) N126(in126,neg126);
   negate #(6) N127(in127,neg127);
   negate #(6) N128(in128,neg128);
   negate #(6) N129(in129,neg129);
   negate #(6) N130(in130,neg130);
   negate #(6) N131(in131,neg131);
   negate #(6) N132(in132,neg132);
   negate #(6) N133(in133,neg133);
   negate #(6) N134(in134,neg134);
   negate #(6) N135(in135,neg135);
   negate #(6) N136(in136,neg136);
   negate #(6) N137(in137,neg137);
   negate #(6) N138(in138,neg138);
   negate #(6) N139(in139,neg139);
   negate #(6) N140(in140,neg140);
   negate #(6) N141(in141,neg141);
   negate #(6) N142(in142,neg142);
   negate #(6) N143(in143,neg143);
   negate #(6) N144(in144,neg144);
   negate #(6) N145(in145,neg145);
   negate #(6) N146(in146,neg146);
   negate #(6) N147(in147,neg147);
   negate #(6) N148(in148,neg148);
   negate #(6) N149(in149,neg149);
   negate #(6) N150(in150,neg150);
   negate #(6) N151(in151,neg151);
   negate #(6) N152(in152,neg152);
   negate #(6) N153(in153,neg153);
   negate #(6) N154(in154,neg154);
   negate #(6) N155(in155,neg155);
   negate #(6) N156(in156,neg156);
   negate #(6) N157(in157,neg157);
   negate #(6) N158(in158,neg158);
   negate #(6) N159(in159,neg159);
   negate #(6) N160(in160,neg160);
   negate #(6) N161(in161,neg161);
   negate #(6) N162(in162,neg162);
   negate #(6) N163(in163,neg163);
   negate #(6) N164(in164,neg164);
   negate #(6) N165(in165,neg165);
   negate #(6) N166(in166,neg166);
   negate #(6) N167(in167,neg167);
   negate #(6) N168(in168,neg168);
   negate #(6) N169(in169,neg169);
   negate #(6) N170(in170,neg170);
   negate #(6) N171(in171,neg171);
   negate #(6) N172(in172,neg172);
   negate #(6) N173(in173,neg173);
   negate #(6) N174(in174,neg174);
   negate #(6) N175(in175,neg175);
   negate #(6) N176(in176,neg176);
   negate #(6) N177(in177,neg177);
   negate #(6) N178(in178,neg178);
   negate #(6) N179(in179,neg179);
   negate #(6) N180(in180,neg180);
   negate #(6) N181(in181,neg181);
   negate #(6) N182(in182,neg182);
   negate #(6) N183(in183,neg183);
   negate #(6) N184(in184,neg184);
   negate #(6) N185(in185,neg185);
   negate #(6) N186(in186,neg186);
   negate #(6) N187(in187,neg187);
   negate #(6) N188(in188,neg188);
   negate #(6) N189(in189,neg189);
   negate #(6) N190(in190,neg190);
   negate #(6) N191(in191,neg191);
   negate #(6) N192(in192,neg192);
   negate #(6) N193(in193,neg193);
   negate #(6) N194(in194,neg194);
   negate #(6) N195(in195,neg195);
   negate #(6) N196(in196,neg196);
   negate #(6) N197(in197,neg197);
   negate #(6) N198(in198,neg198);
   negate #(6) N199(in199,neg199);
   negate #(6) N200(in200,neg200);
   negate #(6) N201(in201,neg201);
   negate #(6) N202(in202,neg202);
   negate #(6) N203(in203,neg203);
   negate #(6) N204(in204,neg204);
   negate #(6) N205(in205,neg205);
   negate #(6) N206(in206,neg206);
   negate #(6) N207(in207,neg207);
   negate #(6) N208(in208,neg208);
   negate #(6) N209(in209,neg209);
   negate #(6) N210(in210,neg210);
   negate #(6) N211(in211,neg211);
   negate #(6) N212(in212,neg212);
   negate #(6) N213(in213,neg213);
   negate #(6) N214(in214,neg214);
   negate #(6) N215(in215,neg215);
   negate #(6) N216(in216,neg216);
   negate #(6) N217(in217,neg217);
   negate #(6) N218(in218,neg218);
   negate #(6) N219(in219,neg219);
   negate #(6) N220(in220,neg220);
   negate #(6) N221(in221,neg221);
   negate #(6) N222(in222,neg222);
   negate #(6) N223(in223,neg223);
   negate #(6) N224(in224,neg224);
   negate #(6) N225(in225,neg225);
   negate #(6) N226(in226,neg226);
   negate #(6) N227(in227,neg227);
   negate #(6) N228(in228,neg228);
   negate #(6) N229(in229,neg229);
   negate #(6) N230(in230,neg230);
   negate #(6) N231(in231,neg231);
   negate #(6) N232(in232,neg232);
   negate #(6) N233(in233,neg233);
   negate #(6) N234(in234,neg234);
   negate #(6) N235(in235,neg235);
   negate #(6) N236(in236,neg236);
   negate #(6) N237(in237,neg237);
   negate #(6) N238(in238,neg238);
   negate #(6) N239(in239,neg239);
   negate #(6) N240(in240,neg240);
   negate #(6) N241(in241,neg241);
   negate #(6) N242(in242,neg242);
   negate #(6) N243(in243,neg243);
   negate #(6) N244(in244,neg244);
   negate #(6) N245(in245,neg245);
   negate #(6) N246(in246,neg246);
   negate #(6) N247(in247,neg247);
   negate #(6) N248(in248,neg248);
   negate #(6) N249(in249,neg249);
   negate #(6) N250(in250,neg250);
   negate #(6) N251(in251,neg251);
   negate #(6) N252(in252,neg252);
   negate #(6) N253(in253,neg253);
   negate #(6) N254(in254,neg254);
   negate #(6) N255(in255,neg255);
   negate #(6) N256(in256,neg256);
   negate #(6) N257(in257,neg257);
   negate #(6) N258(in258,neg258);
   negate #(6) N259(in259,neg259);
   negate #(6) N260(in260,neg260);
   negate #(6) N261(in261,neg261);
   negate #(6) N262(in262,neg262);
   negate #(6) N263(in263,neg263);
   negate #(6) N264(in264,neg264);
   negate #(6) N265(in265,neg265);
   negate #(6) N266(in266,neg266);
   negate #(6) N267(in267,neg267);
   negate #(6) N268(in268,neg268);
   negate #(6) N269(in269,neg269);
   negate #(6) N270(in270,neg270);
   negate #(6) N271(in271,neg271);
   negate #(6) N272(in272,neg272);
   negate #(6) N273(in273,neg273);
   negate #(6) N274(in274,neg274);
   negate #(6) N275(in275,neg275);
   negate #(6) N276(in276,neg276);
   negate #(6) N277(in277,neg277);
   negate #(6) N278(in278,neg278);
   negate #(6) N279(in279,neg279);
   negate #(6) N280(in280,neg280);
   negate #(6) N281(in281,neg281);
   negate #(6) N282(in282,neg282);
   negate #(6) N283(in283,neg283);
   negate #(6) N284(in284,neg284);
   negate #(6) N285(in285,neg285);
   negate #(6) N286(in286,neg286);
   negate #(6) N287(in287,neg287);
   negate #(6) N288(in288,neg288);
   negate #(6) N289(in289,neg289);
   negate #(6) N290(in290,neg290);
   negate #(6) N291(in291,neg291);
   negate #(6) N292(in292,neg292);
   negate #(6) N293(in293,neg293);
   negate #(6) N294(in294,neg294);
   negate #(6) N295(in295,neg295);
   negate #(6) N296(in296,neg296);
   negate #(6) N297(in297,neg297);
   negate #(6) N298(in298,neg298);
   negate #(6) N299(in299,neg299);
   negate #(6) N300(in300,neg300);
   negate #(6) N301(in301,neg301);
   negate #(6) N302(in302,neg302);
   negate #(6) N303(in303,neg303);
   negate #(6) N304(in304,neg304);
   negate #(6) N305(in305,neg305);
   negate #(6) N306(in306,neg306);
   negate #(6) N307(in307,neg307);
   negate #(6) N308(in308,neg308);
   negate #(6) N309(in309,neg309);
   negate #(6) N310(in310,neg310);
   negate #(6) N311(in311,neg311);
   negate #(6) N312(in312,neg312);
   negate #(6) N313(in313,neg313);
   negate #(6) N314(in314,neg314);
   negate #(6) N315(in315,neg315);
   negate #(6) N316(in316,neg316);
   negate #(6) N317(in317,neg317);
   negate #(6) N318(in318,neg318);
   negate #(6) N319(in319,neg319);
   negate #(6) N320(in320,neg320);
   negate #(6) N321(in321,neg321);
   negate #(6) N322(in322,neg322);
   negate #(6) N323(in323,neg323);
   negate #(6) N324(in324,neg324);
   negate #(6) N325(in325,neg325);
   negate #(6) N326(in326,neg326);
   negate #(6) N327(in327,neg327);
   negate #(6) N328(in328,neg328);
   negate #(6) N329(in329,neg329);
   negate #(6) N330(in330,neg330);
   negate #(6) N331(in331,neg331);
   negate #(6) N332(in332,neg332);
   negate #(6) N333(in333,neg333);
   negate #(6) N334(in334,neg334);
   negate #(6) N335(in335,neg335);
   negate #(6) N336(in336,neg336);
   negate #(6) N337(in337,neg337);
   negate #(6) N338(in338,neg338);
   negate #(6) N339(in339,neg339);
   negate #(6) N340(in340,neg340);
   negate #(6) N341(in341,neg341);
   negate #(6) N342(in342,neg342);
   negate #(6) N343(in343,neg343);
   negate #(6) N344(in344,neg344);
   negate #(6) N345(in345,neg345);
   negate #(6) N346(in346,neg346);
   negate #(6) N347(in347,neg347);
   negate #(6) N348(in348,neg348);
   negate #(6) N349(in349,neg349);
   negate #(6) N350(in350,neg350);
   negate #(6) N351(in351,neg351);
   negate #(6) N352(in352,neg352);
   negate #(6) N353(in353,neg353);
   negate #(6) N354(in354,neg354);
   negate #(6) N355(in355,neg355);
   negate #(6) N356(in356,neg356);
   negate #(6) N357(in357,neg357);
   negate #(6) N358(in358,neg358);
   negate #(6) N359(in359,neg359);
   negate #(6) N360(in360,neg360);
   negate #(6) N361(in361,neg361);
   negate #(6) N362(in362,neg362);
   negate #(6) N363(in363,neg363);
   negate #(6) N364(in364,neg364);
   negate #(6) N365(in365,neg365);
   negate #(6) N366(in366,neg366);
   negate #(6) N367(in367,neg367);
   negate #(6) N368(in368,neg368);
   negate #(6) N369(in369,neg369);
   negate #(6) N370(in370,neg370);
   negate #(6) N371(in371,neg371);
   negate #(6) N372(in372,neg372);
   negate #(6) N373(in373,neg373);
   negate #(6) N374(in374,neg374);
   negate #(6) N375(in375,neg375);
   negate #(6) N376(in376,neg376);
   negate #(6) N377(in377,neg377);
   negate #(6) N378(in378,neg378);
   negate #(6) N379(in379,neg379);
   negate #(6) N380(in380,neg380);
   negate #(6) N381(in381,neg381);

   // m1_1 = W*in
   wire signed [9:0] m1_1;
   assign m1_1 =10'b0;

   // m1_2 = W*in
   wire signed [9:0] m1_2;
   assign m1_2 =10'b0;

   // m1_3 = W*in
   wire signed [9:0] m1_3;
   assign m1_3 =10'b0;

   // m1_4 = W*in
   wire signed [9:0] m1_4;
   assign m1_4 =10'b0;

   // m1_5 = W*in
   wire signed [9:0] m1_5;
   assign m1_5 =10'b0;

   // m1_6 = W*in
   wire signed [9:0] m1_6;
   assign m1_6 =10'b0;

   // m1_7 = W*in
   wire signed [9:0] m1_7;
   assign m1_7 =10'b0;

   // m1_8 = W*in
   wire signed [9:0] m1_8;
   assign m1_8 =10'b0;

   // m1_9 = W*in
   wire signed [9:0] m1_9;
   assign m1_9 =10'b0;

   // m1_10 = W*in
   wire signed [9:0] m1_10;
   assign m1_10 =10'b0;

   // m1_11 = W*in
   wire signed [9:0] m1_11;
   assign m1_11 =10'b0;

   // m1_12 = W*in
   wire signed [9:0] m1_12;
   assign m1_12 =10'b0;

   // m1_13 = W*in
   wire signed [9:0] m1_13;
   assign m1_13 =10'b0;

   // m1_14 = W*in
   wire signed [9:0] m1_14;
   assign m1_14 =10'b0;

   // m1_15 = W*in
   wire signed [9:0] m1_15;
   assign m1_15 =10'b0;

   // m1_16 = W*in
   wire signed [9:0] m1_16;
   assign m1_16 =10'b0;

   // m1_17 = W*in
   wire signed [9:0] m1_17;
   assign m1_17 =10'b0;

   // m1_18 = W*in
   wire signed [9:0] m1_18;
   assign m1_18 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_19 = W*in
   wire signed [9:0] m1_19;
   assign m1_19 =10'b0;

   // m1_20 = W*in
   wire signed [9:0] m1_20;
   assign m1_20 =10'b0;

   // m1_21 = W*in
   wire signed [9:0] m1_21;
   assign m1_21 =10'b0;

   // m1_22 = W*in
   wire signed [9:0] m1_22;
   assign m1_22 =10'b0;

   // m1_23 = W*in
   wire signed [9:0] m1_23;
   assign m1_23 =10'b0;

   // m1_24 = W*in
   wire signed [9:0] m1_24;
   assign m1_24 =10'b0;

   // m1_25 = W*in
   wire signed [9:0] m1_25;
   assign m1_25 =10'b0;

   // m1_26 = W*in
   wire signed [9:0] m1_26;
   assign m1_26 =10'b0;

   // m1_27 = W*in
   wire signed [9:0] m1_27;
   assign m1_27 =10'b0;

   // m1_28 = W*in
   wire signed [9:0] m1_28;
   assign m1_28 =10'b0;

   // m1_29 = W*in
   wire signed [9:0] m1_29;
   assign m1_29 =10'b0;

   // m1_30 = W*in
   wire signed [9:0] m1_30;
   assign m1_30 =10'b0;

   // m1_31 = W*in
   wire signed [9:0] m1_31;
   assign m1_31 ={ {5{in1[5]}} , in1[5:1] };

   // m1_32 = W*in
   wire signed [9:0] m1_32;
   assign m1_32 =10'b0;

   // m1_33 = W*in
   wire signed [9:0] m1_33;
   assign m1_33 =10'b0;

   // m1_34 = W*in
   wire signed [9:0] m1_34;
   assign m1_34 =10'b0;

   // m1_35 = W*in
   wire signed [9:0] m1_35;
   assign m1_35 =10'b0;

   // m1_36 = W*in
   wire signed [9:0] m1_36;
   assign m1_36 =10'b0;

   // m1_37 = W*in
   wire signed [9:0] m1_37;
   assign m1_37 =10'b0;

   // m1_38 = W*in
   wire signed [9:0] m1_38;
   assign m1_38 ={ {4{neg1[5]}} , neg1[5:0] };

   // m1_39 = W*in
   wire signed [9:0] m1_39;
   assign m1_39 =10'b0;

   // m1_40 = W*in
   wire signed [9:0] m1_40;
   assign m1_40 =10'b0;

   // m1_41 = W*in
   wire signed [9:0] m1_41;
   assign m1_41 =10'b0;

   // m1_42 = W*in
   wire signed [9:0] m1_42;
   assign m1_42 =10'b0;

   // m1_43 = W*in
   wire signed [9:0] m1_43;
   assign m1_43 ={ {4{neg1[5]}} , neg1[5:0] };

   // m1_44 = W*in
   wire signed [9:0] m1_44;
   assign m1_44 =10'b0;

   // m1_45 = W*in
   wire signed [9:0] m1_45;
   assign m1_45 =10'b0;

   // m1_46 = W*in
   wire signed [9:0] m1_46;
   assign m1_46 =10'b0;

   // m1_47 = W*in
   wire signed [9:0] m1_47;
   assign m1_47 =10'b0;

   // m1_48 = W*in
   wire signed [9:0] m1_48;
   assign m1_48 =10'b0;

   // m1_49 = W*in
   wire signed [9:0] m1_49;
   assign m1_49 =10'b0;

   // m1_50 = W*in
   wire signed [9:0] m1_50;
   assign m1_50 =10'b0;

   // m1_51 = W*in
   wire signed [9:0] m1_51;
   assign m1_51 ={ {4{in1[5]}} , in1[5:0] };

   // m1_52 = W*in
   wire signed [9:0] m1_52;
   assign m1_52 =10'b0;

   // m1_53 = W*in
   wire signed [9:0] m1_53;
   assign m1_53 =10'b0;

   // m1_54 = W*in
   wire signed [9:0] m1_54;
   assign m1_54 =10'b0;

   // m1_55 = W*in
   wire signed [9:0] m1_55;
   assign m1_55 =10'b0;

   // m1_56 = W*in
   wire signed [9:0] m1_56;
   assign m1_56 =10'b0;

   // m1_57 = W*in
   wire signed [9:0] m1_57;
   assign m1_57 =10'b0;

   // m1_58 = W*in
   wire signed [9:0] m1_58;
   assign m1_58 =10'b0;

   // m1_59 = W*in
   wire signed [9:0] m1_59;
   assign m1_59 =10'b0;

   // m1_60 = W*in
   wire signed [9:0] m1_60;
   assign m1_60 =10'b0;

   // m1_61 = W*in
   wire signed [9:0] m1_61;
   assign m1_61 =10'b0;

   // m1_62 = W*in
   wire signed [9:0] m1_62;
   assign m1_62 =10'b0;

   // m1_63 = W*in
   wire signed [9:0] m1_63;
   assign m1_63 ={ {4{neg1[5]}} , neg1[5:0] };

   // m1_64 = W*in
   wire signed [9:0] m1_64;
   assign m1_64 =10'b0;

   // m1_65 = W*in
   wire signed [9:0] m1_65;
   assign m1_65 =10'b0;

   // m1_66 = W*in
   wire signed [9:0] m1_66;
   assign m1_66 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_67 = W*in
   wire signed [9:0] m1_67;
   assign m1_67 ={ {5{in1[5]}} , in1[5:1] };

   // m1_68 = W*in
   wire signed [9:0] m1_68;
   assign m1_68 =10'b0;

   // m1_69 = W*in
   wire signed [9:0] m1_69;
   assign m1_69 =10'b0;

   // m1_70 = W*in
   wire signed [9:0] m1_70;
   assign m1_70 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_71 = W*in
   wire signed [9:0] m1_71;
   assign m1_71 =10'b0;

   // m1_72 = W*in
   wire signed [9:0] m1_72;
   assign m1_72 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_73 = W*in
   wire signed [9:0] m1_73;
   assign m1_73 ={ {4{in1[5]}} , in1[5:0] };

   // m1_74 = W*in
   wire signed [9:0] m1_74;
   assign m1_74 ={ {4{neg1[5]}} , neg1[5:0] };

   // m1_75 = W*in
   wire signed [9:0] m1_75;
   assign m1_75 =10'b0;

   // m1_76 = W*in
   wire signed [9:0] m1_76;
   assign m1_76 =10'b0;

   // m1_77 = W*in
   wire signed [9:0] m1_77;
   assign m1_77 =10'b0;

   // m1_78 = W*in
   wire signed [9:0] m1_78;
   assign m1_78 =10'b0;

   // m1_79 = W*in
   wire signed [9:0] m1_79;
   assign m1_79 =10'b0;

   // m1_80 = W*in
   wire signed [9:0] m1_80;
   assign m1_80 ={ {4{in1[5]}} , in1[5:0] };

   // m1_81 = W*in
   wire signed [9:0] m1_81;
   assign m1_81 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_82 = W*in
   wire signed [9:0] m1_82;
   assign m1_82 =10'b0;

   // m1_83 = W*in
   wire signed [9:0] m1_83;
   assign m1_83 =10'b0;

   // m1_84 = W*in
   wire signed [9:0] m1_84;
   assign m1_84 =10'b0;

   // m1_85 = W*in
   wire signed [9:0] m1_85;
   assign m1_85 =10'b0;

   // m1_86 = W*in
   wire signed [9:0] m1_86;
   assign m1_86 =10'b0;

   // m1_87 = W*in
   wire signed [9:0] m1_87;
   assign m1_87 =10'b0;

   // m1_88 = W*in
   wire signed [9:0] m1_88;
   assign m1_88 =10'b0;

   // m1_89 = W*in
   wire signed [9:0] m1_89;
   assign m1_89 =10'b0;

   // m1_90 = W*in
   wire signed [9:0] m1_90;
   assign m1_90 =10'b0;

   // m1_91 = W*in
   wire signed [9:0] m1_91;
   assign m1_91 =10'b0;

   // m1_92 = W*in
   wire signed [9:0] m1_92;
   assign m1_92 =10'b0;

   // m1_93 = W*in
   wire signed [9:0] m1_93;
   assign m1_93 =10'b0;

   // m1_94 = W*in
   wire signed [9:0] m1_94;
   assign m1_94 =10'b0;

   // m1_95 = W*in
   wire signed [9:0] m1_95;
   assign m1_95 =10'b0;

   // m1_96 = W*in
   wire signed [9:0] m1_96;
   assign m1_96 =10'b0;

   // m1_97 = W*in
   wire signed [9:0] m1_97;
   assign m1_97 =10'b0;

   // m1_98 = W*in
   wire signed [9:0] m1_98;
   assign m1_98 =10'b0;

   // m1_99 = W*in
   wire signed [9:0] m1_99;
   assign m1_99 =10'b0;

   // m1_100 = W*in
   wire signed [9:0] m1_100;
   assign m1_100 =10'b0;

   // m1_101 = W*in
   wire signed [9:0] m1_101;
   assign m1_101 =10'b0;

   // m1_102 = W*in
   wire signed [9:0] m1_102;
   assign m1_102 =10'b0;

   // m1_103 = W*in
   wire signed [9:0] m1_103;
   assign m1_103 =10'b0;

   // m1_104 = W*in
   wire signed [9:0] m1_104;
   assign m1_104 =10'b0;

   // m1_105 = W*in
   wire signed [9:0] m1_105;
   assign m1_105 =10'b0;

   // m1_106 = W*in
   wire signed [9:0] m1_106;
   assign m1_106 =10'b0;

   // m1_107 = W*in
   wire signed [9:0] m1_107;
   assign m1_107 ={ {5{in1[5]}} , in1[5:1] };

   // m1_108 = W*in
   wire signed [9:0] m1_108;
   assign m1_108 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_109 = W*in
   wire signed [9:0] m1_109;
   assign m1_109 =10'b0;

   // m1_110 = W*in
   wire signed [9:0] m1_110;
   assign m1_110 =10'b0;

   // m1_111 = W*in
   wire signed [9:0] m1_111;
   assign m1_111 =10'b0;

   // m1_112 = W*in
   wire signed [9:0] m1_112;
   assign m1_112 =10'b0;

   // m1_113 = W*in
   wire signed [9:0] m1_113;
   assign m1_113 =10'b0;

   // m1_114 = W*in
   wire signed [9:0] m1_114;
   assign m1_114 =10'b0;

   // m1_115 = W*in
   wire signed [9:0] m1_115;
   assign m1_115 =10'b0;

   // m1_116 = W*in
   wire signed [9:0] m1_116;
   assign m1_116 ={ {5{neg1[5]}} , neg1[5:1] };

   // m1_117 = W*in
   wire signed [9:0] m1_117;
   assign m1_117 =10'b0;

   // m2_1 = W*in
   wire signed [9:0] m2_1;
   assign m2_1 =10'b0;

   // m2_2 = W*in
   wire signed [9:0] m2_2;
   assign m2_2 =10'b0;

   // m2_3 = W*in
   wire signed [9:0] m2_3;
   assign m2_3 =10'b0;

   // m2_4 = W*in
   wire signed [9:0] m2_4;
   assign m2_4 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_5 = W*in
   wire signed [9:0] m2_5;
   assign m2_5 =10'b0;

   // m2_6 = W*in
   wire signed [9:0] m2_6;
   assign m2_6 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_7 = W*in
   wire signed [9:0] m2_7;
   assign m2_7 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_8 = W*in
   wire signed [9:0] m2_8;
   assign m2_8 =10'b0;

   // m2_9 = W*in
   wire signed [9:0] m2_9;
   assign m2_9 =10'b0;

   // m2_10 = W*in
   wire signed [9:0] m2_10;
   assign m2_10 =10'b0;

   // m2_11 = W*in
   wire signed [9:0] m2_11;
   assign m2_11 ={ {4{in2[5]}} , in2[5:0] };

   // m2_12 = W*in
   wire signed [9:0] m2_12;
   assign m2_12 ={ {3{in2[5]}} , in2 , {1{1'b0}} };

   // m2_13 = W*in
   wire signed [9:0] m2_13;
   assign m2_13 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_14 = W*in
   wire signed [9:0] m2_14;
   assign m2_14 =10'b0;

   // m2_15 = W*in
   wire signed [9:0] m2_15;
   assign m2_15 =10'b0;

   // m2_16 = W*in
   wire signed [9:0] m2_16;
   assign m2_16 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_17 = W*in
   wire signed [9:0] m2_17;
   assign m2_17 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_18 = W*in
   wire signed [9:0] m2_18;
   assign m2_18 =10'b0;

   // m2_19 = W*in
   wire signed [9:0] m2_19;
   assign m2_19 ={ {4{in2[5]}} , in2[5:0] };

   // m2_20 = W*in
   wire signed [9:0] m2_20;
   assign m2_20 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_21 = W*in
   wire signed [9:0] m2_21;
   assign m2_21 =10'b0;

   // m2_22 = W*in
   wire signed [9:0] m2_22;
   assign m2_22 =10'b0;

   // m2_23 = W*in
   wire signed [9:0] m2_23;
   assign m2_23 =10'b0;

   // m2_24 = W*in
   wire signed [9:0] m2_24;
   assign m2_24 ={ {4{in2[5]}} , in2[5:0] };

   // m2_25 = W*in
   wire signed [9:0] m2_25;
   assign m2_25 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_26 = W*in
   wire signed [9:0] m2_26;
   assign m2_26 =10'b0;

   // m2_27 = W*in
   wire signed [9:0] m2_27;
   assign m2_27 ={ {5{in2[5]}} , in2[5:1] };

   // m2_28 = W*in
   wire signed [9:0] m2_28;
   assign m2_28 =10'b0;

   // m2_29 = W*in
   wire signed [9:0] m2_29;
   assign m2_29 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_30 = W*in
   wire signed [9:0] m2_30;
   assign m2_30 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_31 = W*in
   wire signed [9:0] m2_31;
   assign m2_31 =10'b0;

   // m2_32 = W*in
   wire signed [9:0] m2_32;
   assign m2_32 =10'b0;

   // m2_33 = W*in
   wire signed [9:0] m2_33;
   assign m2_33 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_34 = W*in
   wire signed [9:0] m2_34;
   assign m2_34 =10'b0;

   // m2_35 = W*in
   wire signed [9:0] m2_35;
   assign m2_35 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_36 = W*in
   wire signed [9:0] m2_36;
   assign m2_36 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_37 = W*in
   wire signed [9:0] m2_37;
   assign m2_37 =10'b0;

   // m2_38 = W*in
   wire signed [9:0] m2_38;
   assign m2_38 ={ {4{in2[5]}} , in2[5:0] };

   // m2_39 = W*in
   wire signed [9:0] m2_39;
   assign m2_39 ={ {4{in2[5]}} , in2[5:0] };

   // m2_40 = W*in
   wire signed [9:0] m2_40;
   assign m2_40 =10'b0;

   // m2_41 = W*in
   wire signed [9:0] m2_41;
   assign m2_41 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_42 = W*in
   wire signed [9:0] m2_42;
   assign m2_42 =10'b0;

   // m2_43 = W*in
   wire signed [9:0] m2_43;
   assign m2_43 =10'b0;

   // m2_44 = W*in
   wire signed [9:0] m2_44;
   assign m2_44 =10'b0;

   // m2_45 = W*in
   wire signed [9:0] m2_45;
   assign m2_45 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_46 = W*in
   wire signed [9:0] m2_46;
   assign m2_46 =10'b0;

   // m2_47 = W*in
   wire signed [9:0] m2_47;
   assign m2_47 =10'b0;

   // m2_48 = W*in
   wire signed [9:0] m2_48;
   assign m2_48 =10'b0;

   // m2_49 = W*in
   wire signed [9:0] m2_49;
   assign m2_49 ={ {4{in2[5]}} , in2[5:0] };

   // m2_50 = W*in
   wire signed [9:0] m2_50;
   assign m2_50 ={ {4{in2[5]}} , in2[5:0] };

   // m2_51 = W*in
   wire signed [9:0] m2_51;
   assign m2_51 =10'b0;

   // m2_52 = W*in
   wire signed [9:0] m2_52;
   assign m2_52 =10'b0;

   // m2_53 = W*in
   wire signed [9:0] m2_53;
   assign m2_53 =10'b0;

   // m2_54 = W*in
   wire signed [9:0] m2_54;
   assign m2_54 =10'b0;

   // m2_55 = W*in
   wire signed [9:0] m2_55;
   assign m2_55 =10'b0;

   // m2_56 = W*in
   wire signed [9:0] m2_56;
   assign m2_56 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_57 = W*in
   wire signed [9:0] m2_57;
   assign m2_57 =10'b0;

   // m2_58 = W*in
   wire signed [9:0] m2_58;
   assign m2_58 ={ {4{in2[5]}} , in2[5:0] };

   // m2_59 = W*in
   wire signed [9:0] m2_59;
   assign m2_59 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_60 = W*in
   wire signed [9:0] m2_60;
   assign m2_60 =10'b0;

   // m2_61 = W*in
   wire signed [9:0] m2_61;
   assign m2_61 =10'b0;

   // m2_62 = W*in
   wire signed [9:0] m2_62;
   assign m2_62 =10'b0;

   // m2_63 = W*in
   wire signed [9:0] m2_63;
   assign m2_63 =10'b0;

   // m2_64 = W*in
   wire signed [9:0] m2_64;
   assign m2_64 =10'b0;

   // m2_65 = W*in
   wire signed [9:0] m2_65;
   assign m2_65 ={ {5{in2[5]}} , in2[5:1] };

   // m2_66 = W*in
   wire signed [9:0] m2_66;
   assign m2_66 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_67 = W*in
   wire signed [9:0] m2_67;
   assign m2_67 =10'b0;

   // m2_68 = W*in
   wire signed [9:0] m2_68;
   assign m2_68 ={ {4{in2[5]}} , in2[5:0] };

   // m2_69 = W*in
   wire signed [9:0] m2_69;
   assign m2_69 =10'b0;

   // m2_70 = W*in
   wire signed [9:0] m2_70;
   assign m2_70 =10'b0;

   // m2_71 = W*in
   wire signed [9:0] m2_71;
   assign m2_71 ={ {4{in2[5]}} , in2[5:0] };

   // m2_72 = W*in
   wire signed [9:0] m2_72;
   assign m2_72 =10'b0;

   // m2_73 = W*in
   wire signed [9:0] m2_73;
   assign m2_73 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_74 = W*in
   wire signed [9:0] m2_74;
   assign m2_74 =10'b0;

   // m2_75 = W*in
   wire signed [9:0] m2_75;
   assign m2_75 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_76 = W*in
   wire signed [9:0] m2_76;
   assign m2_76 =10'b0;

   // m2_77 = W*in
   wire signed [9:0] m2_77;
   assign m2_77 =10'b0;

   // m2_78 = W*in
   wire signed [9:0] m2_78;
   assign m2_78 =10'b0;

   // m2_79 = W*in
   wire signed [9:0] m2_79;
   assign m2_79 =10'b0;

   // m2_80 = W*in
   wire signed [9:0] m2_80;
   assign m2_80 =10'b0;

   // m2_81 = W*in
   wire signed [9:0] m2_81;
   assign m2_81 =10'b0;

   // m2_82 = W*in
   wire signed [9:0] m2_82;
   assign m2_82 ={ {4{in2[5]}} , in2[5:0] };

   // m2_83 = W*in
   wire signed [9:0] m2_83;
   assign m2_83 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_84 = W*in
   wire signed [9:0] m2_84;
   assign m2_84 =10'b0;

   // m2_85 = W*in
   wire signed [9:0] m2_85;
   assign m2_85 =10'b0;

   // m2_86 = W*in
   wire signed [9:0] m2_86;
   assign m2_86 =10'b0;

   // m2_87 = W*in
   wire signed [9:0] m2_87;
   assign m2_87 =10'b0;

   // m2_88 = W*in
   wire signed [9:0] m2_88;
   assign m2_88 =10'b0;

   // m2_89 = W*in
   wire signed [9:0] m2_89;
   assign m2_89 =10'b0;

   // m2_90 = W*in
   wire signed [9:0] m2_90;
   assign m2_90 =10'b0;

   // m2_91 = W*in
   wire signed [9:0] m2_91;
   assign m2_91 =10'b0;

   // m2_92 = W*in
   wire signed [9:0] m2_92;
   assign m2_92 =10'b0;

   // m2_93 = W*in
   wire signed [9:0] m2_93;
   assign m2_93 =10'b0;

   // m2_94 = W*in
   wire signed [9:0] m2_94;
   assign m2_94 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_95 = W*in
   wire signed [9:0] m2_95;
   assign m2_95 ={ {4{in2[5]}} , in2[5:0] };

   // m2_96 = W*in
   wire signed [9:0] m2_96;
   assign m2_96 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_97 = W*in
   wire signed [9:0] m2_97;
   assign m2_97 =10'b0;

   // m2_98 = W*in
   wire signed [9:0] m2_98;
   assign m2_98 =10'b0;

   // m2_99 = W*in
   wire signed [9:0] m2_99;
   assign m2_99 =10'b0;

   // m2_100 = W*in
   wire signed [9:0] m2_100;
   assign m2_100 ={ {3{neg2[5]}} , neg2 , {1{1'b0}} };

   // m2_101 = W*in
   wire signed [9:0] m2_101;
   assign m2_101 =10'b0;

   // m2_102 = W*in
   wire signed [9:0] m2_102;
   assign m2_102 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_103 = W*in
   wire signed [9:0] m2_103;
   assign m2_103 =10'b0;

   // m2_104 = W*in
   wire signed [9:0] m2_104;
   assign m2_104 =10'b0;

   // m2_105 = W*in
   wire signed [9:0] m2_105;
   assign m2_105 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_106 = W*in
   wire signed [9:0] m2_106;
   assign m2_106 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_107 = W*in
   wire signed [9:0] m2_107;
   assign m2_107 =10'b0;

   // m2_108 = W*in
   wire signed [9:0] m2_108;
   assign m2_108 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_109 = W*in
   wire signed [9:0] m2_109;
   assign m2_109 ={ {5{neg2[5]}} , neg2[5:1] };

   // m2_110 = W*in
   wire signed [9:0] m2_110;
   assign m2_110 =10'b0;

   // m2_111 = W*in
   wire signed [9:0] m2_111;
   assign m2_111 =10'b0;

   // m2_112 = W*in
   wire signed [9:0] m2_112;
   assign m2_112 =10'b0;

   // m2_113 = W*in
   wire signed [9:0] m2_113;
   assign m2_113 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_114 = W*in
   wire signed [9:0] m2_114;
   assign m2_114 ={ {5{in2[5]}} , in2[5:1] };

   // m2_115 = W*in
   wire signed [9:0] m2_115;
   assign m2_115 =10'b0;

   // m2_116 = W*in
   wire signed [9:0] m2_116;
   assign m2_116 ={ {4{neg2[5]}} , neg2[5:0] };

   // m2_117 = W*in
   wire signed [9:0] m2_117;
   assign m2_117 =10'b0;

   // m3_1 = W*in
   wire signed [9:0] m3_1;
   assign m3_1 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_2 = W*in
   wire signed [9:0] m3_2;
   assign m3_2 =10'b0;

   // m3_3 = W*in
   wire signed [9:0] m3_3;
   assign m3_3 =10'b0;

   // m3_4 = W*in
   wire signed [9:0] m3_4;
   assign m3_4 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_5 = W*in
   wire signed [9:0] m3_5;
   assign m3_5 =10'b0;

   // m3_6 = W*in
   wire signed [9:0] m3_6;
   assign m3_6 ={ {5{in3[5]}} , in3[5:1] };

   // m3_7 = W*in
   wire signed [9:0] m3_7;
   assign m3_7 =10'b0;

   // m3_8 = W*in
   wire signed [9:0] m3_8;
   assign m3_8 =10'b0;

   // m3_9 = W*in
   wire signed [9:0] m3_9;
   assign m3_9 =10'b0;

   // m3_10 = W*in
   wire signed [9:0] m3_10;
   assign m3_10 =10'b0;

   // m3_11 = W*in
   wire signed [9:0] m3_11;
   assign m3_11 =10'b0;

   // m3_12 = W*in
   wire signed [9:0] m3_12;
   assign m3_12 =10'b0;

   // m3_13 = W*in
   wire signed [9:0] m3_13;
   assign m3_13 =10'b0;

   // m3_14 = W*in
   wire signed [9:0] m3_14;
   assign m3_14 =10'b0;

   // m3_15 = W*in
   wire signed [9:0] m3_15;
   assign m3_15 =10'b0;

   // m3_16 = W*in
   wire signed [9:0] m3_16;
   assign m3_16 ={ {3{neg3[5]}} , neg3 , {1{1'b0}} };

   // m3_17 = W*in
   wire signed [9:0] m3_17;
   assign m3_17 =10'b0;

   // m3_18 = W*in
   wire signed [9:0] m3_18;
   assign m3_18 ={ {5{in3[5]}} , in3[5:1] };

   // m3_19 = W*in
   wire signed [9:0] m3_19;
   assign m3_19 ={ {4{in3[5]}} , in3[5:0] };

   // m3_20 = W*in
   wire signed [9:0] m3_20;
   assign m3_20 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_21 = W*in
   wire signed [9:0] m3_21;
   assign m3_21 ={ {4{in3[5]}} , in3[5:0] };

   // m3_22 = W*in
   wire signed [9:0] m3_22;
   assign m3_22 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_23 = W*in
   wire signed [9:0] m3_23;
   assign m3_23 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_24 = W*in
   wire signed [9:0] m3_24;
   assign m3_24 =10'b0;

   // m3_25 = W*in
   wire signed [9:0] m3_25;
   assign m3_25 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_26 = W*in
   wire signed [9:0] m3_26;
   assign m3_26 =10'b0;

   // m3_27 = W*in
   wire signed [9:0] m3_27;
   assign m3_27 =10'b0;

   // m3_28 = W*in
   wire signed [9:0] m3_28;
   assign m3_28 =10'b0;

   // m3_29 = W*in
   wire signed [9:0] m3_29;
   assign m3_29 =10'b0;

   // m3_30 = W*in
   wire signed [9:0] m3_30;
   assign m3_30 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_31 = W*in
   wire signed [9:0] m3_31;
   assign m3_31 =10'b0;

   // m3_32 = W*in
   wire signed [9:0] m3_32;
   assign m3_32 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_33 = W*in
   wire signed [9:0] m3_33;
   assign m3_33 ={ {3{neg3[5]}} , neg3 , {1{1'b0}} };

   // m3_34 = W*in
   wire signed [9:0] m3_34;
   assign m3_34 ={ {4{in3[5]}} , in3[5:0] };

   // m3_35 = W*in
   wire signed [9:0] m3_35;
   assign m3_35 =10'b0;

   // m3_36 = W*in
   wire signed [9:0] m3_36;
   assign m3_36 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_37 = W*in
   wire signed [9:0] m3_37;
   assign m3_37 ={ {3{neg3[5]}} , neg3 , {1{1'b0}} };

   // m3_38 = W*in
   wire signed [9:0] m3_38;
   assign m3_38 ={ {4{in3[5]}} , in3[5:0] };

   // m3_39 = W*in
   wire signed [9:0] m3_39;
   assign m3_39 =10'b0;

   // m3_40 = W*in
   wire signed [9:0] m3_40;
   assign m3_40 =10'b0;

   // m3_41 = W*in
   wire signed [9:0] m3_41;
   assign m3_41 =10'b0;

   // m3_42 = W*in
   wire signed [9:0] m3_42;
   assign m3_42 =10'b0;

   // m3_43 = W*in
   wire signed [9:0] m3_43;
   assign m3_43 =10'b0;

   // m3_44 = W*in
   wire signed [9:0] m3_44;
   assign m3_44 =10'b0;

   // m3_45 = W*in
   wire signed [9:0] m3_45;
   assign m3_45 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_46 = W*in
   wire signed [9:0] m3_46;
   assign m3_46 =10'b0;

   // m3_47 = W*in
   wire signed [9:0] m3_47;
   assign m3_47 =10'b0;

   // m3_48 = W*in
   wire signed [9:0] m3_48;
   assign m3_48 =10'b0;

   // m3_49 = W*in
   wire signed [9:0] m3_49;
   assign m3_49 =10'b0;

   // m3_50 = W*in
   wire signed [9:0] m3_50;
   assign m3_50 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_51 = W*in
   wire signed [9:0] m3_51;
   assign m3_51 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_52 = W*in
   wire signed [9:0] m3_52;
   assign m3_52 =10'b0;

   // m3_53 = W*in
   wire signed [9:0] m3_53;
   assign m3_53 =10'b0;

   // m3_54 = W*in
   wire signed [9:0] m3_54;
   assign m3_54 =10'b0;

   // m3_55 = W*in
   wire signed [9:0] m3_55;
   assign m3_55 =10'b0;

   // m3_56 = W*in
   wire signed [9:0] m3_56;
   assign m3_56 ={ {3{neg3[5]}} , neg3 , {1{1'b0}} };

   // m3_57 = W*in
   wire signed [9:0] m3_57;
   assign m3_57 =10'b0;

   // m3_58 = W*in
   wire signed [9:0] m3_58;
   assign m3_58 ={ {4{in3[5]}} , in3[5:0] };

   // m3_59 = W*in
   wire signed [9:0] m3_59;
   assign m3_59 =10'b0;

   // m3_60 = W*in
   wire signed [9:0] m3_60;
   assign m3_60 =10'b0;

   // m3_61 = W*in
   wire signed [9:0] m3_61;
   assign m3_61 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_62 = W*in
   wire signed [9:0] m3_62;
   assign m3_62 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_63 = W*in
   wire signed [9:0] m3_63;
   assign m3_63 =10'b0;

   // m3_64 = W*in
   wire signed [9:0] m3_64;
   assign m3_64 =10'b0;

   // m3_65 = W*in
   wire signed [9:0] m3_65;
   assign m3_65 =10'b0;

   // m3_66 = W*in
   wire signed [9:0] m3_66;
   assign m3_66 =10'b0;

   // m3_67 = W*in
   wire signed [9:0] m3_67;
   assign m3_67 =10'b0;

   // m3_68 = W*in
   wire signed [9:0] m3_68;
   assign m3_68 =10'b0;

   // m3_69 = W*in
   wire signed [9:0] m3_69;
   assign m3_69 ={ {5{in3[5]}} , in3[5:1] };

   // m3_70 = W*in
   wire signed [9:0] m3_70;
   assign m3_70 =10'b0;

   // m3_71 = W*in
   wire signed [9:0] m3_71;
   assign m3_71 ={ {4{in3[5]}} , in3[5:0] };

   // m3_72 = W*in
   wire signed [9:0] m3_72;
   assign m3_72 ={ {4{in3[5]}} , in3[5:0] };

   // m3_73 = W*in
   wire signed [9:0] m3_73;
   assign m3_73 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_74 = W*in
   wire signed [9:0] m3_74;
   assign m3_74 ={ {4{in3[5]}} , in3[5:0] };

   // m3_75 = W*in
   wire signed [9:0] m3_75;
   assign m3_75 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_76 = W*in
   wire signed [9:0] m3_76;
   assign m3_76 ={ {4{in3[5]}} , in3[5:0] };

   // m3_77 = W*in
   wire signed [9:0] m3_77;
   assign m3_77 =10'b0;

   // m3_78 = W*in
   wire signed [9:0] m3_78;
   assign m3_78 =10'b0;

   // m3_79 = W*in
   wire signed [9:0] m3_79;
   assign m3_79 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_80 = W*in
   wire signed [9:0] m3_80;
   assign m3_80 =10'b0;

   // m3_81 = W*in
   wire signed [9:0] m3_81;
   assign m3_81 =10'b0;

   // m3_82 = W*in
   wire signed [9:0] m3_82;
   assign m3_82 =10'b0;

   // m3_83 = W*in
   wire signed [9:0] m3_83;
   assign m3_83 ={ {3{neg3[5]}} , neg3 , {1{1'b0}} };

   // m3_84 = W*in
   wire signed [9:0] m3_84;
   assign m3_84 =10'b0;

   // m3_85 = W*in
   wire signed [9:0] m3_85;
   assign m3_85 =10'b0;

   // m3_86 = W*in
   wire signed [9:0] m3_86;
   assign m3_86 =10'b0;

   // m3_87 = W*in
   wire signed [9:0] m3_87;
   assign m3_87 =10'b0;

   // m3_88 = W*in
   wire signed [9:0] m3_88;
   assign m3_88 ={ {4{in3[5]}} , in3[5:0] };

   // m3_89 = W*in
   wire signed [9:0] m3_89;
   assign m3_89 =10'b0;

   // m3_90 = W*in
   wire signed [9:0] m3_90;
   assign m3_90 =10'b0;

   // m3_91 = W*in
   wire signed [9:0] m3_91;
   assign m3_91 ={ {4{in3[5]}} , in3[5:0] };

   // m3_92 = W*in
   wire signed [9:0] m3_92;
   assign m3_92 ={ {3{in3[5]}} , in3 , {1{1'b0}} };

   // m3_93 = W*in
   wire signed [9:0] m3_93;
   assign m3_93 =10'b0;

   // m3_94 = W*in
   wire signed [9:0] m3_94;
   assign m3_94 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_95 = W*in
   wire signed [9:0] m3_95;
   assign m3_95 =10'b0;

   // m3_96 = W*in
   wire signed [9:0] m3_96;
   assign m3_96 =10'b0;

   // m3_97 = W*in
   wire signed [9:0] m3_97;
   assign m3_97 ={ {4{in3[5]}} , in3[5:0] };

   // m3_98 = W*in
   wire signed [9:0] m3_98;
   assign m3_98 =10'b0;

   // m3_99 = W*in
   wire signed [9:0] m3_99;
   assign m3_99 =10'b0;

   // m3_100 = W*in
   wire signed [9:0] m3_100;
   assign m3_100 =10'b0;

   // m3_101 = W*in
   wire signed [9:0] m3_101;
   assign m3_101 =10'b0;

   // m3_102 = W*in
   wire signed [9:0] m3_102;
   assign m3_102 ={ {3{neg3[5]}} , neg3 , {1{1'b0}} };

   // m3_103 = W*in
   wire signed [9:0] m3_103;
   assign m3_103 =10'b0;

   // m3_104 = W*in
   wire signed [9:0] m3_104;
   assign m3_104 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_105 = W*in
   wire signed [9:0] m3_105;
   assign m3_105 =10'b0;

   // m3_106 = W*in
   wire signed [9:0] m3_106;
   assign m3_106 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_107 = W*in
   wire signed [9:0] m3_107;
   assign m3_107 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_108 = W*in
   wire signed [9:0] m3_108;
   assign m3_108 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_109 = W*in
   wire signed [9:0] m3_109;
   assign m3_109 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_110 = W*in
   wire signed [9:0] m3_110;
   assign m3_110 =10'b0;

   // m3_111 = W*in
   wire signed [9:0] m3_111;
   assign m3_111 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_112 = W*in
   wire signed [9:0] m3_112;
   assign m3_112 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_113 = W*in
   wire signed [9:0] m3_113;
   assign m3_113 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_114 = W*in
   wire signed [9:0] m3_114;
   assign m3_114 =10'b0;

   // m3_115 = W*in
   wire signed [9:0] m3_115;
   assign m3_115 ={ {4{neg3[5]}} , neg3[5:0] };

   // m3_116 = W*in
   wire signed [9:0] m3_116;
   assign m3_116 ={ {5{neg3[5]}} , neg3[5:1] };

   // m3_117 = W*in
   wire signed [9:0] m3_117;
   assign m3_117 =10'b0;

   // m4_1 = W*in
   wire signed [9:0] m4_1;
   assign m4_1 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_2 = W*in
   wire signed [9:0] m4_2;
   assign m4_2 =10'b0;

   // m4_3 = W*in
   wire signed [9:0] m4_3;
   assign m4_3 =10'b0;

   // m4_4 = W*in
   wire signed [9:0] m4_4;
   assign m4_4 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_5 = W*in
   wire signed [9:0] m4_5;
   assign m4_5 =10'b0;

   // m4_6 = W*in
   wire signed [9:0] m4_6;
   assign m4_6 =10'b0;

   // m4_7 = W*in
   wire signed [9:0] m4_7;
   assign m4_7 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_8 = W*in
   wire signed [9:0] m4_8;
   assign m4_8 =10'b0;

   // m4_9 = W*in
   wire signed [9:0] m4_9;
   assign m4_9 =10'b0;

   // m4_10 = W*in
   wire signed [9:0] m4_10;
   assign m4_10 =10'b0;

   // m4_11 = W*in
   wire signed [9:0] m4_11;
   assign m4_11 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_12 = W*in
   wire signed [9:0] m4_12;
   assign m4_12 =10'b0;

   // m4_13 = W*in
   wire signed [9:0] m4_13;
   assign m4_13 =10'b0;

   // m4_14 = W*in
   wire signed [9:0] m4_14;
   assign m4_14 =10'b0;

   // m4_15 = W*in
   wire signed [9:0] m4_15;
   assign m4_15 ={ {4{in4[5]}} , in4[5:0] };

   // m4_16 = W*in
   wire signed [9:0] m4_16;
   assign m4_16 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_17 = W*in
   wire signed [9:0] m4_17;
   assign m4_17 =10'b0;

   // m4_18 = W*in
   wire signed [9:0] m4_18;
   assign m4_18 =10'b0;

   // m4_19 = W*in
   wire signed [9:0] m4_19;
   assign m4_19 =10'b0;

   // m4_20 = W*in
   wire signed [9:0] m4_20;
   assign m4_20 =10'b0;

   // m4_21 = W*in
   wire signed [9:0] m4_21;
   assign m4_21 =10'b0;

   // m4_22 = W*in
   wire signed [9:0] m4_22;
   assign m4_22 =10'b0;

   // m4_23 = W*in
   wire signed [9:0] m4_23;
   assign m4_23 =10'b0;

   // m4_24 = W*in
   wire signed [9:0] m4_24;
   assign m4_24 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_25 = W*in
   wire signed [9:0] m4_25;
   assign m4_25 =10'b0;

   // m4_26 = W*in
   wire signed [9:0] m4_26;
   assign m4_26 =10'b0;

   // m4_27 = W*in
   wire signed [9:0] m4_27;
   assign m4_27 =10'b0;

   // m4_28 = W*in
   wire signed [9:0] m4_28;
   assign m4_28 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_29 = W*in
   wire signed [9:0] m4_29;
   assign m4_29 =10'b0;

   // m4_30 = W*in
   wire signed [9:0] m4_30;
   assign m4_30 =10'b0;

   // m4_31 = W*in
   wire signed [9:0] m4_31;
   assign m4_31 =10'b0;

   // m4_32 = W*in
   wire signed [9:0] m4_32;
   assign m4_32 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_33 = W*in
   wire signed [9:0] m4_33;
   assign m4_33 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_34 = W*in
   wire signed [9:0] m4_34;
   assign m4_34 ={ {4{in4[5]}} , in4[5:0] };

   // m4_35 = W*in
   wire signed [9:0] m4_35;
   assign m4_35 =10'b0;

   // m4_36 = W*in
   wire signed [9:0] m4_36;
   assign m4_36 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_37 = W*in
   wire signed [9:0] m4_37;
   assign m4_37 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_38 = W*in
   wire signed [9:0] m4_38;
   assign m4_38 ={ {4{in4[5]}} , in4[5:0] };

   // m4_39 = W*in
   wire signed [9:0] m4_39;
   assign m4_39 =10'b0;

   // m4_40 = W*in
   wire signed [9:0] m4_40;
   assign m4_40 =10'b0;

   // m4_41 = W*in
   wire signed [9:0] m4_41;
   assign m4_41 =10'b0;

   // m4_42 = W*in
   wire signed [9:0] m4_42;
   assign m4_42 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_43 = W*in
   wire signed [9:0] m4_43;
   assign m4_43 =10'b0;

   // m4_44 = W*in
   wire signed [9:0] m4_44;
   assign m4_44 =10'b0;

   // m4_45 = W*in
   wire signed [9:0] m4_45;
   assign m4_45 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_46 = W*in
   wire signed [9:0] m4_46;
   assign m4_46 =10'b0;

   // m4_47 = W*in
   wire signed [9:0] m4_47;
   assign m4_47 =10'b0;

   // m4_48 = W*in
   wire signed [9:0] m4_48;
   assign m4_48 =10'b0;

   // m4_49 = W*in
   wire signed [9:0] m4_49;
   assign m4_49 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_50 = W*in
   wire signed [9:0] m4_50;
   assign m4_50 ={ {4{in4[5]}} , in4[5:0] };

   // m4_51 = W*in
   wire signed [9:0] m4_51;
   assign m4_51 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_52 = W*in
   wire signed [9:0] m4_52;
   assign m4_52 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_53 = W*in
   wire signed [9:0] m4_53;
   assign m4_53 =10'b0;

   // m4_54 = W*in
   wire signed [9:0] m4_54;
   assign m4_54 =10'b0;

   // m4_55 = W*in
   wire signed [9:0] m4_55;
   assign m4_55 =10'b0;

   // m4_56 = W*in
   wire signed [9:0] m4_56;
   assign m4_56 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_57 = W*in
   wire signed [9:0] m4_57;
   assign m4_57 =10'b0;

   // m4_58 = W*in
   wire signed [9:0] m4_58;
   assign m4_58 =10'b0;

   // m4_59 = W*in
   wire signed [9:0] m4_59;
   assign m4_59 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_60 = W*in
   wire signed [9:0] m4_60;
   assign m4_60 =10'b0;

   // m4_61 = W*in
   wire signed [9:0] m4_61;
   assign m4_61 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_62 = W*in
   wire signed [9:0] m4_62;
   assign m4_62 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_63 = W*in
   wire signed [9:0] m4_63;
   assign m4_63 =10'b0;

   // m4_64 = W*in
   wire signed [9:0] m4_64;
   assign m4_64 =10'b0;

   // m4_65 = W*in
   wire signed [9:0] m4_65;
   assign m4_65 =10'b0;

   // m4_66 = W*in
   wire signed [9:0] m4_66;
   assign m4_66 =10'b0;

   // m4_67 = W*in
   wire signed [9:0] m4_67;
   assign m4_67 =10'b0;

   // m4_68 = W*in
   wire signed [9:0] m4_68;
   assign m4_68 =10'b0;

   // m4_69 = W*in
   wire signed [9:0] m4_69;
   assign m4_69 ={ {4{in4[5]}} , in4[5:0] };

   // m4_70 = W*in
   wire signed [9:0] m4_70;
   assign m4_70 ={ {4{in4[5]}} , in4[5:0] };

   // m4_71 = W*in
   wire signed [9:0] m4_71;
   assign m4_71 ={ {4{in4[5]}} , in4[5:0] };

   // m4_72 = W*in
   wire signed [9:0] m4_72;
   assign m4_72 ={ {3{in4[5]}} , in4 , {1{1'b0}} };

   // m4_73 = W*in
   wire signed [9:0] m4_73;
   assign m4_73 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_74 = W*in
   wire signed [9:0] m4_74;
   assign m4_74 ={ {4{in4[5]}} , in4[5:0] };

   // m4_75 = W*in
   wire signed [9:0] m4_75;
   assign m4_75 =10'b0;

   // m4_76 = W*in
   wire signed [9:0] m4_76;
   assign m4_76 ={ {4{in4[5]}} , in4[5:0] };

   // m4_77 = W*in
   wire signed [9:0] m4_77;
   assign m4_77 =10'b0;

   // m4_78 = W*in
   wire signed [9:0] m4_78;
   assign m4_78 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_79 = W*in
   wire signed [9:0] m4_79;
   assign m4_79 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_80 = W*in
   wire signed [9:0] m4_80;
   assign m4_80 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_81 = W*in
   wire signed [9:0] m4_81;
   assign m4_81 =10'b0;

   // m4_82 = W*in
   wire signed [9:0] m4_82;
   assign m4_82 =10'b0;

   // m4_83 = W*in
   wire signed [9:0] m4_83;
   assign m4_83 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_84 = W*in
   wire signed [9:0] m4_84;
   assign m4_84 ={ {4{in4[5]}} , in4[5:0] };

   // m4_85 = W*in
   wire signed [9:0] m4_85;
   assign m4_85 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_86 = W*in
   wire signed [9:0] m4_86;
   assign m4_86 =10'b0;

   // m4_87 = W*in
   wire signed [9:0] m4_87;
   assign m4_87 ={ {4{in4[5]}} , in4[5:0] };

   // m4_88 = W*in
   wire signed [9:0] m4_88;
   assign m4_88 ={ {4{in4[5]}} , in4[5:0] };

   // m4_89 = W*in
   wire signed [9:0] m4_89;
   assign m4_89 =10'b0;

   // m4_90 = W*in
   wire signed [9:0] m4_90;
   assign m4_90 ={ {4{in4[5]}} , in4[5:0] };

   // m4_91 = W*in
   wire signed [9:0] m4_91;
   assign m4_91 =10'b0;

   // m4_92 = W*in
   wire signed [9:0] m4_92;
   assign m4_92 =10'b0;

   // m4_93 = W*in
   wire signed [9:0] m4_93;
   assign m4_93 =10'b0;

   // m4_94 = W*in
   wire signed [9:0] m4_94;
   assign m4_94 =10'b0;

   // m4_95 = W*in
   wire signed [9:0] m4_95;
   assign m4_95 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_96 = W*in
   wire signed [9:0] m4_96;
   assign m4_96 =10'b0;

   // m4_97 = W*in
   wire signed [9:0] m4_97;
   assign m4_97 ={ {4{in4[5]}} , in4[5:0] };

   // m4_98 = W*in
   wire signed [9:0] m4_98;
   assign m4_98 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_99 = W*in
   wire signed [9:0] m4_99;
   assign m4_99 ={ {4{in4[5]}} , in4[5:0] };

   // m4_100 = W*in
   wire signed [9:0] m4_100;
   assign m4_100 =10'b0;

   // m4_101 = W*in
   wire signed [9:0] m4_101;
   assign m4_101 =10'b0;

   // m4_102 = W*in
   wire signed [9:0] m4_102;
   assign m4_102 ={ {3{neg4[5]}} , neg4 , {1{1'b0}} };

   // m4_103 = W*in
   wire signed [9:0] m4_103;
   assign m4_103 ={ {4{in4[5]}} , in4[5:0] };

   // m4_104 = W*in
   wire signed [9:0] m4_104;
   assign m4_104 ={ {4{in4[5]}} , in4[5:0] };

   // m4_105 = W*in
   wire signed [9:0] m4_105;
   assign m4_105 =10'b0;

   // m4_106 = W*in
   wire signed [9:0] m4_106;
   assign m4_106 ={ {4{neg4[5]}} , neg4[5:0] };

   // m4_107 = W*in
   wire signed [9:0] m4_107;
   assign m4_107 =10'b0;

   // m4_108 = W*in
   wire signed [9:0] m4_108;
   assign m4_108 =10'b0;

   // m4_109 = W*in
   wire signed [9:0] m4_109;
   assign m4_109 =10'b0;

   // m4_110 = W*in
   wire signed [9:0] m4_110;
   assign m4_110 ={ {5{neg4[5]}} , neg4[5:1] };

   // m4_111 = W*in
   wire signed [9:0] m4_111;
   assign m4_111 =10'b0;

   // m4_112 = W*in
   wire signed [9:0] m4_112;
   assign m4_112 ={ {5{neg4[5]}} , neg4[5:1] };

   // m4_113 = W*in
   wire signed [9:0] m4_113;
   assign m4_113 ={ {5{neg4[5]}} , neg4[5:1] };

   // m4_114 = W*in
   wire signed [9:0] m4_114;
   assign m4_114 ={ {4{in4[5]}} , in4[5:0] };

   // m4_115 = W*in
   wire signed [9:0] m4_115;
   assign m4_115 =10'b0;

   // m4_116 = W*in
   wire signed [9:0] m4_116;
   assign m4_116 =10'b0;

   // m4_117 = W*in
   wire signed [9:0] m4_117;
   assign m4_117 =10'b0;

   // m5_1 = W*in
   wire signed [9:0] m5_1;
   assign m5_1 =10'b0;

   // m5_2 = W*in
   wire signed [9:0] m5_2;
   assign m5_2 =10'b0;

   // m5_3 = W*in
   wire signed [9:0] m5_3;
   assign m5_3 =10'b0;

   // m5_4 = W*in
   wire signed [9:0] m5_4;
   assign m5_4 =10'b0;

   // m5_5 = W*in
   wire signed [9:0] m5_5;
   assign m5_5 =10'b0;

   // m5_6 = W*in
   wire signed [9:0] m5_6;
   assign m5_6 =10'b0;

   // m5_7 = W*in
   wire signed [9:0] m5_7;
   assign m5_7 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_8 = W*in
   wire signed [9:0] m5_8;
   assign m5_8 =10'b0;

   // m5_9 = W*in
   wire signed [9:0] m5_9;
   assign m5_9 =10'b0;

   // m5_10 = W*in
   wire signed [9:0] m5_10;
   assign m5_10 =10'b0;

   // m5_11 = W*in
   wire signed [9:0] m5_11;
   assign m5_11 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_12 = W*in
   wire signed [9:0] m5_12;
   assign m5_12 =10'b0;

   // m5_13 = W*in
   wire signed [9:0] m5_13;
   assign m5_13 =10'b0;

   // m5_14 = W*in
   wire signed [9:0] m5_14;
   assign m5_14 =10'b0;

   // m5_15 = W*in
   wire signed [9:0] m5_15;
   assign m5_15 =10'b0;

   // m5_16 = W*in
   wire signed [9:0] m5_16;
   assign m5_16 =10'b0;

   // m5_17 = W*in
   wire signed [9:0] m5_17;
   assign m5_17 =10'b0;

   // m5_18 = W*in
   wire signed [9:0] m5_18;
   assign m5_18 =10'b0;

   // m5_19 = W*in
   wire signed [9:0] m5_19;
   assign m5_19 =10'b0;

   // m5_20 = W*in
   wire signed [9:0] m5_20;
   assign m5_20 =10'b0;

   // m5_21 = W*in
   wire signed [9:0] m5_21;
   assign m5_21 =10'b0;

   // m5_22 = W*in
   wire signed [9:0] m5_22;
   assign m5_22 =10'b0;

   // m5_23 = W*in
   wire signed [9:0] m5_23;
   assign m5_23 ={ {4{in5[5]}} , in5[5:0] };

   // m5_24 = W*in
   wire signed [9:0] m5_24;
   assign m5_24 =10'b0;

   // m5_25 = W*in
   wire signed [9:0] m5_25;
   assign m5_25 =10'b0;

   // m5_26 = W*in
   wire signed [9:0] m5_26;
   assign m5_26 =10'b0;

   // m5_27 = W*in
   wire signed [9:0] m5_27;
   assign m5_27 =10'b0;

   // m5_28 = W*in
   wire signed [9:0] m5_28;
   assign m5_28 =10'b0;

   // m5_29 = W*in
   wire signed [9:0] m5_29;
   assign m5_29 =10'b0;

   // m5_30 = W*in
   wire signed [9:0] m5_30;
   assign m5_30 =10'b0;

   // m5_31 = W*in
   wire signed [9:0] m5_31;
   assign m5_31 =10'b0;

   // m5_32 = W*in
   wire signed [9:0] m5_32;
   assign m5_32 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_33 = W*in
   wire signed [9:0] m5_33;
   assign m5_33 =10'b0;

   // m5_34 = W*in
   wire signed [9:0] m5_34;
   assign m5_34 =10'b0;

   // m5_35 = W*in
   wire signed [9:0] m5_35;
   assign m5_35 =10'b0;

   // m5_36 = W*in
   wire signed [9:0] m5_36;
   assign m5_36 ={ {5{neg5[5]}} , neg5[5:1] };

   // m5_37 = W*in
   wire signed [9:0] m5_37;
   assign m5_37 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_38 = W*in
   wire signed [9:0] m5_38;
   assign m5_38 =10'b0;

   // m5_39 = W*in
   wire signed [9:0] m5_39;
   assign m5_39 =10'b0;

   // m5_40 = W*in
   wire signed [9:0] m5_40;
   assign m5_40 =10'b0;

   // m5_41 = W*in
   wire signed [9:0] m5_41;
   assign m5_41 =10'b0;

   // m5_42 = W*in
   wire signed [9:0] m5_42;
   assign m5_42 =10'b0;

   // m5_43 = W*in
   wire signed [9:0] m5_43;
   assign m5_43 =10'b0;

   // m5_44 = W*in
   wire signed [9:0] m5_44;
   assign m5_44 =10'b0;

   // m5_45 = W*in
   wire signed [9:0] m5_45;
   assign m5_45 =10'b0;

   // m5_46 = W*in
   wire signed [9:0] m5_46;
   assign m5_46 =10'b0;

   // m5_47 = W*in
   wire signed [9:0] m5_47;
   assign m5_47 =10'b0;

   // m5_48 = W*in
   wire signed [9:0] m5_48;
   assign m5_48 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_49 = W*in
   wire signed [9:0] m5_49;
   assign m5_49 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_50 = W*in
   wire signed [9:0] m5_50;
   assign m5_50 =10'b0;

   // m5_51 = W*in
   wire signed [9:0] m5_51;
   assign m5_51 =10'b0;

   // m5_52 = W*in
   wire signed [9:0] m5_52;
   assign m5_52 =10'b0;

   // m5_53 = W*in
   wire signed [9:0] m5_53;
   assign m5_53 =10'b0;

   // m5_54 = W*in
   wire signed [9:0] m5_54;
   assign m5_54 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_55 = W*in
   wire signed [9:0] m5_55;
   assign m5_55 =10'b0;

   // m5_56 = W*in
   wire signed [9:0] m5_56;
   assign m5_56 =10'b0;

   // m5_57 = W*in
   wire signed [9:0] m5_57;
   assign m5_57 =10'b0;

   // m5_58 = W*in
   wire signed [9:0] m5_58;
   assign m5_58 =10'b0;

   // m5_59 = W*in
   wire signed [9:0] m5_59;
   assign m5_59 =10'b0;

   // m5_60 = W*in
   wire signed [9:0] m5_60;
   assign m5_60 =10'b0;

   // m5_61 = W*in
   wire signed [9:0] m5_61;
   assign m5_61 ={ {3{neg5[5]}} , neg5 , {1{1'b0}} };

   // m5_62 = W*in
   wire signed [9:0] m5_62;
   assign m5_62 =10'b0;

   // m5_63 = W*in
   wire signed [9:0] m5_63;
   assign m5_63 =10'b0;

   // m5_64 = W*in
   wire signed [9:0] m5_64;
   assign m5_64 ={ {4{in5[5]}} , in5[5:0] };

   // m5_65 = W*in
   wire signed [9:0] m5_65;
   assign m5_65 ={ {4{in5[5]}} , in5[5:0] };

   // m5_66 = W*in
   wire signed [9:0] m5_66;
   assign m5_66 =10'b0;

   // m5_67 = W*in
   wire signed [9:0] m5_67;
   assign m5_67 =10'b0;

   // m5_68 = W*in
   wire signed [9:0] m5_68;
   assign m5_68 =10'b0;

   // m5_69 = W*in
   wire signed [9:0] m5_69;
   assign m5_69 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_70 = W*in
   wire signed [9:0] m5_70;
   assign m5_70 =10'b0;

   // m5_71 = W*in
   wire signed [9:0] m5_71;
   assign m5_71 =10'b0;

   // m5_72 = W*in
   wire signed [9:0] m5_72;
   assign m5_72 ={ {5{neg5[5]}} , neg5[5:1] };

   // m5_73 = W*in
   wire signed [9:0] m5_73;
   assign m5_73 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_74 = W*in
   wire signed [9:0] m5_74;
   assign m5_74 =10'b0;

   // m5_75 = W*in
   wire signed [9:0] m5_75;
   assign m5_75 =10'b0;

   // m5_76 = W*in
   wire signed [9:0] m5_76;
   assign m5_76 =10'b0;

   // m5_77 = W*in
   wire signed [9:0] m5_77;
   assign m5_77 =10'b0;

   // m5_78 = W*in
   wire signed [9:0] m5_78;
   assign m5_78 =10'b0;

   // m5_79 = W*in
   wire signed [9:0] m5_79;
   assign m5_79 =10'b0;

   // m5_80 = W*in
   wire signed [9:0] m5_80;
   assign m5_80 =10'b0;

   // m5_81 = W*in
   wire signed [9:0] m5_81;
   assign m5_81 ={ {4{in5[5]}} , in5[5:0] };

   // m5_82 = W*in
   wire signed [9:0] m5_82;
   assign m5_82 =10'b0;

   // m5_83 = W*in
   wire signed [9:0] m5_83;
   assign m5_83 =10'b0;

   // m5_84 = W*in
   wire signed [9:0] m5_84;
   assign m5_84 =10'b0;

   // m5_85 = W*in
   wire signed [9:0] m5_85;
   assign m5_85 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_86 = W*in
   wire signed [9:0] m5_86;
   assign m5_86 =10'b0;

   // m5_87 = W*in
   wire signed [9:0] m5_87;
   assign m5_87 =10'b0;

   // m5_88 = W*in
   wire signed [9:0] m5_88;
   assign m5_88 =10'b0;

   // m5_89 = W*in
   wire signed [9:0] m5_89;
   assign m5_89 =10'b0;

   // m5_90 = W*in
   wire signed [9:0] m5_90;
   assign m5_90 =10'b0;

   // m5_91 = W*in
   wire signed [9:0] m5_91;
   assign m5_91 =10'b0;

   // m5_92 = W*in
   wire signed [9:0] m5_92;
   assign m5_92 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_93 = W*in
   wire signed [9:0] m5_93;
   assign m5_93 =10'b0;

   // m5_94 = W*in
   wire signed [9:0] m5_94;
   assign m5_94 =10'b0;

   // m5_95 = W*in
   wire signed [9:0] m5_95;
   assign m5_95 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_96 = W*in
   wire signed [9:0] m5_96;
   assign m5_96 =10'b0;

   // m5_97 = W*in
   wire signed [9:0] m5_97;
   assign m5_97 ={ {4{neg5[5]}} , neg5[5:0] };

   // m5_98 = W*in
   wire signed [9:0] m5_98;
   assign m5_98 =10'b0;

   // m5_99 = W*in
   wire signed [9:0] m5_99;
   assign m5_99 =10'b0;

   // m5_100 = W*in
   wire signed [9:0] m5_100;
   assign m5_100 =10'b0;

   // m5_101 = W*in
   wire signed [9:0] m5_101;
   assign m5_101 =10'b0;

   // m5_102 = W*in
   wire signed [9:0] m5_102;
   assign m5_102 =10'b0;

   // m5_103 = W*in
   wire signed [9:0] m5_103;
   assign m5_103 =10'b0;

   // m5_104 = W*in
   wire signed [9:0] m5_104;
   assign m5_104 =10'b0;

   // m5_105 = W*in
   wire signed [9:0] m5_105;
   assign m5_105 =10'b0;

   // m5_106 = W*in
   wire signed [9:0] m5_106;
   assign m5_106 =10'b0;

   // m5_107 = W*in
   wire signed [9:0] m5_107;
   assign m5_107 =10'b0;

   // m5_108 = W*in
   wire signed [9:0] m5_108;
   assign m5_108 =10'b0;

   // m5_109 = W*in
   wire signed [9:0] m5_109;
   assign m5_109 =10'b0;

   // m5_110 = W*in
   wire signed [9:0] m5_110;
   assign m5_110 =10'b0;

   // m5_111 = W*in
   wire signed [9:0] m5_111;
   assign m5_111 =10'b0;

   // m5_112 = W*in
   wire signed [9:0] m5_112;
   assign m5_112 ={ {4{in5[5]}} , in5[5:0] };

   // m5_113 = W*in
   wire signed [9:0] m5_113;
   assign m5_113 =10'b0;

   // m5_114 = W*in
   wire signed [9:0] m5_114;
   assign m5_114 =10'b0;

   // m5_115 = W*in
   wire signed [9:0] m5_115;
   assign m5_115 =10'b0;

   // m5_116 = W*in
   wire signed [9:0] m5_116;
   assign m5_116 =10'b0;

   // m5_117 = W*in
   wire signed [9:0] m5_117;
   assign m5_117 ={ {4{neg5[5]}} , neg5[5:0] };

   // m6_1 = W*in
   wire signed [9:0] m6_1;
   assign m6_1 =10'b0;

   // m6_2 = W*in
   wire signed [9:0] m6_2;
   assign m6_2 ={ {4{in6[5]}} , in6[5:0] };

   // m6_3 = W*in
   wire signed [9:0] m6_3;
   assign m6_3 =10'b0;

   // m6_4 = W*in
   wire signed [9:0] m6_4;
   assign m6_4 =10'b0;

   // m6_5 = W*in
   wire signed [9:0] m6_5;
   assign m6_5 =10'b0;

   // m6_6 = W*in
   wire signed [9:0] m6_6;
   assign m6_6 =10'b0;

   // m6_7 = W*in
   wire signed [9:0] m6_7;
   assign m6_7 =10'b0;

   // m6_8 = W*in
   wire signed [9:0] m6_8;
   assign m6_8 ={ {4{in6[5]}} , in6[5:0] };

   // m6_9 = W*in
   wire signed [9:0] m6_9;
   assign m6_9 =10'b0;

   // m6_10 = W*in
   wire signed [9:0] m6_10;
   assign m6_10 =10'b0;

   // m6_11 = W*in
   wire signed [9:0] m6_11;
   assign m6_11 =10'b0;

   // m6_12 = W*in
   wire signed [9:0] m6_12;
   assign m6_12 =10'b0;

   // m6_13 = W*in
   wire signed [9:0] m6_13;
   assign m6_13 =10'b0;

   // m6_14 = W*in
   wire signed [9:0] m6_14;
   assign m6_14 =10'b0;

   // m6_15 = W*in
   wire signed [9:0] m6_15;
   assign m6_15 =10'b0;

   // m6_16 = W*in
   wire signed [9:0] m6_16;
   assign m6_16 =10'b0;

   // m6_17 = W*in
   wire signed [9:0] m6_17;
   assign m6_17 ={ {5{in6[5]}} , in6[5:1] };

   // m6_18 = W*in
   wire signed [9:0] m6_18;
   assign m6_18 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_19 = W*in
   wire signed [9:0] m6_19;
   assign m6_19 =10'b0;

   // m6_20 = W*in
   wire signed [9:0] m6_20;
   assign m6_20 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_21 = W*in
   wire signed [9:0] m6_21;
   assign m6_21 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_22 = W*in
   wire signed [9:0] m6_22;
   assign m6_22 =10'b0;

   // m6_23 = W*in
   wire signed [9:0] m6_23;
   assign m6_23 =10'b0;

   // m6_24 = W*in
   wire signed [9:0] m6_24;
   assign m6_24 =10'b0;

   // m6_25 = W*in
   wire signed [9:0] m6_25;
   assign m6_25 ={ {4{in6[5]}} , in6[5:0] };

   // m6_26 = W*in
   wire signed [9:0] m6_26;
   assign m6_26 ={ {4{neg6[5]}} , neg6[5:0] };

   // m6_27 = W*in
   wire signed [9:0] m6_27;
   assign m6_27 ={ {5{in6[5]}} , in6[5:1] };

   // m6_28 = W*in
   wire signed [9:0] m6_28;
   assign m6_28 =10'b0;

   // m6_29 = W*in
   wire signed [9:0] m6_29;
   assign m6_29 =10'b0;

   // m6_30 = W*in
   wire signed [9:0] m6_30;
   assign m6_30 =10'b0;

   // m6_31 = W*in
   wire signed [9:0] m6_31;
   assign m6_31 ={ {4{in6[5]}} , in6[5:0] };

   // m6_32 = W*in
   wire signed [9:0] m6_32;
   assign m6_32 =10'b0;

   // m6_33 = W*in
   wire signed [9:0] m6_33;
   assign m6_33 =10'b0;

   // m6_34 = W*in
   wire signed [9:0] m6_34;
   assign m6_34 =10'b0;

   // m6_35 = W*in
   wire signed [9:0] m6_35;
   assign m6_35 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_36 = W*in
   wire signed [9:0] m6_36;
   assign m6_36 ={ {4{in6[5]}} , in6[5:0] };

   // m6_37 = W*in
   wire signed [9:0] m6_37;
   assign m6_37 =10'b0;

   // m6_38 = W*in
   wire signed [9:0] m6_38;
   assign m6_38 =10'b0;

   // m6_39 = W*in
   wire signed [9:0] m6_39;
   assign m6_39 =10'b0;

   // m6_40 = W*in
   wire signed [9:0] m6_40;
   assign m6_40 =10'b0;

   // m6_41 = W*in
   wire signed [9:0] m6_41;
   assign m6_41 ={ {4{neg6[5]}} , neg6[5:0] };

   // m6_42 = W*in
   wire signed [9:0] m6_42;
   assign m6_42 =10'b0;

   // m6_43 = W*in
   wire signed [9:0] m6_43;
   assign m6_43 =10'b0;

   // m6_44 = W*in
   wire signed [9:0] m6_44;
   assign m6_44 =10'b0;

   // m6_45 = W*in
   wire signed [9:0] m6_45;
   assign m6_45 =10'b0;

   // m6_46 = W*in
   wire signed [9:0] m6_46;
   assign m6_46 =10'b0;

   // m6_47 = W*in
   wire signed [9:0] m6_47;
   assign m6_47 =10'b0;

   // m6_48 = W*in
   wire signed [9:0] m6_48;
   assign m6_48 =10'b0;

   // m6_49 = W*in
   wire signed [9:0] m6_49;
   assign m6_49 =10'b0;

   // m6_50 = W*in
   wire signed [9:0] m6_50;
   assign m6_50 =10'b0;

   // m6_51 = W*in
   wire signed [9:0] m6_51;
   assign m6_51 =10'b0;

   // m6_52 = W*in
   wire signed [9:0] m6_52;
   assign m6_52 ={ {4{in6[5]}} , in6[5:0] };

   // m6_53 = W*in
   wire signed [9:0] m6_53;
   assign m6_53 ={ {4{in6[5]}} , in6[5:0] };

   // m6_54 = W*in
   wire signed [9:0] m6_54;
   assign m6_54 =10'b0;

   // m6_55 = W*in
   wire signed [9:0] m6_55;
   assign m6_55 =10'b0;

   // m6_56 = W*in
   wire signed [9:0] m6_56;
   assign m6_56 =10'b0;

   // m6_57 = W*in
   wire signed [9:0] m6_57;
   assign m6_57 =10'b0;

   // m6_58 = W*in
   wire signed [9:0] m6_58;
   assign m6_58 =10'b0;

   // m6_59 = W*in
   wire signed [9:0] m6_59;
   assign m6_59 ={ {4{in6[5]}} , in6[5:0] };

   // m6_60 = W*in
   wire signed [9:0] m6_60;
   assign m6_60 =10'b0;

   // m6_61 = W*in
   wire signed [9:0] m6_61;
   assign m6_61 =10'b0;

   // m6_62 = W*in
   wire signed [9:0] m6_62;
   assign m6_62 =10'b0;

   // m6_63 = W*in
   wire signed [9:0] m6_63;
   assign m6_63 =10'b0;

   // m6_64 = W*in
   wire signed [9:0] m6_64;
   assign m6_64 =10'b0;

   // m6_65 = W*in
   wire signed [9:0] m6_65;
   assign m6_65 =10'b0;

   // m6_66 = W*in
   wire signed [9:0] m6_66;
   assign m6_66 =10'b0;

   // m6_67 = W*in
   wire signed [9:0] m6_67;
   assign m6_67 =10'b0;

   // m6_68 = W*in
   wire signed [9:0] m6_68;
   assign m6_68 ={ {4{in6[5]}} , in6[5:0] };

   // m6_69 = W*in
   wire signed [9:0] m6_69;
   assign m6_69 =10'b0;

   // m6_70 = W*in
   wire signed [9:0] m6_70;
   assign m6_70 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_71 = W*in
   wire signed [9:0] m6_71;
   assign m6_71 =10'b0;

   // m6_72 = W*in
   wire signed [9:0] m6_72;
   assign m6_72 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_73 = W*in
   wire signed [9:0] m6_73;
   assign m6_73 ={ {4{in6[5]}} , in6[5:0] };

   // m6_74 = W*in
   wire signed [9:0] m6_74;
   assign m6_74 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_75 = W*in
   wire signed [9:0] m6_75;
   assign m6_75 =10'b0;

   // m6_76 = W*in
   wire signed [9:0] m6_76;
   assign m6_76 =10'b0;

   // m6_77 = W*in
   wire signed [9:0] m6_77;
   assign m6_77 =10'b0;

   // m6_78 = W*in
   wire signed [9:0] m6_78;
   assign m6_78 =10'b0;

   // m6_79 = W*in
   wire signed [9:0] m6_79;
   assign m6_79 =10'b0;

   // m6_80 = W*in
   wire signed [9:0] m6_80;
   assign m6_80 ={ {4{in6[5]}} , in6[5:0] };

   // m6_81 = W*in
   wire signed [9:0] m6_81;
   assign m6_81 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_82 = W*in
   wire signed [9:0] m6_82;
   assign m6_82 =10'b0;

   // m6_83 = W*in
   wire signed [9:0] m6_83;
   assign m6_83 =10'b0;

   // m6_84 = W*in
   wire signed [9:0] m6_84;
   assign m6_84 =10'b0;

   // m6_85 = W*in
   wire signed [9:0] m6_85;
   assign m6_85 =10'b0;

   // m6_86 = W*in
   wire signed [9:0] m6_86;
   assign m6_86 =10'b0;

   // m6_87 = W*in
   wire signed [9:0] m6_87;
   assign m6_87 =10'b0;

   // m6_88 = W*in
   wire signed [9:0] m6_88;
   assign m6_88 =10'b0;

   // m6_89 = W*in
   wire signed [9:0] m6_89;
   assign m6_89 =10'b0;

   // m6_90 = W*in
   wire signed [9:0] m6_90;
   assign m6_90 =10'b0;

   // m6_91 = W*in
   wire signed [9:0] m6_91;
   assign m6_91 =10'b0;

   // m6_92 = W*in
   wire signed [9:0] m6_92;
   assign m6_92 =10'b0;

   // m6_93 = W*in
   wire signed [9:0] m6_93;
   assign m6_93 =10'b0;

   // m6_94 = W*in
   wire signed [9:0] m6_94;
   assign m6_94 =10'b0;

   // m6_95 = W*in
   wire signed [9:0] m6_95;
   assign m6_95 =10'b0;

   // m6_96 = W*in
   wire signed [9:0] m6_96;
   assign m6_96 =10'b0;

   // m6_97 = W*in
   wire signed [9:0] m6_97;
   assign m6_97 =10'b0;

   // m6_98 = W*in
   wire signed [9:0] m6_98;
   assign m6_98 ={ {4{in6[5]}} , in6[5:0] };

   // m6_99 = W*in
   wire signed [9:0] m6_99;
   assign m6_99 =10'b0;

   // m6_100 = W*in
   wire signed [9:0] m6_100;
   assign m6_100 =10'b0;

   // m6_101 = W*in
   wire signed [9:0] m6_101;
   assign m6_101 =10'b0;

   // m6_102 = W*in
   wire signed [9:0] m6_102;
   assign m6_102 =10'b0;

   // m6_103 = W*in
   wire signed [9:0] m6_103;
   assign m6_103 =10'b0;

   // m6_104 = W*in
   wire signed [9:0] m6_104;
   assign m6_104 =10'b0;

   // m6_105 = W*in
   wire signed [9:0] m6_105;
   assign m6_105 ={ {4{in6[5]}} , in6[5:0] };

   // m6_106 = W*in
   wire signed [9:0] m6_106;
   assign m6_106 =10'b0;

   // m6_107 = W*in
   wire signed [9:0] m6_107;
   assign m6_107 =10'b0;

   // m6_108 = W*in
   wire signed [9:0] m6_108;
   assign m6_108 ={ {4{neg6[5]}} , neg6[5:0] };

   // m6_109 = W*in
   wire signed [9:0] m6_109;
   assign m6_109 =10'b0;

   // m6_110 = W*in
   wire signed [9:0] m6_110;
   assign m6_110 =10'b0;

   // m6_111 = W*in
   wire signed [9:0] m6_111;
   assign m6_111 =10'b0;

   // m6_112 = W*in
   wire signed [9:0] m6_112;
   assign m6_112 =10'b0;

   // m6_113 = W*in
   wire signed [9:0] m6_113;
   assign m6_113 =10'b0;

   // m6_114 = W*in
   wire signed [9:0] m6_114;
   assign m6_114 =10'b0;

   // m6_115 = W*in
   wire signed [9:0] m6_115;
   assign m6_115 =10'b0;

   // m6_116 = W*in
   wire signed [9:0] m6_116;
   assign m6_116 ={ {5{neg6[5]}} , neg6[5:1] };

   // m6_117 = W*in
   wire signed [9:0] m6_117;
   assign m6_117 =10'b0;

   // m7_1 = W*in
   wire signed [9:0] m7_1;
   assign m7_1 =10'b0;

   // m7_2 = W*in
   wire signed [9:0] m7_2;
   assign m7_2 =10'b0;

   // m7_3 = W*in
   wire signed [9:0] m7_3;
   assign m7_3 =10'b0;

   // m7_4 = W*in
   wire signed [9:0] m7_4;
   assign m7_4 =10'b0;

   // m7_5 = W*in
   wire signed [9:0] m7_5;
   assign m7_5 =10'b0;

   // m7_6 = W*in
   wire signed [9:0] m7_6;
   assign m7_6 =10'b0;

   // m7_7 = W*in
   wire signed [9:0] m7_7;
   assign m7_7 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_8 = W*in
   wire signed [9:0] m7_8;
   assign m7_8 ={ {4{in7[5]}} , in7[5:0] };

   // m7_9 = W*in
   wire signed [9:0] m7_9;
   assign m7_9 =10'b0;

   // m7_10 = W*in
   wire signed [9:0] m7_10;
   assign m7_10 =10'b0;

   // m7_11 = W*in
   wire signed [9:0] m7_11;
   assign m7_11 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_12 = W*in
   wire signed [9:0] m7_12;
   assign m7_12 =10'b0;

   // m7_13 = W*in
   wire signed [9:0] m7_13;
   assign m7_13 =10'b0;

   // m7_14 = W*in
   wire signed [9:0] m7_14;
   assign m7_14 =10'b0;

   // m7_15 = W*in
   wire signed [9:0] m7_15;
   assign m7_15 ={ {4{in7[5]}} , in7[5:0] };

   // m7_16 = W*in
   wire signed [9:0] m7_16;
   assign m7_16 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_17 = W*in
   wire signed [9:0] m7_17;
   assign m7_17 ={ {5{in7[5]}} , in7[5:1] };

   // m7_18 = W*in
   wire signed [9:0] m7_18;
   assign m7_18 =10'b0;

   // m7_19 = W*in
   wire signed [9:0] m7_19;
   assign m7_19 =10'b0;

   // m7_20 = W*in
   wire signed [9:0] m7_20;
   assign m7_20 ={ {5{neg7[5]}} , neg7[5:1] };

   // m7_21 = W*in
   wire signed [9:0] m7_21;
   assign m7_21 ={ {5{neg7[5]}} , neg7[5:1] };

   // m7_22 = W*in
   wire signed [9:0] m7_22;
   assign m7_22 =10'b0;

   // m7_23 = W*in
   wire signed [9:0] m7_23;
   assign m7_23 =10'b0;

   // m7_24 = W*in
   wire signed [9:0] m7_24;
   assign m7_24 =10'b0;

   // m7_25 = W*in
   wire signed [9:0] m7_25;
   assign m7_25 =10'b0;

   // m7_26 = W*in
   wire signed [9:0] m7_26;
   assign m7_26 ={ {5{neg7[5]}} , neg7[5:1] };

   // m7_27 = W*in
   wire signed [9:0] m7_27;
   assign m7_27 =10'b0;

   // m7_28 = W*in
   wire signed [9:0] m7_28;
   assign m7_28 =10'b0;

   // m7_29 = W*in
   wire signed [9:0] m7_29;
   assign m7_29 =10'b0;

   // m7_30 = W*in
   wire signed [9:0] m7_30;
   assign m7_30 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_31 = W*in
   wire signed [9:0] m7_31;
   assign m7_31 ={ {4{in7[5]}} , in7[5:0] };

   // m7_32 = W*in
   wire signed [9:0] m7_32;
   assign m7_32 =10'b0;

   // m7_33 = W*in
   wire signed [9:0] m7_33;
   assign m7_33 =10'b0;

   // m7_34 = W*in
   wire signed [9:0] m7_34;
   assign m7_34 ={ {4{in7[5]}} , in7[5:0] };

   // m7_35 = W*in
   wire signed [9:0] m7_35;
   assign m7_35 ={ {5{neg7[5]}} , neg7[5:1] };

   // m7_36 = W*in
   wire signed [9:0] m7_36;
   assign m7_36 =10'b0;

   // m7_37 = W*in
   wire signed [9:0] m7_37;
   assign m7_37 =10'b0;

   // m7_38 = W*in
   wire signed [9:0] m7_38;
   assign m7_38 ={ {4{in7[5]}} , in7[5:0] };

   // m7_39 = W*in
   wire signed [9:0] m7_39;
   assign m7_39 =10'b0;

   // m7_40 = W*in
   wire signed [9:0] m7_40;
   assign m7_40 =10'b0;

   // m7_41 = W*in
   wire signed [9:0] m7_41;
   assign m7_41 =10'b0;

   // m7_42 = W*in
   wire signed [9:0] m7_42;
   assign m7_42 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_43 = W*in
   wire signed [9:0] m7_43;
   assign m7_43 =10'b0;

   // m7_44 = W*in
   wire signed [9:0] m7_44;
   assign m7_44 =10'b0;

   // m7_45 = W*in
   wire signed [9:0] m7_45;
   assign m7_45 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_46 = W*in
   wire signed [9:0] m7_46;
   assign m7_46 =10'b0;

   // m7_47 = W*in
   wire signed [9:0] m7_47;
   assign m7_47 =10'b0;

   // m7_48 = W*in
   wire signed [9:0] m7_48;
   assign m7_48 =10'b0;

   // m7_49 = W*in
   wire signed [9:0] m7_49;
   assign m7_49 =10'b0;

   // m7_50 = W*in
   wire signed [9:0] m7_50;
   assign m7_50 =10'b0;

   // m7_51 = W*in
   wire signed [9:0] m7_51;
   assign m7_51 =10'b0;

   // m7_52 = W*in
   wire signed [9:0] m7_52;
   assign m7_52 ={ {4{in7[5]}} , in7[5:0] };

   // m7_53 = W*in
   wire signed [9:0] m7_53;
   assign m7_53 ={ {4{in7[5]}} , in7[5:0] };

   // m7_54 = W*in
   wire signed [9:0] m7_54;
   assign m7_54 =10'b0;

   // m7_55 = W*in
   wire signed [9:0] m7_55;
   assign m7_55 ={ {5{neg7[5]}} , neg7[5:1] };

   // m7_56 = W*in
   wire signed [9:0] m7_56;
   assign m7_56 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_57 = W*in
   wire signed [9:0] m7_57;
   assign m7_57 =10'b0;

   // m7_58 = W*in
   wire signed [9:0] m7_58;
   assign m7_58 =10'b0;

   // m7_59 = W*in
   wire signed [9:0] m7_59;
   assign m7_59 =10'b0;

   // m7_60 = W*in
   wire signed [9:0] m7_60;
   assign m7_60 ={ {4{in7[5]}} , in7[5:0] };

   // m7_61 = W*in
   wire signed [9:0] m7_61;
   assign m7_61 =10'b0;

   // m7_62 = W*in
   wire signed [9:0] m7_62;
   assign m7_62 =10'b0;

   // m7_63 = W*in
   wire signed [9:0] m7_63;
   assign m7_63 =10'b0;

   // m7_64 = W*in
   wire signed [9:0] m7_64;
   assign m7_64 =10'b0;

   // m7_65 = W*in
   wire signed [9:0] m7_65;
   assign m7_65 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_66 = W*in
   wire signed [9:0] m7_66;
   assign m7_66 =10'b0;

   // m7_67 = W*in
   wire signed [9:0] m7_67;
   assign m7_67 =10'b0;

   // m7_68 = W*in
   wire signed [9:0] m7_68;
   assign m7_68 =10'b0;

   // m7_69 = W*in
   wire signed [9:0] m7_69;
   assign m7_69 =10'b0;

   // m7_70 = W*in
   wire signed [9:0] m7_70;
   assign m7_70 =10'b0;

   // m7_71 = W*in
   wire signed [9:0] m7_71;
   assign m7_71 ={ {4{in7[5]}} , in7[5:0] };

   // m7_72 = W*in
   wire signed [9:0] m7_72;
   assign m7_72 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_73 = W*in
   wire signed [9:0] m7_73;
   assign m7_73 ={ {4{in7[5]}} , in7[5:0] };

   // m7_74 = W*in
   wire signed [9:0] m7_74;
   assign m7_74 =10'b0;

   // m7_75 = W*in
   wire signed [9:0] m7_75;
   assign m7_75 =10'b0;

   // m7_76 = W*in
   wire signed [9:0] m7_76;
   assign m7_76 =10'b0;

   // m7_77 = W*in
   wire signed [9:0] m7_77;
   assign m7_77 =10'b0;

   // m7_78 = W*in
   wire signed [9:0] m7_78;
   assign m7_78 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_79 = W*in
   wire signed [9:0] m7_79;
   assign m7_79 =10'b0;

   // m7_80 = W*in
   wire signed [9:0] m7_80;
   assign m7_80 ={ {4{in7[5]}} , in7[5:0] };

   // m7_81 = W*in
   wire signed [9:0] m7_81;
   assign m7_81 =10'b0;

   // m7_82 = W*in
   wire signed [9:0] m7_82;
   assign m7_82 =10'b0;

   // m7_83 = W*in
   wire signed [9:0] m7_83;
   assign m7_83 =10'b0;

   // m7_84 = W*in
   wire signed [9:0] m7_84;
   assign m7_84 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_85 = W*in
   wire signed [9:0] m7_85;
   assign m7_85 =10'b0;

   // m7_86 = W*in
   wire signed [9:0] m7_86;
   assign m7_86 =10'b0;

   // m7_87 = W*in
   wire signed [9:0] m7_87;
   assign m7_87 =10'b0;

   // m7_88 = W*in
   wire signed [9:0] m7_88;
   assign m7_88 ={ {4{in7[5]}} , in7[5:0] };

   // m7_89 = W*in
   wire signed [9:0] m7_89;
   assign m7_89 =10'b0;

   // m7_90 = W*in
   wire signed [9:0] m7_90;
   assign m7_90 =10'b0;

   // m7_91 = W*in
   wire signed [9:0] m7_91;
   assign m7_91 =10'b0;

   // m7_92 = W*in
   wire signed [9:0] m7_92;
   assign m7_92 =10'b0;

   // m7_93 = W*in
   wire signed [9:0] m7_93;
   assign m7_93 =10'b0;

   // m7_94 = W*in
   wire signed [9:0] m7_94;
   assign m7_94 =10'b0;

   // m7_95 = W*in
   wire signed [9:0] m7_95;
   assign m7_95 =10'b0;

   // m7_96 = W*in
   wire signed [9:0] m7_96;
   assign m7_96 =10'b0;

   // m7_97 = W*in
   wire signed [9:0] m7_97;
   assign m7_97 ={ {3{in7[5]}} , in7 , {1{1'b0}} };

   // m7_98 = W*in
   wire signed [9:0] m7_98;
   assign m7_98 ={ {4{in7[5]}} , in7[5:0] };

   // m7_99 = W*in
   wire signed [9:0] m7_99;
   assign m7_99 ={ {4{in7[5]}} , in7[5:0] };

   // m7_100 = W*in
   wire signed [9:0] m7_100;
   assign m7_100 =10'b0;

   // m7_101 = W*in
   wire signed [9:0] m7_101;
   assign m7_101 =10'b0;

   // m7_102 = W*in
   wire signed [9:0] m7_102;
   assign m7_102 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_103 = W*in
   wire signed [9:0] m7_103;
   assign m7_103 =10'b0;

   // m7_104 = W*in
   wire signed [9:0] m7_104;
   assign m7_104 =10'b0;

   // m7_105 = W*in
   wire signed [9:0] m7_105;
   assign m7_105 ={ {4{in7[5]}} , in7[5:0] };

   // m7_106 = W*in
   wire signed [9:0] m7_106;
   assign m7_106 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_107 = W*in
   wire signed [9:0] m7_107;
   assign m7_107 =10'b0;

   // m7_108 = W*in
   wire signed [9:0] m7_108;
   assign m7_108 ={ {5{neg7[5]}} , neg7[5:1] };

   // m7_109 = W*in
   wire signed [9:0] m7_109;
   assign m7_109 =10'b0;

   // m7_110 = W*in
   wire signed [9:0] m7_110;
   assign m7_110 ={ {4{in7[5]}} , in7[5:0] };

   // m7_111 = W*in
   wire signed [9:0] m7_111;
   assign m7_111 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_112 = W*in
   wire signed [9:0] m7_112;
   assign m7_112 =10'b0;

   // m7_113 = W*in
   wire signed [9:0] m7_113;
   assign m7_113 =10'b0;

   // m7_114 = W*in
   wire signed [9:0] m7_114;
   assign m7_114 =10'b0;

   // m7_115 = W*in
   wire signed [9:0] m7_115;
   assign m7_115 =10'b0;

   // m7_116 = W*in
   wire signed [9:0] m7_116;
   assign m7_116 ={ {4{neg7[5]}} , neg7[5:0] };

   // m7_117 = W*in
   wire signed [9:0] m7_117;
   assign m7_117 =10'b0;

   // m8_1 = W*in
   wire signed [9:0] m8_1;
   assign m8_1 =10'b0;

   // m8_2 = W*in
   wire signed [9:0] m8_2;
   assign m8_2 =10'b0;

   // m8_3 = W*in
   wire signed [9:0] m8_3;
   assign m8_3 =10'b0;

   // m8_4 = W*in
   wire signed [9:0] m8_4;
   assign m8_4 =10'b0;

   // m8_5 = W*in
   wire signed [9:0] m8_5;
   assign m8_5 =10'b0;

   // m8_6 = W*in
   wire signed [9:0] m8_6;
   assign m8_6 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_7 = W*in
   wire signed [9:0] m8_7;
   assign m8_7 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_8 = W*in
   wire signed [9:0] m8_8;
   assign m8_8 =10'b0;

   // m8_9 = W*in
   wire signed [9:0] m8_9;
   assign m8_9 =10'b0;

   // m8_10 = W*in
   wire signed [9:0] m8_10;
   assign m8_10 =10'b0;

   // m8_11 = W*in
   wire signed [9:0] m8_11;
   assign m8_11 =10'b0;

   // m8_12 = W*in
   wire signed [9:0] m8_12;
   assign m8_12 ={ {4{in8[5]}} , in8[5:0] };

   // m8_13 = W*in
   wire signed [9:0] m8_13;
   assign m8_13 =10'b0;

   // m8_14 = W*in
   wire signed [9:0] m8_14;
   assign m8_14 =10'b0;

   // m8_15 = W*in
   wire signed [9:0] m8_15;
   assign m8_15 ={ {5{in8[5]}} , in8[5:1] };

   // m8_16 = W*in
   wire signed [9:0] m8_16;
   assign m8_16 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_17 = W*in
   wire signed [9:0] m8_17;
   assign m8_17 =10'b0;

   // m8_18 = W*in
   wire signed [9:0] m8_18;
   assign m8_18 =10'b0;

   // m8_19 = W*in
   wire signed [9:0] m8_19;
   assign m8_19 =10'b0;

   // m8_20 = W*in
   wire signed [9:0] m8_20;
   assign m8_20 =10'b0;

   // m8_21 = W*in
   wire signed [9:0] m8_21;
   assign m8_21 =10'b0;

   // m8_22 = W*in
   wire signed [9:0] m8_22;
   assign m8_22 ={ {5{neg8[5]}} , neg8[5:1] };

   // m8_23 = W*in
   wire signed [9:0] m8_23;
   assign m8_23 ={ {4{in8[5]}} , in8[5:0] };

   // m8_24 = W*in
   wire signed [9:0] m8_24;
   assign m8_24 =10'b0;

   // m8_25 = W*in
   wire signed [9:0] m8_25;
   assign m8_25 =10'b0;

   // m8_26 = W*in
   wire signed [9:0] m8_26;
   assign m8_26 =10'b0;

   // m8_27 = W*in
   wire signed [9:0] m8_27;
   assign m8_27 ={ {4{in8[5]}} , in8[5:0] };

   // m8_28 = W*in
   wire signed [9:0] m8_28;
   assign m8_28 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_29 = W*in
   wire signed [9:0] m8_29;
   assign m8_29 ={ {5{neg8[5]}} , neg8[5:1] };

   // m8_30 = W*in
   wire signed [9:0] m8_30;
   assign m8_30 =10'b0;

   // m8_31 = W*in
   wire signed [9:0] m8_31;
   assign m8_31 ={ {4{in8[5]}} , in8[5:0] };

   // m8_32 = W*in
   wire signed [9:0] m8_32;
   assign m8_32 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_33 = W*in
   wire signed [9:0] m8_33;
   assign m8_33 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_34 = W*in
   wire signed [9:0] m8_34;
   assign m8_34 =10'b0;

   // m8_35 = W*in
   wire signed [9:0] m8_35;
   assign m8_35 ={ {4{in8[5]}} , in8[5:0] };

   // m8_36 = W*in
   wire signed [9:0] m8_36;
   assign m8_36 =10'b0;

   // m8_37 = W*in
   wire signed [9:0] m8_37;
   assign m8_37 =10'b0;

   // m8_38 = W*in
   wire signed [9:0] m8_38;
   assign m8_38 =10'b0;

   // m8_39 = W*in
   wire signed [9:0] m8_39;
   assign m8_39 =10'b0;

   // m8_40 = W*in
   wire signed [9:0] m8_40;
   assign m8_40 =10'b0;

   // m8_41 = W*in
   wire signed [9:0] m8_41;
   assign m8_41 =10'b0;

   // m8_42 = W*in
   wire signed [9:0] m8_42;
   assign m8_42 =10'b0;

   // m8_43 = W*in
   wire signed [9:0] m8_43;
   assign m8_43 =10'b0;

   // m8_44 = W*in
   wire signed [9:0] m8_44;
   assign m8_44 =10'b0;

   // m8_45 = W*in
   wire signed [9:0] m8_45;
   assign m8_45 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_46 = W*in
   wire signed [9:0] m8_46;
   assign m8_46 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_47 = W*in
   wire signed [9:0] m8_47;
   assign m8_47 =10'b0;

   // m8_48 = W*in
   wire signed [9:0] m8_48;
   assign m8_48 =10'b0;

   // m8_49 = W*in
   wire signed [9:0] m8_49;
   assign m8_49 =10'b0;

   // m8_50 = W*in
   wire signed [9:0] m8_50;
   assign m8_50 =10'b0;

   // m8_51 = W*in
   wire signed [9:0] m8_51;
   assign m8_51 =10'b0;

   // m8_52 = W*in
   wire signed [9:0] m8_52;
   assign m8_52 ={ {4{in8[5]}} , in8[5:0] };

   // m8_53 = W*in
   wire signed [9:0] m8_53;
   assign m8_53 =10'b0;

   // m8_54 = W*in
   wire signed [9:0] m8_54;
   assign m8_54 =10'b0;

   // m8_55 = W*in
   wire signed [9:0] m8_55;
   assign m8_55 =10'b0;

   // m8_56 = W*in
   wire signed [9:0] m8_56;
   assign m8_56 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_57 = W*in
   wire signed [9:0] m8_57;
   assign m8_57 =10'b0;

   // m8_58 = W*in
   wire signed [9:0] m8_58;
   assign m8_58 =10'b0;

   // m8_59 = W*in
   wire signed [9:0] m8_59;
   assign m8_59 =10'b0;

   // m8_60 = W*in
   wire signed [9:0] m8_60;
   assign m8_60 =10'b0;

   // m8_61 = W*in
   wire signed [9:0] m8_61;
   assign m8_61 =10'b0;

   // m8_62 = W*in
   wire signed [9:0] m8_62;
   assign m8_62 =10'b0;

   // m8_63 = W*in
   wire signed [9:0] m8_63;
   assign m8_63 =10'b0;

   // m8_64 = W*in
   wire signed [9:0] m8_64;
   assign m8_64 =10'b0;

   // m8_65 = W*in
   wire signed [9:0] m8_65;
   assign m8_65 =10'b0;

   // m8_66 = W*in
   wire signed [9:0] m8_66;
   assign m8_66 =10'b0;

   // m8_67 = W*in
   wire signed [9:0] m8_67;
   assign m8_67 ={ {5{neg8[5]}} , neg8[5:1] };

   // m8_68 = W*in
   wire signed [9:0] m8_68;
   assign m8_68 =10'b0;

   // m8_69 = W*in
   wire signed [9:0] m8_69;
   assign m8_69 =10'b0;

   // m8_70 = W*in
   wire signed [9:0] m8_70;
   assign m8_70 =10'b0;

   // m8_71 = W*in
   wire signed [9:0] m8_71;
   assign m8_71 ={ {5{in8[5]}} , in8[5:1] };

   // m8_72 = W*in
   wire signed [9:0] m8_72;
   assign m8_72 =10'b0;

   // m8_73 = W*in
   wire signed [9:0] m8_73;
   assign m8_73 =10'b0;

   // m8_74 = W*in
   wire signed [9:0] m8_74;
   assign m8_74 =10'b0;

   // m8_75 = W*in
   wire signed [9:0] m8_75;
   assign m8_75 =10'b0;

   // m8_76 = W*in
   wire signed [9:0] m8_76;
   assign m8_76 =10'b0;

   // m8_77 = W*in
   wire signed [9:0] m8_77;
   assign m8_77 =10'b0;

   // m8_78 = W*in
   wire signed [9:0] m8_78;
   assign m8_78 =10'b0;

   // m8_79 = W*in
   wire signed [9:0] m8_79;
   assign m8_79 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_80 = W*in
   wire signed [9:0] m8_80;
   assign m8_80 =10'b0;

   // m8_81 = W*in
   wire signed [9:0] m8_81;
   assign m8_81 =10'b0;

   // m8_82 = W*in
   wire signed [9:0] m8_82;
   assign m8_82 ={ {4{in8[5]}} , in8[5:0] };

   // m8_83 = W*in
   wire signed [9:0] m8_83;
   assign m8_83 =10'b0;

   // m8_84 = W*in
   wire signed [9:0] m8_84;
   assign m8_84 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_85 = W*in
   wire signed [9:0] m8_85;
   assign m8_85 =10'b0;

   // m8_86 = W*in
   wire signed [9:0] m8_86;
   assign m8_86 =10'b0;

   // m8_87 = W*in
   wire signed [9:0] m8_87;
   assign m8_87 =10'b0;

   // m8_88 = W*in
   wire signed [9:0] m8_88;
   assign m8_88 ={ {4{in8[5]}} , in8[5:0] };

   // m8_89 = W*in
   wire signed [9:0] m8_89;
   assign m8_89 =10'b0;

   // m8_90 = W*in
   wire signed [9:0] m8_90;
   assign m8_90 =10'b0;

   // m8_91 = W*in
   wire signed [9:0] m8_91;
   assign m8_91 =10'b0;

   // m8_92 = W*in
   wire signed [9:0] m8_92;
   assign m8_92 =10'b0;

   // m8_93 = W*in
   wire signed [9:0] m8_93;
   assign m8_93 =10'b0;

   // m8_94 = W*in
   wire signed [9:0] m8_94;
   assign m8_94 =10'b0;

   // m8_95 = W*in
   wire signed [9:0] m8_95;
   assign m8_95 =10'b0;

   // m8_96 = W*in
   wire signed [9:0] m8_96;
   assign m8_96 =10'b0;

   // m8_97 = W*in
   wire signed [9:0] m8_97;
   assign m8_97 ={ {5{in8[5]}} , in8[5:1] };

   // m8_98 = W*in
   wire signed [9:0] m8_98;
   assign m8_98 ={ {4{in8[5]}} , in8[5:0] };

   // m8_99 = W*in
   wire signed [9:0] m8_99;
   assign m8_99 =10'b0;

   // m8_100 = W*in
   wire signed [9:0] m8_100;
   assign m8_100 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_101 = W*in
   wire signed [9:0] m8_101;
   assign m8_101 =10'b0;

   // m8_102 = W*in
   wire signed [9:0] m8_102;
   assign m8_102 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_103 = W*in
   wire signed [9:0] m8_103;
   assign m8_103 =10'b0;

   // m8_104 = W*in
   wire signed [9:0] m8_104;
   assign m8_104 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_105 = W*in
   wire signed [9:0] m8_105;
   assign m8_105 =10'b0;

   // m8_106 = W*in
   wire signed [9:0] m8_106;
   assign m8_106 ={ {4{neg8[5]}} , neg8[5:0] };

   // m8_107 = W*in
   wire signed [9:0] m8_107;
   assign m8_107 =10'b0;

   // m8_108 = W*in
   wire signed [9:0] m8_108;
   assign m8_108 =10'b0;

   // m8_109 = W*in
   wire signed [9:0] m8_109;
   assign m8_109 ={ {4{in8[5]}} , in8[5:0] };

   // m8_110 = W*in
   wire signed [9:0] m8_110;
   assign m8_110 =10'b0;

   // m8_111 = W*in
   wire signed [9:0] m8_111;
   assign m8_111 =10'b0;

   // m8_112 = W*in
   wire signed [9:0] m8_112;
   assign m8_112 =10'b0;

   // m8_113 = W*in
   wire signed [9:0] m8_113;
   assign m8_113 =10'b0;

   // m8_114 = W*in
   wire signed [9:0] m8_114;
   assign m8_114 =10'b0;

   // m8_115 = W*in
   wire signed [9:0] m8_115;
   assign m8_115 =10'b0;

   // m8_116 = W*in
   wire signed [9:0] m8_116;
   assign m8_116 =10'b0;

   // m8_117 = W*in
   wire signed [9:0] m8_117;
   assign m8_117 ={ {5{in8[5]}} , in8[5:1] };

   // m9_1 = W*in
   wire signed [9:0] m9_1;
   assign m9_1 =10'b0;

   // m9_2 = W*in
   wire signed [9:0] m9_2;
   assign m9_2 ={ {4{in9[5]}} , in9[5:0] };

   // m9_3 = W*in
   wire signed [9:0] m9_3;
   assign m9_3 =10'b0;

   // m9_4 = W*in
   wire signed [9:0] m9_4;
   assign m9_4 =10'b0;

   // m9_5 = W*in
   wire signed [9:0] m9_5;
   assign m9_5 =10'b0;

   // m9_6 = W*in
   wire signed [9:0] m9_6;
   assign m9_6 =10'b0;

   // m9_7 = W*in
   wire signed [9:0] m9_7;
   assign m9_7 =10'b0;

   // m9_8 = W*in
   wire signed [9:0] m9_8;
   assign m9_8 ={ {4{in9[5]}} , in9[5:0] };

   // m9_9 = W*in
   wire signed [9:0] m9_9;
   assign m9_9 =10'b0;

   // m9_10 = W*in
   wire signed [9:0] m9_10;
   assign m9_10 =10'b0;

   // m9_11 = W*in
   wire signed [9:0] m9_11;
   assign m9_11 ={ {4{in9[5]}} , in9[5:0] };

   // m9_12 = W*in
   wire signed [9:0] m9_12;
   assign m9_12 =10'b0;

   // m9_13 = W*in
   wire signed [9:0] m9_13;
   assign m9_13 =10'b0;

   // m9_14 = W*in
   wire signed [9:0] m9_14;
   assign m9_14 =10'b0;

   // m9_15 = W*in
   wire signed [9:0] m9_15;
   assign m9_15 ={ {5{in9[5]}} , in9[5:1] };

   // m9_16 = W*in
   wire signed [9:0] m9_16;
   assign m9_16 ={ {4{in9[5]}} , in9[5:0] };

   // m9_17 = W*in
   wire signed [9:0] m9_17;
   assign m9_17 =10'b0;

   // m9_18 = W*in
   wire signed [9:0] m9_18;
   assign m9_18 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_19 = W*in
   wire signed [9:0] m9_19;
   assign m9_19 =10'b0;

   // m9_20 = W*in
   wire signed [9:0] m9_20;
   assign m9_20 ={ {4{in9[5]}} , in9[5:0] };

   // m9_21 = W*in
   wire signed [9:0] m9_21;
   assign m9_21 =10'b0;

   // m9_22 = W*in
   wire signed [9:0] m9_22;
   assign m9_22 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_23 = W*in
   wire signed [9:0] m9_23;
   assign m9_23 =10'b0;

   // m9_24 = W*in
   wire signed [9:0] m9_24;
   assign m9_24 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_25 = W*in
   wire signed [9:0] m9_25;
   assign m9_25 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_26 = W*in
   wire signed [9:0] m9_26;
   assign m9_26 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_27 = W*in
   wire signed [9:0] m9_27;
   assign m9_27 =10'b0;

   // m9_28 = W*in
   wire signed [9:0] m9_28;
   assign m9_28 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_29 = W*in
   wire signed [9:0] m9_29;
   assign m9_29 =10'b0;

   // m9_30 = W*in
   wire signed [9:0] m9_30;
   assign m9_30 ={ {3{in9[5]}} , in9 , {1{1'b0}} };

   // m9_31 = W*in
   wire signed [9:0] m9_31;
   assign m9_31 ={ {4{in9[5]}} , in9[5:0] };

   // m9_32 = W*in
   wire signed [9:0] m9_32;
   assign m9_32 =10'b0;

   // m9_33 = W*in
   wire signed [9:0] m9_33;
   assign m9_33 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_34 = W*in
   wire signed [9:0] m9_34;
   assign m9_34 =10'b0;

   // m9_35 = W*in
   wire signed [9:0] m9_35;
   assign m9_35 ={ {4{in9[5]}} , in9[5:0] };

   // m9_36 = W*in
   wire signed [9:0] m9_36;
   assign m9_36 =10'b0;

   // m9_37 = W*in
   wire signed [9:0] m9_37;
   assign m9_37 =10'b0;

   // m9_38 = W*in
   wire signed [9:0] m9_38;
   assign m9_38 =10'b0;

   // m9_39 = W*in
   wire signed [9:0] m9_39;
   assign m9_39 =10'b0;

   // m9_40 = W*in
   wire signed [9:0] m9_40;
   assign m9_40 =10'b0;

   // m9_41 = W*in
   wire signed [9:0] m9_41;
   assign m9_41 ={ {4{in9[5]}} , in9[5:0] };

   // m9_42 = W*in
   wire signed [9:0] m9_42;
   assign m9_42 =10'b0;

   // m9_43 = W*in
   wire signed [9:0] m9_43;
   assign m9_43 =10'b0;

   // m9_44 = W*in
   wire signed [9:0] m9_44;
   assign m9_44 =10'b0;

   // m9_45 = W*in
   wire signed [9:0] m9_45;
   assign m9_45 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_46 = W*in
   wire signed [9:0] m9_46;
   assign m9_46 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_47 = W*in
   wire signed [9:0] m9_47;
   assign m9_47 =10'b0;

   // m9_48 = W*in
   wire signed [9:0] m9_48;
   assign m9_48 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_49 = W*in
   wire signed [9:0] m9_49;
   assign m9_49 =10'b0;

   // m9_50 = W*in
   wire signed [9:0] m9_50;
   assign m9_50 =10'b0;

   // m9_51 = W*in
   wire signed [9:0] m9_51;
   assign m9_51 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_52 = W*in
   wire signed [9:0] m9_52;
   assign m9_52 ={ {4{in9[5]}} , in9[5:0] };

   // m9_53 = W*in
   wire signed [9:0] m9_53;
   assign m9_53 ={ {4{in9[5]}} , in9[5:0] };

   // m9_54 = W*in
   wire signed [9:0] m9_54;
   assign m9_54 =10'b0;

   // m9_55 = W*in
   wire signed [9:0] m9_55;
   assign m9_55 =10'b0;

   // m9_56 = W*in
   wire signed [9:0] m9_56;
   assign m9_56 =10'b0;

   // m9_57 = W*in
   wire signed [9:0] m9_57;
   assign m9_57 =10'b0;

   // m9_58 = W*in
   wire signed [9:0] m9_58;
   assign m9_58 =10'b0;

   // m9_59 = W*in
   wire signed [9:0] m9_59;
   assign m9_59 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_60 = W*in
   wire signed [9:0] m9_60;
   assign m9_60 =10'b0;

   // m9_61 = W*in
   wire signed [9:0] m9_61;
   assign m9_61 =10'b0;

   // m9_62 = W*in
   wire signed [9:0] m9_62;
   assign m9_62 =10'b0;

   // m9_63 = W*in
   wire signed [9:0] m9_63;
   assign m9_63 =10'b0;

   // m9_64 = W*in
   wire signed [9:0] m9_64;
   assign m9_64 =10'b0;

   // m9_65 = W*in
   wire signed [9:0] m9_65;
   assign m9_65 =10'b0;

   // m9_66 = W*in
   wire signed [9:0] m9_66;
   assign m9_66 ={ {4{in9[5]}} , in9[5:0] };

   // m9_67 = W*in
   wire signed [9:0] m9_67;
   assign m9_67 =10'b0;

   // m9_68 = W*in
   wire signed [9:0] m9_68;
   assign m9_68 =10'b0;

   // m9_69 = W*in
   wire signed [9:0] m9_69;
   assign m9_69 =10'b0;

   // m9_70 = W*in
   wire signed [9:0] m9_70;
   assign m9_70 =10'b0;

   // m9_71 = W*in
   wire signed [9:0] m9_71;
   assign m9_71 =10'b0;

   // m9_72 = W*in
   wire signed [9:0] m9_72;
   assign m9_72 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_73 = W*in
   wire signed [9:0] m9_73;
   assign m9_73 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_74 = W*in
   wire signed [9:0] m9_74;
   assign m9_74 =10'b0;

   // m9_75 = W*in
   wire signed [9:0] m9_75;
   assign m9_75 =10'b0;

   // m9_76 = W*in
   wire signed [9:0] m9_76;
   assign m9_76 =10'b0;

   // m9_77 = W*in
   wire signed [9:0] m9_77;
   assign m9_77 =10'b0;

   // m9_78 = W*in
   wire signed [9:0] m9_78;
   assign m9_78 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_79 = W*in
   wire signed [9:0] m9_79;
   assign m9_79 ={ {4{in9[5]}} , in9[5:0] };

   // m9_80 = W*in
   wire signed [9:0] m9_80;
   assign m9_80 =10'b0;

   // m9_81 = W*in
   wire signed [9:0] m9_81;
   assign m9_81 =10'b0;

   // m9_82 = W*in
   wire signed [9:0] m9_82;
   assign m9_82 =10'b0;

   // m9_83 = W*in
   wire signed [9:0] m9_83;
   assign m9_83 =10'b0;

   // m9_84 = W*in
   wire signed [9:0] m9_84;
   assign m9_84 =10'b0;

   // m9_85 = W*in
   wire signed [9:0] m9_85;
   assign m9_85 =10'b0;

   // m9_86 = W*in
   wire signed [9:0] m9_86;
   assign m9_86 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_87 = W*in
   wire signed [9:0] m9_87;
   assign m9_87 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_88 = W*in
   wire signed [9:0] m9_88;
   assign m9_88 ={ {4{in9[5]}} , in9[5:0] };

   // m9_89 = W*in
   wire signed [9:0] m9_89;
   assign m9_89 =10'b0;

   // m9_90 = W*in
   wire signed [9:0] m9_90;
   assign m9_90 =10'b0;

   // m9_91 = W*in
   wire signed [9:0] m9_91;
   assign m9_91 =10'b0;

   // m9_92 = W*in
   wire signed [9:0] m9_92;
   assign m9_92 =10'b0;

   // m9_93 = W*in
   wire signed [9:0] m9_93;
   assign m9_93 =10'b0;

   // m9_94 = W*in
   wire signed [9:0] m9_94;
   assign m9_94 ={ {4{in9[5]}} , in9[5:0] };

   // m9_95 = W*in
   wire signed [9:0] m9_95;
   assign m9_95 =10'b0;

   // m9_96 = W*in
   wire signed [9:0] m9_96;
   assign m9_96 =10'b0;

   // m9_97 = W*in
   wire signed [9:0] m9_97;
   assign m9_97 =10'b0;

   // m9_98 = W*in
   wire signed [9:0] m9_98;
   assign m9_98 ={ {4{in9[5]}} , in9[5:0] };

   // m9_99 = W*in
   wire signed [9:0] m9_99;
   assign m9_99 =10'b0;

   // m9_100 = W*in
   wire signed [9:0] m9_100;
   assign m9_100 =10'b0;

   // m9_101 = W*in
   wire signed [9:0] m9_101;
   assign m9_101 =10'b0;

   // m9_102 = W*in
   wire signed [9:0] m9_102;
   assign m9_102 =10'b0;

   // m9_103 = W*in
   wire signed [9:0] m9_103;
   assign m9_103 =10'b0;

   // m9_104 = W*in
   wire signed [9:0] m9_104;
   assign m9_104 =10'b0;

   // m9_105 = W*in
   wire signed [9:0] m9_105;
   assign m9_105 ={ {4{in9[5]}} , in9[5:0] };

   // m9_106 = W*in
   wire signed [9:0] m9_106;
   assign m9_106 ={ {4{in9[5]}} , in9[5:0] };

   // m9_107 = W*in
   wire signed [9:0] m9_107;
   assign m9_107 ={ {5{neg9[5]}} , neg9[5:1] };

   // m9_108 = W*in
   wire signed [9:0] m9_108;
   assign m9_108 ={ {4{in9[5]}} , in9[5:0] };

   // m9_109 = W*in
   wire signed [9:0] m9_109;
   assign m9_109 ={ {4{in9[5]}} , in9[5:0] };

   // m9_110 = W*in
   wire signed [9:0] m9_110;
   assign m9_110 =10'b0;

   // m9_111 = W*in
   wire signed [9:0] m9_111;
   assign m9_111 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_112 = W*in
   wire signed [9:0] m9_112;
   assign m9_112 =10'b0;

   // m9_113 = W*in
   wire signed [9:0] m9_113;
   assign m9_113 =10'b0;

   // m9_114 = W*in
   wire signed [9:0] m9_114;
   assign m9_114 ={ {4{neg9[5]}} , neg9[5:0] };

   // m9_115 = W*in
   wire signed [9:0] m9_115;
   assign m9_115 ={ {4{in9[5]}} , in9[5:0] };

   // m9_116 = W*in
   wire signed [9:0] m9_116;
   assign m9_116 ={ {4{in9[5]}} , in9[5:0] };

   // m9_117 = W*in
   wire signed [9:0] m9_117;
   assign m9_117 ={ {4{in9[5]}} , in9[5:0] };

   // m10_1 = W*in
   wire signed [9:0] m10_1;
   assign m10_1 =10'b0;

   // m10_2 = W*in
   wire signed [9:0] m10_2;
   assign m10_2 =10'b0;

   // m10_3 = W*in
   wire signed [9:0] m10_3;
   assign m10_3 =10'b0;

   // m10_4 = W*in
   wire signed [9:0] m10_4;
   assign m10_4 =10'b0;

   // m10_5 = W*in
   wire signed [9:0] m10_5;
   assign m10_5 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_6 = W*in
   wire signed [9:0] m10_6;
   assign m10_6 =10'b0;

   // m10_7 = W*in
   wire signed [9:0] m10_7;
   assign m10_7 =10'b0;

   // m10_8 = W*in
   wire signed [9:0] m10_8;
   assign m10_8 =10'b0;

   // m10_9 = W*in
   wire signed [9:0] m10_9;
   assign m10_9 =10'b0;

   // m10_10 = W*in
   wire signed [9:0] m10_10;
   assign m10_10 =10'b0;

   // m10_11 = W*in
   wire signed [9:0] m10_11;
   assign m10_11 =10'b0;

   // m10_12 = W*in
   wire signed [9:0] m10_12;
   assign m10_12 =10'b0;

   // m10_13 = W*in
   wire signed [9:0] m10_13;
   assign m10_13 ={ {4{in10[5]}} , in10[5:0] };

   // m10_14 = W*in
   wire signed [9:0] m10_14;
   assign m10_14 =10'b0;

   // m10_15 = W*in
   wire signed [9:0] m10_15;
   assign m10_15 =10'b0;

   // m10_16 = W*in
   wire signed [9:0] m10_16;
   assign m10_16 ={ {4{in10[5]}} , in10[5:0] };

   // m10_17 = W*in
   wire signed [9:0] m10_17;
   assign m10_17 =10'b0;

   // m10_18 = W*in
   wire signed [9:0] m10_18;
   assign m10_18 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_19 = W*in
   wire signed [9:0] m10_19;
   assign m10_19 =10'b0;

   // m10_20 = W*in
   wire signed [9:0] m10_20;
   assign m10_20 =10'b0;

   // m10_21 = W*in
   wire signed [9:0] m10_21;
   assign m10_21 =10'b0;

   // m10_22 = W*in
   wire signed [9:0] m10_22;
   assign m10_22 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_23 = W*in
   wire signed [9:0] m10_23;
   assign m10_23 =10'b0;

   // m10_24 = W*in
   wire signed [9:0] m10_24;
   assign m10_24 =10'b0;

   // m10_25 = W*in
   wire signed [9:0] m10_25;
   assign m10_25 =10'b0;

   // m10_26 = W*in
   wire signed [9:0] m10_26;
   assign m10_26 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_27 = W*in
   wire signed [9:0] m10_27;
   assign m10_27 =10'b0;

   // m10_28 = W*in
   wire signed [9:0] m10_28;
   assign m10_28 =10'b0;

   // m10_29 = W*in
   wire signed [9:0] m10_29;
   assign m10_29 =10'b0;

   // m10_30 = W*in
   wire signed [9:0] m10_30;
   assign m10_30 ={ {4{in10[5]}} , in10[5:0] };

   // m10_31 = W*in
   wire signed [9:0] m10_31;
   assign m10_31 =10'b0;

   // m10_32 = W*in
   wire signed [9:0] m10_32;
   assign m10_32 =10'b0;

   // m10_33 = W*in
   wire signed [9:0] m10_33;
   assign m10_33 =10'b0;

   // m10_34 = W*in
   wire signed [9:0] m10_34;
   assign m10_34 =10'b0;

   // m10_35 = W*in
   wire signed [9:0] m10_35;
   assign m10_35 ={ {4{in10[5]}} , in10[5:0] };

   // m10_36 = W*in
   wire signed [9:0] m10_36;
   assign m10_36 =10'b0;

   // m10_37 = W*in
   wire signed [9:0] m10_37;
   assign m10_37 =10'b0;

   // m10_38 = W*in
   wire signed [9:0] m10_38;
   assign m10_38 =10'b0;

   // m10_39 = W*in
   wire signed [9:0] m10_39;
   assign m10_39 =10'b0;

   // m10_40 = W*in
   wire signed [9:0] m10_40;
   assign m10_40 =10'b0;

   // m10_41 = W*in
   wire signed [9:0] m10_41;
   assign m10_41 ={ {4{in10[5]}} , in10[5:0] };

   // m10_42 = W*in
   wire signed [9:0] m10_42;
   assign m10_42 ={ {5{in10[5]}} , in10[5:1] };

   // m10_43 = W*in
   wire signed [9:0] m10_43;
   assign m10_43 =10'b0;

   // m10_44 = W*in
   wire signed [9:0] m10_44;
   assign m10_44 =10'b0;

   // m10_45 = W*in
   wire signed [9:0] m10_45;
   assign m10_45 =10'b0;

   // m10_46 = W*in
   wire signed [9:0] m10_46;
   assign m10_46 =10'b0;

   // m10_47 = W*in
   wire signed [9:0] m10_47;
   assign m10_47 =10'b0;

   // m10_48 = W*in
   wire signed [9:0] m10_48;
   assign m10_48 =10'b0;

   // m10_49 = W*in
   wire signed [9:0] m10_49;
   assign m10_49 =10'b0;

   // m10_50 = W*in
   wire signed [9:0] m10_50;
   assign m10_50 =10'b0;

   // m10_51 = W*in
   wire signed [9:0] m10_51;
   assign m10_51 =10'b0;

   // m10_52 = W*in
   wire signed [9:0] m10_52;
   assign m10_52 ={ {4{in10[5]}} , in10[5:0] };

   // m10_53 = W*in
   wire signed [9:0] m10_53;
   assign m10_53 =10'b0;

   // m10_54 = W*in
   wire signed [9:0] m10_54;
   assign m10_54 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_55 = W*in
   wire signed [9:0] m10_55;
   assign m10_55 =10'b0;

   // m10_56 = W*in
   wire signed [9:0] m10_56;
   assign m10_56 ={ {4{in10[5]}} , in10[5:0] };

   // m10_57 = W*in
   wire signed [9:0] m10_57;
   assign m10_57 =10'b0;

   // m10_58 = W*in
   wire signed [9:0] m10_58;
   assign m10_58 =10'b0;

   // m10_59 = W*in
   wire signed [9:0] m10_59;
   assign m10_59 =10'b0;

   // m10_60 = W*in
   wire signed [9:0] m10_60;
   assign m10_60 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_61 = W*in
   wire signed [9:0] m10_61;
   assign m10_61 =10'b0;

   // m10_62 = W*in
   wire signed [9:0] m10_62;
   assign m10_62 =10'b0;

   // m10_63 = W*in
   wire signed [9:0] m10_63;
   assign m10_63 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_64 = W*in
   wire signed [9:0] m10_64;
   assign m10_64 =10'b0;

   // m10_65 = W*in
   wire signed [9:0] m10_65;
   assign m10_65 =10'b0;

   // m10_66 = W*in
   wire signed [9:0] m10_66;
   assign m10_66 ={ {5{in10[5]}} , in10[5:1] };

   // m10_67 = W*in
   wire signed [9:0] m10_67;
   assign m10_67 =10'b0;

   // m10_68 = W*in
   wire signed [9:0] m10_68;
   assign m10_68 =10'b0;

   // m10_69 = W*in
   wire signed [9:0] m10_69;
   assign m10_69 =10'b0;

   // m10_70 = W*in
   wire signed [9:0] m10_70;
   assign m10_70 =10'b0;

   // m10_71 = W*in
   wire signed [9:0] m10_71;
   assign m10_71 ={ {5{neg10[5]}} , neg10[5:1] };

   // m10_72 = W*in
   wire signed [9:0] m10_72;
   assign m10_72 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_73 = W*in
   wire signed [9:0] m10_73;
   assign m10_73 =10'b0;

   // m10_74 = W*in
   wire signed [9:0] m10_74;
   assign m10_74 =10'b0;

   // m10_75 = W*in
   wire signed [9:0] m10_75;
   assign m10_75 ={ {5{neg10[5]}} , neg10[5:1] };

   // m10_76 = W*in
   wire signed [9:0] m10_76;
   assign m10_76 =10'b0;

   // m10_77 = W*in
   wire signed [9:0] m10_77;
   assign m10_77 =10'b0;

   // m10_78 = W*in
   wire signed [9:0] m10_78;
   assign m10_78 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_79 = W*in
   wire signed [9:0] m10_79;
   assign m10_79 ={ {4{in10[5]}} , in10[5:0] };

   // m10_80 = W*in
   wire signed [9:0] m10_80;
   assign m10_80 ={ {4{in10[5]}} , in10[5:0] };

   // m10_81 = W*in
   wire signed [9:0] m10_81;
   assign m10_81 =10'b0;

   // m10_82 = W*in
   wire signed [9:0] m10_82;
   assign m10_82 =10'b0;

   // m10_83 = W*in
   wire signed [9:0] m10_83;
   assign m10_83 =10'b0;

   // m10_84 = W*in
   wire signed [9:0] m10_84;
   assign m10_84 =10'b0;

   // m10_85 = W*in
   wire signed [9:0] m10_85;
   assign m10_85 =10'b0;

   // m10_86 = W*in
   wire signed [9:0] m10_86;
   assign m10_86 =10'b0;

   // m10_87 = W*in
   wire signed [9:0] m10_87;
   assign m10_87 ={ {4{neg10[5]}} , neg10[5:0] };

   // m10_88 = W*in
   wire signed [9:0] m10_88;
   assign m10_88 =10'b0;

   // m10_89 = W*in
   wire signed [9:0] m10_89;
   assign m10_89 =10'b0;

   // m10_90 = W*in
   wire signed [9:0] m10_90;
   assign m10_90 =10'b0;

   // m10_91 = W*in
   wire signed [9:0] m10_91;
   assign m10_91 =10'b0;

   // m10_92 = W*in
   wire signed [9:0] m10_92;
   assign m10_92 =10'b0;

   // m10_93 = W*in
   wire signed [9:0] m10_93;
   assign m10_93 =10'b0;

   // m10_94 = W*in
   wire signed [9:0] m10_94;
   assign m10_94 ={ {4{in10[5]}} , in10[5:0] };

   // m10_95 = W*in
   wire signed [9:0] m10_95;
   assign m10_95 =10'b0;

   // m10_96 = W*in
   wire signed [9:0] m10_96;
   assign m10_96 ={ {5{in10[5]}} , in10[5:1] };

   // m10_97 = W*in
   wire signed [9:0] m10_97;
   assign m10_97 ={ {4{in10[5]}} , in10[5:0] };

   // m10_98 = W*in
   wire signed [9:0] m10_98;
   assign m10_98 =10'b0;

   // m10_99 = W*in
   wire signed [9:0] m10_99;
   assign m10_99 =10'b0;

   // m10_100 = W*in
   wire signed [9:0] m10_100;
   assign m10_100 ={ {5{in10[5]}} , in10[5:1] };

   // m10_101 = W*in
   wire signed [9:0] m10_101;
   assign m10_101 =10'b0;

   // m10_102 = W*in
   wire signed [9:0] m10_102;
   assign m10_102 =10'b0;

   // m10_103 = W*in
   wire signed [9:0] m10_103;
   assign m10_103 =10'b0;

   // m10_104 = W*in
   wire signed [9:0] m10_104;
   assign m10_104 =10'b0;

   // m10_105 = W*in
   wire signed [9:0] m10_105;
   assign m10_105 =10'b0;

   // m10_106 = W*in
   wire signed [9:0] m10_106;
   assign m10_106 =10'b0;

   // m10_107 = W*in
   wire signed [9:0] m10_107;
   assign m10_107 =10'b0;

   // m10_108 = W*in
   wire signed [9:0] m10_108;
   assign m10_108 ={ {4{in10[5]}} , in10[5:0] };

   // m10_109 = W*in
   wire signed [9:0] m10_109;
   assign m10_109 ={ {4{in10[5]}} , in10[5:0] };

   // m10_110 = W*in
   wire signed [9:0] m10_110;
   assign m10_110 =10'b0;

   // m10_111 = W*in
   wire signed [9:0] m10_111;
   assign m10_111 =10'b0;

   // m10_112 = W*in
   wire signed [9:0] m10_112;
   assign m10_112 =10'b0;

   // m10_113 = W*in
   wire signed [9:0] m10_113;
   assign m10_113 =10'b0;

   // m10_114 = W*in
   wire signed [9:0] m10_114;
   assign m10_114 =10'b0;

   // m10_115 = W*in
   wire signed [9:0] m10_115;
   assign m10_115 =10'b0;

   // m10_116 = W*in
   wire signed [9:0] m10_116;
   assign m10_116 ={ {3{in10[5]}} , in10 , {1{1'b0}} };

   // m10_117 = W*in
   wire signed [9:0] m10_117;
   assign m10_117 =10'b0;

   // m11_1 = W*in
   wire signed [9:0] m11_1;
   assign m11_1 =10'b0;

   // m11_2 = W*in
   wire signed [9:0] m11_2;
   assign m11_2 =10'b0;

   // m11_3 = W*in
   wire signed [9:0] m11_3;
   assign m11_3 =10'b0;

   // m11_4 = W*in
   wire signed [9:0] m11_4;
   assign m11_4 =10'b0;

   // m11_5 = W*in
   wire signed [9:0] m11_5;
   assign m11_5 =10'b0;

   // m11_6 = W*in
   wire signed [9:0] m11_6;
   assign m11_6 =10'b0;

   // m11_7 = W*in
   wire signed [9:0] m11_7;
   assign m11_7 =10'b0;

   // m11_8 = W*in
   wire signed [9:0] m11_8;
   assign m11_8 =10'b0;

   // m11_9 = W*in
   wire signed [9:0] m11_9;
   assign m11_9 =10'b0;

   // m11_10 = W*in
   wire signed [9:0] m11_10;
   assign m11_10 =10'b0;

   // m11_11 = W*in
   wire signed [9:0] m11_11;
   assign m11_11 =10'b0;

   // m11_12 = W*in
   wire signed [9:0] m11_12;
   assign m11_12 ={ {4{in11[5]}} , in11[5:0] };

   // m11_13 = W*in
   wire signed [9:0] m11_13;
   assign m11_13 =10'b0;

   // m11_14 = W*in
   wire signed [9:0] m11_14;
   assign m11_14 =10'b0;

   // m11_15 = W*in
   wire signed [9:0] m11_15;
   assign m11_15 =10'b0;

   // m11_16 = W*in
   wire signed [9:0] m11_16;
   assign m11_16 =10'b0;

   // m11_17 = W*in
   wire signed [9:0] m11_17;
   assign m11_17 ={ {4{in11[5]}} , in11[5:0] };

   // m11_18 = W*in
   wire signed [9:0] m11_18;
   assign m11_18 =10'b0;

   // m11_19 = W*in
   wire signed [9:0] m11_19;
   assign m11_19 ={ {5{in11[5]}} , in11[5:1] };

   // m11_20 = W*in
   wire signed [9:0] m11_20;
   assign m11_20 ={ {4{neg11[5]}} , neg11[5:0] };

   // m11_21 = W*in
   wire signed [9:0] m11_21;
   assign m11_21 =10'b0;

   // m11_22 = W*in
   wire signed [9:0] m11_22;
   assign m11_22 ={ {5{neg11[5]}} , neg11[5:1] };

   // m11_23 = W*in
   wire signed [9:0] m11_23;
   assign m11_23 =10'b0;

   // m11_24 = W*in
   wire signed [9:0] m11_24;
   assign m11_24 =10'b0;

   // m11_25 = W*in
   wire signed [9:0] m11_25;
   assign m11_25 ={ {4{in11[5]}} , in11[5:0] };

   // m11_26 = W*in
   wire signed [9:0] m11_26;
   assign m11_26 ={ {5{neg11[5]}} , neg11[5:1] };

   // m11_27 = W*in
   wire signed [9:0] m11_27;
   assign m11_27 =10'b0;

   // m11_28 = W*in
   wire signed [9:0] m11_28;
   assign m11_28 =10'b0;

   // m11_29 = W*in
   wire signed [9:0] m11_29;
   assign m11_29 ={ {5{in11[5]}} , in11[5:1] };

   // m11_30 = W*in
   wire signed [9:0] m11_30;
   assign m11_30 =10'b0;

   // m11_31 = W*in
   wire signed [9:0] m11_31;
   assign m11_31 =10'b0;

   // m11_32 = W*in
   wire signed [9:0] m11_32;
   assign m11_32 =10'b0;

   // m11_33 = W*in
   wire signed [9:0] m11_33;
   assign m11_33 =10'b0;

   // m11_34 = W*in
   wire signed [9:0] m11_34;
   assign m11_34 =10'b0;

   // m11_35 = W*in
   wire signed [9:0] m11_35;
   assign m11_35 ={ {5{neg11[5]}} , neg11[5:1] };

   // m11_36 = W*in
   wire signed [9:0] m11_36;
   assign m11_36 ={ {5{in11[5]}} , in11[5:1] };

   // m11_37 = W*in
   wire signed [9:0] m11_37;
   assign m11_37 =10'b0;

   // m11_38 = W*in
   wire signed [9:0] m11_38;
   assign m11_38 =10'b0;

   // m11_39 = W*in
   wire signed [9:0] m11_39;
   assign m11_39 =10'b0;

   // m11_40 = W*in
   wire signed [9:0] m11_40;
   assign m11_40 =10'b0;

   // m11_41 = W*in
   wire signed [9:0] m11_41;
   assign m11_41 =10'b0;

   // m11_42 = W*in
   wire signed [9:0] m11_42;
   assign m11_42 =10'b0;

   // m11_43 = W*in
   wire signed [9:0] m11_43;
   assign m11_43 =10'b0;

   // m11_44 = W*in
   wire signed [9:0] m11_44;
   assign m11_44 ={ {4{in11[5]}} , in11[5:0] };

   // m11_45 = W*in
   wire signed [9:0] m11_45;
   assign m11_45 =10'b0;

   // m11_46 = W*in
   wire signed [9:0] m11_46;
   assign m11_46 =10'b0;

   // m11_47 = W*in
   wire signed [9:0] m11_47;
   assign m11_47 =10'b0;

   // m11_48 = W*in
   wire signed [9:0] m11_48;
   assign m11_48 =10'b0;

   // m11_49 = W*in
   wire signed [9:0] m11_49;
   assign m11_49 ={ {4{in11[5]}} , in11[5:0] };

   // m11_50 = W*in
   wire signed [9:0] m11_50;
   assign m11_50 =10'b0;

   // m11_51 = W*in
   wire signed [9:0] m11_51;
   assign m11_51 =10'b0;

   // m11_52 = W*in
   wire signed [9:0] m11_52;
   assign m11_52 =10'b0;

   // m11_53 = W*in
   wire signed [9:0] m11_53;
   assign m11_53 =10'b0;

   // m11_54 = W*in
   wire signed [9:0] m11_54;
   assign m11_54 ={ {4{in11[5]}} , in11[5:0] };

   // m11_55 = W*in
   wire signed [9:0] m11_55;
   assign m11_55 =10'b0;

   // m11_56 = W*in
   wire signed [9:0] m11_56;
   assign m11_56 =10'b0;

   // m11_57 = W*in
   wire signed [9:0] m11_57;
   assign m11_57 =10'b0;

   // m11_58 = W*in
   wire signed [9:0] m11_58;
   assign m11_58 =10'b0;

   // m11_59 = W*in
   wire signed [9:0] m11_59;
   assign m11_59 =10'b0;

   // m11_60 = W*in
   wire signed [9:0] m11_60;
   assign m11_60 =10'b0;

   // m11_61 = W*in
   wire signed [9:0] m11_61;
   assign m11_61 =10'b0;

   // m11_62 = W*in
   wire signed [9:0] m11_62;
   assign m11_62 =10'b0;

   // m11_63 = W*in
   wire signed [9:0] m11_63;
   assign m11_63 =10'b0;

   // m11_64 = W*in
   wire signed [9:0] m11_64;
   assign m11_64 ={ {4{neg11[5]}} , neg11[5:0] };

   // m11_65 = W*in
   wire signed [9:0] m11_65;
   assign m11_65 =10'b0;

   // m11_66 = W*in
   wire signed [9:0] m11_66;
   assign m11_66 ={ {4{in11[5]}} , in11[5:0] };

   // m11_67 = W*in
   wire signed [9:0] m11_67;
   assign m11_67 =10'b0;

   // m11_68 = W*in
   wire signed [9:0] m11_68;
   assign m11_68 =10'b0;

   // m11_69 = W*in
   wire signed [9:0] m11_69;
   assign m11_69 =10'b0;

   // m11_70 = W*in
   wire signed [9:0] m11_70;
   assign m11_70 =10'b0;

   // m11_71 = W*in
   wire signed [9:0] m11_71;
   assign m11_71 =10'b0;

   // m11_72 = W*in
   wire signed [9:0] m11_72;
   assign m11_72 ={ {5{neg11[5]}} , neg11[5:1] };

   // m11_73 = W*in
   wire signed [9:0] m11_73;
   assign m11_73 =10'b0;

   // m11_74 = W*in
   wire signed [9:0] m11_74;
   assign m11_74 ={ {5{neg11[5]}} , neg11[5:1] };

   // m11_75 = W*in
   wire signed [9:0] m11_75;
   assign m11_75 =10'b0;

   // m11_76 = W*in
   wire signed [9:0] m11_76;
   assign m11_76 =10'b0;

   // m11_77 = W*in
   wire signed [9:0] m11_77;
   assign m11_77 =10'b0;

   // m11_78 = W*in
   wire signed [9:0] m11_78;
   assign m11_78 =10'b0;

   // m11_79 = W*in
   wire signed [9:0] m11_79;
   assign m11_79 =10'b0;

   // m11_80 = W*in
   wire signed [9:0] m11_80;
   assign m11_80 =10'b0;

   // m11_81 = W*in
   wire signed [9:0] m11_81;
   assign m11_81 ={ {5{neg11[5]}} , neg11[5:1] };

   // m11_82 = W*in
   wire signed [9:0] m11_82;
   assign m11_82 ={ {4{neg11[5]}} , neg11[5:0] };

   // m11_83 = W*in
   wire signed [9:0] m11_83;
   assign m11_83 =10'b0;

   // m11_84 = W*in
   wire signed [9:0] m11_84;
   assign m11_84 =10'b0;

   // m11_85 = W*in
   wire signed [9:0] m11_85;
   assign m11_85 ={ {4{in11[5]}} , in11[5:0] };

   // m11_86 = W*in
   wire signed [9:0] m11_86;
   assign m11_86 =10'b0;

   // m11_87 = W*in
   wire signed [9:0] m11_87;
   assign m11_87 =10'b0;

   // m11_88 = W*in
   wire signed [9:0] m11_88;
   assign m11_88 =10'b0;

   // m11_89 = W*in
   wire signed [9:0] m11_89;
   assign m11_89 =10'b0;

   // m11_90 = W*in
   wire signed [9:0] m11_90;
   assign m11_90 =10'b0;

   // m11_91 = W*in
   wire signed [9:0] m11_91;
   assign m11_91 =10'b0;

   // m11_92 = W*in
   wire signed [9:0] m11_92;
   assign m11_92 =10'b0;

   // m11_93 = W*in
   wire signed [9:0] m11_93;
   assign m11_93 =10'b0;

   // m11_94 = W*in
   wire signed [9:0] m11_94;
   assign m11_94 =10'b0;

   // m11_95 = W*in
   wire signed [9:0] m11_95;
   assign m11_95 ={ {4{in11[5]}} , in11[5:0] };

   // m11_96 = W*in
   wire signed [9:0] m11_96;
   assign m11_96 =10'b0;

   // m11_97 = W*in
   wire signed [9:0] m11_97;
   assign m11_97 ={ {4{in11[5]}} , in11[5:0] };

   // m11_98 = W*in
   wire signed [9:0] m11_98;
   assign m11_98 =10'b0;

   // m11_99 = W*in
   wire signed [9:0] m11_99;
   assign m11_99 =10'b0;

   // m11_100 = W*in
   wire signed [9:0] m11_100;
   assign m11_100 =10'b0;

   // m11_101 = W*in
   wire signed [9:0] m11_101;
   assign m11_101 =10'b0;

   // m11_102 = W*in
   wire signed [9:0] m11_102;
   assign m11_102 =10'b0;

   // m11_103 = W*in
   wire signed [9:0] m11_103;
   assign m11_103 =10'b0;

   // m11_104 = W*in
   wire signed [9:0] m11_104;
   assign m11_104 =10'b0;

   // m11_105 = W*in
   wire signed [9:0] m11_105;
   assign m11_105 =10'b0;

   // m11_106 = W*in
   wire signed [9:0] m11_106;
   assign m11_106 =10'b0;

   // m11_107 = W*in
   wire signed [9:0] m11_107;
   assign m11_107 ={ {5{in11[5]}} , in11[5:1] };

   // m11_108 = W*in
   wire signed [9:0] m11_108;
   assign m11_108 =10'b0;

   // m11_109 = W*in
   wire signed [9:0] m11_109;
   assign m11_109 =10'b0;

   // m11_110 = W*in
   wire signed [9:0] m11_110;
   assign m11_110 =10'b0;

   // m11_111 = W*in
   wire signed [9:0] m11_111;
   assign m11_111 =10'b0;

   // m11_112 = W*in
   wire signed [9:0] m11_112;
   assign m11_112 =10'b0;

   // m11_113 = W*in
   wire signed [9:0] m11_113;
   assign m11_113 =10'b0;

   // m11_114 = W*in
   wire signed [9:0] m11_114;
   assign m11_114 =10'b0;

   // m11_115 = W*in
   wire signed [9:0] m11_115;
   assign m11_115 ={ {4{neg11[5]}} , neg11[5:0] };

   // m11_116 = W*in
   wire signed [9:0] m11_116;
   assign m11_116 =10'b0;

   // m11_117 = W*in
   wire signed [9:0] m11_117;
   assign m11_117 =10'b0;

   // m12_1 = W*in
   wire signed [9:0] m12_1;
   assign m12_1 =10'b0;

   // m12_2 = W*in
   wire signed [9:0] m12_2;
   assign m12_2 =10'b0;

   // m12_3 = W*in
   wire signed [9:0] m12_3;
   assign m12_3 ={ {4{in12[5]}} , in12[5:0] };

   // m12_4 = W*in
   wire signed [9:0] m12_4;
   assign m12_4 =10'b0;

   // m12_5 = W*in
   wire signed [9:0] m12_5;
   assign m12_5 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_6 = W*in
   wire signed [9:0] m12_6;
   assign m12_6 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_7 = W*in
   wire signed [9:0] m12_7;
   assign m12_7 =10'b0;

   // m12_8 = W*in
   wire signed [9:0] m12_8;
   assign m12_8 =10'b0;

   // m12_9 = W*in
   wire signed [9:0] m12_9;
   assign m12_9 =10'b0;

   // m12_10 = W*in
   wire signed [9:0] m12_10;
   assign m12_10 =10'b0;

   // m12_11 = W*in
   wire signed [9:0] m12_11;
   assign m12_11 =10'b0;

   // m12_12 = W*in
   wire signed [9:0] m12_12;
   assign m12_12 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_13 = W*in
   wire signed [9:0] m12_13;
   assign m12_13 ={ {4{in12[5]}} , in12[5:0] };

   // m12_14 = W*in
   wire signed [9:0] m12_14;
   assign m12_14 =10'b0;

   // m12_15 = W*in
   wire signed [9:0] m12_15;
   assign m12_15 =10'b0;

   // m12_16 = W*in
   wire signed [9:0] m12_16;
   assign m12_16 =10'b0;

   // m12_17 = W*in
   wire signed [9:0] m12_17;
   assign m12_17 ={ {4{in12[5]}} , in12[5:0] };

   // m12_18 = W*in
   wire signed [9:0] m12_18;
   assign m12_18 ={ {5{in12[5]}} , in12[5:1] };

   // m12_19 = W*in
   wire signed [9:0] m12_19;
   assign m12_19 =10'b0;

   // m12_20 = W*in
   wire signed [9:0] m12_20;
   assign m12_20 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_21 = W*in
   wire signed [9:0] m12_21;
   assign m12_21 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_22 = W*in
   wire signed [9:0] m12_22;
   assign m12_22 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_23 = W*in
   wire signed [9:0] m12_23;
   assign m12_23 =10'b0;

   // m12_24 = W*in
   wire signed [9:0] m12_24;
   assign m12_24 =10'b0;

   // m12_25 = W*in
   wire signed [9:0] m12_25;
   assign m12_25 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_26 = W*in
   wire signed [9:0] m12_26;
   assign m12_26 =10'b0;

   // m12_27 = W*in
   wire signed [9:0] m12_27;
   assign m12_27 =10'b0;

   // m12_28 = W*in
   wire signed [9:0] m12_28;
   assign m12_28 =10'b0;

   // m12_29 = W*in
   wire signed [9:0] m12_29;
   assign m12_29 =10'b0;

   // m12_30 = W*in
   wire signed [9:0] m12_30;
   assign m12_30 =10'b0;

   // m12_31 = W*in
   wire signed [9:0] m12_31;
   assign m12_31 ={ {5{in12[5]}} , in12[5:1] };

   // m12_32 = W*in
   wire signed [9:0] m12_32;
   assign m12_32 =10'b0;

   // m12_33 = W*in
   wire signed [9:0] m12_33;
   assign m12_33 =10'b0;

   // m12_34 = W*in
   wire signed [9:0] m12_34;
   assign m12_34 =10'b0;

   // m12_35 = W*in
   wire signed [9:0] m12_35;
   assign m12_35 =10'b0;

   // m12_36 = W*in
   wire signed [9:0] m12_36;
   assign m12_36 ={ {4{in12[5]}} , in12[5:0] };

   // m12_37 = W*in
   wire signed [9:0] m12_37;
   assign m12_37 =10'b0;

   // m12_38 = W*in
   wire signed [9:0] m12_38;
   assign m12_38 =10'b0;

   // m12_39 = W*in
   wire signed [9:0] m12_39;
   assign m12_39 =10'b0;

   // m12_40 = W*in
   wire signed [9:0] m12_40;
   assign m12_40 =10'b0;

   // m12_41 = W*in
   wire signed [9:0] m12_41;
   assign m12_41 =10'b0;

   // m12_42 = W*in
   wire signed [9:0] m12_42;
   assign m12_42 =10'b0;

   // m12_43 = W*in
   wire signed [9:0] m12_43;
   assign m12_43 =10'b0;

   // m12_44 = W*in
   wire signed [9:0] m12_44;
   assign m12_44 =10'b0;

   // m12_45 = W*in
   wire signed [9:0] m12_45;
   assign m12_45 =10'b0;

   // m12_46 = W*in
   wire signed [9:0] m12_46;
   assign m12_46 =10'b0;

   // m12_47 = W*in
   wire signed [9:0] m12_47;
   assign m12_47 =10'b0;

   // m12_48 = W*in
   wire signed [9:0] m12_48;
   assign m12_48 =10'b0;

   // m12_49 = W*in
   wire signed [9:0] m12_49;
   assign m12_49 =10'b0;

   // m12_50 = W*in
   wire signed [9:0] m12_50;
   assign m12_50 =10'b0;

   // m12_51 = W*in
   wire signed [9:0] m12_51;
   assign m12_51 =10'b0;

   // m12_52 = W*in
   wire signed [9:0] m12_52;
   assign m12_52 =10'b0;

   // m12_53 = W*in
   wire signed [9:0] m12_53;
   assign m12_53 =10'b0;

   // m12_54 = W*in
   wire signed [9:0] m12_54;
   assign m12_54 =10'b0;

   // m12_55 = W*in
   wire signed [9:0] m12_55;
   assign m12_55 =10'b0;

   // m12_56 = W*in
   wire signed [9:0] m12_56;
   assign m12_56 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_57 = W*in
   wire signed [9:0] m12_57;
   assign m12_57 =10'b0;

   // m12_58 = W*in
   wire signed [9:0] m12_58;
   assign m12_58 =10'b0;

   // m12_59 = W*in
   wire signed [9:0] m12_59;
   assign m12_59 ={ {4{in12[5]}} , in12[5:0] };

   // m12_60 = W*in
   wire signed [9:0] m12_60;
   assign m12_60 ={ {4{in12[5]}} , in12[5:0] };

   // m12_61 = W*in
   wire signed [9:0] m12_61;
   assign m12_61 =10'b0;

   // m12_62 = W*in
   wire signed [9:0] m12_62;
   assign m12_62 =10'b0;

   // m12_63 = W*in
   wire signed [9:0] m12_63;
   assign m12_63 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_64 = W*in
   wire signed [9:0] m12_64;
   assign m12_64 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_65 = W*in
   wire signed [9:0] m12_65;
   assign m12_65 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_66 = W*in
   wire signed [9:0] m12_66;
   assign m12_66 ={ {4{in12[5]}} , in12[5:0] };

   // m12_67 = W*in
   wire signed [9:0] m12_67;
   assign m12_67 =10'b0;

   // m12_68 = W*in
   wire signed [9:0] m12_68;
   assign m12_68 =10'b0;

   // m12_69 = W*in
   wire signed [9:0] m12_69;
   assign m12_69 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_70 = W*in
   wire signed [9:0] m12_70;
   assign m12_70 =10'b0;

   // m12_71 = W*in
   wire signed [9:0] m12_71;
   assign m12_71 =10'b0;

   // m12_72 = W*in
   wire signed [9:0] m12_72;
   assign m12_72 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_73 = W*in
   wire signed [9:0] m12_73;
   assign m12_73 =10'b0;

   // m12_74 = W*in
   wire signed [9:0] m12_74;
   assign m12_74 ={ {5{neg12[5]}} , neg12[5:1] };

   // m12_75 = W*in
   wire signed [9:0] m12_75;
   assign m12_75 ={ {5{in12[5]}} , in12[5:1] };

   // m12_76 = W*in
   wire signed [9:0] m12_76;
   assign m12_76 =10'b0;

   // m12_77 = W*in
   wire signed [9:0] m12_77;
   assign m12_77 =10'b0;

   // m12_78 = W*in
   wire signed [9:0] m12_78;
   assign m12_78 =10'b0;

   // m12_79 = W*in
   wire signed [9:0] m12_79;
   assign m12_79 =10'b0;

   // m12_80 = W*in
   wire signed [9:0] m12_80;
   assign m12_80 =10'b0;

   // m12_81 = W*in
   wire signed [9:0] m12_81;
   assign m12_81 =10'b0;

   // m12_82 = W*in
   wire signed [9:0] m12_82;
   assign m12_82 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_83 = W*in
   wire signed [9:0] m12_83;
   assign m12_83 =10'b0;

   // m12_84 = W*in
   wire signed [9:0] m12_84;
   assign m12_84 =10'b0;

   // m12_85 = W*in
   wire signed [9:0] m12_85;
   assign m12_85 =10'b0;

   // m12_86 = W*in
   wire signed [9:0] m12_86;
   assign m12_86 =10'b0;

   // m12_87 = W*in
   wire signed [9:0] m12_87;
   assign m12_87 =10'b0;

   // m12_88 = W*in
   wire signed [9:0] m12_88;
   assign m12_88 =10'b0;

   // m12_89 = W*in
   wire signed [9:0] m12_89;
   assign m12_89 =10'b0;

   // m12_90 = W*in
   wire signed [9:0] m12_90;
   assign m12_90 =10'b0;

   // m12_91 = W*in
   wire signed [9:0] m12_91;
   assign m12_91 =10'b0;

   // m12_92 = W*in
   wire signed [9:0] m12_92;
   assign m12_92 =10'b0;

   // m12_93 = W*in
   wire signed [9:0] m12_93;
   assign m12_93 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_94 = W*in
   wire signed [9:0] m12_94;
   assign m12_94 =10'b0;

   // m12_95 = W*in
   wire signed [9:0] m12_95;
   assign m12_95 =10'b0;

   // m12_96 = W*in
   wire signed [9:0] m12_96;
   assign m12_96 =10'b0;

   // m12_97 = W*in
   wire signed [9:0] m12_97;
   assign m12_97 =10'b0;

   // m12_98 = W*in
   wire signed [9:0] m12_98;
   assign m12_98 =10'b0;

   // m12_99 = W*in
   wire signed [9:0] m12_99;
   assign m12_99 =10'b0;

   // m12_100 = W*in
   wire signed [9:0] m12_100;
   assign m12_100 ={ {3{in12[5]}} , in12 , {1{1'b0}} };

   // m12_101 = W*in
   wire signed [9:0] m12_101;
   assign m12_101 =10'b0;

   // m12_102 = W*in
   wire signed [9:0] m12_102;
   assign m12_102 =10'b0;

   // m12_103 = W*in
   wire signed [9:0] m12_103;
   assign m12_103 ={ {4{in12[5]}} , in12[5:0] };

   // m12_104 = W*in
   wire signed [9:0] m12_104;
   assign m12_104 ={ {4{in12[5]}} , in12[5:0] };

   // m12_105 = W*in
   wire signed [9:0] m12_105;
   assign m12_105 =10'b0;

   // m12_106 = W*in
   wire signed [9:0] m12_106;
   assign m12_106 =10'b0;

   // m12_107 = W*in
   wire signed [9:0] m12_107;
   assign m12_107 ={ {4{in12[5]}} , in12[5:0] };

   // m12_108 = W*in
   wire signed [9:0] m12_108;
   assign m12_108 =10'b0;

   // m12_109 = W*in
   wire signed [9:0] m12_109;
   assign m12_109 =10'b0;

   // m12_110 = W*in
   wire signed [9:0] m12_110;
   assign m12_110 =10'b0;

   // m12_111 = W*in
   wire signed [9:0] m12_111;
   assign m12_111 =10'b0;

   // m12_112 = W*in
   wire signed [9:0] m12_112;
   assign m12_112 ={ {4{in12[5]}} , in12[5:0] };

   // m12_113 = W*in
   wire signed [9:0] m12_113;
   assign m12_113 ={ {4{neg12[5]}} , neg12[5:0] };

   // m12_114 = W*in
   wire signed [9:0] m12_114;
   assign m12_114 =10'b0;

   // m12_115 = W*in
   wire signed [9:0] m12_115;
   assign m12_115 =10'b0;

   // m12_116 = W*in
   wire signed [9:0] m12_116;
   assign m12_116 ={ {4{in12[5]}} , in12[5:0] };

   // m12_117 = W*in
   wire signed [9:0] m12_117;
   assign m12_117 =10'b0;

   // m13_1 = W*in
   wire signed [9:0] m13_1;
   assign m13_1 =10'b0;

   // m13_2 = W*in
   wire signed [9:0] m13_2;
   assign m13_2 =10'b0;

   // m13_3 = W*in
   wire signed [9:0] m13_3;
   assign m13_3 =10'b0;

   // m13_4 = W*in
   wire signed [9:0] m13_4;
   assign m13_4 =10'b0;

   // m13_5 = W*in
   wire signed [9:0] m13_5;
   assign m13_5 =10'b0;

   // m13_6 = W*in
   wire signed [9:0] m13_6;
   assign m13_6 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_7 = W*in
   wire signed [9:0] m13_7;
   assign m13_7 =10'b0;

   // m13_8 = W*in
   wire signed [9:0] m13_8;
   assign m13_8 =10'b0;

   // m13_9 = W*in
   wire signed [9:0] m13_9;
   assign m13_9 =10'b0;

   // m13_10 = W*in
   wire signed [9:0] m13_10;
   assign m13_10 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_11 = W*in
   wire signed [9:0] m13_11;
   assign m13_11 =10'b0;

   // m13_12 = W*in
   wire signed [9:0] m13_12;
   assign m13_12 =10'b0;

   // m13_13 = W*in
   wire signed [9:0] m13_13;
   assign m13_13 ={ {4{in13[5]}} , in13[5:0] };

   // m13_14 = W*in
   wire signed [9:0] m13_14;
   assign m13_14 =10'b0;

   // m13_15 = W*in
   wire signed [9:0] m13_15;
   assign m13_15 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_16 = W*in
   wire signed [9:0] m13_16;
   assign m13_16 =10'b0;

   // m13_17 = W*in
   wire signed [9:0] m13_17;
   assign m13_17 =10'b0;

   // m13_18 = W*in
   wire signed [9:0] m13_18;
   assign m13_18 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_19 = W*in
   wire signed [9:0] m13_19;
   assign m13_19 =10'b0;

   // m13_20 = W*in
   wire signed [9:0] m13_20;
   assign m13_20 =10'b0;

   // m13_21 = W*in
   wire signed [9:0] m13_21;
   assign m13_21 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_22 = W*in
   wire signed [9:0] m13_22;
   assign m13_22 ={ {5{neg13[5]}} , neg13[5:1] };

   // m13_23 = W*in
   wire signed [9:0] m13_23;
   assign m13_23 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_24 = W*in
   wire signed [9:0] m13_24;
   assign m13_24 =10'b0;

   // m13_25 = W*in
   wire signed [9:0] m13_25;
   assign m13_25 =10'b0;

   // m13_26 = W*in
   wire signed [9:0] m13_26;
   assign m13_26 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_27 = W*in
   wire signed [9:0] m13_27;
   assign m13_27 ={ {5{in13[5]}} , in13[5:1] };

   // m13_28 = W*in
   wire signed [9:0] m13_28;
   assign m13_28 ={ {5{in13[5]}} , in13[5:1] };

   // m13_29 = W*in
   wire signed [9:0] m13_29;
   assign m13_29 =10'b0;

   // m13_30 = W*in
   wire signed [9:0] m13_30;
   assign m13_30 =10'b0;

   // m13_31 = W*in
   wire signed [9:0] m13_31;
   assign m13_31 ={ {5{neg13[5]}} , neg13[5:1] };

   // m13_32 = W*in
   wire signed [9:0] m13_32;
   assign m13_32 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_33 = W*in
   wire signed [9:0] m13_33;
   assign m13_33 =10'b0;

   // m13_34 = W*in
   wire signed [9:0] m13_34;
   assign m13_34 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_35 = W*in
   wire signed [9:0] m13_35;
   assign m13_35 =10'b0;

   // m13_36 = W*in
   wire signed [9:0] m13_36;
   assign m13_36 ={ {5{in13[5]}} , in13[5:1] };

   // m13_37 = W*in
   wire signed [9:0] m13_37;
   assign m13_37 =10'b0;

   // m13_38 = W*in
   wire signed [9:0] m13_38;
   assign m13_38 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_39 = W*in
   wire signed [9:0] m13_39;
   assign m13_39 =10'b0;

   // m13_40 = W*in
   wire signed [9:0] m13_40;
   assign m13_40 =10'b0;

   // m13_41 = W*in
   wire signed [9:0] m13_41;
   assign m13_41 ={ {4{in13[5]}} , in13[5:0] };

   // m13_42 = W*in
   wire signed [9:0] m13_42;
   assign m13_42 =10'b0;

   // m13_43 = W*in
   wire signed [9:0] m13_43;
   assign m13_43 =10'b0;

   // m13_44 = W*in
   wire signed [9:0] m13_44;
   assign m13_44 ={ {4{in13[5]}} , in13[5:0] };

   // m13_45 = W*in
   wire signed [9:0] m13_45;
   assign m13_45 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_46 = W*in
   wire signed [9:0] m13_46;
   assign m13_46 =10'b0;

   // m13_47 = W*in
   wire signed [9:0] m13_47;
   assign m13_47 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_48 = W*in
   wire signed [9:0] m13_48;
   assign m13_48 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_49 = W*in
   wire signed [9:0] m13_49;
   assign m13_49 ={ {4{in13[5]}} , in13[5:0] };

   // m13_50 = W*in
   wire signed [9:0] m13_50;
   assign m13_50 =10'b0;

   // m13_51 = W*in
   wire signed [9:0] m13_51;
   assign m13_51 =10'b0;

   // m13_52 = W*in
   wire signed [9:0] m13_52;
   assign m13_52 =10'b0;

   // m13_53 = W*in
   wire signed [9:0] m13_53;
   assign m13_53 =10'b0;

   // m13_54 = W*in
   wire signed [9:0] m13_54;
   assign m13_54 ={ {4{in13[5]}} , in13[5:0] };

   // m13_55 = W*in
   wire signed [9:0] m13_55;
   assign m13_55 =10'b0;

   // m13_56 = W*in
   wire signed [9:0] m13_56;
   assign m13_56 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_57 = W*in
   wire signed [9:0] m13_57;
   assign m13_57 =10'b0;

   // m13_58 = W*in
   wire signed [9:0] m13_58;
   assign m13_58 =10'b0;

   // m13_59 = W*in
   wire signed [9:0] m13_59;
   assign m13_59 ={ {4{in13[5]}} , in13[5:0] };

   // m13_60 = W*in
   wire signed [9:0] m13_60;
   assign m13_60 ={ {4{in13[5]}} , in13[5:0] };

   // m13_61 = W*in
   wire signed [9:0] m13_61;
   assign m13_61 =10'b0;

   // m13_62 = W*in
   wire signed [9:0] m13_62;
   assign m13_62 =10'b0;

   // m13_63 = W*in
   wire signed [9:0] m13_63;
   assign m13_63 =10'b0;

   // m13_64 = W*in
   wire signed [9:0] m13_64;
   assign m13_64 ={ {5{neg13[5]}} , neg13[5:1] };

   // m13_65 = W*in
   wire signed [9:0] m13_65;
   assign m13_65 ={ {4{in13[5]}} , in13[5:0] };

   // m13_66 = W*in
   wire signed [9:0] m13_66;
   assign m13_66 ={ {4{in13[5]}} , in13[5:0] };

   // m13_67 = W*in
   wire signed [9:0] m13_67;
   assign m13_67 =10'b0;

   // m13_68 = W*in
   wire signed [9:0] m13_68;
   assign m13_68 =10'b0;

   // m13_69 = W*in
   wire signed [9:0] m13_69;
   assign m13_69 ={ {5{neg13[5]}} , neg13[5:1] };

   // m13_70 = W*in
   wire signed [9:0] m13_70;
   assign m13_70 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_71 = W*in
   wire signed [9:0] m13_71;
   assign m13_71 =10'b0;

   // m13_72 = W*in
   wire signed [9:0] m13_72;
   assign m13_72 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_73 = W*in
   wire signed [9:0] m13_73;
   assign m13_73 =10'b0;

   // m13_74 = W*in
   wire signed [9:0] m13_74;
   assign m13_74 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_75 = W*in
   wire signed [9:0] m13_75;
   assign m13_75 ={ {4{in13[5]}} , in13[5:0] };

   // m13_76 = W*in
   wire signed [9:0] m13_76;
   assign m13_76 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_77 = W*in
   wire signed [9:0] m13_77;
   assign m13_77 =10'b0;

   // m13_78 = W*in
   wire signed [9:0] m13_78;
   assign m13_78 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_79 = W*in
   wire signed [9:0] m13_79;
   assign m13_79 ={ {4{in13[5]}} , in13[5:0] };

   // m13_80 = W*in
   wire signed [9:0] m13_80;
   assign m13_80 =10'b0;

   // m13_81 = W*in
   wire signed [9:0] m13_81;
   assign m13_81 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_82 = W*in
   wire signed [9:0] m13_82;
   assign m13_82 =10'b0;

   // m13_83 = W*in
   wire signed [9:0] m13_83;
   assign m13_83 =10'b0;

   // m13_84 = W*in
   wire signed [9:0] m13_84;
   assign m13_84 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_85 = W*in
   wire signed [9:0] m13_85;
   assign m13_85 =10'b0;

   // m13_86 = W*in
   wire signed [9:0] m13_86;
   assign m13_86 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_87 = W*in
   wire signed [9:0] m13_87;
   assign m13_87 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_88 = W*in
   wire signed [9:0] m13_88;
   assign m13_88 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_89 = W*in
   wire signed [9:0] m13_89;
   assign m13_89 =10'b0;

   // m13_90 = W*in
   wire signed [9:0] m13_90;
   assign m13_90 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_91 = W*in
   wire signed [9:0] m13_91;
   assign m13_91 ={ {5{neg13[5]}} , neg13[5:1] };

   // m13_92 = W*in
   wire signed [9:0] m13_92;
   assign m13_92 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_93 = W*in
   wire signed [9:0] m13_93;
   assign m13_93 =10'b0;

   // m13_94 = W*in
   wire signed [9:0] m13_94;
   assign m13_94 =10'b0;

   // m13_95 = W*in
   wire signed [9:0] m13_95;
   assign m13_95 =10'b0;

   // m13_96 = W*in
   wire signed [9:0] m13_96;
   assign m13_96 =10'b0;

   // m13_97 = W*in
   wire signed [9:0] m13_97;
   assign m13_97 =10'b0;

   // m13_98 = W*in
   wire signed [9:0] m13_98;
   assign m13_98 =10'b0;

   // m13_99 = W*in
   wire signed [9:0] m13_99;
   assign m13_99 ={ {3{neg13[5]}} , neg13 , {1{1'b0}} };

   // m13_100 = W*in
   wire signed [9:0] m13_100;
   assign m13_100 ={ {4{in13[5]}} , in13[5:0] };

   // m13_101 = W*in
   wire signed [9:0] m13_101;
   assign m13_101 ={ {4{in13[5]}} , in13[5:0] };

   // m13_102 = W*in
   wire signed [9:0] m13_102;
   assign m13_102 =10'b0;

   // m13_103 = W*in
   wire signed [9:0] m13_103;
   assign m13_103 ={ {4{in13[5]}} , in13[5:0] };

   // m13_104 = W*in
   wire signed [9:0] m13_104;
   assign m13_104 ={ {4{in13[5]}} , in13[5:0] };

   // m13_105 = W*in
   wire signed [9:0] m13_105;
   assign m13_105 =10'b0;

   // m13_106 = W*in
   wire signed [9:0] m13_106;
   assign m13_106 =10'b0;

   // m13_107 = W*in
   wire signed [9:0] m13_107;
   assign m13_107 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_108 = W*in
   wire signed [9:0] m13_108;
   assign m13_108 ={ {4{in13[5]}} , in13[5:0] };

   // m13_109 = W*in
   wire signed [9:0] m13_109;
   assign m13_109 ={ {4{in13[5]}} , in13[5:0] };

   // m13_110 = W*in
   wire signed [9:0] m13_110;
   assign m13_110 =10'b0;

   // m13_111 = W*in
   wire signed [9:0] m13_111;
   assign m13_111 =10'b0;

   // m13_112 = W*in
   wire signed [9:0] m13_112;
   assign m13_112 =10'b0;

   // m13_113 = W*in
   wire signed [9:0] m13_113;
   assign m13_113 =10'b0;

   // m13_114 = W*in
   wire signed [9:0] m13_114;
   assign m13_114 ={ {4{neg13[5]}} , neg13[5:0] };

   // m13_115 = W*in
   wire signed [9:0] m13_115;
   assign m13_115 =10'b0;

   // m13_116 = W*in
   wire signed [9:0] m13_116;
   assign m13_116 ={ {4{in13[5]}} , in13[5:0] };

   // m13_117 = W*in
   wire signed [9:0] m13_117;
   assign m13_117 ={ {4{in13[5]}} , in13[5:0] };

   // m14_1 = W*in
   wire signed [9:0] m14_1;
   assign m14_1 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_2 = W*in
   wire signed [9:0] m14_2;
   assign m14_2 =10'b0;

   // m14_3 = W*in
   wire signed [9:0] m14_3;
   assign m14_3 =10'b0;

   // m14_4 = W*in
   wire signed [9:0] m14_4;
   assign m14_4 =10'b0;

   // m14_5 = W*in
   wire signed [9:0] m14_5;
   assign m14_5 =10'b0;

   // m14_6 = W*in
   wire signed [9:0] m14_6;
   assign m14_6 =10'b0;

   // m14_7 = W*in
   wire signed [9:0] m14_7;
   assign m14_7 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_8 = W*in
   wire signed [9:0] m14_8;
   assign m14_8 =10'b0;

   // m14_9 = W*in
   wire signed [9:0] m14_9;
   assign m14_9 =10'b0;

   // m14_10 = W*in
   wire signed [9:0] m14_10;
   assign m14_10 =10'b0;

   // m14_11 = W*in
   wire signed [9:0] m14_11;
   assign m14_11 ={ {4{in14[5]}} , in14[5:0] };

   // m14_12 = W*in
   wire signed [9:0] m14_12;
   assign m14_12 ={ {5{in14[5]}} , in14[5:1] };

   // m14_13 = W*in
   wire signed [9:0] m14_13;
   assign m14_13 =10'b0;

   // m14_14 = W*in
   wire signed [9:0] m14_14;
   assign m14_14 =10'b0;

   // m14_15 = W*in
   wire signed [9:0] m14_15;
   assign m14_15 =10'b0;

   // m14_16 = W*in
   wire signed [9:0] m14_16;
   assign m14_16 ={ {4{in14[5]}} , in14[5:0] };

   // m14_17 = W*in
   wire signed [9:0] m14_17;
   assign m14_17 =10'b0;

   // m14_18 = W*in
   wire signed [9:0] m14_18;
   assign m14_18 ={ {5{neg14[5]}} , neg14[5:1] };

   // m14_19 = W*in
   wire signed [9:0] m14_19;
   assign m14_19 ={ {4{in14[5]}} , in14[5:0] };

   // m14_20 = W*in
   wire signed [9:0] m14_20;
   assign m14_20 ={ {4{in14[5]}} , in14[5:0] };

   // m14_21 = W*in
   wire signed [9:0] m14_21;
   assign m14_21 ={ {4{in14[5]}} , in14[5:0] };

   // m14_22 = W*in
   wire signed [9:0] m14_22;
   assign m14_22 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_23 = W*in
   wire signed [9:0] m14_23;
   assign m14_23 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_24 = W*in
   wire signed [9:0] m14_24;
   assign m14_24 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_25 = W*in
   wire signed [9:0] m14_25;
   assign m14_25 =10'b0;

   // m14_26 = W*in
   wire signed [9:0] m14_26;
   assign m14_26 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_27 = W*in
   wire signed [9:0] m14_27;
   assign m14_27 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_28 = W*in
   wire signed [9:0] m14_28;
   assign m14_28 =10'b0;

   // m14_29 = W*in
   wire signed [9:0] m14_29;
   assign m14_29 =10'b0;

   // m14_30 = W*in
   wire signed [9:0] m14_30;
   assign m14_30 ={ {4{in14[5]}} , in14[5:0] };

   // m14_31 = W*in
   wire signed [9:0] m14_31;
   assign m14_31 =10'b0;

   // m14_32 = W*in
   wire signed [9:0] m14_32;
   assign m14_32 =10'b0;

   // m14_33 = W*in
   wire signed [9:0] m14_33;
   assign m14_33 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_34 = W*in
   wire signed [9:0] m14_34;
   assign m14_34 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_35 = W*in
   wire signed [9:0] m14_35;
   assign m14_35 ={ {4{in14[5]}} , in14[5:0] };

   // m14_36 = W*in
   wire signed [9:0] m14_36;
   assign m14_36 =10'b0;

   // m14_37 = W*in
   wire signed [9:0] m14_37;
   assign m14_37 =10'b0;

   // m14_38 = W*in
   wire signed [9:0] m14_38;
   assign m14_38 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_39 = W*in
   wire signed [9:0] m14_39;
   assign m14_39 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_40 = W*in
   wire signed [9:0] m14_40;
   assign m14_40 ={ {4{in14[5]}} , in14[5:0] };

   // m14_41 = W*in
   wire signed [9:0] m14_41;
   assign m14_41 ={ {4{in14[5]}} , in14[5:0] };

   // m14_42 = W*in
   wire signed [9:0] m14_42;
   assign m14_42 =10'b0;

   // m14_43 = W*in
   wire signed [9:0] m14_43;
   assign m14_43 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_44 = W*in
   wire signed [9:0] m14_44;
   assign m14_44 ={ {4{in14[5]}} , in14[5:0] };

   // m14_45 = W*in
   wire signed [9:0] m14_45;
   assign m14_45 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_46 = W*in
   wire signed [9:0] m14_46;
   assign m14_46 =10'b0;

   // m14_47 = W*in
   wire signed [9:0] m14_47;
   assign m14_47 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_48 = W*in
   wire signed [9:0] m14_48;
   assign m14_48 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_49 = W*in
   wire signed [9:0] m14_49;
   assign m14_49 ={ {4{in14[5]}} , in14[5:0] };

   // m14_50 = W*in
   wire signed [9:0] m14_50;
   assign m14_50 =10'b0;

   // m14_51 = W*in
   wire signed [9:0] m14_51;
   assign m14_51 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_52 = W*in
   wire signed [9:0] m14_52;
   assign m14_52 =10'b0;

   // m14_53 = W*in
   wire signed [9:0] m14_53;
   assign m14_53 ={ {4{in14[5]}} , in14[5:0] };

   // m14_54 = W*in
   wire signed [9:0] m14_54;
   assign m14_54 ={ {4{in14[5]}} , in14[5:0] };

   // m14_55 = W*in
   wire signed [9:0] m14_55;
   assign m14_55 =10'b0;

   // m14_56 = W*in
   wire signed [9:0] m14_56;
   assign m14_56 =10'b0;

   // m14_57 = W*in
   wire signed [9:0] m14_57;
   assign m14_57 =10'b0;

   // m14_58 = W*in
   wire signed [9:0] m14_58;
   assign m14_58 =10'b0;

   // m14_59 = W*in
   wire signed [9:0] m14_59;
   assign m14_59 =10'b0;

   // m14_60 = W*in
   wire signed [9:0] m14_60;
   assign m14_60 ={ {5{in14[5]}} , in14[5:1] };

   // m14_61 = W*in
   wire signed [9:0] m14_61;
   assign m14_61 ={ {4{in14[5]}} , in14[5:0] };

   // m14_62 = W*in
   wire signed [9:0] m14_62;
   assign m14_62 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_63 = W*in
   wire signed [9:0] m14_63;
   assign m14_63 =10'b0;

   // m14_64 = W*in
   wire signed [9:0] m14_64;
   assign m14_64 =10'b0;

   // m14_65 = W*in
   wire signed [9:0] m14_65;
   assign m14_65 ={ {4{in14[5]}} , in14[5:0] };

   // m14_66 = W*in
   wire signed [9:0] m14_66;
   assign m14_66 ={ {4{in14[5]}} , in14[5:0] };

   // m14_67 = W*in
   wire signed [9:0] m14_67;
   assign m14_67 ={ {4{in14[5]}} , in14[5:0] };

   // m14_68 = W*in
   wire signed [9:0] m14_68;
   assign m14_68 =10'b0;

   // m14_69 = W*in
   wire signed [9:0] m14_69;
   assign m14_69 =10'b0;

   // m14_70 = W*in
   wire signed [9:0] m14_70;
   assign m14_70 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_71 = W*in
   wire signed [9:0] m14_71;
   assign m14_71 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_72 = W*in
   wire signed [9:0] m14_72;
   assign m14_72 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_73 = W*in
   wire signed [9:0] m14_73;
   assign m14_73 =10'b0;

   // m14_74 = W*in
   wire signed [9:0] m14_74;
   assign m14_74 =10'b0;

   // m14_75 = W*in
   wire signed [9:0] m14_75;
   assign m14_75 ={ {5{in14[5]}} , in14[5:1] };

   // m14_76 = W*in
   wire signed [9:0] m14_76;
   assign m14_76 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_77 = W*in
   wire signed [9:0] m14_77;
   assign m14_77 =10'b0;

   // m14_78 = W*in
   wire signed [9:0] m14_78;
   assign m14_78 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_79 = W*in
   wire signed [9:0] m14_79;
   assign m14_79 ={ {3{in14[5]}} , in14 , {1{1'b0}} };

   // m14_80 = W*in
   wire signed [9:0] m14_80;
   assign m14_80 =10'b0;

   // m14_81 = W*in
   wire signed [9:0] m14_81;
   assign m14_81 =10'b0;

   // m14_82 = W*in
   wire signed [9:0] m14_82;
   assign m14_82 ={ {4{in14[5]}} , in14[5:0] };

   // m14_83 = W*in
   wire signed [9:0] m14_83;
   assign m14_83 =10'b0;

   // m14_84 = W*in
   wire signed [9:0] m14_84;
   assign m14_84 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_85 = W*in
   wire signed [9:0] m14_85;
   assign m14_85 =10'b0;

   // m14_86 = W*in
   wire signed [9:0] m14_86;
   assign m14_86 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_87 = W*in
   wire signed [9:0] m14_87;
   assign m14_87 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_88 = W*in
   wire signed [9:0] m14_88;
   assign m14_88 =10'b0;

   // m14_89 = W*in
   wire signed [9:0] m14_89;
   assign m14_89 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_90 = W*in
   wire signed [9:0] m14_90;
   assign m14_90 =10'b0;

   // m14_91 = W*in
   wire signed [9:0] m14_91;
   assign m14_91 ={ {4{in14[5]}} , in14[5:0] };

   // m14_92 = W*in
   wire signed [9:0] m14_92;
   assign m14_92 =10'b0;

   // m14_93 = W*in
   wire signed [9:0] m14_93;
   assign m14_93 =10'b0;

   // m14_94 = W*in
   wire signed [9:0] m14_94;
   assign m14_94 ={ {4{in14[5]}} , in14[5:0] };

   // m14_95 = W*in
   wire signed [9:0] m14_95;
   assign m14_95 =10'b0;

   // m14_96 = W*in
   wire signed [9:0] m14_96;
   assign m14_96 =10'b0;

   // m14_97 = W*in
   wire signed [9:0] m14_97;
   assign m14_97 =10'b0;

   // m14_98 = W*in
   wire signed [9:0] m14_98;
   assign m14_98 =10'b0;

   // m14_99 = W*in
   wire signed [9:0] m14_99;
   assign m14_99 ={ {3{neg14[5]}} , neg14 , {1{1'b0}} };

   // m14_100 = W*in
   wire signed [9:0] m14_100;
   assign m14_100 =10'b0;

   // m14_101 = W*in
   wire signed [9:0] m14_101;
   assign m14_101 =10'b0;

   // m14_102 = W*in
   wire signed [9:0] m14_102;
   assign m14_102 ={ {4{in14[5]}} , in14[5:0] };

   // m14_103 = W*in
   wire signed [9:0] m14_103;
   assign m14_103 =10'b0;

   // m14_104 = W*in
   wire signed [9:0] m14_104;
   assign m14_104 =10'b0;

   // m14_105 = W*in
   wire signed [9:0] m14_105;
   assign m14_105 =10'b0;

   // m14_106 = W*in
   wire signed [9:0] m14_106;
   assign m14_106 ={ {4{in14[5]}} , in14[5:0] };

   // m14_107 = W*in
   wire signed [9:0] m14_107;
   assign m14_107 =10'b0;

   // m14_108 = W*in
   wire signed [9:0] m14_108;
   assign m14_108 ={ {4{in14[5]}} , in14[5:0] };

   // m14_109 = W*in
   wire signed [9:0] m14_109;
   assign m14_109 =10'b0;

   // m14_110 = W*in
   wire signed [9:0] m14_110;
   assign m14_110 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_111 = W*in
   wire signed [9:0] m14_111;
   assign m14_111 =10'b0;

   // m14_112 = W*in
   wire signed [9:0] m14_112;
   assign m14_112 =10'b0;

   // m14_113 = W*in
   wire signed [9:0] m14_113;
   assign m14_113 =10'b0;

   // m14_114 = W*in
   wire signed [9:0] m14_114;
   assign m14_114 ={ {4{neg14[5]}} , neg14[5:0] };

   // m14_115 = W*in
   wire signed [9:0] m14_115;
   assign m14_115 =10'b0;

   // m14_116 = W*in
   wire signed [9:0] m14_116;
   assign m14_116 ={ {4{in14[5]}} , in14[5:0] };

   // m14_117 = W*in
   wire signed [9:0] m14_117;
   assign m14_117 ={ {4{in14[5]}} , in14[5:0] };

   // m15_1 = W*in
   wire signed [9:0] m15_1;
   assign m15_1 =10'b0;

   // m15_2 = W*in
   wire signed [9:0] m15_2;
   assign m15_2 =10'b0;

   // m15_3 = W*in
   wire signed [9:0] m15_3;
   assign m15_3 =10'b0;

   // m15_4 = W*in
   wire signed [9:0] m15_4;
   assign m15_4 =10'b0;

   // m15_5 = W*in
   wire signed [9:0] m15_5;
   assign m15_5 =10'b0;

   // m15_6 = W*in
   wire signed [9:0] m15_6;
   assign m15_6 =10'b0;

   // m15_7 = W*in
   wire signed [9:0] m15_7;
   assign m15_7 ={ {4{in15[5]}} , in15[5:0] };

   // m15_8 = W*in
   wire signed [9:0] m15_8;
   assign m15_8 =10'b0;

   // m15_9 = W*in
   wire signed [9:0] m15_9;
   assign m15_9 =10'b0;

   // m15_10 = W*in
   wire signed [9:0] m15_10;
   assign m15_10 =10'b0;

   // m15_11 = W*in
   wire signed [9:0] m15_11;
   assign m15_11 ={ {4{in15[5]}} , in15[5:0] };

   // m15_12 = W*in
   wire signed [9:0] m15_12;
   assign m15_12 =10'b0;

   // m15_13 = W*in
   wire signed [9:0] m15_13;
   assign m15_13 =10'b0;

   // m15_14 = W*in
   wire signed [9:0] m15_14;
   assign m15_14 =10'b0;

   // m15_15 = W*in
   wire signed [9:0] m15_15;
   assign m15_15 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_16 = W*in
   wire signed [9:0] m15_16;
   assign m15_16 ={ {4{in15[5]}} , in15[5:0] };

   // m15_17 = W*in
   wire signed [9:0] m15_17;
   assign m15_17 =10'b0;

   // m15_18 = W*in
   wire signed [9:0] m15_18;
   assign m15_18 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_19 = W*in
   wire signed [9:0] m15_19;
   assign m15_19 ={ {5{in15[5]}} , in15[5:1] };

   // m15_20 = W*in
   wire signed [9:0] m15_20;
   assign m15_20 =10'b0;

   // m15_21 = W*in
   wire signed [9:0] m15_21;
   assign m15_21 =10'b0;

   // m15_22 = W*in
   wire signed [9:0] m15_22;
   assign m15_22 ={ {5{neg15[5]}} , neg15[5:1] };

   // m15_23 = W*in
   wire signed [9:0] m15_23;
   assign m15_23 =10'b0;

   // m15_24 = W*in
   wire signed [9:0] m15_24;
   assign m15_24 =10'b0;

   // m15_25 = W*in
   wire signed [9:0] m15_25;
   assign m15_25 ={ {4{in15[5]}} , in15[5:0] };

   // m15_26 = W*in
   wire signed [9:0] m15_26;
   assign m15_26 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_27 = W*in
   wire signed [9:0] m15_27;
   assign m15_27 ={ {5{neg15[5]}} , neg15[5:1] };

   // m15_28 = W*in
   wire signed [9:0] m15_28;
   assign m15_28 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_29 = W*in
   wire signed [9:0] m15_29;
   assign m15_29 =10'b0;

   // m15_30 = W*in
   wire signed [9:0] m15_30;
   assign m15_30 =10'b0;

   // m15_31 = W*in
   wire signed [9:0] m15_31;
   assign m15_31 =10'b0;

   // m15_32 = W*in
   wire signed [9:0] m15_32;
   assign m15_32 =10'b0;

   // m15_33 = W*in
   wire signed [9:0] m15_33;
   assign m15_33 =10'b0;

   // m15_34 = W*in
   wire signed [9:0] m15_34;
   assign m15_34 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_35 = W*in
   wire signed [9:0] m15_35;
   assign m15_35 =10'b0;

   // m15_36 = W*in
   wire signed [9:0] m15_36;
   assign m15_36 ={ {4{in15[5]}} , in15[5:0] };

   // m15_37 = W*in
   wire signed [9:0] m15_37;
   assign m15_37 =10'b0;

   // m15_38 = W*in
   wire signed [9:0] m15_38;
   assign m15_38 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_39 = W*in
   wire signed [9:0] m15_39;
   assign m15_39 =10'b0;

   // m15_40 = W*in
   wire signed [9:0] m15_40;
   assign m15_40 =10'b0;

   // m15_41 = W*in
   wire signed [9:0] m15_41;
   assign m15_41 ={ {4{in15[5]}} , in15[5:0] };

   // m15_42 = W*in
   wire signed [9:0] m15_42;
   assign m15_42 =10'b0;

   // m15_43 = W*in
   wire signed [9:0] m15_43;
   assign m15_43 =10'b0;

   // m15_44 = W*in
   wire signed [9:0] m15_44;
   assign m15_44 =10'b0;

   // m15_45 = W*in
   wire signed [9:0] m15_45;
   assign m15_45 =10'b0;

   // m15_46 = W*in
   wire signed [9:0] m15_46;
   assign m15_46 =10'b0;

   // m15_47 = W*in
   wire signed [9:0] m15_47;
   assign m15_47 =10'b0;

   // m15_48 = W*in
   wire signed [9:0] m15_48;
   assign m15_48 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_49 = W*in
   wire signed [9:0] m15_49;
   assign m15_49 ={ {4{in15[5]}} , in15[5:0] };

   // m15_50 = W*in
   wire signed [9:0] m15_50;
   assign m15_50 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_51 = W*in
   wire signed [9:0] m15_51;
   assign m15_51 =10'b0;

   // m15_52 = W*in
   wire signed [9:0] m15_52;
   assign m15_52 =10'b0;

   // m15_53 = W*in
   wire signed [9:0] m15_53;
   assign m15_53 ={ {4{in15[5]}} , in15[5:0] };

   // m15_54 = W*in
   wire signed [9:0] m15_54;
   assign m15_54 =10'b0;

   // m15_55 = W*in
   wire signed [9:0] m15_55;
   assign m15_55 =10'b0;

   // m15_56 = W*in
   wire signed [9:0] m15_56;
   assign m15_56 ={ {4{in15[5]}} , in15[5:0] };

   // m15_57 = W*in
   wire signed [9:0] m15_57;
   assign m15_57 =10'b0;

   // m15_58 = W*in
   wire signed [9:0] m15_58;
   assign m15_58 =10'b0;

   // m15_59 = W*in
   wire signed [9:0] m15_59;
   assign m15_59 =10'b0;

   // m15_60 = W*in
   wire signed [9:0] m15_60;
   assign m15_60 =10'b0;

   // m15_61 = W*in
   wire signed [9:0] m15_61;
   assign m15_61 =10'b0;

   // m15_62 = W*in
   wire signed [9:0] m15_62;
   assign m15_62 =10'b0;

   // m15_63 = W*in
   wire signed [9:0] m15_63;
   assign m15_63 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_64 = W*in
   wire signed [9:0] m15_64;
   assign m15_64 ={ {5{neg15[5]}} , neg15[5:1] };

   // m15_65 = W*in
   wire signed [9:0] m15_65;
   assign m15_65 ={ {5{in15[5]}} , in15[5:1] };

   // m15_66 = W*in
   wire signed [9:0] m15_66;
   assign m15_66 ={ {4{in15[5]}} , in15[5:0] };

   // m15_67 = W*in
   wire signed [9:0] m15_67;
   assign m15_67 =10'b0;

   // m15_68 = W*in
   wire signed [9:0] m15_68;
   assign m15_68 =10'b0;

   // m15_69 = W*in
   wire signed [9:0] m15_69;
   assign m15_69 =10'b0;

   // m15_70 = W*in
   wire signed [9:0] m15_70;
   assign m15_70 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_71 = W*in
   wire signed [9:0] m15_71;
   assign m15_71 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_72 = W*in
   wire signed [9:0] m15_72;
   assign m15_72 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_73 = W*in
   wire signed [9:0] m15_73;
   assign m15_73 ={ {4{in15[5]}} , in15[5:0] };

   // m15_74 = W*in
   wire signed [9:0] m15_74;
   assign m15_74 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_75 = W*in
   wire signed [9:0] m15_75;
   assign m15_75 =10'b0;

   // m15_76 = W*in
   wire signed [9:0] m15_76;
   assign m15_76 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_77 = W*in
   wire signed [9:0] m15_77;
   assign m15_77 =10'b0;

   // m15_78 = W*in
   wire signed [9:0] m15_78;
   assign m15_78 =10'b0;

   // m15_79 = W*in
   wire signed [9:0] m15_79;
   assign m15_79 ={ {4{in15[5]}} , in15[5:0] };

   // m15_80 = W*in
   wire signed [9:0] m15_80;
   assign m15_80 =10'b0;

   // m15_81 = W*in
   wire signed [9:0] m15_81;
   assign m15_81 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_82 = W*in
   wire signed [9:0] m15_82;
   assign m15_82 =10'b0;

   // m15_83 = W*in
   wire signed [9:0] m15_83;
   assign m15_83 =10'b0;

   // m15_84 = W*in
   wire signed [9:0] m15_84;
   assign m15_84 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_85 = W*in
   wire signed [9:0] m15_85;
   assign m15_85 =10'b0;

   // m15_86 = W*in
   wire signed [9:0] m15_86;
   assign m15_86 ={ {5{neg15[5]}} , neg15[5:1] };

   // m15_87 = W*in
   wire signed [9:0] m15_87;
   assign m15_87 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_88 = W*in
   wire signed [9:0] m15_88;
   assign m15_88 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_89 = W*in
   wire signed [9:0] m15_89;
   assign m15_89 =10'b0;

   // m15_90 = W*in
   wire signed [9:0] m15_90;
   assign m15_90 =10'b0;

   // m15_91 = W*in
   wire signed [9:0] m15_91;
   assign m15_91 ={ {4{in15[5]}} , in15[5:0] };

   // m15_92 = W*in
   wire signed [9:0] m15_92;
   assign m15_92 ={ {4{neg15[5]}} , neg15[5:0] };

   // m15_93 = W*in
   wire signed [9:0] m15_93;
   assign m15_93 =10'b0;

   // m15_94 = W*in
   wire signed [9:0] m15_94;
   assign m15_94 ={ {4{in15[5]}} , in15[5:0] };

   // m15_95 = W*in
   wire signed [9:0] m15_95;
   assign m15_95 =10'b0;

   // m15_96 = W*in
   wire signed [9:0] m15_96;
   assign m15_96 =10'b0;

   // m15_97 = W*in
   wire signed [9:0] m15_97;
   assign m15_97 ={ {4{in15[5]}} , in15[5:0] };

   // m15_98 = W*in
   wire signed [9:0] m15_98;
   assign m15_98 =10'b0;

   // m15_99 = W*in
   wire signed [9:0] m15_99;
   assign m15_99 ={ {3{neg15[5]}} , neg15 , {1{1'b0}} };

   // m15_100 = W*in
   wire signed [9:0] m15_100;
   assign m15_100 =10'b0;

   // m15_101 = W*in
   wire signed [9:0] m15_101;
   assign m15_101 =10'b0;

   // m15_102 = W*in
   wire signed [9:0] m15_102;
   assign m15_102 ={ {3{in15[5]}} , in15 , {1{1'b0}} };

   // m15_103 = W*in
   wire signed [9:0] m15_103;
   assign m15_103 =10'b0;

   // m15_104 = W*in
   wire signed [9:0] m15_104;
   assign m15_104 =10'b0;

   // m15_105 = W*in
   wire signed [9:0] m15_105;
   assign m15_105 =10'b0;

   // m15_106 = W*in
   wire signed [9:0] m15_106;
   assign m15_106 ={ {4{in15[5]}} , in15[5:0] };

   // m15_107 = W*in
   wire signed [9:0] m15_107;
   assign m15_107 =10'b0;

   // m15_108 = W*in
   wire signed [9:0] m15_108;
   assign m15_108 =10'b0;

   // m15_109 = W*in
   wire signed [9:0] m15_109;
   assign m15_109 =10'b0;

   // m15_110 = W*in
   wire signed [9:0] m15_110;
   assign m15_110 =10'b0;

   // m15_111 = W*in
   wire signed [9:0] m15_111;
   assign m15_111 =10'b0;

   // m15_112 = W*in
   wire signed [9:0] m15_112;
   assign m15_112 =10'b0;

   // m15_113 = W*in
   wire signed [9:0] m15_113;
   assign m15_113 =10'b0;

   // m15_114 = W*in
   wire signed [9:0] m15_114;
   assign m15_114 =10'b0;

   // m15_115 = W*in
   wire signed [9:0] m15_115;
   assign m15_115 =10'b0;

   // m15_116 = W*in
   wire signed [9:0] m15_116;
   assign m15_116 =10'b0;

   // m15_117 = W*in
   wire signed [9:0] m15_117;
   assign m15_117 =10'b0;

   // m16_1 = W*in
   wire signed [9:0] m16_1;
   assign m16_1 =10'b0;

   // m16_2 = W*in
   wire signed [9:0] m16_2;
   assign m16_2 =10'b0;

   // m16_3 = W*in
   wire signed [9:0] m16_3;
   assign m16_3 =10'b0;

   // m16_4 = W*in
   wire signed [9:0] m16_4;
   assign m16_4 =10'b0;

   // m16_5 = W*in
   wire signed [9:0] m16_5;
   assign m16_5 =10'b0;

   // m16_6 = W*in
   wire signed [9:0] m16_6;
   assign m16_6 =10'b0;

   // m16_7 = W*in
   wire signed [9:0] m16_7;
   assign m16_7 =10'b0;

   // m16_8 = W*in
   wire signed [9:0] m16_8;
   assign m16_8 =10'b0;

   // m16_9 = W*in
   wire signed [9:0] m16_9;
   assign m16_9 =10'b0;

   // m16_10 = W*in
   wire signed [9:0] m16_10;
   assign m16_10 ={ {4{in16[5]}} , in16[5:0] };

   // m16_11 = W*in
   wire signed [9:0] m16_11;
   assign m16_11 =10'b0;

   // m16_12 = W*in
   wire signed [9:0] m16_12;
   assign m16_12 =10'b0;

   // m16_13 = W*in
   wire signed [9:0] m16_13;
   assign m16_13 =10'b0;

   // m16_14 = W*in
   wire signed [9:0] m16_14;
   assign m16_14 =10'b0;

   // m16_15 = W*in
   wire signed [9:0] m16_15;
   assign m16_15 =10'b0;

   // m16_16 = W*in
   wire signed [9:0] m16_16;
   assign m16_16 =10'b0;

   // m16_17 = W*in
   wire signed [9:0] m16_17;
   assign m16_17 =10'b0;

   // m16_18 = W*in
   wire signed [9:0] m16_18;
   assign m16_18 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_19 = W*in
   wire signed [9:0] m16_19;
   assign m16_19 ={ {4{in16[5]}} , in16[5:0] };

   // m16_20 = W*in
   wire signed [9:0] m16_20;
   assign m16_20 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_21 = W*in
   wire signed [9:0] m16_21;
   assign m16_21 ={ {4{in16[5]}} , in16[5:0] };

   // m16_22 = W*in
   wire signed [9:0] m16_22;
   assign m16_22 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_23 = W*in
   wire signed [9:0] m16_23;
   assign m16_23 =10'b0;

   // m16_24 = W*in
   wire signed [9:0] m16_24;
   assign m16_24 =10'b0;

   // m16_25 = W*in
   wire signed [9:0] m16_25;
   assign m16_25 =10'b0;

   // m16_26 = W*in
   wire signed [9:0] m16_26;
   assign m16_26 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_27 = W*in
   wire signed [9:0] m16_27;
   assign m16_27 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_28 = W*in
   wire signed [9:0] m16_28;
   assign m16_28 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_29 = W*in
   wire signed [9:0] m16_29;
   assign m16_29 ={ {4{in16[5]}} , in16[5:0] };

   // m16_30 = W*in
   wire signed [9:0] m16_30;
   assign m16_30 =10'b0;

   // m16_31 = W*in
   wire signed [9:0] m16_31;
   assign m16_31 =10'b0;

   // m16_32 = W*in
   wire signed [9:0] m16_32;
   assign m16_32 =10'b0;

   // m16_33 = W*in
   wire signed [9:0] m16_33;
   assign m16_33 =10'b0;

   // m16_34 = W*in
   wire signed [9:0] m16_34;
   assign m16_34 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_35 = W*in
   wire signed [9:0] m16_35;
   assign m16_35 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_36 = W*in
   wire signed [9:0] m16_36;
   assign m16_36 =10'b0;

   // m16_37 = W*in
   wire signed [9:0] m16_37;
   assign m16_37 ={ {4{in16[5]}} , in16[5:0] };

   // m16_38 = W*in
   wire signed [9:0] m16_38;
   assign m16_38 =10'b0;

   // m16_39 = W*in
   wire signed [9:0] m16_39;
   assign m16_39 =10'b0;

   // m16_40 = W*in
   wire signed [9:0] m16_40;
   assign m16_40 =10'b0;

   // m16_41 = W*in
   wire signed [9:0] m16_41;
   assign m16_41 =10'b0;

   // m16_42 = W*in
   wire signed [9:0] m16_42;
   assign m16_42 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_43 = W*in
   wire signed [9:0] m16_43;
   assign m16_43 =10'b0;

   // m16_44 = W*in
   wire signed [9:0] m16_44;
   assign m16_44 ={ {4{in16[5]}} , in16[5:0] };

   // m16_45 = W*in
   wire signed [9:0] m16_45;
   assign m16_45 =10'b0;

   // m16_46 = W*in
   wire signed [9:0] m16_46;
   assign m16_46 =10'b0;

   // m16_47 = W*in
   wire signed [9:0] m16_47;
   assign m16_47 =10'b0;

   // m16_48 = W*in
   wire signed [9:0] m16_48;
   assign m16_48 =10'b0;

   // m16_49 = W*in
   wire signed [9:0] m16_49;
   assign m16_49 =10'b0;

   // m16_50 = W*in
   wire signed [9:0] m16_50;
   assign m16_50 =10'b0;

   // m16_51 = W*in
   wire signed [9:0] m16_51;
   assign m16_51 =10'b0;

   // m16_52 = W*in
   wire signed [9:0] m16_52;
   assign m16_52 =10'b0;

   // m16_53 = W*in
   wire signed [9:0] m16_53;
   assign m16_53 =10'b0;

   // m16_54 = W*in
   wire signed [9:0] m16_54;
   assign m16_54 ={ {4{in16[5]}} , in16[5:0] };

   // m16_55 = W*in
   wire signed [9:0] m16_55;
   assign m16_55 =10'b0;

   // m16_56 = W*in
   wire signed [9:0] m16_56;
   assign m16_56 =10'b0;

   // m16_57 = W*in
   wire signed [9:0] m16_57;
   assign m16_57 =10'b0;

   // m16_58 = W*in
   wire signed [9:0] m16_58;
   assign m16_58 =10'b0;

   // m16_59 = W*in
   wire signed [9:0] m16_59;
   assign m16_59 =10'b0;

   // m16_60 = W*in
   wire signed [9:0] m16_60;
   assign m16_60 =10'b0;

   // m16_61 = W*in
   wire signed [9:0] m16_61;
   assign m16_61 =10'b0;

   // m16_62 = W*in
   wire signed [9:0] m16_62;
   assign m16_62 =10'b0;

   // m16_63 = W*in
   wire signed [9:0] m16_63;
   assign m16_63 ={ {4{in16[5]}} , in16[5:0] };

   // m16_64 = W*in
   wire signed [9:0] m16_64;
   assign m16_64 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_65 = W*in
   wire signed [9:0] m16_65;
   assign m16_65 ={ {5{in16[5]}} , in16[5:1] };

   // m16_66 = W*in
   wire signed [9:0] m16_66;
   assign m16_66 =10'b0;

   // m16_67 = W*in
   wire signed [9:0] m16_67;
   assign m16_67 ={ {4{in16[5]}} , in16[5:0] };

   // m16_68 = W*in
   wire signed [9:0] m16_68;
   assign m16_68 =10'b0;

   // m16_69 = W*in
   wire signed [9:0] m16_69;
   assign m16_69 ={ {4{in16[5]}} , in16[5:0] };

   // m16_70 = W*in
   wire signed [9:0] m16_70;
   assign m16_70 ={ {4{in16[5]}} , in16[5:0] };

   // m16_71 = W*in
   wire signed [9:0] m16_71;
   assign m16_71 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_72 = W*in
   wire signed [9:0] m16_72;
   assign m16_72 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_73 = W*in
   wire signed [9:0] m16_73;
   assign m16_73 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_74 = W*in
   wire signed [9:0] m16_74;
   assign m16_74 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_75 = W*in
   wire signed [9:0] m16_75;
   assign m16_75 ={ {5{neg16[5]}} , neg16[5:1] };

   // m16_76 = W*in
   wire signed [9:0] m16_76;
   assign m16_76 =10'b0;

   // m16_77 = W*in
   wire signed [9:0] m16_77;
   assign m16_77 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_78 = W*in
   wire signed [9:0] m16_78;
   assign m16_78 =10'b0;

   // m16_79 = W*in
   wire signed [9:0] m16_79;
   assign m16_79 ={ {4{in16[5]}} , in16[5:0] };

   // m16_80 = W*in
   wire signed [9:0] m16_80;
   assign m16_80 =10'b0;

   // m16_81 = W*in
   wire signed [9:0] m16_81;
   assign m16_81 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_82 = W*in
   wire signed [9:0] m16_82;
   assign m16_82 =10'b0;

   // m16_83 = W*in
   wire signed [9:0] m16_83;
   assign m16_83 =10'b0;

   // m16_84 = W*in
   wire signed [9:0] m16_84;
   assign m16_84 =10'b0;

   // m16_85 = W*in
   wire signed [9:0] m16_85;
   assign m16_85 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_86 = W*in
   wire signed [9:0] m16_86;
   assign m16_86 =10'b0;

   // m16_87 = W*in
   wire signed [9:0] m16_87;
   assign m16_87 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_88 = W*in
   wire signed [9:0] m16_88;
   assign m16_88 =10'b0;

   // m16_89 = W*in
   wire signed [9:0] m16_89;
   assign m16_89 =10'b0;

   // m16_90 = W*in
   wire signed [9:0] m16_90;
   assign m16_90 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_91 = W*in
   wire signed [9:0] m16_91;
   assign m16_91 =10'b0;

   // m16_92 = W*in
   wire signed [9:0] m16_92;
   assign m16_92 =10'b0;

   // m16_93 = W*in
   wire signed [9:0] m16_93;
   assign m16_93 ={ {3{in16[5]}} , in16 , {1{1'b0}} };

   // m16_94 = W*in
   wire signed [9:0] m16_94;
   assign m16_94 =10'b0;

   // m16_95 = W*in
   wire signed [9:0] m16_95;
   assign m16_95 ={ {4{in16[5]}} , in16[5:0] };

   // m16_96 = W*in
   wire signed [9:0] m16_96;
   assign m16_96 ={ {4{in16[5]}} , in16[5:0] };

   // m16_97 = W*in
   wire signed [9:0] m16_97;
   assign m16_97 =10'b0;

   // m16_98 = W*in
   wire signed [9:0] m16_98;
   assign m16_98 =10'b0;

   // m16_99 = W*in
   wire signed [9:0] m16_99;
   assign m16_99 =10'b0;

   // m16_100 = W*in
   wire signed [9:0] m16_100;
   assign m16_100 ={ {4{neg16[5]}} , neg16[5:0] };

   // m16_101 = W*in
   wire signed [9:0] m16_101;
   assign m16_101 =10'b0;

   // m16_102 = W*in
   wire signed [9:0] m16_102;
   assign m16_102 =10'b0;

   // m16_103 = W*in
   wire signed [9:0] m16_103;
   assign m16_103 =10'b0;

   // m16_104 = W*in
   wire signed [9:0] m16_104;
   assign m16_104 =10'b0;

   // m16_105 = W*in
   wire signed [9:0] m16_105;
   assign m16_105 =10'b0;

   // m16_106 = W*in
   wire signed [9:0] m16_106;
   assign m16_106 =10'b0;

   // m16_107 = W*in
   wire signed [9:0] m16_107;
   assign m16_107 =10'b0;

   // m16_108 = W*in
   wire signed [9:0] m16_108;
   assign m16_108 ={ {5{in16[5]}} , in16[5:1] };

   // m16_109 = W*in
   wire signed [9:0] m16_109;
   assign m16_109 =10'b0;

   // m16_110 = W*in
   wire signed [9:0] m16_110;
   assign m16_110 =10'b0;

   // m16_111 = W*in
   wire signed [9:0] m16_111;
   assign m16_111 =10'b0;

   // m16_112 = W*in
   wire signed [9:0] m16_112;
   assign m16_112 =10'b0;

   // m16_113 = W*in
   wire signed [9:0] m16_113;
   assign m16_113 =10'b0;

   // m16_114 = W*in
   wire signed [9:0] m16_114;
   assign m16_114 =10'b0;

   // m16_115 = W*in
   wire signed [9:0] m16_115;
   assign m16_115 =10'b0;

   // m16_116 = W*in
   wire signed [9:0] m16_116;
   assign m16_116 ={ {4{in16[5]}} , in16[5:0] };

   // m16_117 = W*in
   wire signed [9:0] m16_117;
   assign m16_117 ={ {4{neg16[5]}} , neg16[5:0] };

   // m17_1 = W*in
   wire signed [9:0] m17_1;
   assign m17_1 =10'b0;

   // m17_2 = W*in
   wire signed [9:0] m17_2;
   assign m17_2 =10'b0;

   // m17_3 = W*in
   wire signed [9:0] m17_3;
   assign m17_3 =10'b0;

   // m17_4 = W*in
   wire signed [9:0] m17_4;
   assign m17_4 =10'b0;

   // m17_5 = W*in
   wire signed [9:0] m17_5;
   assign m17_5 =10'b0;

   // m17_6 = W*in
   wire signed [9:0] m17_6;
   assign m17_6 =10'b0;

   // m17_7 = W*in
   wire signed [9:0] m17_7;
   assign m17_7 =10'b0;

   // m17_8 = W*in
   wire signed [9:0] m17_8;
   assign m17_8 =10'b0;

   // m17_9 = W*in
   wire signed [9:0] m17_9;
   assign m17_9 =10'b0;

   // m17_10 = W*in
   wire signed [9:0] m17_10;
   assign m17_10 =10'b0;

   // m17_11 = W*in
   wire signed [9:0] m17_11;
   assign m17_11 =10'b0;

   // m17_12 = W*in
   wire signed [9:0] m17_12;
   assign m17_12 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_13 = W*in
   wire signed [9:0] m17_13;
   assign m17_13 =10'b0;

   // m17_14 = W*in
   wire signed [9:0] m17_14;
   assign m17_14 =10'b0;

   // m17_15 = W*in
   wire signed [9:0] m17_15;
   assign m17_15 =10'b0;

   // m17_16 = W*in
   wire signed [9:0] m17_16;
   assign m17_16 =10'b0;

   // m17_17 = W*in
   wire signed [9:0] m17_17;
   assign m17_17 ={ {4{in17[5]}} , in17[5:0] };

   // m17_18 = W*in
   wire signed [9:0] m17_18;
   assign m17_18 ={ {5{neg17[5]}} , neg17[5:1] };

   // m17_19 = W*in
   wire signed [9:0] m17_19;
   assign m17_19 =10'b0;

   // m17_20 = W*in
   wire signed [9:0] m17_20;
   assign m17_20 =10'b0;

   // m17_21 = W*in
   wire signed [9:0] m17_21;
   assign m17_21 =10'b0;

   // m17_22 = W*in
   wire signed [9:0] m17_22;
   assign m17_22 =10'b0;

   // m17_23 = W*in
   wire signed [9:0] m17_23;
   assign m17_23 =10'b0;

   // m17_24 = W*in
   wire signed [9:0] m17_24;
   assign m17_24 =10'b0;

   // m17_25 = W*in
   wire signed [9:0] m17_25;
   assign m17_25 =10'b0;

   // m17_26 = W*in
   wire signed [9:0] m17_26;
   assign m17_26 ={ {5{neg17[5]}} , neg17[5:1] };

   // m17_27 = W*in
   wire signed [9:0] m17_27;
   assign m17_27 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_28 = W*in
   wire signed [9:0] m17_28;
   assign m17_28 =10'b0;

   // m17_29 = W*in
   wire signed [9:0] m17_29;
   assign m17_29 =10'b0;

   // m17_30 = W*in
   wire signed [9:0] m17_30;
   assign m17_30 =10'b0;

   // m17_31 = W*in
   wire signed [9:0] m17_31;
   assign m17_31 ={ {5{neg17[5]}} , neg17[5:1] };

   // m17_32 = W*in
   wire signed [9:0] m17_32;
   assign m17_32 ={ {5{in17[5]}} , in17[5:1] };

   // m17_33 = W*in
   wire signed [9:0] m17_33;
   assign m17_33 =10'b0;

   // m17_34 = W*in
   wire signed [9:0] m17_34;
   assign m17_34 =10'b0;

   // m17_35 = W*in
   wire signed [9:0] m17_35;
   assign m17_35 =10'b0;

   // m17_36 = W*in
   wire signed [9:0] m17_36;
   assign m17_36 ={ {5{in17[5]}} , in17[5:1] };

   // m17_37 = W*in
   wire signed [9:0] m17_37;
   assign m17_37 ={ {4{in17[5]}} , in17[5:0] };

   // m17_38 = W*in
   wire signed [9:0] m17_38;
   assign m17_38 =10'b0;

   // m17_39 = W*in
   wire signed [9:0] m17_39;
   assign m17_39 =10'b0;

   // m17_40 = W*in
   wire signed [9:0] m17_40;
   assign m17_40 =10'b0;

   // m17_41 = W*in
   wire signed [9:0] m17_41;
   assign m17_41 =10'b0;

   // m17_42 = W*in
   wire signed [9:0] m17_42;
   assign m17_42 =10'b0;

   // m17_43 = W*in
   wire signed [9:0] m17_43;
   assign m17_43 =10'b0;

   // m17_44 = W*in
   wire signed [9:0] m17_44;
   assign m17_44 =10'b0;

   // m17_45 = W*in
   wire signed [9:0] m17_45;
   assign m17_45 ={ {4{in17[5]}} , in17[5:0] };

   // m17_46 = W*in
   wire signed [9:0] m17_46;
   assign m17_46 =10'b0;

   // m17_47 = W*in
   wire signed [9:0] m17_47;
   assign m17_47 ={ {4{in17[5]}} , in17[5:0] };

   // m17_48 = W*in
   wire signed [9:0] m17_48;
   assign m17_48 =10'b0;

   // m17_49 = W*in
   wire signed [9:0] m17_49;
   assign m17_49 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_50 = W*in
   wire signed [9:0] m17_50;
   assign m17_50 =10'b0;

   // m17_51 = W*in
   wire signed [9:0] m17_51;
   assign m17_51 ={ {4{in17[5]}} , in17[5:0] };

   // m17_52 = W*in
   wire signed [9:0] m17_52;
   assign m17_52 =10'b0;

   // m17_53 = W*in
   wire signed [9:0] m17_53;
   assign m17_53 =10'b0;

   // m17_54 = W*in
   wire signed [9:0] m17_54;
   assign m17_54 =10'b0;

   // m17_55 = W*in
   wire signed [9:0] m17_55;
   assign m17_55 =10'b0;

   // m17_56 = W*in
   wire signed [9:0] m17_56;
   assign m17_56 =10'b0;

   // m17_57 = W*in
   wire signed [9:0] m17_57;
   assign m17_57 ={ {4{in17[5]}} , in17[5:0] };

   // m17_58 = W*in
   wire signed [9:0] m17_58;
   assign m17_58 =10'b0;

   // m17_59 = W*in
   wire signed [9:0] m17_59;
   assign m17_59 =10'b0;

   // m17_60 = W*in
   wire signed [9:0] m17_60;
   assign m17_60 =10'b0;

   // m17_61 = W*in
   wire signed [9:0] m17_61;
   assign m17_61 =10'b0;

   // m17_62 = W*in
   wire signed [9:0] m17_62;
   assign m17_62 =10'b0;

   // m17_63 = W*in
   wire signed [9:0] m17_63;
   assign m17_63 ={ {4{in17[5]}} , in17[5:0] };

   // m17_64 = W*in
   wire signed [9:0] m17_64;
   assign m17_64 =10'b0;

   // m17_65 = W*in
   wire signed [9:0] m17_65;
   assign m17_65 =10'b0;

   // m17_66 = W*in
   wire signed [9:0] m17_66;
   assign m17_66 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_67 = W*in
   wire signed [9:0] m17_67;
   assign m17_67 ={ {4{in17[5]}} , in17[5:0] };

   // m17_68 = W*in
   wire signed [9:0] m17_68;
   assign m17_68 =10'b0;

   // m17_69 = W*in
   wire signed [9:0] m17_69;
   assign m17_69 =10'b0;

   // m17_70 = W*in
   wire signed [9:0] m17_70;
   assign m17_70 =10'b0;

   // m17_71 = W*in
   wire signed [9:0] m17_71;
   assign m17_71 ={ {5{neg17[5]}} , neg17[5:1] };

   // m17_72 = W*in
   wire signed [9:0] m17_72;
   assign m17_72 =10'b0;

   // m17_73 = W*in
   wire signed [9:0] m17_73;
   assign m17_73 =10'b0;

   // m17_74 = W*in
   wire signed [9:0] m17_74;
   assign m17_74 =10'b0;

   // m17_75 = W*in
   wire signed [9:0] m17_75;
   assign m17_75 =10'b0;

   // m17_76 = W*in
   wire signed [9:0] m17_76;
   assign m17_76 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_77 = W*in
   wire signed [9:0] m17_77;
   assign m17_77 =10'b0;

   // m17_78 = W*in
   wire signed [9:0] m17_78;
   assign m17_78 =10'b0;

   // m17_79 = W*in
   wire signed [9:0] m17_79;
   assign m17_79 =10'b0;

   // m17_80 = W*in
   wire signed [9:0] m17_80;
   assign m17_80 =10'b0;

   // m17_81 = W*in
   wire signed [9:0] m17_81;
   assign m17_81 ={ {5{neg17[5]}} , neg17[5:1] };

   // m17_82 = W*in
   wire signed [9:0] m17_82;
   assign m17_82 =10'b0;

   // m17_83 = W*in
   wire signed [9:0] m17_83;
   assign m17_83 =10'b0;

   // m17_84 = W*in
   wire signed [9:0] m17_84;
   assign m17_84 =10'b0;

   // m17_85 = W*in
   wire signed [9:0] m17_85;
   assign m17_85 =10'b0;

   // m17_86 = W*in
   wire signed [9:0] m17_86;
   assign m17_86 =10'b0;

   // m17_87 = W*in
   wire signed [9:0] m17_87;
   assign m17_87 =10'b0;

   // m17_88 = W*in
   wire signed [9:0] m17_88;
   assign m17_88 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_89 = W*in
   wire signed [9:0] m17_89;
   assign m17_89 =10'b0;

   // m17_90 = W*in
   wire signed [9:0] m17_90;
   assign m17_90 =10'b0;

   // m17_91 = W*in
   wire signed [9:0] m17_91;
   assign m17_91 =10'b0;

   // m17_92 = W*in
   wire signed [9:0] m17_92;
   assign m17_92 =10'b0;

   // m17_93 = W*in
   wire signed [9:0] m17_93;
   assign m17_93 =10'b0;

   // m17_94 = W*in
   wire signed [9:0] m17_94;
   assign m17_94 =10'b0;

   // m17_95 = W*in
   wire signed [9:0] m17_95;
   assign m17_95 =10'b0;

   // m17_96 = W*in
   wire signed [9:0] m17_96;
   assign m17_96 =10'b0;

   // m17_97 = W*in
   wire signed [9:0] m17_97;
   assign m17_97 =10'b0;

   // m17_98 = W*in
   wire signed [9:0] m17_98;
   assign m17_98 =10'b0;

   // m17_99 = W*in
   wire signed [9:0] m17_99;
   assign m17_99 =10'b0;

   // m17_100 = W*in
   wire signed [9:0] m17_100;
   assign m17_100 ={ {4{neg17[5]}} , neg17[5:0] };

   // m17_101 = W*in
   wire signed [9:0] m17_101;
   assign m17_101 =10'b0;

   // m17_102 = W*in
   wire signed [9:0] m17_102;
   assign m17_102 =10'b0;

   // m17_103 = W*in
   wire signed [9:0] m17_103;
   assign m17_103 =10'b0;

   // m17_104 = W*in
   wire signed [9:0] m17_104;
   assign m17_104 =10'b0;

   // m17_105 = W*in
   wire signed [9:0] m17_105;
   assign m17_105 =10'b0;

   // m17_106 = W*in
   wire signed [9:0] m17_106;
   assign m17_106 =10'b0;

   // m17_107 = W*in
   wire signed [9:0] m17_107;
   assign m17_107 =10'b0;

   // m17_108 = W*in
   wire signed [9:0] m17_108;
   assign m17_108 =10'b0;

   // m17_109 = W*in
   wire signed [9:0] m17_109;
   assign m17_109 =10'b0;

   // m17_110 = W*in
   wire signed [9:0] m17_110;
   assign m17_110 =10'b0;

   // m17_111 = W*in
   wire signed [9:0] m17_111;
   assign m17_111 =10'b0;

   // m17_112 = W*in
   wire signed [9:0] m17_112;
   assign m17_112 =10'b0;

   // m17_113 = W*in
   wire signed [9:0] m17_113;
   assign m17_113 =10'b0;

   // m17_114 = W*in
   wire signed [9:0] m17_114;
   assign m17_114 =10'b0;

   // m17_115 = W*in
   wire signed [9:0] m17_115;
   assign m17_115 ={ {4{in17[5]}} , in17[5:0] };

   // m17_116 = W*in
   wire signed [9:0] m17_116;
   assign m17_116 =10'b0;

   // m17_117 = W*in
   wire signed [9:0] m17_117;
   assign m17_117 =10'b0;

   // m18_1 = W*in
   wire signed [9:0] m18_1;
   assign m18_1 =10'b0;

   // m18_2 = W*in
   wire signed [9:0] m18_2;
   assign m18_2 =10'b0;

   // m18_3 = W*in
   wire signed [9:0] m18_3;
   assign m18_3 ={ {4{in18[5]}} , in18[5:0] };

   // m18_4 = W*in
   wire signed [9:0] m18_4;
   assign m18_4 =10'b0;

   // m18_5 = W*in
   wire signed [9:0] m18_5;
   assign m18_5 =10'b0;

   // m18_6 = W*in
   wire signed [9:0] m18_6;
   assign m18_6 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_7 = W*in
   wire signed [9:0] m18_7;
   assign m18_7 =10'b0;

   // m18_8 = W*in
   wire signed [9:0] m18_8;
   assign m18_8 =10'b0;

   // m18_9 = W*in
   wire signed [9:0] m18_9;
   assign m18_9 =10'b0;

   // m18_10 = W*in
   wire signed [9:0] m18_10;
   assign m18_10 =10'b0;

   // m18_11 = W*in
   wire signed [9:0] m18_11;
   assign m18_11 =10'b0;

   // m18_12 = W*in
   wire signed [9:0] m18_12;
   assign m18_12 ={ {5{neg18[5]}} , neg18[5:1] };

   // m18_13 = W*in
   wire signed [9:0] m18_13;
   assign m18_13 ={ {4{in18[5]}} , in18[5:0] };

   // m18_14 = W*in
   wire signed [9:0] m18_14;
   assign m18_14 =10'b0;

   // m18_15 = W*in
   wire signed [9:0] m18_15;
   assign m18_15 =10'b0;

   // m18_16 = W*in
   wire signed [9:0] m18_16;
   assign m18_16 =10'b0;

   // m18_17 = W*in
   wire signed [9:0] m18_17;
   assign m18_17 =10'b0;

   // m18_18 = W*in
   wire signed [9:0] m18_18;
   assign m18_18 =10'b0;

   // m18_19 = W*in
   wire signed [9:0] m18_19;
   assign m18_19 =10'b0;

   // m18_20 = W*in
   wire signed [9:0] m18_20;
   assign m18_20 =10'b0;

   // m18_21 = W*in
   wire signed [9:0] m18_21;
   assign m18_21 =10'b0;

   // m18_22 = W*in
   wire signed [9:0] m18_22;
   assign m18_22 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_23 = W*in
   wire signed [9:0] m18_23;
   assign m18_23 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_24 = W*in
   wire signed [9:0] m18_24;
   assign m18_24 =10'b0;

   // m18_25 = W*in
   wire signed [9:0] m18_25;
   assign m18_25 =10'b0;

   // m18_26 = W*in
   wire signed [9:0] m18_26;
   assign m18_26 =10'b0;

   // m18_27 = W*in
   wire signed [9:0] m18_27;
   assign m18_27 =10'b0;

   // m18_28 = W*in
   wire signed [9:0] m18_28;
   assign m18_28 =10'b0;

   // m18_29 = W*in
   wire signed [9:0] m18_29;
   assign m18_29 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_30 = W*in
   wire signed [9:0] m18_30;
   assign m18_30 =10'b0;

   // m18_31 = W*in
   wire signed [9:0] m18_31;
   assign m18_31 ={ {5{neg18[5]}} , neg18[5:1] };

   // m18_32 = W*in
   wire signed [9:0] m18_32;
   assign m18_32 =10'b0;

   // m18_33 = W*in
   wire signed [9:0] m18_33;
   assign m18_33 =10'b0;

   // m18_34 = W*in
   wire signed [9:0] m18_34;
   assign m18_34 =10'b0;

   // m18_35 = W*in
   wire signed [9:0] m18_35;
   assign m18_35 ={ {5{in18[5]}} , in18[5:1] };

   // m18_36 = W*in
   wire signed [9:0] m18_36;
   assign m18_36 ={ {5{in18[5]}} , in18[5:1] };

   // m18_37 = W*in
   wire signed [9:0] m18_37;
   assign m18_37 =10'b0;

   // m18_38 = W*in
   wire signed [9:0] m18_38;
   assign m18_38 =10'b0;

   // m18_39 = W*in
   wire signed [9:0] m18_39;
   assign m18_39 =10'b0;

   // m18_40 = W*in
   wire signed [9:0] m18_40;
   assign m18_40 =10'b0;

   // m18_41 = W*in
   wire signed [9:0] m18_41;
   assign m18_41 =10'b0;

   // m18_42 = W*in
   wire signed [9:0] m18_42;
   assign m18_42 =10'b0;

   // m18_43 = W*in
   wire signed [9:0] m18_43;
   assign m18_43 =10'b0;

   // m18_44 = W*in
   wire signed [9:0] m18_44;
   assign m18_44 =10'b0;

   // m18_45 = W*in
   wire signed [9:0] m18_45;
   assign m18_45 =10'b0;

   // m18_46 = W*in
   wire signed [9:0] m18_46;
   assign m18_46 ={ {4{in18[5]}} , in18[5:0] };

   // m18_47 = W*in
   wire signed [9:0] m18_47;
   assign m18_47 =10'b0;

   // m18_48 = W*in
   wire signed [9:0] m18_48;
   assign m18_48 =10'b0;

   // m18_49 = W*in
   wire signed [9:0] m18_49;
   assign m18_49 =10'b0;

   // m18_50 = W*in
   wire signed [9:0] m18_50;
   assign m18_50 =10'b0;

   // m18_51 = W*in
   wire signed [9:0] m18_51;
   assign m18_51 =10'b0;

   // m18_52 = W*in
   wire signed [9:0] m18_52;
   assign m18_52 =10'b0;

   // m18_53 = W*in
   wire signed [9:0] m18_53;
   assign m18_53 =10'b0;

   // m18_54 = W*in
   wire signed [9:0] m18_54;
   assign m18_54 =10'b0;

   // m18_55 = W*in
   wire signed [9:0] m18_55;
   assign m18_55 =10'b0;

   // m18_56 = W*in
   wire signed [9:0] m18_56;
   assign m18_56 ={ {5{neg18[5]}} , neg18[5:1] };

   // m18_57 = W*in
   wire signed [9:0] m18_57;
   assign m18_57 ={ {4{in18[5]}} , in18[5:0] };

   // m18_58 = W*in
   wire signed [9:0] m18_58;
   assign m18_58 =10'b0;

   // m18_59 = W*in
   wire signed [9:0] m18_59;
   assign m18_59 =10'b0;

   // m18_60 = W*in
   wire signed [9:0] m18_60;
   assign m18_60 ={ {4{in18[5]}} , in18[5:0] };

   // m18_61 = W*in
   wire signed [9:0] m18_61;
   assign m18_61 =10'b0;

   // m18_62 = W*in
   wire signed [9:0] m18_62;
   assign m18_62 =10'b0;

   // m18_63 = W*in
   wire signed [9:0] m18_63;
   assign m18_63 =10'b0;

   // m18_64 = W*in
   wire signed [9:0] m18_64;
   assign m18_64 =10'b0;

   // m18_65 = W*in
   wire signed [9:0] m18_65;
   assign m18_65 ={ {4{in18[5]}} , in18[5:0] };

   // m18_66 = W*in
   wire signed [9:0] m18_66;
   assign m18_66 ={ {4{in18[5]}} , in18[5:0] };

   // m18_67 = W*in
   wire signed [9:0] m18_67;
   assign m18_67 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_68 = W*in
   wire signed [9:0] m18_68;
   assign m18_68 =10'b0;

   // m18_69 = W*in
   wire signed [9:0] m18_69;
   assign m18_69 =10'b0;

   // m18_70 = W*in
   wire signed [9:0] m18_70;
   assign m18_70 =10'b0;

   // m18_71 = W*in
   wire signed [9:0] m18_71;
   assign m18_71 =10'b0;

   // m18_72 = W*in
   wire signed [9:0] m18_72;
   assign m18_72 =10'b0;

   // m18_73 = W*in
   wire signed [9:0] m18_73;
   assign m18_73 =10'b0;

   // m18_74 = W*in
   wire signed [9:0] m18_74;
   assign m18_74 =10'b0;

   // m18_75 = W*in
   wire signed [9:0] m18_75;
   assign m18_75 =10'b0;

   // m18_76 = W*in
   wire signed [9:0] m18_76;
   assign m18_76 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_77 = W*in
   wire signed [9:0] m18_77;
   assign m18_77 =10'b0;

   // m18_78 = W*in
   wire signed [9:0] m18_78;
   assign m18_78 =10'b0;

   // m18_79 = W*in
   wire signed [9:0] m18_79;
   assign m18_79 =10'b0;

   // m18_80 = W*in
   wire signed [9:0] m18_80;
   assign m18_80 =10'b0;

   // m18_81 = W*in
   wire signed [9:0] m18_81;
   assign m18_81 ={ {5{neg18[5]}} , neg18[5:1] };

   // m18_82 = W*in
   wire signed [9:0] m18_82;
   assign m18_82 =10'b0;

   // m18_83 = W*in
   wire signed [9:0] m18_83;
   assign m18_83 =10'b0;

   // m18_84 = W*in
   wire signed [9:0] m18_84;
   assign m18_84 =10'b0;

   // m18_85 = W*in
   wire signed [9:0] m18_85;
   assign m18_85 =10'b0;

   // m18_86 = W*in
   wire signed [9:0] m18_86;
   assign m18_86 =10'b0;

   // m18_87 = W*in
   wire signed [9:0] m18_87;
   assign m18_87 =10'b0;

   // m18_88 = W*in
   wire signed [9:0] m18_88;
   assign m18_88 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_89 = W*in
   wire signed [9:0] m18_89;
   assign m18_89 =10'b0;

   // m18_90 = W*in
   wire signed [9:0] m18_90;
   assign m18_90 =10'b0;

   // m18_91 = W*in
   wire signed [9:0] m18_91;
   assign m18_91 ={ {5{in18[5]}} , in18[5:1] };

   // m18_92 = W*in
   wire signed [9:0] m18_92;
   assign m18_92 =10'b0;

   // m18_93 = W*in
   wire signed [9:0] m18_93;
   assign m18_93 =10'b0;

   // m18_94 = W*in
   wire signed [9:0] m18_94;
   assign m18_94 ={ {4{in18[5]}} , in18[5:0] };

   // m18_95 = W*in
   wire signed [9:0] m18_95;
   assign m18_95 =10'b0;

   // m18_96 = W*in
   wire signed [9:0] m18_96;
   assign m18_96 =10'b0;

   // m18_97 = W*in
   wire signed [9:0] m18_97;
   assign m18_97 ={ {5{in18[5]}} , in18[5:1] };

   // m18_98 = W*in
   wire signed [9:0] m18_98;
   assign m18_98 ={ {4{neg18[5]}} , neg18[5:0] };

   // m18_99 = W*in
   wire signed [9:0] m18_99;
   assign m18_99 =10'b0;

   // m18_100 = W*in
   wire signed [9:0] m18_100;
   assign m18_100 =10'b0;

   // m18_101 = W*in
   wire signed [9:0] m18_101;
   assign m18_101 =10'b0;

   // m18_102 = W*in
   wire signed [9:0] m18_102;
   assign m18_102 =10'b0;

   // m18_103 = W*in
   wire signed [9:0] m18_103;
   assign m18_103 =10'b0;

   // m18_104 = W*in
   wire signed [9:0] m18_104;
   assign m18_104 ={ {4{in18[5]}} , in18[5:0] };

   // m18_105 = W*in
   wire signed [9:0] m18_105;
   assign m18_105 =10'b0;

   // m18_106 = W*in
   wire signed [9:0] m18_106;
   assign m18_106 ={ {4{in18[5]}} , in18[5:0] };

   // m18_107 = W*in
   wire signed [9:0] m18_107;
   assign m18_107 =10'b0;

   // m18_108 = W*in
   wire signed [9:0] m18_108;
   assign m18_108 =10'b0;

   // m18_109 = W*in
   wire signed [9:0] m18_109;
   assign m18_109 =10'b0;

   // m18_110 = W*in
   wire signed [9:0] m18_110;
   assign m18_110 =10'b0;

   // m18_111 = W*in
   wire signed [9:0] m18_111;
   assign m18_111 =10'b0;

   // m18_112 = W*in
   wire signed [9:0] m18_112;
   assign m18_112 ={ {4{in18[5]}} , in18[5:0] };

   // m18_113 = W*in
   wire signed [9:0] m18_113;
   assign m18_113 =10'b0;

   // m18_114 = W*in
   wire signed [9:0] m18_114;
   assign m18_114 =10'b0;

   // m18_115 = W*in
   wire signed [9:0] m18_115;
   assign m18_115 =10'b0;

   // m18_116 = W*in
   wire signed [9:0] m18_116;
   assign m18_116 =10'b0;

   // m18_117 = W*in
   wire signed [9:0] m18_117;
   assign m18_117 =10'b0;

   // m19_1 = W*in
   wire signed [9:0] m19_1;
   assign m19_1 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_2 = W*in
   wire signed [9:0] m19_2;
   assign m19_2 =10'b0;

   // m19_3 = W*in
   wire signed [9:0] m19_3;
   assign m19_3 =10'b0;

   // m19_4 = W*in
   wire signed [9:0] m19_4;
   assign m19_4 =10'b0;

   // m19_5 = W*in
   wire signed [9:0] m19_5;
   assign m19_5 =10'b0;

   // m19_6 = W*in
   wire signed [9:0] m19_6;
   assign m19_6 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_7 = W*in
   wire signed [9:0] m19_7;
   assign m19_7 =10'b0;

   // m19_8 = W*in
   wire signed [9:0] m19_8;
   assign m19_8 =10'b0;

   // m19_9 = W*in
   wire signed [9:0] m19_9;
   assign m19_9 =10'b0;

   // m19_10 = W*in
   wire signed [9:0] m19_10;
   assign m19_10 =10'b0;

   // m19_11 = W*in
   wire signed [9:0] m19_11;
   assign m19_11 ={ {5{in19[5]}} , in19[5:1] };

   // m19_12 = W*in
   wire signed [9:0] m19_12;
   assign m19_12 =10'b0;

   // m19_13 = W*in
   wire signed [9:0] m19_13;
   assign m19_13 =10'b0;

   // m19_14 = W*in
   wire signed [9:0] m19_14;
   assign m19_14 =10'b0;

   // m19_15 = W*in
   wire signed [9:0] m19_15;
   assign m19_15 =10'b0;

   // m19_16 = W*in
   wire signed [9:0] m19_16;
   assign m19_16 =10'b0;

   // m19_17 = W*in
   wire signed [9:0] m19_17;
   assign m19_17 =10'b0;

   // m19_18 = W*in
   wire signed [9:0] m19_18;
   assign m19_18 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_19 = W*in
   wire signed [9:0] m19_19;
   assign m19_19 =10'b0;

   // m19_20 = W*in
   wire signed [9:0] m19_20;
   assign m19_20 =10'b0;

   // m19_21 = W*in
   wire signed [9:0] m19_21;
   assign m19_21 ={ {5{in19[5]}} , in19[5:1] };

   // m19_22 = W*in
   wire signed [9:0] m19_22;
   assign m19_22 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_23 = W*in
   wire signed [9:0] m19_23;
   assign m19_23 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_24 = W*in
   wire signed [9:0] m19_24;
   assign m19_24 =10'b0;

   // m19_25 = W*in
   wire signed [9:0] m19_25;
   assign m19_25 =10'b0;

   // m19_26 = W*in
   wire signed [9:0] m19_26;
   assign m19_26 =10'b0;

   // m19_27 = W*in
   wire signed [9:0] m19_27;
   assign m19_27 ={ {4{in19[5]}} , in19[5:0] };

   // m19_28 = W*in
   wire signed [9:0] m19_28;
   assign m19_28 ={ {4{in19[5]}} , in19[5:0] };

   // m19_29 = W*in
   wire signed [9:0] m19_29;
   assign m19_29 ={ {5{neg19[5]}} , neg19[5:1] };

   // m19_30 = W*in
   wire signed [9:0] m19_30;
   assign m19_30 ={ {5{in19[5]}} , in19[5:1] };

   // m19_31 = W*in
   wire signed [9:0] m19_31;
   assign m19_31 =10'b0;

   // m19_32 = W*in
   wire signed [9:0] m19_32;
   assign m19_32 =10'b0;

   // m19_33 = W*in
   wire signed [9:0] m19_33;
   assign m19_33 =10'b0;

   // m19_34 = W*in
   wire signed [9:0] m19_34;
   assign m19_34 =10'b0;

   // m19_35 = W*in
   wire signed [9:0] m19_35;
   assign m19_35 =10'b0;

   // m19_36 = W*in
   wire signed [9:0] m19_36;
   assign m19_36 =10'b0;

   // m19_37 = W*in
   wire signed [9:0] m19_37;
   assign m19_37 =10'b0;

   // m19_38 = W*in
   wire signed [9:0] m19_38;
   assign m19_38 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_39 = W*in
   wire signed [9:0] m19_39;
   assign m19_39 =10'b0;

   // m19_40 = W*in
   wire signed [9:0] m19_40;
   assign m19_40 =10'b0;

   // m19_41 = W*in
   wire signed [9:0] m19_41;
   assign m19_41 =10'b0;

   // m19_42 = W*in
   wire signed [9:0] m19_42;
   assign m19_42 =10'b0;

   // m19_43 = W*in
   wire signed [9:0] m19_43;
   assign m19_43 =10'b0;

   // m19_44 = W*in
   wire signed [9:0] m19_44;
   assign m19_44 =10'b0;

   // m19_45 = W*in
   wire signed [9:0] m19_45;
   assign m19_45 =10'b0;

   // m19_46 = W*in
   wire signed [9:0] m19_46;
   assign m19_46 ={ {4{in19[5]}} , in19[5:0] };

   // m19_47 = W*in
   wire signed [9:0] m19_47;
   assign m19_47 =10'b0;

   // m19_48 = W*in
   wire signed [9:0] m19_48;
   assign m19_48 =10'b0;

   // m19_49 = W*in
   wire signed [9:0] m19_49;
   assign m19_49 =10'b0;

   // m19_50 = W*in
   wire signed [9:0] m19_50;
   assign m19_50 =10'b0;

   // m19_51 = W*in
   wire signed [9:0] m19_51;
   assign m19_51 =10'b0;

   // m19_52 = W*in
   wire signed [9:0] m19_52;
   assign m19_52 =10'b0;

   // m19_53 = W*in
   wire signed [9:0] m19_53;
   assign m19_53 =10'b0;

   // m19_54 = W*in
   wire signed [9:0] m19_54;
   assign m19_54 =10'b0;

   // m19_55 = W*in
   wire signed [9:0] m19_55;
   assign m19_55 =10'b0;

   // m19_56 = W*in
   wire signed [9:0] m19_56;
   assign m19_56 =10'b0;

   // m19_57 = W*in
   wire signed [9:0] m19_57;
   assign m19_57 =10'b0;

   // m19_58 = W*in
   wire signed [9:0] m19_58;
   assign m19_58 =10'b0;

   // m19_59 = W*in
   wire signed [9:0] m19_59;
   assign m19_59 =10'b0;

   // m19_60 = W*in
   wire signed [9:0] m19_60;
   assign m19_60 =10'b0;

   // m19_61 = W*in
   wire signed [9:0] m19_61;
   assign m19_61 =10'b0;

   // m19_62 = W*in
   wire signed [9:0] m19_62;
   assign m19_62 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_63 = W*in
   wire signed [9:0] m19_63;
   assign m19_63 =10'b0;

   // m19_64 = W*in
   wire signed [9:0] m19_64;
   assign m19_64 =10'b0;

   // m19_65 = W*in
   wire signed [9:0] m19_65;
   assign m19_65 ={ {4{in19[5]}} , in19[5:0] };

   // m19_66 = W*in
   wire signed [9:0] m19_66;
   assign m19_66 ={ {4{in19[5]}} , in19[5:0] };

   // m19_67 = W*in
   wire signed [9:0] m19_67;
   assign m19_67 =10'b0;

   // m19_68 = W*in
   wire signed [9:0] m19_68;
   assign m19_68 ={ {4{in19[5]}} , in19[5:0] };

   // m19_69 = W*in
   wire signed [9:0] m19_69;
   assign m19_69 =10'b0;

   // m19_70 = W*in
   wire signed [9:0] m19_70;
   assign m19_70 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_71 = W*in
   wire signed [9:0] m19_71;
   assign m19_71 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_72 = W*in
   wire signed [9:0] m19_72;
   assign m19_72 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_73 = W*in
   wire signed [9:0] m19_73;
   assign m19_73 =10'b0;

   // m19_74 = W*in
   wire signed [9:0] m19_74;
   assign m19_74 =10'b0;

   // m19_75 = W*in
   wire signed [9:0] m19_75;
   assign m19_75 =10'b0;

   // m19_76 = W*in
   wire signed [9:0] m19_76;
   assign m19_76 ={ {3{neg19[5]}} , neg19 , {1{1'b0}} };

   // m19_77 = W*in
   wire signed [9:0] m19_77;
   assign m19_77 ={ {4{in19[5]}} , in19[5:0] };

   // m19_78 = W*in
   wire signed [9:0] m19_78;
   assign m19_78 =10'b0;

   // m19_79 = W*in
   wire signed [9:0] m19_79;
   assign m19_79 =10'b0;

   // m19_80 = W*in
   wire signed [9:0] m19_80;
   assign m19_80 =10'b0;

   // m19_81 = W*in
   wire signed [9:0] m19_81;
   assign m19_81 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_82 = W*in
   wire signed [9:0] m19_82;
   assign m19_82 ={ {4{in19[5]}} , in19[5:0] };

   // m19_83 = W*in
   wire signed [9:0] m19_83;
   assign m19_83 =10'b0;

   // m19_84 = W*in
   wire signed [9:0] m19_84;
   assign m19_84 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_85 = W*in
   wire signed [9:0] m19_85;
   assign m19_85 ={ {5{in19[5]}} , in19[5:1] };

   // m19_86 = W*in
   wire signed [9:0] m19_86;
   assign m19_86 =10'b0;

   // m19_87 = W*in
   wire signed [9:0] m19_87;
   assign m19_87 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_88 = W*in
   wire signed [9:0] m19_88;
   assign m19_88 =10'b0;

   // m19_89 = W*in
   wire signed [9:0] m19_89;
   assign m19_89 =10'b0;

   // m19_90 = W*in
   wire signed [9:0] m19_90;
   assign m19_90 =10'b0;

   // m19_91 = W*in
   wire signed [9:0] m19_91;
   assign m19_91 =10'b0;

   // m19_92 = W*in
   wire signed [9:0] m19_92;
   assign m19_92 =10'b0;

   // m19_93 = W*in
   wire signed [9:0] m19_93;
   assign m19_93 =10'b0;

   // m19_94 = W*in
   wire signed [9:0] m19_94;
   assign m19_94 =10'b0;

   // m19_95 = W*in
   wire signed [9:0] m19_95;
   assign m19_95 =10'b0;

   // m19_96 = W*in
   wire signed [9:0] m19_96;
   assign m19_96 =10'b0;

   // m19_97 = W*in
   wire signed [9:0] m19_97;
   assign m19_97 ={ {5{in19[5]}} , in19[5:1] };

   // m19_98 = W*in
   wire signed [9:0] m19_98;
   assign m19_98 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_99 = W*in
   wire signed [9:0] m19_99;
   assign m19_99 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_100 = W*in
   wire signed [9:0] m19_100;
   assign m19_100 =10'b0;

   // m19_101 = W*in
   wire signed [9:0] m19_101;
   assign m19_101 =10'b0;

   // m19_102 = W*in
   wire signed [9:0] m19_102;
   assign m19_102 =10'b0;

   // m19_103 = W*in
   wire signed [9:0] m19_103;
   assign m19_103 =10'b0;

   // m19_104 = W*in
   wire signed [9:0] m19_104;
   assign m19_104 =10'b0;

   // m19_105 = W*in
   wire signed [9:0] m19_105;
   assign m19_105 =10'b0;

   // m19_106 = W*in
   wire signed [9:0] m19_106;
   assign m19_106 =10'b0;

   // m19_107 = W*in
   wire signed [9:0] m19_107;
   assign m19_107 ={ {5{neg19[5]}} , neg19[5:1] };

   // m19_108 = W*in
   wire signed [9:0] m19_108;
   assign m19_108 =10'b0;

   // m19_109 = W*in
   wire signed [9:0] m19_109;
   assign m19_109 =10'b0;

   // m19_110 = W*in
   wire signed [9:0] m19_110;
   assign m19_110 =10'b0;

   // m19_111 = W*in
   wire signed [9:0] m19_111;
   assign m19_111 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_112 = W*in
   wire signed [9:0] m19_112;
   assign m19_112 ={ {4{in19[5]}} , in19[5:0] };

   // m19_113 = W*in
   wire signed [9:0] m19_113;
   assign m19_113 ={ {4{neg19[5]}} , neg19[5:0] };

   // m19_114 = W*in
   wire signed [9:0] m19_114;
   assign m19_114 =10'b0;

   // m19_115 = W*in
   wire signed [9:0] m19_115;
   assign m19_115 ={ {4{in19[5]}} , in19[5:0] };

   // m19_116 = W*in
   wire signed [9:0] m19_116;
   assign m19_116 =10'b0;

   // m19_117 = W*in
   wire signed [9:0] m19_117;
   assign m19_117 ={ {4{in19[5]}} , in19[5:0] };

   // m20_1 = W*in
   wire signed [9:0] m20_1;
   assign m20_1 =10'b0;

   // m20_2 = W*in
   wire signed [9:0] m20_2;
   assign m20_2 =10'b0;

   // m20_3 = W*in
   wire signed [9:0] m20_3;
   assign m20_3 =10'b0;

   // m20_4 = W*in
   wire signed [9:0] m20_4;
   assign m20_4 =10'b0;

   // m20_5 = W*in
   wire signed [9:0] m20_5;
   assign m20_5 =10'b0;

   // m20_6 = W*in
   wire signed [9:0] m20_6;
   assign m20_6 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_7 = W*in
   wire signed [9:0] m20_7;
   assign m20_7 ={ {4{in20[5]}} , in20[5:0] };

   // m20_8 = W*in
   wire signed [9:0] m20_8;
   assign m20_8 =10'b0;

   // m20_9 = W*in
   wire signed [9:0] m20_9;
   assign m20_9 =10'b0;

   // m20_10 = W*in
   wire signed [9:0] m20_10;
   assign m20_10 =10'b0;

   // m20_11 = W*in
   wire signed [9:0] m20_11;
   assign m20_11 ={ {4{in20[5]}} , in20[5:0] };

   // m20_12 = W*in
   wire signed [9:0] m20_12;
   assign m20_12 =10'b0;

   // m20_13 = W*in
   wire signed [9:0] m20_13;
   assign m20_13 =10'b0;

   // m20_14 = W*in
   wire signed [9:0] m20_14;
   assign m20_14 =10'b0;

   // m20_15 = W*in
   wire signed [9:0] m20_15;
   assign m20_15 =10'b0;

   // m20_16 = W*in
   wire signed [9:0] m20_16;
   assign m20_16 =10'b0;

   // m20_17 = W*in
   wire signed [9:0] m20_17;
   assign m20_17 ={ {5{in20[5]}} , in20[5:1] };

   // m20_18 = W*in
   wire signed [9:0] m20_18;
   assign m20_18 =10'b0;

   // m20_19 = W*in
   wire signed [9:0] m20_19;
   assign m20_19 ={ {5{neg20[5]}} , neg20[5:1] };

   // m20_20 = W*in
   wire signed [9:0] m20_20;
   assign m20_20 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_21 = W*in
   wire signed [9:0] m20_21;
   assign m20_21 =10'b0;

   // m20_22 = W*in
   wire signed [9:0] m20_22;
   assign m20_22 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_23 = W*in
   wire signed [9:0] m20_23;
   assign m20_23 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_24 = W*in
   wire signed [9:0] m20_24;
   assign m20_24 =10'b0;

   // m20_25 = W*in
   wire signed [9:0] m20_25;
   assign m20_25 =10'b0;

   // m20_26 = W*in
   wire signed [9:0] m20_26;
   assign m20_26 =10'b0;

   // m20_27 = W*in
   wire signed [9:0] m20_27;
   assign m20_27 ={ {4{in20[5]}} , in20[5:0] };

   // m20_28 = W*in
   wire signed [9:0] m20_28;
   assign m20_28 ={ {4{in20[5]}} , in20[5:0] };

   // m20_29 = W*in
   wire signed [9:0] m20_29;
   assign m20_29 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_30 = W*in
   wire signed [9:0] m20_30;
   assign m20_30 =10'b0;

   // m20_31 = W*in
   wire signed [9:0] m20_31;
   assign m20_31 =10'b0;

   // m20_32 = W*in
   wire signed [9:0] m20_32;
   assign m20_32 =10'b0;

   // m20_33 = W*in
   wire signed [9:0] m20_33;
   assign m20_33 =10'b0;

   // m20_34 = W*in
   wire signed [9:0] m20_34;
   assign m20_34 =10'b0;

   // m20_35 = W*in
   wire signed [9:0] m20_35;
   assign m20_35 =10'b0;

   // m20_36 = W*in
   wire signed [9:0] m20_36;
   assign m20_36 =10'b0;

   // m20_37 = W*in
   wire signed [9:0] m20_37;
   assign m20_37 ={ {4{in20[5]}} , in20[5:0] };

   // m20_38 = W*in
   wire signed [9:0] m20_38;
   assign m20_38 =10'b0;

   // m20_39 = W*in
   wire signed [9:0] m20_39;
   assign m20_39 =10'b0;

   // m20_40 = W*in
   wire signed [9:0] m20_40;
   assign m20_40 ={ {4{in20[5]}} , in20[5:0] };

   // m20_41 = W*in
   wire signed [9:0] m20_41;
   assign m20_41 =10'b0;

   // m20_42 = W*in
   wire signed [9:0] m20_42;
   assign m20_42 =10'b0;

   // m20_43 = W*in
   wire signed [9:0] m20_43;
   assign m20_43 =10'b0;

   // m20_44 = W*in
   wire signed [9:0] m20_44;
   assign m20_44 =10'b0;

   // m20_45 = W*in
   wire signed [9:0] m20_45;
   assign m20_45 ={ {4{in20[5]}} , in20[5:0] };

   // m20_46 = W*in
   wire signed [9:0] m20_46;
   assign m20_46 ={ {4{in20[5]}} , in20[5:0] };

   // m20_47 = W*in
   wire signed [9:0] m20_47;
   assign m20_47 =10'b0;

   // m20_48 = W*in
   wire signed [9:0] m20_48;
   assign m20_48 =10'b0;

   // m20_49 = W*in
   wire signed [9:0] m20_49;
   assign m20_49 =10'b0;

   // m20_50 = W*in
   wire signed [9:0] m20_50;
   assign m20_50 =10'b0;

   // m20_51 = W*in
   wire signed [9:0] m20_51;
   assign m20_51 ={ {4{in20[5]}} , in20[5:0] };

   // m20_52 = W*in
   wire signed [9:0] m20_52;
   assign m20_52 =10'b0;

   // m20_53 = W*in
   wire signed [9:0] m20_53;
   assign m20_53 =10'b0;

   // m20_54 = W*in
   wire signed [9:0] m20_54;
   assign m20_54 ={ {4{in20[5]}} , in20[5:0] };

   // m20_55 = W*in
   wire signed [9:0] m20_55;
   assign m20_55 =10'b0;

   // m20_56 = W*in
   wire signed [9:0] m20_56;
   assign m20_56 =10'b0;

   // m20_57 = W*in
   wire signed [9:0] m20_57;
   assign m20_57 =10'b0;

   // m20_58 = W*in
   wire signed [9:0] m20_58;
   assign m20_58 =10'b0;

   // m20_59 = W*in
   wire signed [9:0] m20_59;
   assign m20_59 ={ {4{in20[5]}} , in20[5:0] };

   // m20_60 = W*in
   wire signed [9:0] m20_60;
   assign m20_60 =10'b0;

   // m20_61 = W*in
   wire signed [9:0] m20_61;
   assign m20_61 =10'b0;

   // m20_62 = W*in
   wire signed [9:0] m20_62;
   assign m20_62 =10'b0;

   // m20_63 = W*in
   wire signed [9:0] m20_63;
   assign m20_63 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_64 = W*in
   wire signed [9:0] m20_64;
   assign m20_64 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_65 = W*in
   wire signed [9:0] m20_65;
   assign m20_65 =10'b0;

   // m20_66 = W*in
   wire signed [9:0] m20_66;
   assign m20_66 ={ {4{in20[5]}} , in20[5:0] };

   // m20_67 = W*in
   wire signed [9:0] m20_67;
   assign m20_67 =10'b0;

   // m20_68 = W*in
   wire signed [9:0] m20_68;
   assign m20_68 =10'b0;

   // m20_69 = W*in
   wire signed [9:0] m20_69;
   assign m20_69 =10'b0;

   // m20_70 = W*in
   wire signed [9:0] m20_70;
   assign m20_70 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_71 = W*in
   wire signed [9:0] m20_71;
   assign m20_71 ={ {5{in20[5]}} , in20[5:1] };

   // m20_72 = W*in
   wire signed [9:0] m20_72;
   assign m20_72 ={ {5{neg20[5]}} , neg20[5:1] };

   // m20_73 = W*in
   wire signed [9:0] m20_73;
   assign m20_73 ={ {5{in20[5]}} , in20[5:1] };

   // m20_74 = W*in
   wire signed [9:0] m20_74;
   assign m20_74 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_75 = W*in
   wire signed [9:0] m20_75;
   assign m20_75 =10'b0;

   // m20_76 = W*in
   wire signed [9:0] m20_76;
   assign m20_76 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_77 = W*in
   wire signed [9:0] m20_77;
   assign m20_77 ={ {3{in20[5]}} , in20 , {1{1'b0}} };

   // m20_78 = W*in
   wire signed [9:0] m20_78;
   assign m20_78 =10'b0;

   // m20_79 = W*in
   wire signed [9:0] m20_79;
   assign m20_79 =10'b0;

   // m20_80 = W*in
   wire signed [9:0] m20_80;
   assign m20_80 =10'b0;

   // m20_81 = W*in
   wire signed [9:0] m20_81;
   assign m20_81 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_82 = W*in
   wire signed [9:0] m20_82;
   assign m20_82 =10'b0;

   // m20_83 = W*in
   wire signed [9:0] m20_83;
   assign m20_83 =10'b0;

   // m20_84 = W*in
   wire signed [9:0] m20_84;
   assign m20_84 =10'b0;

   // m20_85 = W*in
   wire signed [9:0] m20_85;
   assign m20_85 ={ {4{in20[5]}} , in20[5:0] };

   // m20_86 = W*in
   wire signed [9:0] m20_86;
   assign m20_86 =10'b0;

   // m20_87 = W*in
   wire signed [9:0] m20_87;
   assign m20_87 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_88 = W*in
   wire signed [9:0] m20_88;
   assign m20_88 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_89 = W*in
   wire signed [9:0] m20_89;
   assign m20_89 =10'b0;

   // m20_90 = W*in
   wire signed [9:0] m20_90;
   assign m20_90 =10'b0;

   // m20_91 = W*in
   wire signed [9:0] m20_91;
   assign m20_91 =10'b0;

   // m20_92 = W*in
   wire signed [9:0] m20_92;
   assign m20_92 =10'b0;

   // m20_93 = W*in
   wire signed [9:0] m20_93;
   assign m20_93 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_94 = W*in
   wire signed [9:0] m20_94;
   assign m20_94 =10'b0;

   // m20_95 = W*in
   wire signed [9:0] m20_95;
   assign m20_95 ={ {4{in20[5]}} , in20[5:0] };

   // m20_96 = W*in
   wire signed [9:0] m20_96;
   assign m20_96 =10'b0;

   // m20_97 = W*in
   wire signed [9:0] m20_97;
   assign m20_97 ={ {5{in20[5]}} , in20[5:1] };

   // m20_98 = W*in
   wire signed [9:0] m20_98;
   assign m20_98 =10'b0;

   // m20_99 = W*in
   wire signed [9:0] m20_99;
   assign m20_99 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_100 = W*in
   wire signed [9:0] m20_100;
   assign m20_100 =10'b0;

   // m20_101 = W*in
   wire signed [9:0] m20_101;
   assign m20_101 =10'b0;

   // m20_102 = W*in
   wire signed [9:0] m20_102;
   assign m20_102 =10'b0;

   // m20_103 = W*in
   wire signed [9:0] m20_103;
   assign m20_103 =10'b0;

   // m20_104 = W*in
   wire signed [9:0] m20_104;
   assign m20_104 =10'b0;

   // m20_105 = W*in
   wire signed [9:0] m20_105;
   assign m20_105 =10'b0;

   // m20_106 = W*in
   wire signed [9:0] m20_106;
   assign m20_106 =10'b0;

   // m20_107 = W*in
   wire signed [9:0] m20_107;
   assign m20_107 ={ {4{in20[5]}} , in20[5:0] };

   // m20_108 = W*in
   wire signed [9:0] m20_108;
   assign m20_108 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_109 = W*in
   wire signed [9:0] m20_109;
   assign m20_109 =10'b0;

   // m20_110 = W*in
   wire signed [9:0] m20_110;
   assign m20_110 =10'b0;

   // m20_111 = W*in
   wire signed [9:0] m20_111;
   assign m20_111 =10'b0;

   // m20_112 = W*in
   wire signed [9:0] m20_112;
   assign m20_112 =10'b0;

   // m20_113 = W*in
   wire signed [9:0] m20_113;
   assign m20_113 =10'b0;

   // m20_114 = W*in
   wire signed [9:0] m20_114;
   assign m20_114 ={ {4{neg20[5]}} , neg20[5:0] };

   // m20_115 = W*in
   wire signed [9:0] m20_115;
   assign m20_115 =10'b0;

   // m20_116 = W*in
   wire signed [9:0] m20_116;
   assign m20_116 =10'b0;

   // m20_117 = W*in
   wire signed [9:0] m20_117;
   assign m20_117 =10'b0;

   // m21_1 = W*in
   wire signed [9:0] m21_1;
   assign m21_1 =10'b0;

   // m21_2 = W*in
   wire signed [9:0] m21_2;
   assign m21_2 =10'b0;

   // m21_3 = W*in
   wire signed [9:0] m21_3;
   assign m21_3 =10'b0;

   // m21_4 = W*in
   wire signed [9:0] m21_4;
   assign m21_4 =10'b0;

   // m21_5 = W*in
   wire signed [9:0] m21_5;
   assign m21_5 ={ {4{in21[5]}} , in21[5:0] };

   // m21_6 = W*in
   wire signed [9:0] m21_6;
   assign m21_6 ={ {4{in21[5]}} , in21[5:0] };

   // m21_7 = W*in
   wire signed [9:0] m21_7;
   assign m21_7 =10'b0;

   // m21_8 = W*in
   wire signed [9:0] m21_8;
   assign m21_8 =10'b0;

   // m21_9 = W*in
   wire signed [9:0] m21_9;
   assign m21_9 =10'b0;

   // m21_10 = W*in
   wire signed [9:0] m21_10;
   assign m21_10 =10'b0;

   // m21_11 = W*in
   wire signed [9:0] m21_11;
   assign m21_11 =10'b0;

   // m21_12 = W*in
   wire signed [9:0] m21_12;
   assign m21_12 ={ {4{neg21[5]}} , neg21[5:0] };

   // m21_13 = W*in
   wire signed [9:0] m21_13;
   assign m21_13 =10'b0;

   // m21_14 = W*in
   wire signed [9:0] m21_14;
   assign m21_14 =10'b0;

   // m21_15 = W*in
   wire signed [9:0] m21_15;
   assign m21_15 =10'b0;

   // m21_16 = W*in
   wire signed [9:0] m21_16;
   assign m21_16 =10'b0;

   // m21_17 = W*in
   wire signed [9:0] m21_17;
   assign m21_17 =10'b0;

   // m21_18 = W*in
   wire signed [9:0] m21_18;
   assign m21_18 ={ {5{neg21[5]}} , neg21[5:1] };

   // m21_19 = W*in
   wire signed [9:0] m21_19;
   assign m21_19 =10'b0;

   // m21_20 = W*in
   wire signed [9:0] m21_20;
   assign m21_20 =10'b0;

   // m21_21 = W*in
   wire signed [9:0] m21_21;
   assign m21_21 ={ {5{in21[5]}} , in21[5:1] };

   // m21_22 = W*in
   wire signed [9:0] m21_22;
   assign m21_22 =10'b0;

   // m21_23 = W*in
   wire signed [9:0] m21_23;
   assign m21_23 =10'b0;

   // m21_24 = W*in
   wire signed [9:0] m21_24;
   assign m21_24 =10'b0;

   // m21_25 = W*in
   wire signed [9:0] m21_25;
   assign m21_25 =10'b0;

   // m21_26 = W*in
   wire signed [9:0] m21_26;
   assign m21_26 =10'b0;

   // m21_27 = W*in
   wire signed [9:0] m21_27;
   assign m21_27 ={ {5{neg21[5]}} , neg21[5:1] };

   // m21_28 = W*in
   wire signed [9:0] m21_28;
   assign m21_28 =10'b0;

   // m21_29 = W*in
   wire signed [9:0] m21_29;
   assign m21_29 ={ {5{in21[5]}} , in21[5:1] };

   // m21_30 = W*in
   wire signed [9:0] m21_30;
   assign m21_30 =10'b0;

   // m21_31 = W*in
   wire signed [9:0] m21_31;
   assign m21_31 =10'b0;

   // m21_32 = W*in
   wire signed [9:0] m21_32;
   assign m21_32 =10'b0;

   // m21_33 = W*in
   wire signed [9:0] m21_33;
   assign m21_33 =10'b0;

   // m21_34 = W*in
   wire signed [9:0] m21_34;
   assign m21_34 =10'b0;

   // m21_35 = W*in
   wire signed [9:0] m21_35;
   assign m21_35 =10'b0;

   // m21_36 = W*in
   wire signed [9:0] m21_36;
   assign m21_36 =10'b0;

   // m21_37 = W*in
   wire signed [9:0] m21_37;
   assign m21_37 ={ {4{in21[5]}} , in21[5:0] };

   // m21_38 = W*in
   wire signed [9:0] m21_38;
   assign m21_38 =10'b0;

   // m21_39 = W*in
   wire signed [9:0] m21_39;
   assign m21_39 =10'b0;

   // m21_40 = W*in
   wire signed [9:0] m21_40;
   assign m21_40 =10'b0;

   // m21_41 = W*in
   wire signed [9:0] m21_41;
   assign m21_41 ={ {4{in21[5]}} , in21[5:0] };

   // m21_42 = W*in
   wire signed [9:0] m21_42;
   assign m21_42 =10'b0;

   // m21_43 = W*in
   wire signed [9:0] m21_43;
   assign m21_43 =10'b0;

   // m21_44 = W*in
   wire signed [9:0] m21_44;
   assign m21_44 =10'b0;

   // m21_45 = W*in
   wire signed [9:0] m21_45;
   assign m21_45 =10'b0;

   // m21_46 = W*in
   wire signed [9:0] m21_46;
   assign m21_46 =10'b0;

   // m21_47 = W*in
   wire signed [9:0] m21_47;
   assign m21_47 =10'b0;

   // m21_48 = W*in
   wire signed [9:0] m21_48;
   assign m21_48 =10'b0;

   // m21_49 = W*in
   wire signed [9:0] m21_49;
   assign m21_49 =10'b0;

   // m21_50 = W*in
   wire signed [9:0] m21_50;
   assign m21_50 =10'b0;

   // m21_51 = W*in
   wire signed [9:0] m21_51;
   assign m21_51 =10'b0;

   // m21_52 = W*in
   wire signed [9:0] m21_52;
   assign m21_52 =10'b0;

   // m21_53 = W*in
   wire signed [9:0] m21_53;
   assign m21_53 =10'b0;

   // m21_54 = W*in
   wire signed [9:0] m21_54;
   assign m21_54 =10'b0;

   // m21_55 = W*in
   wire signed [9:0] m21_55;
   assign m21_55 =10'b0;

   // m21_56 = W*in
   wire signed [9:0] m21_56;
   assign m21_56 =10'b0;

   // m21_57 = W*in
   wire signed [9:0] m21_57;
   assign m21_57 =10'b0;

   // m21_58 = W*in
   wire signed [9:0] m21_58;
   assign m21_58 =10'b0;

   // m21_59 = W*in
   wire signed [9:0] m21_59;
   assign m21_59 =10'b0;

   // m21_60 = W*in
   wire signed [9:0] m21_60;
   assign m21_60 =10'b0;

   // m21_61 = W*in
   wire signed [9:0] m21_61;
   assign m21_61 =10'b0;

   // m21_62 = W*in
   wire signed [9:0] m21_62;
   assign m21_62 =10'b0;

   // m21_63 = W*in
   wire signed [9:0] m21_63;
   assign m21_63 ={ {4{in21[5]}} , in21[5:0] };

   // m21_64 = W*in
   wire signed [9:0] m21_64;
   assign m21_64 ={ {4{neg21[5]}} , neg21[5:0] };

   // m21_65 = W*in
   wire signed [9:0] m21_65;
   assign m21_65 ={ {5{in21[5]}} , in21[5:1] };

   // m21_66 = W*in
   wire signed [9:0] m21_66;
   assign m21_66 =10'b0;

   // m21_67 = W*in
   wire signed [9:0] m21_67;
   assign m21_67 =10'b0;

   // m21_68 = W*in
   wire signed [9:0] m21_68;
   assign m21_68 ={ {4{neg21[5]}} , neg21[5:0] };

   // m21_69 = W*in
   wire signed [9:0] m21_69;
   assign m21_69 ={ {5{in21[5]}} , in21[5:1] };

   // m21_70 = W*in
   wire signed [9:0] m21_70;
   assign m21_70 ={ {5{in21[5]}} , in21[5:1] };

   // m21_71 = W*in
   wire signed [9:0] m21_71;
   assign m21_71 ={ {5{neg21[5]}} , neg21[5:1] };

   // m21_72 = W*in
   wire signed [9:0] m21_72;
   assign m21_72 =10'b0;

   // m21_73 = W*in
   wire signed [9:0] m21_73;
   assign m21_73 =10'b0;

   // m21_74 = W*in
   wire signed [9:0] m21_74;
   assign m21_74 =10'b0;

   // m21_75 = W*in
   wire signed [9:0] m21_75;
   assign m21_75 =10'b0;

   // m21_76 = W*in
   wire signed [9:0] m21_76;
   assign m21_76 =10'b0;

   // m21_77 = W*in
   wire signed [9:0] m21_77;
   assign m21_77 =10'b0;

   // m21_78 = W*in
   wire signed [9:0] m21_78;
   assign m21_78 =10'b0;

   // m21_79 = W*in
   wire signed [9:0] m21_79;
   assign m21_79 =10'b0;

   // m21_80 = W*in
   wire signed [9:0] m21_80;
   assign m21_80 =10'b0;

   // m21_81 = W*in
   wire signed [9:0] m21_81;
   assign m21_81 ={ {5{neg21[5]}} , neg21[5:1] };

   // m21_82 = W*in
   wire signed [9:0] m21_82;
   assign m21_82 ={ {5{in21[5]}} , in21[5:1] };

   // m21_83 = W*in
   wire signed [9:0] m21_83;
   assign m21_83 =10'b0;

   // m21_84 = W*in
   wire signed [9:0] m21_84;
   assign m21_84 =10'b0;

   // m21_85 = W*in
   wire signed [9:0] m21_85;
   assign m21_85 ={ {4{in21[5]}} , in21[5:0] };

   // m21_86 = W*in
   wire signed [9:0] m21_86;
   assign m21_86 =10'b0;

   // m21_87 = W*in
   wire signed [9:0] m21_87;
   assign m21_87 =10'b0;

   // m21_88 = W*in
   wire signed [9:0] m21_88;
   assign m21_88 =10'b0;

   // m21_89 = W*in
   wire signed [9:0] m21_89;
   assign m21_89 =10'b0;

   // m21_90 = W*in
   wire signed [9:0] m21_90;
   assign m21_90 =10'b0;

   // m21_91 = W*in
   wire signed [9:0] m21_91;
   assign m21_91 =10'b0;

   // m21_92 = W*in
   wire signed [9:0] m21_92;
   assign m21_92 =10'b0;

   // m21_93 = W*in
   wire signed [9:0] m21_93;
   assign m21_93 ={ {4{in21[5]}} , in21[5:0] };

   // m21_94 = W*in
   wire signed [9:0] m21_94;
   assign m21_94 =10'b0;

   // m21_95 = W*in
   wire signed [9:0] m21_95;
   assign m21_95 =10'b0;

   // m21_96 = W*in
   wire signed [9:0] m21_96;
   assign m21_96 =10'b0;

   // m21_97 = W*in
   wire signed [9:0] m21_97;
   assign m21_97 =10'b0;

   // m21_98 = W*in
   wire signed [9:0] m21_98;
   assign m21_98 =10'b0;

   // m21_99 = W*in
   wire signed [9:0] m21_99;
   assign m21_99 =10'b0;

   // m21_100 = W*in
   wire signed [9:0] m21_100;
   assign m21_100 =10'b0;

   // m21_101 = W*in
   wire signed [9:0] m21_101;
   assign m21_101 =10'b0;

   // m21_102 = W*in
   wire signed [9:0] m21_102;
   assign m21_102 =10'b0;

   // m21_103 = W*in
   wire signed [9:0] m21_103;
   assign m21_103 =10'b0;

   // m21_104 = W*in
   wire signed [9:0] m21_104;
   assign m21_104 =10'b0;

   // m21_105 = W*in
   wire signed [9:0] m21_105;
   assign m21_105 =10'b0;

   // m21_106 = W*in
   wire signed [9:0] m21_106;
   assign m21_106 =10'b0;

   // m21_107 = W*in
   wire signed [9:0] m21_107;
   assign m21_107 =10'b0;

   // m21_108 = W*in
   wire signed [9:0] m21_108;
   assign m21_108 ={ {4{in21[5]}} , in21[5:0] };

   // m21_109 = W*in
   wire signed [9:0] m21_109;
   assign m21_109 =10'b0;

   // m21_110 = W*in
   wire signed [9:0] m21_110;
   assign m21_110 =10'b0;

   // m21_111 = W*in
   wire signed [9:0] m21_111;
   assign m21_111 =10'b0;

   // m21_112 = W*in
   wire signed [9:0] m21_112;
   assign m21_112 =10'b0;

   // m21_113 = W*in
   wire signed [9:0] m21_113;
   assign m21_113 =10'b0;

   // m21_114 = W*in
   wire signed [9:0] m21_114;
   assign m21_114 =10'b0;

   // m21_115 = W*in
   wire signed [9:0] m21_115;
   assign m21_115 =10'b0;

   // m21_116 = W*in
   wire signed [9:0] m21_116;
   assign m21_116 =10'b0;

   // m21_117 = W*in
   wire signed [9:0] m21_117;
   assign m21_117 =10'b0;

   // m22_1 = W*in
   wire signed [9:0] m22_1;
   assign m22_1 =10'b0;

   // m22_2 = W*in
   wire signed [9:0] m22_2;
   assign m22_2 =10'b0;

   // m22_3 = W*in
   wire signed [9:0] m22_3;
   assign m22_3 =10'b0;

   // m22_4 = W*in
   wire signed [9:0] m22_4;
   assign m22_4 =10'b0;

   // m22_5 = W*in
   wire signed [9:0] m22_5;
   assign m22_5 =10'b0;

   // m22_6 = W*in
   wire signed [9:0] m22_6;
   assign m22_6 ={ {5{in22[5]}} , in22[5:1] };

   // m22_7 = W*in
   wire signed [9:0] m22_7;
   assign m22_7 =10'b0;

   // m22_8 = W*in
   wire signed [9:0] m22_8;
   assign m22_8 =10'b0;

   // m22_9 = W*in
   wire signed [9:0] m22_9;
   assign m22_9 =10'b0;

   // m22_10 = W*in
   wire signed [9:0] m22_10;
   assign m22_10 =10'b0;

   // m22_11 = W*in
   wire signed [9:0] m22_11;
   assign m22_11 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_12 = W*in
   wire signed [9:0] m22_12;
   assign m22_12 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_13 = W*in
   wire signed [9:0] m22_13;
   assign m22_13 =10'b0;

   // m22_14 = W*in
   wire signed [9:0] m22_14;
   assign m22_14 =10'b0;

   // m22_15 = W*in
   wire signed [9:0] m22_15;
   assign m22_15 =10'b0;

   // m22_16 = W*in
   wire signed [9:0] m22_16;
   assign m22_16 =10'b0;

   // m22_17 = W*in
   wire signed [9:0] m22_17;
   assign m22_17 =10'b0;

   // m22_18 = W*in
   wire signed [9:0] m22_18;
   assign m22_18 =10'b0;

   // m22_19 = W*in
   wire signed [9:0] m22_19;
   assign m22_19 =10'b0;

   // m22_20 = W*in
   wire signed [9:0] m22_20;
   assign m22_20 =10'b0;

   // m22_21 = W*in
   wire signed [9:0] m22_21;
   assign m22_21 =10'b0;

   // m22_22 = W*in
   wire signed [9:0] m22_22;
   assign m22_22 =10'b0;

   // m22_23 = W*in
   wire signed [9:0] m22_23;
   assign m22_23 =10'b0;

   // m22_24 = W*in
   wire signed [9:0] m22_24;
   assign m22_24 =10'b0;

   // m22_25 = W*in
   wire signed [9:0] m22_25;
   assign m22_25 =10'b0;

   // m22_26 = W*in
   wire signed [9:0] m22_26;
   assign m22_26 ={ {5{neg22[5]}} , neg22[5:1] };

   // m22_27 = W*in
   wire signed [9:0] m22_27;
   assign m22_27 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_28 = W*in
   wire signed [9:0] m22_28;
   assign m22_28 ={ {5{neg22[5]}} , neg22[5:1] };

   // m22_29 = W*in
   wire signed [9:0] m22_29;
   assign m22_29 =10'b0;

   // m22_30 = W*in
   wire signed [9:0] m22_30;
   assign m22_30 =10'b0;

   // m22_31 = W*in
   wire signed [9:0] m22_31;
   assign m22_31 ={ {5{neg22[5]}} , neg22[5:1] };

   // m22_32 = W*in
   wire signed [9:0] m22_32;
   assign m22_32 ={ {5{in22[5]}} , in22[5:1] };

   // m22_33 = W*in
   wire signed [9:0] m22_33;
   assign m22_33 =10'b0;

   // m22_34 = W*in
   wire signed [9:0] m22_34;
   assign m22_34 =10'b0;

   // m22_35 = W*in
   wire signed [9:0] m22_35;
   assign m22_35 =10'b0;

   // m22_36 = W*in
   wire signed [9:0] m22_36;
   assign m22_36 =10'b0;

   // m22_37 = W*in
   wire signed [9:0] m22_37;
   assign m22_37 ={ {4{in22[5]}} , in22[5:0] };

   // m22_38 = W*in
   wire signed [9:0] m22_38;
   assign m22_38 =10'b0;

   // m22_39 = W*in
   wire signed [9:0] m22_39;
   assign m22_39 =10'b0;

   // m22_40 = W*in
   wire signed [9:0] m22_40;
   assign m22_40 =10'b0;

   // m22_41 = W*in
   wire signed [9:0] m22_41;
   assign m22_41 =10'b0;

   // m22_42 = W*in
   wire signed [9:0] m22_42;
   assign m22_42 =10'b0;

   // m22_43 = W*in
   wire signed [9:0] m22_43;
   assign m22_43 =10'b0;

   // m22_44 = W*in
   wire signed [9:0] m22_44;
   assign m22_44 =10'b0;

   // m22_45 = W*in
   wire signed [9:0] m22_45;
   assign m22_45 ={ {4{in22[5]}} , in22[5:0] };

   // m22_46 = W*in
   wire signed [9:0] m22_46;
   assign m22_46 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_47 = W*in
   wire signed [9:0] m22_47;
   assign m22_47 =10'b0;

   // m22_48 = W*in
   wire signed [9:0] m22_48;
   assign m22_48 ={ {4{in22[5]}} , in22[5:0] };

   // m22_49 = W*in
   wire signed [9:0] m22_49;
   assign m22_49 =10'b0;

   // m22_50 = W*in
   wire signed [9:0] m22_50;
   assign m22_50 =10'b0;

   // m22_51 = W*in
   wire signed [9:0] m22_51;
   assign m22_51 =10'b0;

   // m22_52 = W*in
   wire signed [9:0] m22_52;
   assign m22_52 =10'b0;

   // m22_53 = W*in
   wire signed [9:0] m22_53;
   assign m22_53 =10'b0;

   // m22_54 = W*in
   wire signed [9:0] m22_54;
   assign m22_54 =10'b0;

   // m22_55 = W*in
   wire signed [9:0] m22_55;
   assign m22_55 =10'b0;

   // m22_56 = W*in
   wire signed [9:0] m22_56;
   assign m22_56 =10'b0;

   // m22_57 = W*in
   wire signed [9:0] m22_57;
   assign m22_57 =10'b0;

   // m22_58 = W*in
   wire signed [9:0] m22_58;
   assign m22_58 =10'b0;

   // m22_59 = W*in
   wire signed [9:0] m22_59;
   assign m22_59 =10'b0;

   // m22_60 = W*in
   wire signed [9:0] m22_60;
   assign m22_60 =10'b0;

   // m22_61 = W*in
   wire signed [9:0] m22_61;
   assign m22_61 =10'b0;

   // m22_62 = W*in
   wire signed [9:0] m22_62;
   assign m22_62 =10'b0;

   // m22_63 = W*in
   wire signed [9:0] m22_63;
   assign m22_63 =10'b0;

   // m22_64 = W*in
   wire signed [9:0] m22_64;
   assign m22_64 =10'b0;

   // m22_65 = W*in
   wire signed [9:0] m22_65;
   assign m22_65 ={ {5{in22[5]}} , in22[5:1] };

   // m22_66 = W*in
   wire signed [9:0] m22_66;
   assign m22_66 ={ {5{neg22[5]}} , neg22[5:1] };

   // m22_67 = W*in
   wire signed [9:0] m22_67;
   assign m22_67 =10'b0;

   // m22_68 = W*in
   wire signed [9:0] m22_68;
   assign m22_68 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_69 = W*in
   wire signed [9:0] m22_69;
   assign m22_69 ={ {4{in22[5]}} , in22[5:0] };

   // m22_70 = W*in
   wire signed [9:0] m22_70;
   assign m22_70 ={ {5{in22[5]}} , in22[5:1] };

   // m22_71 = W*in
   wire signed [9:0] m22_71;
   assign m22_71 =10'b0;

   // m22_72 = W*in
   wire signed [9:0] m22_72;
   assign m22_72 ={ {5{in22[5]}} , in22[5:1] };

   // m22_73 = W*in
   wire signed [9:0] m22_73;
   assign m22_73 =10'b0;

   // m22_74 = W*in
   wire signed [9:0] m22_74;
   assign m22_74 =10'b0;

   // m22_75 = W*in
   wire signed [9:0] m22_75;
   assign m22_75 =10'b0;

   // m22_76 = W*in
   wire signed [9:0] m22_76;
   assign m22_76 =10'b0;

   // m22_77 = W*in
   wire signed [9:0] m22_77;
   assign m22_77 =10'b0;

   // m22_78 = W*in
   wire signed [9:0] m22_78;
   assign m22_78 =10'b0;

   // m22_79 = W*in
   wire signed [9:0] m22_79;
   assign m22_79 =10'b0;

   // m22_80 = W*in
   wire signed [9:0] m22_80;
   assign m22_80 =10'b0;

   // m22_81 = W*in
   wire signed [9:0] m22_81;
   assign m22_81 =10'b0;

   // m22_82 = W*in
   wire signed [9:0] m22_82;
   assign m22_82 =10'b0;

   // m22_83 = W*in
   wire signed [9:0] m22_83;
   assign m22_83 =10'b0;

   // m22_84 = W*in
   wire signed [9:0] m22_84;
   assign m22_84 =10'b0;

   // m22_85 = W*in
   wire signed [9:0] m22_85;
   assign m22_85 =10'b0;

   // m22_86 = W*in
   wire signed [9:0] m22_86;
   assign m22_86 =10'b0;

   // m22_87 = W*in
   wire signed [9:0] m22_87;
   assign m22_87 =10'b0;

   // m22_88 = W*in
   wire signed [9:0] m22_88;
   assign m22_88 =10'b0;

   // m22_89 = W*in
   wire signed [9:0] m22_89;
   assign m22_89 =10'b0;

   // m22_90 = W*in
   wire signed [9:0] m22_90;
   assign m22_90 =10'b0;

   // m22_91 = W*in
   wire signed [9:0] m22_91;
   assign m22_91 =10'b0;

   // m22_92 = W*in
   wire signed [9:0] m22_92;
   assign m22_92 =10'b0;

   // m22_93 = W*in
   wire signed [9:0] m22_93;
   assign m22_93 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_94 = W*in
   wire signed [9:0] m22_94;
   assign m22_94 =10'b0;

   // m22_95 = W*in
   wire signed [9:0] m22_95;
   assign m22_95 =10'b0;

   // m22_96 = W*in
   wire signed [9:0] m22_96;
   assign m22_96 =10'b0;

   // m22_97 = W*in
   wire signed [9:0] m22_97;
   assign m22_97 =10'b0;

   // m22_98 = W*in
   wire signed [9:0] m22_98;
   assign m22_98 =10'b0;

   // m22_99 = W*in
   wire signed [9:0] m22_99;
   assign m22_99 ={ {4{in22[5]}} , in22[5:0] };

   // m22_100 = W*in
   wire signed [9:0] m22_100;
   assign m22_100 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_101 = W*in
   wire signed [9:0] m22_101;
   assign m22_101 =10'b0;

   // m22_102 = W*in
   wire signed [9:0] m22_102;
   assign m22_102 =10'b0;

   // m22_103 = W*in
   wire signed [9:0] m22_103;
   assign m22_103 =10'b0;

   // m22_104 = W*in
   wire signed [9:0] m22_104;
   assign m22_104 ={ {4{neg22[5]}} , neg22[5:0] };

   // m22_105 = W*in
   wire signed [9:0] m22_105;
   assign m22_105 =10'b0;

   // m22_106 = W*in
   wire signed [9:0] m22_106;
   assign m22_106 =10'b0;

   // m22_107 = W*in
   wire signed [9:0] m22_107;
   assign m22_107 =10'b0;

   // m22_108 = W*in
   wire signed [9:0] m22_108;
   assign m22_108 =10'b0;

   // m22_109 = W*in
   wire signed [9:0] m22_109;
   assign m22_109 =10'b0;

   // m22_110 = W*in
   wire signed [9:0] m22_110;
   assign m22_110 =10'b0;

   // m22_111 = W*in
   wire signed [9:0] m22_111;
   assign m22_111 =10'b0;

   // m22_112 = W*in
   wire signed [9:0] m22_112;
   assign m22_112 =10'b0;

   // m22_113 = W*in
   wire signed [9:0] m22_113;
   assign m22_113 =10'b0;

   // m22_114 = W*in
   wire signed [9:0] m22_114;
   assign m22_114 =10'b0;

   // m22_115 = W*in
   wire signed [9:0] m22_115;
   assign m22_115 =10'b0;

   // m22_116 = W*in
   wire signed [9:0] m22_116;
   assign m22_116 =10'b0;

   // m22_117 = W*in
   wire signed [9:0] m22_117;
   assign m22_117 =10'b0;

   // m23_1 = W*in
   wire signed [9:0] m23_1;
   assign m23_1 =10'b0;

   // m23_2 = W*in
   wire signed [9:0] m23_2;
   assign m23_2 =10'b0;

   // m23_3 = W*in
   wire signed [9:0] m23_3;
   assign m23_3 ={ {4{in23[5]}} , in23[5:0] };

   // m23_4 = W*in
   wire signed [9:0] m23_4;
   assign m23_4 =10'b0;

   // m23_5 = W*in
   wire signed [9:0] m23_5;
   assign m23_5 =10'b0;

   // m23_6 = W*in
   wire signed [9:0] m23_6;
   assign m23_6 =10'b0;

   // m23_7 = W*in
   wire signed [9:0] m23_7;
   assign m23_7 =10'b0;

   // m23_8 = W*in
   wire signed [9:0] m23_8;
   assign m23_8 =10'b0;

   // m23_9 = W*in
   wire signed [9:0] m23_9;
   assign m23_9 =10'b0;

   // m23_10 = W*in
   wire signed [9:0] m23_10;
   assign m23_10 =10'b0;

   // m23_11 = W*in
   wire signed [9:0] m23_11;
   assign m23_11 =10'b0;

   // m23_12 = W*in
   wire signed [9:0] m23_12;
   assign m23_12 =10'b0;

   // m23_13 = W*in
   wire signed [9:0] m23_13;
   assign m23_13 =10'b0;

   // m23_14 = W*in
   wire signed [9:0] m23_14;
   assign m23_14 =10'b0;

   // m23_15 = W*in
   wire signed [9:0] m23_15;
   assign m23_15 =10'b0;

   // m23_16 = W*in
   wire signed [9:0] m23_16;
   assign m23_16 =10'b0;

   // m23_17 = W*in
   wire signed [9:0] m23_17;
   assign m23_17 =10'b0;

   // m23_18 = W*in
   wire signed [9:0] m23_18;
   assign m23_18 =10'b0;

   // m23_19 = W*in
   wire signed [9:0] m23_19;
   assign m23_19 ={ {4{in23[5]}} , in23[5:0] };

   // m23_20 = W*in
   wire signed [9:0] m23_20;
   assign m23_20 =10'b0;

   // m23_21 = W*in
   wire signed [9:0] m23_21;
   assign m23_21 =10'b0;

   // m23_22 = W*in
   wire signed [9:0] m23_22;
   assign m23_22 =10'b0;

   // m23_23 = W*in
   wire signed [9:0] m23_23;
   assign m23_23 =10'b0;

   // m23_24 = W*in
   wire signed [9:0] m23_24;
   assign m23_24 =10'b0;

   // m23_25 = W*in
   wire signed [9:0] m23_25;
   assign m23_25 =10'b0;

   // m23_26 = W*in
   wire signed [9:0] m23_26;
   assign m23_26 =10'b0;

   // m23_27 = W*in
   wire signed [9:0] m23_27;
   assign m23_27 =10'b0;

   // m23_28 = W*in
   wire signed [9:0] m23_28;
   assign m23_28 ={ {5{neg23[5]}} , neg23[5:1] };

   // m23_29 = W*in
   wire signed [9:0] m23_29;
   assign m23_29 =10'b0;

   // m23_30 = W*in
   wire signed [9:0] m23_30;
   assign m23_30 =10'b0;

   // m23_31 = W*in
   wire signed [9:0] m23_31;
   assign m23_31 =10'b0;

   // m23_32 = W*in
   wire signed [9:0] m23_32;
   assign m23_32 =10'b0;

   // m23_33 = W*in
   wire signed [9:0] m23_33;
   assign m23_33 =10'b0;

   // m23_34 = W*in
   wire signed [9:0] m23_34;
   assign m23_34 =10'b0;

   // m23_35 = W*in
   wire signed [9:0] m23_35;
   assign m23_35 =10'b0;

   // m23_36 = W*in
   wire signed [9:0] m23_36;
   assign m23_36 =10'b0;

   // m23_37 = W*in
   wire signed [9:0] m23_37;
   assign m23_37 =10'b0;

   // m23_38 = W*in
   wire signed [9:0] m23_38;
   assign m23_38 =10'b0;

   // m23_39 = W*in
   wire signed [9:0] m23_39;
   assign m23_39 =10'b0;

   // m23_40 = W*in
   wire signed [9:0] m23_40;
   assign m23_40 =10'b0;

   // m23_41 = W*in
   wire signed [9:0] m23_41;
   assign m23_41 =10'b0;

   // m23_42 = W*in
   wire signed [9:0] m23_42;
   assign m23_42 =10'b0;

   // m23_43 = W*in
   wire signed [9:0] m23_43;
   assign m23_43 =10'b0;

   // m23_44 = W*in
   wire signed [9:0] m23_44;
   assign m23_44 =10'b0;

   // m23_45 = W*in
   wire signed [9:0] m23_45;
   assign m23_45 =10'b0;

   // m23_46 = W*in
   wire signed [9:0] m23_46;
   assign m23_46 =10'b0;

   // m23_47 = W*in
   wire signed [9:0] m23_47;
   assign m23_47 =10'b0;

   // m23_48 = W*in
   wire signed [9:0] m23_48;
   assign m23_48 =10'b0;

   // m23_49 = W*in
   wire signed [9:0] m23_49;
   assign m23_49 =10'b0;

   // m23_50 = W*in
   wire signed [9:0] m23_50;
   assign m23_50 =10'b0;

   // m23_51 = W*in
   wire signed [9:0] m23_51;
   assign m23_51 =10'b0;

   // m23_52 = W*in
   wire signed [9:0] m23_52;
   assign m23_52 =10'b0;

   // m23_53 = W*in
   wire signed [9:0] m23_53;
   assign m23_53 =10'b0;

   // m23_54 = W*in
   wire signed [9:0] m23_54;
   assign m23_54 =10'b0;

   // m23_55 = W*in
   wire signed [9:0] m23_55;
   assign m23_55 =10'b0;

   // m23_56 = W*in
   wire signed [9:0] m23_56;
   assign m23_56 =10'b0;

   // m23_57 = W*in
   wire signed [9:0] m23_57;
   assign m23_57 =10'b0;

   // m23_58 = W*in
   wire signed [9:0] m23_58;
   assign m23_58 =10'b0;

   // m23_59 = W*in
   wire signed [9:0] m23_59;
   assign m23_59 =10'b0;

   // m23_60 = W*in
   wire signed [9:0] m23_60;
   assign m23_60 ={ {4{in23[5]}} , in23[5:0] };

   // m23_61 = W*in
   wire signed [9:0] m23_61;
   assign m23_61 =10'b0;

   // m23_62 = W*in
   wire signed [9:0] m23_62;
   assign m23_62 =10'b0;

   // m23_63 = W*in
   wire signed [9:0] m23_63;
   assign m23_63 =10'b0;

   // m23_64 = W*in
   wire signed [9:0] m23_64;
   assign m23_64 ={ {5{neg23[5]}} , neg23[5:1] };

   // m23_65 = W*in
   wire signed [9:0] m23_65;
   assign m23_65 ={ {5{neg23[5]}} , neg23[5:1] };

   // m23_66 = W*in
   wire signed [9:0] m23_66;
   assign m23_66 =10'b0;

   // m23_67 = W*in
   wire signed [9:0] m23_67;
   assign m23_67 =10'b0;

   // m23_68 = W*in
   wire signed [9:0] m23_68;
   assign m23_68 =10'b0;

   // m23_69 = W*in
   wire signed [9:0] m23_69;
   assign m23_69 =10'b0;

   // m23_70 = W*in
   wire signed [9:0] m23_70;
   assign m23_70 =10'b0;

   // m23_71 = W*in
   wire signed [9:0] m23_71;
   assign m23_71 =10'b0;

   // m23_72 = W*in
   wire signed [9:0] m23_72;
   assign m23_72 =10'b0;

   // m23_73 = W*in
   wire signed [9:0] m23_73;
   assign m23_73 =10'b0;

   // m23_74 = W*in
   wire signed [9:0] m23_74;
   assign m23_74 =10'b0;

   // m23_75 = W*in
   wire signed [9:0] m23_75;
   assign m23_75 =10'b0;

   // m23_76 = W*in
   wire signed [9:0] m23_76;
   assign m23_76 ={ {4{neg23[5]}} , neg23[5:0] };

   // m23_77 = W*in
   wire signed [9:0] m23_77;
   assign m23_77 =10'b0;

   // m23_78 = W*in
   wire signed [9:0] m23_78;
   assign m23_78 =10'b0;

   // m23_79 = W*in
   wire signed [9:0] m23_79;
   assign m23_79 =10'b0;

   // m23_80 = W*in
   wire signed [9:0] m23_80;
   assign m23_80 =10'b0;

   // m23_81 = W*in
   wire signed [9:0] m23_81;
   assign m23_81 =10'b0;

   // m23_82 = W*in
   wire signed [9:0] m23_82;
   assign m23_82 =10'b0;

   // m23_83 = W*in
   wire signed [9:0] m23_83;
   assign m23_83 =10'b0;

   // m23_84 = W*in
   wire signed [9:0] m23_84;
   assign m23_84 =10'b0;

   // m23_85 = W*in
   wire signed [9:0] m23_85;
   assign m23_85 =10'b0;

   // m23_86 = W*in
   wire signed [9:0] m23_86;
   assign m23_86 =10'b0;

   // m23_87 = W*in
   wire signed [9:0] m23_87;
   assign m23_87 =10'b0;

   // m23_88 = W*in
   wire signed [9:0] m23_88;
   assign m23_88 =10'b0;

   // m23_89 = W*in
   wire signed [9:0] m23_89;
   assign m23_89 =10'b0;

   // m23_90 = W*in
   wire signed [9:0] m23_90;
   assign m23_90 =10'b0;

   // m23_91 = W*in
   wire signed [9:0] m23_91;
   assign m23_91 =10'b0;

   // m23_92 = W*in
   wire signed [9:0] m23_92;
   assign m23_92 =10'b0;

   // m23_93 = W*in
   wire signed [9:0] m23_93;
   assign m23_93 =10'b0;

   // m23_94 = W*in
   wire signed [9:0] m23_94;
   assign m23_94 =10'b0;

   // m23_95 = W*in
   wire signed [9:0] m23_95;
   assign m23_95 =10'b0;

   // m23_96 = W*in
   wire signed [9:0] m23_96;
   assign m23_96 =10'b0;

   // m23_97 = W*in
   wire signed [9:0] m23_97;
   assign m23_97 ={ {4{neg23[5]}} , neg23[5:0] };

   // m23_98 = W*in
   wire signed [9:0] m23_98;
   assign m23_98 =10'b0;

   // m23_99 = W*in
   wire signed [9:0] m23_99;
   assign m23_99 =10'b0;

   // m23_100 = W*in
   wire signed [9:0] m23_100;
   assign m23_100 =10'b0;

   // m23_101 = W*in
   wire signed [9:0] m23_101;
   assign m23_101 =10'b0;

   // m23_102 = W*in
   wire signed [9:0] m23_102;
   assign m23_102 =10'b0;

   // m23_103 = W*in
   wire signed [9:0] m23_103;
   assign m23_103 ={ {4{in23[5]}} , in23[5:0] };

   // m23_104 = W*in
   wire signed [9:0] m23_104;
   assign m23_104 =10'b0;

   // m23_105 = W*in
   wire signed [9:0] m23_105;
   assign m23_105 =10'b0;

   // m23_106 = W*in
   wire signed [9:0] m23_106;
   assign m23_106 =10'b0;

   // m23_107 = W*in
   wire signed [9:0] m23_107;
   assign m23_107 ={ {4{in23[5]}} , in23[5:0] };

   // m23_108 = W*in
   wire signed [9:0] m23_108;
   assign m23_108 =10'b0;

   // m23_109 = W*in
   wire signed [9:0] m23_109;
   assign m23_109 =10'b0;

   // m23_110 = W*in
   wire signed [9:0] m23_110;
   assign m23_110 =10'b0;

   // m23_111 = W*in
   wire signed [9:0] m23_111;
   assign m23_111 =10'b0;

   // m23_112 = W*in
   wire signed [9:0] m23_112;
   assign m23_112 =10'b0;

   // m23_113 = W*in
   wire signed [9:0] m23_113;
   assign m23_113 =10'b0;

   // m23_114 = W*in
   wire signed [9:0] m23_114;
   assign m23_114 =10'b0;

   // m23_115 = W*in
   wire signed [9:0] m23_115;
   assign m23_115 =10'b0;

   // m23_116 = W*in
   wire signed [9:0] m23_116;
   assign m23_116 ={ {4{in23[5]}} , in23[5:0] };

   // m23_117 = W*in
   wire signed [9:0] m23_117;
   assign m23_117 =10'b0;

   // m24_1 = W*in
   wire signed [9:0] m24_1;
   assign m24_1 =10'b0;

   // m24_2 = W*in
   wire signed [9:0] m24_2;
   assign m24_2 =10'b0;

   // m24_3 = W*in
   wire signed [9:0] m24_3;
   assign m24_3 =10'b0;

   // m24_4 = W*in
   wire signed [9:0] m24_4;
   assign m24_4 =10'b0;

   // m24_5 = W*in
   wire signed [9:0] m24_5;
   assign m24_5 =10'b0;

   // m24_6 = W*in
   wire signed [9:0] m24_6;
   assign m24_6 =10'b0;

   // m24_7 = W*in
   wire signed [9:0] m24_7;
   assign m24_7 =10'b0;

   // m24_8 = W*in
   wire signed [9:0] m24_8;
   assign m24_8 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_9 = W*in
   wire signed [9:0] m24_9;
   assign m24_9 =10'b0;

   // m24_10 = W*in
   wire signed [9:0] m24_10;
   assign m24_10 =10'b0;

   // m24_11 = W*in
   wire signed [9:0] m24_11;
   assign m24_11 ={ {4{in24[5]}} , in24[5:0] };

   // m24_12 = W*in
   wire signed [9:0] m24_12;
   assign m24_12 =10'b0;

   // m24_13 = W*in
   wire signed [9:0] m24_13;
   assign m24_13 =10'b0;

   // m24_14 = W*in
   wire signed [9:0] m24_14;
   assign m24_14 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_15 = W*in
   wire signed [9:0] m24_15;
   assign m24_15 =10'b0;

   // m24_16 = W*in
   wire signed [9:0] m24_16;
   assign m24_16 =10'b0;

   // m24_17 = W*in
   wire signed [9:0] m24_17;
   assign m24_17 ={ {5{in24[5]}} , in24[5:1] };

   // m24_18 = W*in
   wire signed [9:0] m24_18;
   assign m24_18 =10'b0;

   // m24_19 = W*in
   wire signed [9:0] m24_19;
   assign m24_19 =10'b0;

   // m24_20 = W*in
   wire signed [9:0] m24_20;
   assign m24_20 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_21 = W*in
   wire signed [9:0] m24_21;
   assign m24_21 =10'b0;

   // m24_22 = W*in
   wire signed [9:0] m24_22;
   assign m24_22 =10'b0;

   // m24_23 = W*in
   wire signed [9:0] m24_23;
   assign m24_23 =10'b0;

   // m24_24 = W*in
   wire signed [9:0] m24_24;
   assign m24_24 =10'b0;

   // m24_25 = W*in
   wire signed [9:0] m24_25;
   assign m24_25 =10'b0;

   // m24_26 = W*in
   wire signed [9:0] m24_26;
   assign m24_26 =10'b0;

   // m24_27 = W*in
   wire signed [9:0] m24_27;
   assign m24_27 ={ {5{in24[5]}} , in24[5:1] };

   // m24_28 = W*in
   wire signed [9:0] m24_28;
   assign m24_28 =10'b0;

   // m24_29 = W*in
   wire signed [9:0] m24_29;
   assign m24_29 =10'b0;

   // m24_30 = W*in
   wire signed [9:0] m24_30;
   assign m24_30 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_31 = W*in
   wire signed [9:0] m24_31;
   assign m24_31 ={ {5{neg24[5]}} , neg24[5:1] };

   // m24_32 = W*in
   wire signed [9:0] m24_32;
   assign m24_32 =10'b0;

   // m24_33 = W*in
   wire signed [9:0] m24_33;
   assign m24_33 =10'b0;

   // m24_34 = W*in
   wire signed [9:0] m24_34;
   assign m24_34 =10'b0;

   // m24_35 = W*in
   wire signed [9:0] m24_35;
   assign m24_35 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_36 = W*in
   wire signed [9:0] m24_36;
   assign m24_36 =10'b0;

   // m24_37 = W*in
   wire signed [9:0] m24_37;
   assign m24_37 ={ {4{in24[5]}} , in24[5:0] };

   // m24_38 = W*in
   wire signed [9:0] m24_38;
   assign m24_38 =10'b0;

   // m24_39 = W*in
   wire signed [9:0] m24_39;
   assign m24_39 ={ {4{in24[5]}} , in24[5:0] };

   // m24_40 = W*in
   wire signed [9:0] m24_40;
   assign m24_40 =10'b0;

   // m24_41 = W*in
   wire signed [9:0] m24_41;
   assign m24_41 =10'b0;

   // m24_42 = W*in
   wire signed [9:0] m24_42;
   assign m24_42 =10'b0;

   // m24_43 = W*in
   wire signed [9:0] m24_43;
   assign m24_43 =10'b0;

   // m24_44 = W*in
   wire signed [9:0] m24_44;
   assign m24_44 =10'b0;

   // m24_45 = W*in
   wire signed [9:0] m24_45;
   assign m24_45 =10'b0;

   // m24_46 = W*in
   wire signed [9:0] m24_46;
   assign m24_46 ={ {4{in24[5]}} , in24[5:0] };

   // m24_47 = W*in
   wire signed [9:0] m24_47;
   assign m24_47 =10'b0;

   // m24_48 = W*in
   wire signed [9:0] m24_48;
   assign m24_48 =10'b0;

   // m24_49 = W*in
   wire signed [9:0] m24_49;
   assign m24_49 =10'b0;

   // m24_50 = W*in
   wire signed [9:0] m24_50;
   assign m24_50 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_51 = W*in
   wire signed [9:0] m24_51;
   assign m24_51 =10'b0;

   // m24_52 = W*in
   wire signed [9:0] m24_52;
   assign m24_52 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_53 = W*in
   wire signed [9:0] m24_53;
   assign m24_53 =10'b0;

   // m24_54 = W*in
   wire signed [9:0] m24_54;
   assign m24_54 =10'b0;

   // m24_55 = W*in
   wire signed [9:0] m24_55;
   assign m24_55 =10'b0;

   // m24_56 = W*in
   wire signed [9:0] m24_56;
   assign m24_56 ={ {4{in24[5]}} , in24[5:0] };

   // m24_57 = W*in
   wire signed [9:0] m24_57;
   assign m24_57 =10'b0;

   // m24_58 = W*in
   wire signed [9:0] m24_58;
   assign m24_58 =10'b0;

   // m24_59 = W*in
   wire signed [9:0] m24_59;
   assign m24_59 =10'b0;

   // m24_60 = W*in
   wire signed [9:0] m24_60;
   assign m24_60 =10'b0;

   // m24_61 = W*in
   wire signed [9:0] m24_61;
   assign m24_61 =10'b0;

   // m24_62 = W*in
   wire signed [9:0] m24_62;
   assign m24_62 =10'b0;

   // m24_63 = W*in
   wire signed [9:0] m24_63;
   assign m24_63 =10'b0;

   // m24_64 = W*in
   wire signed [9:0] m24_64;
   assign m24_64 ={ {5{neg24[5]}} , neg24[5:1] };

   // m24_65 = W*in
   wire signed [9:0] m24_65;
   assign m24_65 ={ {5{neg24[5]}} , neg24[5:1] };

   // m24_66 = W*in
   wire signed [9:0] m24_66;
   assign m24_66 =10'b0;

   // m24_67 = W*in
   wire signed [9:0] m24_67;
   assign m24_67 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_68 = W*in
   wire signed [9:0] m24_68;
   assign m24_68 ={ {5{neg24[5]}} , neg24[5:1] };

   // m24_69 = W*in
   wire signed [9:0] m24_69;
   assign m24_69 =10'b0;

   // m24_70 = W*in
   wire signed [9:0] m24_70;
   assign m24_70 ={ {5{neg24[5]}} , neg24[5:1] };

   // m24_71 = W*in
   wire signed [9:0] m24_71;
   assign m24_71 =10'b0;

   // m24_72 = W*in
   wire signed [9:0] m24_72;
   assign m24_72 =10'b0;

   // m24_73 = W*in
   wire signed [9:0] m24_73;
   assign m24_73 =10'b0;

   // m24_74 = W*in
   wire signed [9:0] m24_74;
   assign m24_74 =10'b0;

   // m24_75 = W*in
   wire signed [9:0] m24_75;
   assign m24_75 =10'b0;

   // m24_76 = W*in
   wire signed [9:0] m24_76;
   assign m24_76 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_77 = W*in
   wire signed [9:0] m24_77;
   assign m24_77 =10'b0;

   // m24_78 = W*in
   wire signed [9:0] m24_78;
   assign m24_78 =10'b0;

   // m24_79 = W*in
   wire signed [9:0] m24_79;
   assign m24_79 =10'b0;

   // m24_80 = W*in
   wire signed [9:0] m24_80;
   assign m24_80 =10'b0;

   // m24_81 = W*in
   wire signed [9:0] m24_81;
   assign m24_81 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_82 = W*in
   wire signed [9:0] m24_82;
   assign m24_82 =10'b0;

   // m24_83 = W*in
   wire signed [9:0] m24_83;
   assign m24_83 ={ {4{in24[5]}} , in24[5:0] };

   // m24_84 = W*in
   wire signed [9:0] m24_84;
   assign m24_84 =10'b0;

   // m24_85 = W*in
   wire signed [9:0] m24_85;
   assign m24_85 ={ {4{in24[5]}} , in24[5:0] };

   // m24_86 = W*in
   wire signed [9:0] m24_86;
   assign m24_86 =10'b0;

   // m24_87 = W*in
   wire signed [9:0] m24_87;
   assign m24_87 =10'b0;

   // m24_88 = W*in
   wire signed [9:0] m24_88;
   assign m24_88 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_89 = W*in
   wire signed [9:0] m24_89;
   assign m24_89 =10'b0;

   // m24_90 = W*in
   wire signed [9:0] m24_90;
   assign m24_90 =10'b0;

   // m24_91 = W*in
   wire signed [9:0] m24_91;
   assign m24_91 =10'b0;

   // m24_92 = W*in
   wire signed [9:0] m24_92;
   assign m24_92 =10'b0;

   // m24_93 = W*in
   wire signed [9:0] m24_93;
   assign m24_93 =10'b0;

   // m24_94 = W*in
   wire signed [9:0] m24_94;
   assign m24_94 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_95 = W*in
   wire signed [9:0] m24_95;
   assign m24_95 ={ {4{in24[5]}} , in24[5:0] };

   // m24_96 = W*in
   wire signed [9:0] m24_96;
   assign m24_96 =10'b0;

   // m24_97 = W*in
   wire signed [9:0] m24_97;
   assign m24_97 =10'b0;

   // m24_98 = W*in
   wire signed [9:0] m24_98;
   assign m24_98 =10'b0;

   // m24_99 = W*in
   wire signed [9:0] m24_99;
   assign m24_99 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_100 = W*in
   wire signed [9:0] m24_100;
   assign m24_100 =10'b0;

   // m24_101 = W*in
   wire signed [9:0] m24_101;
   assign m24_101 ={ {4{in24[5]}} , in24[5:0] };

   // m24_102 = W*in
   wire signed [9:0] m24_102;
   assign m24_102 =10'b0;

   // m24_103 = W*in
   wire signed [9:0] m24_103;
   assign m24_103 =10'b0;

   // m24_104 = W*in
   wire signed [9:0] m24_104;
   assign m24_104 ={ {4{in24[5]}} , in24[5:0] };

   // m24_105 = W*in
   wire signed [9:0] m24_105;
   assign m24_105 =10'b0;

   // m24_106 = W*in
   wire signed [9:0] m24_106;
   assign m24_106 =10'b0;

   // m24_107 = W*in
   wire signed [9:0] m24_107;
   assign m24_107 ={ {4{in24[5]}} , in24[5:0] };

   // m24_108 = W*in
   wire signed [9:0] m24_108;
   assign m24_108 ={ {4{neg24[5]}} , neg24[5:0] };

   // m24_109 = W*in
   wire signed [9:0] m24_109;
   assign m24_109 =10'b0;

   // m24_110 = W*in
   wire signed [9:0] m24_110;
   assign m24_110 =10'b0;

   // m24_111 = W*in
   wire signed [9:0] m24_111;
   assign m24_111 =10'b0;

   // m24_112 = W*in
   wire signed [9:0] m24_112;
   assign m24_112 =10'b0;

   // m24_113 = W*in
   wire signed [9:0] m24_113;
   assign m24_113 =10'b0;

   // m24_114 = W*in
   wire signed [9:0] m24_114;
   assign m24_114 =10'b0;

   // m24_115 = W*in
   wire signed [9:0] m24_115;
   assign m24_115 =10'b0;

   // m24_116 = W*in
   wire signed [9:0] m24_116;
   assign m24_116 =10'b0;

   // m24_117 = W*in
   wire signed [9:0] m24_117;
   assign m24_117 ={ {4{neg24[5]}} , neg24[5:0] };

   // m25_1 = W*in
   wire signed [9:0] m25_1;
   assign m25_1 =10'b0;

   // m25_2 = W*in
   wire signed [9:0] m25_2;
   assign m25_2 =10'b0;

   // m25_3 = W*in
   wire signed [9:0] m25_3;
   assign m25_3 =10'b0;

   // m25_4 = W*in
   wire signed [9:0] m25_4;
   assign m25_4 =10'b0;

   // m25_5 = W*in
   wire signed [9:0] m25_5;
   assign m25_5 =10'b0;

   // m25_6 = W*in
   wire signed [9:0] m25_6;
   assign m25_6 =10'b0;

   // m25_7 = W*in
   wire signed [9:0] m25_7;
   assign m25_7 =10'b0;

   // m25_8 = W*in
   wire signed [9:0] m25_8;
   assign m25_8 ={ {4{neg25[5]}} , neg25[5:0] };

   // m25_9 = W*in
   wire signed [9:0] m25_9;
   assign m25_9 =10'b0;

   // m25_10 = W*in
   wire signed [9:0] m25_10;
   assign m25_10 =10'b0;

   // m25_11 = W*in
   wire signed [9:0] m25_11;
   assign m25_11 =10'b0;

   // m25_12 = W*in
   wire signed [9:0] m25_12;
   assign m25_12 =10'b0;

   // m25_13 = W*in
   wire signed [9:0] m25_13;
   assign m25_13 =10'b0;

   // m25_14 = W*in
   wire signed [9:0] m25_14;
   assign m25_14 ={ {4{neg25[5]}} , neg25[5:0] };

   // m25_15 = W*in
   wire signed [9:0] m25_15;
   assign m25_15 =10'b0;

   // m25_16 = W*in
   wire signed [9:0] m25_16;
   assign m25_16 =10'b0;

   // m25_17 = W*in
   wire signed [9:0] m25_17;
   assign m25_17 ={ {5{in25[5]}} , in25[5:1] };

   // m25_18 = W*in
   wire signed [9:0] m25_18;
   assign m25_18 =10'b0;

   // m25_19 = W*in
   wire signed [9:0] m25_19;
   assign m25_19 =10'b0;

   // m25_20 = W*in
   wire signed [9:0] m25_20;
   assign m25_20 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_21 = W*in
   wire signed [9:0] m25_21;
   assign m25_21 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_22 = W*in
   wire signed [9:0] m25_22;
   assign m25_22 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_23 = W*in
   wire signed [9:0] m25_23;
   assign m25_23 =10'b0;

   // m25_24 = W*in
   wire signed [9:0] m25_24;
   assign m25_24 =10'b0;

   // m25_25 = W*in
   wire signed [9:0] m25_25;
   assign m25_25 =10'b0;

   // m25_26 = W*in
   wire signed [9:0] m25_26;
   assign m25_26 =10'b0;

   // m25_27 = W*in
   wire signed [9:0] m25_27;
   assign m25_27 ={ {5{in25[5]}} , in25[5:1] };

   // m25_28 = W*in
   wire signed [9:0] m25_28;
   assign m25_28 =10'b0;

   // m25_29 = W*in
   wire signed [9:0] m25_29;
   assign m25_29 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_30 = W*in
   wire signed [9:0] m25_30;
   assign m25_30 =10'b0;

   // m25_31 = W*in
   wire signed [9:0] m25_31;
   assign m25_31 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_32 = W*in
   wire signed [9:0] m25_32;
   assign m25_32 =10'b0;

   // m25_33 = W*in
   wire signed [9:0] m25_33;
   assign m25_33 =10'b0;

   // m25_34 = W*in
   wire signed [9:0] m25_34;
   assign m25_34 =10'b0;

   // m25_35 = W*in
   wire signed [9:0] m25_35;
   assign m25_35 =10'b0;

   // m25_36 = W*in
   wire signed [9:0] m25_36;
   assign m25_36 =10'b0;

   // m25_37 = W*in
   wire signed [9:0] m25_37;
   assign m25_37 =10'b0;

   // m25_38 = W*in
   wire signed [9:0] m25_38;
   assign m25_38 =10'b0;

   // m25_39 = W*in
   wire signed [9:0] m25_39;
   assign m25_39 =10'b0;

   // m25_40 = W*in
   wire signed [9:0] m25_40;
   assign m25_40 =10'b0;

   // m25_41 = W*in
   wire signed [9:0] m25_41;
   assign m25_41 =10'b0;

   // m25_42 = W*in
   wire signed [9:0] m25_42;
   assign m25_42 =10'b0;

   // m25_43 = W*in
   wire signed [9:0] m25_43;
   assign m25_43 =10'b0;

   // m25_44 = W*in
   wire signed [9:0] m25_44;
   assign m25_44 =10'b0;

   // m25_45 = W*in
   wire signed [9:0] m25_45;
   assign m25_45 =10'b0;

   // m25_46 = W*in
   wire signed [9:0] m25_46;
   assign m25_46 =10'b0;

   // m25_47 = W*in
   wire signed [9:0] m25_47;
   assign m25_47 =10'b0;

   // m25_48 = W*in
   wire signed [9:0] m25_48;
   assign m25_48 =10'b0;

   // m25_49 = W*in
   wire signed [9:0] m25_49;
   assign m25_49 =10'b0;

   // m25_50 = W*in
   wire signed [9:0] m25_50;
   assign m25_50 ={ {4{neg25[5]}} , neg25[5:0] };

   // m25_51 = W*in
   wire signed [9:0] m25_51;
   assign m25_51 =10'b0;

   // m25_52 = W*in
   wire signed [9:0] m25_52;
   assign m25_52 =10'b0;

   // m25_53 = W*in
   wire signed [9:0] m25_53;
   assign m25_53 =10'b0;

   // m25_54 = W*in
   wire signed [9:0] m25_54;
   assign m25_54 =10'b0;

   // m25_55 = W*in
   wire signed [9:0] m25_55;
   assign m25_55 =10'b0;

   // m25_56 = W*in
   wire signed [9:0] m25_56;
   assign m25_56 =10'b0;

   // m25_57 = W*in
   wire signed [9:0] m25_57;
   assign m25_57 =10'b0;

   // m25_58 = W*in
   wire signed [9:0] m25_58;
   assign m25_58 =10'b0;

   // m25_59 = W*in
   wire signed [9:0] m25_59;
   assign m25_59 =10'b0;

   // m25_60 = W*in
   wire signed [9:0] m25_60;
   assign m25_60 =10'b0;

   // m25_61 = W*in
   wire signed [9:0] m25_61;
   assign m25_61 ={ {4{in25[5]}} , in25[5:0] };

   // m25_62 = W*in
   wire signed [9:0] m25_62;
   assign m25_62 =10'b0;

   // m25_63 = W*in
   wire signed [9:0] m25_63;
   assign m25_63 =10'b0;

   // m25_64 = W*in
   wire signed [9:0] m25_64;
   assign m25_64 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_65 = W*in
   wire signed [9:0] m25_65;
   assign m25_65 ={ {4{neg25[5]}} , neg25[5:0] };

   // m25_66 = W*in
   wire signed [9:0] m25_66;
   assign m25_66 =10'b0;

   // m25_67 = W*in
   wire signed [9:0] m25_67;
   assign m25_67 ={ {4{neg25[5]}} , neg25[5:0] };

   // m25_68 = W*in
   wire signed [9:0] m25_68;
   assign m25_68 =10'b0;

   // m25_69 = W*in
   wire signed [9:0] m25_69;
   assign m25_69 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_70 = W*in
   wire signed [9:0] m25_70;
   assign m25_70 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_71 = W*in
   wire signed [9:0] m25_71;
   assign m25_71 ={ {5{in25[5]}} , in25[5:1] };

   // m25_72 = W*in
   wire signed [9:0] m25_72;
   assign m25_72 =10'b0;

   // m25_73 = W*in
   wire signed [9:0] m25_73;
   assign m25_73 =10'b0;

   // m25_74 = W*in
   wire signed [9:0] m25_74;
   assign m25_74 =10'b0;

   // m25_75 = W*in
   wire signed [9:0] m25_75;
   assign m25_75 =10'b0;

   // m25_76 = W*in
   wire signed [9:0] m25_76;
   assign m25_76 =10'b0;

   // m25_77 = W*in
   wire signed [9:0] m25_77;
   assign m25_77 =10'b0;

   // m25_78 = W*in
   wire signed [9:0] m25_78;
   assign m25_78 =10'b0;

   // m25_79 = W*in
   wire signed [9:0] m25_79;
   assign m25_79 =10'b0;

   // m25_80 = W*in
   wire signed [9:0] m25_80;
   assign m25_80 =10'b0;

   // m25_81 = W*in
   wire signed [9:0] m25_81;
   assign m25_81 ={ {4{neg25[5]}} , neg25[5:0] };

   // m25_82 = W*in
   wire signed [9:0] m25_82;
   assign m25_82 ={ {5{neg25[5]}} , neg25[5:1] };

   // m25_83 = W*in
   wire signed [9:0] m25_83;
   assign m25_83 ={ {4{in25[5]}} , in25[5:0] };

   // m25_84 = W*in
   wire signed [9:0] m25_84;
   assign m25_84 =10'b0;

   // m25_85 = W*in
   wire signed [9:0] m25_85;
   assign m25_85 =10'b0;

   // m25_86 = W*in
   wire signed [9:0] m25_86;
   assign m25_86 =10'b0;

   // m25_87 = W*in
   wire signed [9:0] m25_87;
   assign m25_87 =10'b0;

   // m25_88 = W*in
   wire signed [9:0] m25_88;
   assign m25_88 =10'b0;

   // m25_89 = W*in
   wire signed [9:0] m25_89;
   assign m25_89 =10'b0;

   // m25_90 = W*in
   wire signed [9:0] m25_90;
   assign m25_90 =10'b0;

   // m25_91 = W*in
   wire signed [9:0] m25_91;
   assign m25_91 =10'b0;

   // m25_92 = W*in
   wire signed [9:0] m25_92;
   assign m25_92 =10'b0;

   // m25_93 = W*in
   wire signed [9:0] m25_93;
   assign m25_93 =10'b0;

   // m25_94 = W*in
   wire signed [9:0] m25_94;
   assign m25_94 =10'b0;

   // m25_95 = W*in
   wire signed [9:0] m25_95;
   assign m25_95 ={ {4{in25[5]}} , in25[5:0] };

   // m25_96 = W*in
   wire signed [9:0] m25_96;
   assign m25_96 =10'b0;

   // m25_97 = W*in
   wire signed [9:0] m25_97;
   assign m25_97 =10'b0;

   // m25_98 = W*in
   wire signed [9:0] m25_98;
   assign m25_98 =10'b0;

   // m25_99 = W*in
   wire signed [9:0] m25_99;
   assign m25_99 =10'b0;

   // m25_100 = W*in
   wire signed [9:0] m25_100;
   assign m25_100 =10'b0;

   // m25_101 = W*in
   wire signed [9:0] m25_101;
   assign m25_101 =10'b0;

   // m25_102 = W*in
   wire signed [9:0] m25_102;
   assign m25_102 =10'b0;

   // m25_103 = W*in
   wire signed [9:0] m25_103;
   assign m25_103 ={ {4{in25[5]}} , in25[5:0] };

   // m25_104 = W*in
   wire signed [9:0] m25_104;
   assign m25_104 ={ {4{in25[5]}} , in25[5:0] };

   // m25_105 = W*in
   wire signed [9:0] m25_105;
   assign m25_105 =10'b0;

   // m25_106 = W*in
   wire signed [9:0] m25_106;
   assign m25_106 =10'b0;

   // m25_107 = W*in
   wire signed [9:0] m25_107;
   assign m25_107 ={ {4{in25[5]}} , in25[5:0] };

   // m25_108 = W*in
   wire signed [9:0] m25_108;
   assign m25_108 =10'b0;

   // m25_109 = W*in
   wire signed [9:0] m25_109;
   assign m25_109 =10'b0;

   // m25_110 = W*in
   wire signed [9:0] m25_110;
   assign m25_110 =10'b0;

   // m25_111 = W*in
   wire signed [9:0] m25_111;
   assign m25_111 =10'b0;

   // m25_112 = W*in
   wire signed [9:0] m25_112;
   assign m25_112 =10'b0;

   // m25_113 = W*in
   wire signed [9:0] m25_113;
   assign m25_113 =10'b0;

   // m25_114 = W*in
   wire signed [9:0] m25_114;
   assign m25_114 =10'b0;

   // m25_115 = W*in
   wire signed [9:0] m25_115;
   assign m25_115 =10'b0;

   // m25_116 = W*in
   wire signed [9:0] m25_116;
   assign m25_116 =10'b0;

   // m25_117 = W*in
   wire signed [9:0] m25_117;
   assign m25_117 =10'b0;

   // m26_1 = W*in
   wire signed [9:0] m26_1;
   assign m26_1 =10'b0;

   // m26_2 = W*in
   wire signed [9:0] m26_2;
   assign m26_2 =10'b0;

   // m26_3 = W*in
   wire signed [9:0] m26_3;
   assign m26_3 =10'b0;

   // m26_4 = W*in
   wire signed [9:0] m26_4;
   assign m26_4 =10'b0;

   // m26_5 = W*in
   wire signed [9:0] m26_5;
   assign m26_5 =10'b0;

   // m26_6 = W*in
   wire signed [9:0] m26_6;
   assign m26_6 =10'b0;

   // m26_7 = W*in
   wire signed [9:0] m26_7;
   assign m26_7 =10'b0;

   // m26_8 = W*in
   wire signed [9:0] m26_8;
   assign m26_8 =10'b0;

   // m26_9 = W*in
   wire signed [9:0] m26_9;
   assign m26_9 =10'b0;

   // m26_10 = W*in
   wire signed [9:0] m26_10;
   assign m26_10 =10'b0;

   // m26_11 = W*in
   wire signed [9:0] m26_11;
   assign m26_11 =10'b0;

   // m26_12 = W*in
   wire signed [9:0] m26_12;
   assign m26_12 =10'b0;

   // m26_13 = W*in
   wire signed [9:0] m26_13;
   assign m26_13 =10'b0;

   // m26_14 = W*in
   wire signed [9:0] m26_14;
   assign m26_14 =10'b0;

   // m26_15 = W*in
   wire signed [9:0] m26_15;
   assign m26_15 =10'b0;

   // m26_16 = W*in
   wire signed [9:0] m26_16;
   assign m26_16 =10'b0;

   // m26_17 = W*in
   wire signed [9:0] m26_17;
   assign m26_17 =10'b0;

   // m26_18 = W*in
   wire signed [9:0] m26_18;
   assign m26_18 =10'b0;

   // m26_19 = W*in
   wire signed [9:0] m26_19;
   assign m26_19 =10'b0;

   // m26_20 = W*in
   wire signed [9:0] m26_20;
   assign m26_20 ={ {5{in26[5]}} , in26[5:1] };

   // m26_21 = W*in
   wire signed [9:0] m26_21;
   assign m26_21 =10'b0;

   // m26_22 = W*in
   wire signed [9:0] m26_22;
   assign m26_22 =10'b0;

   // m26_23 = W*in
   wire signed [9:0] m26_23;
   assign m26_23 =10'b0;

   // m26_24 = W*in
   wire signed [9:0] m26_24;
   assign m26_24 =10'b0;

   // m26_25 = W*in
   wire signed [9:0] m26_25;
   assign m26_25 =10'b0;

   // m26_26 = W*in
   wire signed [9:0] m26_26;
   assign m26_26 =10'b0;

   // m26_27 = W*in
   wire signed [9:0] m26_27;
   assign m26_27 =10'b0;

   // m26_28 = W*in
   wire signed [9:0] m26_28;
   assign m26_28 =10'b0;

   // m26_29 = W*in
   wire signed [9:0] m26_29;
   assign m26_29 =10'b0;

   // m26_30 = W*in
   wire signed [9:0] m26_30;
   assign m26_30 =10'b0;

   // m26_31 = W*in
   wire signed [9:0] m26_31;
   assign m26_31 =10'b0;

   // m26_32 = W*in
   wire signed [9:0] m26_32;
   assign m26_32 =10'b0;

   // m26_33 = W*in
   wire signed [9:0] m26_33;
   assign m26_33 =10'b0;

   // m26_34 = W*in
   wire signed [9:0] m26_34;
   assign m26_34 =10'b0;

   // m26_35 = W*in
   wire signed [9:0] m26_35;
   assign m26_35 =10'b0;

   // m26_36 = W*in
   wire signed [9:0] m26_36;
   assign m26_36 =10'b0;

   // m26_37 = W*in
   wire signed [9:0] m26_37;
   assign m26_37 =10'b0;

   // m26_38 = W*in
   wire signed [9:0] m26_38;
   assign m26_38 =10'b0;

   // m26_39 = W*in
   wire signed [9:0] m26_39;
   assign m26_39 =10'b0;

   // m26_40 = W*in
   wire signed [9:0] m26_40;
   assign m26_40 =10'b0;

   // m26_41 = W*in
   wire signed [9:0] m26_41;
   assign m26_41 =10'b0;

   // m26_42 = W*in
   wire signed [9:0] m26_42;
   assign m26_42 =10'b0;

   // m26_43 = W*in
   wire signed [9:0] m26_43;
   assign m26_43 =10'b0;

   // m26_44 = W*in
   wire signed [9:0] m26_44;
   assign m26_44 =10'b0;

   // m26_45 = W*in
   wire signed [9:0] m26_45;
   assign m26_45 =10'b0;

   // m26_46 = W*in
   wire signed [9:0] m26_46;
   assign m26_46 =10'b0;

   // m26_47 = W*in
   wire signed [9:0] m26_47;
   assign m26_47 =10'b0;

   // m26_48 = W*in
   wire signed [9:0] m26_48;
   assign m26_48 =10'b0;

   // m26_49 = W*in
   wire signed [9:0] m26_49;
   assign m26_49 =10'b0;

   // m26_50 = W*in
   wire signed [9:0] m26_50;
   assign m26_50 =10'b0;

   // m26_51 = W*in
   wire signed [9:0] m26_51;
   assign m26_51 =10'b0;

   // m26_52 = W*in
   wire signed [9:0] m26_52;
   assign m26_52 =10'b0;

   // m26_53 = W*in
   wire signed [9:0] m26_53;
   assign m26_53 =10'b0;

   // m26_54 = W*in
   wire signed [9:0] m26_54;
   assign m26_54 =10'b0;

   // m26_55 = W*in
   wire signed [9:0] m26_55;
   assign m26_55 =10'b0;

   // m26_56 = W*in
   wire signed [9:0] m26_56;
   assign m26_56 =10'b0;

   // m26_57 = W*in
   wire signed [9:0] m26_57;
   assign m26_57 =10'b0;

   // m26_58 = W*in
   wire signed [9:0] m26_58;
   assign m26_58 =10'b0;

   // m26_59 = W*in
   wire signed [9:0] m26_59;
   assign m26_59 =10'b0;

   // m26_60 = W*in
   wire signed [9:0] m26_60;
   assign m26_60 =10'b0;

   // m26_61 = W*in
   wire signed [9:0] m26_61;
   assign m26_61 =10'b0;

   // m26_62 = W*in
   wire signed [9:0] m26_62;
   assign m26_62 =10'b0;

   // m26_63 = W*in
   wire signed [9:0] m26_63;
   assign m26_63 =10'b0;

   // m26_64 = W*in
   wire signed [9:0] m26_64;
   assign m26_64 =10'b0;

   // m26_65 = W*in
   wire signed [9:0] m26_65;
   assign m26_65 =10'b0;

   // m26_66 = W*in
   wire signed [9:0] m26_66;
   assign m26_66 =10'b0;

   // m26_67 = W*in
   wire signed [9:0] m26_67;
   assign m26_67 =10'b0;

   // m26_68 = W*in
   wire signed [9:0] m26_68;
   assign m26_68 =10'b0;

   // m26_69 = W*in
   wire signed [9:0] m26_69;
   assign m26_69 =10'b0;

   // m26_70 = W*in
   wire signed [9:0] m26_70;
   assign m26_70 =10'b0;

   // m26_71 = W*in
   wire signed [9:0] m26_71;
   assign m26_71 =10'b0;

   // m26_72 = W*in
   wire signed [9:0] m26_72;
   assign m26_72 =10'b0;

   // m26_73 = W*in
   wire signed [9:0] m26_73;
   assign m26_73 =10'b0;

   // m26_74 = W*in
   wire signed [9:0] m26_74;
   assign m26_74 =10'b0;

   // m26_75 = W*in
   wire signed [9:0] m26_75;
   assign m26_75 =10'b0;

   // m26_76 = W*in
   wire signed [9:0] m26_76;
   assign m26_76 =10'b0;

   // m26_77 = W*in
   wire signed [9:0] m26_77;
   assign m26_77 =10'b0;

   // m26_78 = W*in
   wire signed [9:0] m26_78;
   assign m26_78 =10'b0;

   // m26_79 = W*in
   wire signed [9:0] m26_79;
   assign m26_79 =10'b0;

   // m26_80 = W*in
   wire signed [9:0] m26_80;
   assign m26_80 =10'b0;

   // m26_81 = W*in
   wire signed [9:0] m26_81;
   assign m26_81 =10'b0;

   // m26_82 = W*in
   wire signed [9:0] m26_82;
   assign m26_82 =10'b0;

   // m26_83 = W*in
   wire signed [9:0] m26_83;
   assign m26_83 =10'b0;

   // m26_84 = W*in
   wire signed [9:0] m26_84;
   assign m26_84 =10'b0;

   // m26_85 = W*in
   wire signed [9:0] m26_85;
   assign m26_85 =10'b0;

   // m26_86 = W*in
   wire signed [9:0] m26_86;
   assign m26_86 =10'b0;

   // m26_87 = W*in
   wire signed [9:0] m26_87;
   assign m26_87 =10'b0;

   // m26_88 = W*in
   wire signed [9:0] m26_88;
   assign m26_88 =10'b0;

   // m26_89 = W*in
   wire signed [9:0] m26_89;
   assign m26_89 =10'b0;

   // m26_90 = W*in
   wire signed [9:0] m26_90;
   assign m26_90 =10'b0;

   // m26_91 = W*in
   wire signed [9:0] m26_91;
   assign m26_91 =10'b0;

   // m26_92 = W*in
   wire signed [9:0] m26_92;
   assign m26_92 =10'b0;

   // m26_93 = W*in
   wire signed [9:0] m26_93;
   assign m26_93 =10'b0;

   // m26_94 = W*in
   wire signed [9:0] m26_94;
   assign m26_94 =10'b0;

   // m26_95 = W*in
   wire signed [9:0] m26_95;
   assign m26_95 =10'b0;

   // m26_96 = W*in
   wire signed [9:0] m26_96;
   assign m26_96 =10'b0;

   // m26_97 = W*in
   wire signed [9:0] m26_97;
   assign m26_97 =10'b0;

   // m26_98 = W*in
   wire signed [9:0] m26_98;
   assign m26_98 =10'b0;

   // m26_99 = W*in
   wire signed [9:0] m26_99;
   assign m26_99 =10'b0;

   // m26_100 = W*in
   wire signed [9:0] m26_100;
   assign m26_100 =10'b0;

   // m26_101 = W*in
   wire signed [9:0] m26_101;
   assign m26_101 =10'b0;

   // m26_102 = W*in
   wire signed [9:0] m26_102;
   assign m26_102 =10'b0;

   // m26_103 = W*in
   wire signed [9:0] m26_103;
   assign m26_103 =10'b0;

   // m26_104 = W*in
   wire signed [9:0] m26_104;
   assign m26_104 =10'b0;

   // m26_105 = W*in
   wire signed [9:0] m26_105;
   assign m26_105 =10'b0;

   // m26_106 = W*in
   wire signed [9:0] m26_106;
   assign m26_106 =10'b0;

   // m26_107 = W*in
   wire signed [9:0] m26_107;
   assign m26_107 =10'b0;

   // m26_108 = W*in
   wire signed [9:0] m26_108;
   assign m26_108 ={ {5{in26[5]}} , in26[5:1] };

   // m26_109 = W*in
   wire signed [9:0] m26_109;
   assign m26_109 =10'b0;

   // m26_110 = W*in
   wire signed [9:0] m26_110;
   assign m26_110 =10'b0;

   // m26_111 = W*in
   wire signed [9:0] m26_111;
   assign m26_111 =10'b0;

   // m26_112 = W*in
   wire signed [9:0] m26_112;
   assign m26_112 =10'b0;

   // m26_113 = W*in
   wire signed [9:0] m26_113;
   assign m26_113 =10'b0;

   // m26_114 = W*in
   wire signed [9:0] m26_114;
   assign m26_114 =10'b0;

   // m26_115 = W*in
   wire signed [9:0] m26_115;
   assign m26_115 =10'b0;

   // m26_116 = W*in
   wire signed [9:0] m26_116;
   assign m26_116 ={ {5{in26[5]}} , in26[5:1] };

   // m26_117 = W*in
   wire signed [9:0] m26_117;
   assign m26_117 =10'b0;

   // m27_1 = W*in
   wire signed [9:0] m27_1;
   assign m27_1 =10'b0;

   // m27_2 = W*in
   wire signed [9:0] m27_2;
   assign m27_2 =10'b0;

   // m27_3 = W*in
   wire signed [9:0] m27_3;
   assign m27_3 =10'b0;

   // m27_4 = W*in
   wire signed [9:0] m27_4;
   assign m27_4 =10'b0;

   // m27_5 = W*in
   wire signed [9:0] m27_5;
   assign m27_5 =10'b0;

   // m27_6 = W*in
   wire signed [9:0] m27_6;
   assign m27_6 =10'b0;

   // m27_7 = W*in
   wire signed [9:0] m27_7;
   assign m27_7 =10'b0;

   // m27_8 = W*in
   wire signed [9:0] m27_8;
   assign m27_8 =10'b0;

   // m27_9 = W*in
   wire signed [9:0] m27_9;
   assign m27_9 =10'b0;

   // m27_10 = W*in
   wire signed [9:0] m27_10;
   assign m27_10 =10'b0;

   // m27_11 = W*in
   wire signed [9:0] m27_11;
   assign m27_11 =10'b0;

   // m27_12 = W*in
   wire signed [9:0] m27_12;
   assign m27_12 =10'b0;

   // m27_13 = W*in
   wire signed [9:0] m27_13;
   assign m27_13 =10'b0;

   // m27_14 = W*in
   wire signed [9:0] m27_14;
   assign m27_14 =10'b0;

   // m27_15 = W*in
   wire signed [9:0] m27_15;
   assign m27_15 =10'b0;

   // m27_16 = W*in
   wire signed [9:0] m27_16;
   assign m27_16 =10'b0;

   // m27_17 = W*in
   wire signed [9:0] m27_17;
   assign m27_17 =10'b0;

   // m27_18 = W*in
   wire signed [9:0] m27_18;
   assign m27_18 =10'b0;

   // m27_19 = W*in
   wire signed [9:0] m27_19;
   assign m27_19 =10'b0;

   // m27_20 = W*in
   wire signed [9:0] m27_20;
   assign m27_20 =10'b0;

   // m27_21 = W*in
   wire signed [9:0] m27_21;
   assign m27_21 =10'b0;

   // m27_22 = W*in
   wire signed [9:0] m27_22;
   assign m27_22 =10'b0;

   // m27_23 = W*in
   wire signed [9:0] m27_23;
   assign m27_23 =10'b0;

   // m27_24 = W*in
   wire signed [9:0] m27_24;
   assign m27_24 =10'b0;

   // m27_25 = W*in
   wire signed [9:0] m27_25;
   assign m27_25 =10'b0;

   // m27_26 = W*in
   wire signed [9:0] m27_26;
   assign m27_26 =10'b0;

   // m27_27 = W*in
   wire signed [9:0] m27_27;
   assign m27_27 =10'b0;

   // m27_28 = W*in
   wire signed [9:0] m27_28;
   assign m27_28 =10'b0;

   // m27_29 = W*in
   wire signed [9:0] m27_29;
   assign m27_29 ={ {5{in27[5]}} , in27[5:1] };

   // m27_30 = W*in
   wire signed [9:0] m27_30;
   assign m27_30 =10'b0;

   // m27_31 = W*in
   wire signed [9:0] m27_31;
   assign m27_31 =10'b0;

   // m27_32 = W*in
   wire signed [9:0] m27_32;
   assign m27_32 =10'b0;

   // m27_33 = W*in
   wire signed [9:0] m27_33;
   assign m27_33 =10'b0;

   // m27_34 = W*in
   wire signed [9:0] m27_34;
   assign m27_34 =10'b0;

   // m27_35 = W*in
   wire signed [9:0] m27_35;
   assign m27_35 =10'b0;

   // m27_36 = W*in
   wire signed [9:0] m27_36;
   assign m27_36 =10'b0;

   // m27_37 = W*in
   wire signed [9:0] m27_37;
   assign m27_37 =10'b0;

   // m27_38 = W*in
   wire signed [9:0] m27_38;
   assign m27_38 =10'b0;

   // m27_39 = W*in
   wire signed [9:0] m27_39;
   assign m27_39 =10'b0;

   // m27_40 = W*in
   wire signed [9:0] m27_40;
   assign m27_40 =10'b0;

   // m27_41 = W*in
   wire signed [9:0] m27_41;
   assign m27_41 =10'b0;

   // m27_42 = W*in
   wire signed [9:0] m27_42;
   assign m27_42 =10'b0;

   // m27_43 = W*in
   wire signed [9:0] m27_43;
   assign m27_43 =10'b0;

   // m27_44 = W*in
   wire signed [9:0] m27_44;
   assign m27_44 =10'b0;

   // m27_45 = W*in
   wire signed [9:0] m27_45;
   assign m27_45 =10'b0;

   // m27_46 = W*in
   wire signed [9:0] m27_46;
   assign m27_46 =10'b0;

   // m27_47 = W*in
   wire signed [9:0] m27_47;
   assign m27_47 =10'b0;

   // m27_48 = W*in
   wire signed [9:0] m27_48;
   assign m27_48 =10'b0;

   // m27_49 = W*in
   wire signed [9:0] m27_49;
   assign m27_49 =10'b0;

   // m27_50 = W*in
   wire signed [9:0] m27_50;
   assign m27_50 =10'b0;

   // m27_51 = W*in
   wire signed [9:0] m27_51;
   assign m27_51 =10'b0;

   // m27_52 = W*in
   wire signed [9:0] m27_52;
   assign m27_52 =10'b0;

   // m27_53 = W*in
   wire signed [9:0] m27_53;
   assign m27_53 =10'b0;

   // m27_54 = W*in
   wire signed [9:0] m27_54;
   assign m27_54 =10'b0;

   // m27_55 = W*in
   wire signed [9:0] m27_55;
   assign m27_55 =10'b0;

   // m27_56 = W*in
   wire signed [9:0] m27_56;
   assign m27_56 =10'b0;

   // m27_57 = W*in
   wire signed [9:0] m27_57;
   assign m27_57 =10'b0;

   // m27_58 = W*in
   wire signed [9:0] m27_58;
   assign m27_58 =10'b0;

   // m27_59 = W*in
   wire signed [9:0] m27_59;
   assign m27_59 =10'b0;

   // m27_60 = W*in
   wire signed [9:0] m27_60;
   assign m27_60 =10'b0;

   // m27_61 = W*in
   wire signed [9:0] m27_61;
   assign m27_61 =10'b0;

   // m27_62 = W*in
   wire signed [9:0] m27_62;
   assign m27_62 =10'b0;

   // m27_63 = W*in
   wire signed [9:0] m27_63;
   assign m27_63 =10'b0;

   // m27_64 = W*in
   wire signed [9:0] m27_64;
   assign m27_64 =10'b0;

   // m27_65 = W*in
   wire signed [9:0] m27_65;
   assign m27_65 =10'b0;

   // m27_66 = W*in
   wire signed [9:0] m27_66;
   assign m27_66 =10'b0;

   // m27_67 = W*in
   wire signed [9:0] m27_67;
   assign m27_67 =10'b0;

   // m27_68 = W*in
   wire signed [9:0] m27_68;
   assign m27_68 =10'b0;

   // m27_69 = W*in
   wire signed [9:0] m27_69;
   assign m27_69 =10'b0;

   // m27_70 = W*in
   wire signed [9:0] m27_70;
   assign m27_70 ={ {5{in27[5]}} , in27[5:1] };

   // m27_71 = W*in
   wire signed [9:0] m27_71;
   assign m27_71 =10'b0;

   // m27_72 = W*in
   wire signed [9:0] m27_72;
   assign m27_72 =10'b0;

   // m27_73 = W*in
   wire signed [9:0] m27_73;
   assign m27_73 =10'b0;

   // m27_74 = W*in
   wire signed [9:0] m27_74;
   assign m27_74 =10'b0;

   // m27_75 = W*in
   wire signed [9:0] m27_75;
   assign m27_75 =10'b0;

   // m27_76 = W*in
   wire signed [9:0] m27_76;
   assign m27_76 =10'b0;

   // m27_77 = W*in
   wire signed [9:0] m27_77;
   assign m27_77 =10'b0;

   // m27_78 = W*in
   wire signed [9:0] m27_78;
   assign m27_78 =10'b0;

   // m27_79 = W*in
   wire signed [9:0] m27_79;
   assign m27_79 =10'b0;

   // m27_80 = W*in
   wire signed [9:0] m27_80;
   assign m27_80 =10'b0;

   // m27_81 = W*in
   wire signed [9:0] m27_81;
   assign m27_81 ={ {5{neg27[5]}} , neg27[5:1] };

   // m27_82 = W*in
   wire signed [9:0] m27_82;
   assign m27_82 =10'b0;

   // m27_83 = W*in
   wire signed [9:0] m27_83;
   assign m27_83 =10'b0;

   // m27_84 = W*in
   wire signed [9:0] m27_84;
   assign m27_84 =10'b0;

   // m27_85 = W*in
   wire signed [9:0] m27_85;
   assign m27_85 =10'b0;

   // m27_86 = W*in
   wire signed [9:0] m27_86;
   assign m27_86 =10'b0;

   // m27_87 = W*in
   wire signed [9:0] m27_87;
   assign m27_87 =10'b0;

   // m27_88 = W*in
   wire signed [9:0] m27_88;
   assign m27_88 =10'b0;

   // m27_89 = W*in
   wire signed [9:0] m27_89;
   assign m27_89 =10'b0;

   // m27_90 = W*in
   wire signed [9:0] m27_90;
   assign m27_90 =10'b0;

   // m27_91 = W*in
   wire signed [9:0] m27_91;
   assign m27_91 =10'b0;

   // m27_92 = W*in
   wire signed [9:0] m27_92;
   assign m27_92 =10'b0;

   // m27_93 = W*in
   wire signed [9:0] m27_93;
   assign m27_93 =10'b0;

   // m27_94 = W*in
   wire signed [9:0] m27_94;
   assign m27_94 =10'b0;

   // m27_95 = W*in
   wire signed [9:0] m27_95;
   assign m27_95 =10'b0;

   // m27_96 = W*in
   wire signed [9:0] m27_96;
   assign m27_96 =10'b0;

   // m27_97 = W*in
   wire signed [9:0] m27_97;
   assign m27_97 =10'b0;

   // m27_98 = W*in
   wire signed [9:0] m27_98;
   assign m27_98 =10'b0;

   // m27_99 = W*in
   wire signed [9:0] m27_99;
   assign m27_99 =10'b0;

   // m27_100 = W*in
   wire signed [9:0] m27_100;
   assign m27_100 =10'b0;

   // m27_101 = W*in
   wire signed [9:0] m27_101;
   assign m27_101 =10'b0;

   // m27_102 = W*in
   wire signed [9:0] m27_102;
   assign m27_102 =10'b0;

   // m27_103 = W*in
   wire signed [9:0] m27_103;
   assign m27_103 =10'b0;

   // m27_104 = W*in
   wire signed [9:0] m27_104;
   assign m27_104 =10'b0;

   // m27_105 = W*in
   wire signed [9:0] m27_105;
   assign m27_105 =10'b0;

   // m27_106 = W*in
   wire signed [9:0] m27_106;
   assign m27_106 =10'b0;

   // m27_107 = W*in
   wire signed [9:0] m27_107;
   assign m27_107 =10'b0;

   // m27_108 = W*in
   wire signed [9:0] m27_108;
   assign m27_108 =10'b0;

   // m27_109 = W*in
   wire signed [9:0] m27_109;
   assign m27_109 =10'b0;

   // m27_110 = W*in
   wire signed [9:0] m27_110;
   assign m27_110 =10'b0;

   // m27_111 = W*in
   wire signed [9:0] m27_111;
   assign m27_111 =10'b0;

   // m27_112 = W*in
   wire signed [9:0] m27_112;
   assign m27_112 =10'b0;

   // m27_113 = W*in
   wire signed [9:0] m27_113;
   assign m27_113 =10'b0;

   // m27_114 = W*in
   wire signed [9:0] m27_114;
   assign m27_114 =10'b0;

   // m27_115 = W*in
   wire signed [9:0] m27_115;
   assign m27_115 =10'b0;

   // m27_116 = W*in
   wire signed [9:0] m27_116;
   assign m27_116 =10'b0;

   // m27_117 = W*in
   wire signed [9:0] m27_117;
   assign m27_117 =10'b0;

   // m28_1 = W*in
   wire signed [9:0] m28_1;
   assign m28_1 =10'b0;

   // m28_2 = W*in
   wire signed [9:0] m28_2;
   assign m28_2 =10'b0;

   // m28_3 = W*in
   wire signed [9:0] m28_3;
   assign m28_3 =10'b0;

   // m28_4 = W*in
   wire signed [9:0] m28_4;
   assign m28_4 =10'b0;

   // m28_5 = W*in
   wire signed [9:0] m28_5;
   assign m28_5 =10'b0;

   // m28_6 = W*in
   wire signed [9:0] m28_6;
   assign m28_6 =10'b0;

   // m28_7 = W*in
   wire signed [9:0] m28_7;
   assign m28_7 =10'b0;

   // m28_8 = W*in
   wire signed [9:0] m28_8;
   assign m28_8 =10'b0;

   // m28_9 = W*in
   wire signed [9:0] m28_9;
   assign m28_9 =10'b0;

   // m28_10 = W*in
   wire signed [9:0] m28_10;
   assign m28_10 =10'b0;

   // m28_11 = W*in
   wire signed [9:0] m28_11;
   assign m28_11 =10'b0;

   // m28_12 = W*in
   wire signed [9:0] m28_12;
   assign m28_12 =10'b0;

   // m28_13 = W*in
   wire signed [9:0] m28_13;
   assign m28_13 =10'b0;

   // m28_14 = W*in
   wire signed [9:0] m28_14;
   assign m28_14 =10'b0;

   // m28_15 = W*in
   wire signed [9:0] m28_15;
   assign m28_15 =10'b0;

   // m28_16 = W*in
   wire signed [9:0] m28_16;
   assign m28_16 =10'b0;

   // m28_17 = W*in
   wire signed [9:0] m28_17;
   assign m28_17 =10'b0;

   // m28_18 = W*in
   wire signed [9:0] m28_18;
   assign m28_18 =10'b0;

   // m28_19 = W*in
   wire signed [9:0] m28_19;
   assign m28_19 =10'b0;

   // m28_20 = W*in
   wire signed [9:0] m28_20;
   assign m28_20 ={ {5{neg28[5]}} , neg28[5:1] };

   // m28_21 = W*in
   wire signed [9:0] m28_21;
   assign m28_21 =10'b0;

   // m28_22 = W*in
   wire signed [9:0] m28_22;
   assign m28_22 =10'b0;

   // m28_23 = W*in
   wire signed [9:0] m28_23;
   assign m28_23 =10'b0;

   // m28_24 = W*in
   wire signed [9:0] m28_24;
   assign m28_24 =10'b0;

   // m28_25 = W*in
   wire signed [9:0] m28_25;
   assign m28_25 =10'b0;

   // m28_26 = W*in
   wire signed [9:0] m28_26;
   assign m28_26 =10'b0;

   // m28_27 = W*in
   wire signed [9:0] m28_27;
   assign m28_27 =10'b0;

   // m28_28 = W*in
   wire signed [9:0] m28_28;
   assign m28_28 =10'b0;

   // m28_29 = W*in
   wire signed [9:0] m28_29;
   assign m28_29 ={ {5{in28[5]}} , in28[5:1] };

   // m28_30 = W*in
   wire signed [9:0] m28_30;
   assign m28_30 =10'b0;

   // m28_31 = W*in
   wire signed [9:0] m28_31;
   assign m28_31 =10'b0;

   // m28_32 = W*in
   wire signed [9:0] m28_32;
   assign m28_32 =10'b0;

   // m28_33 = W*in
   wire signed [9:0] m28_33;
   assign m28_33 =10'b0;

   // m28_34 = W*in
   wire signed [9:0] m28_34;
   assign m28_34 =10'b0;

   // m28_35 = W*in
   wire signed [9:0] m28_35;
   assign m28_35 =10'b0;

   // m28_36 = W*in
   wire signed [9:0] m28_36;
   assign m28_36 =10'b0;

   // m28_37 = W*in
   wire signed [9:0] m28_37;
   assign m28_37 =10'b0;

   // m28_38 = W*in
   wire signed [9:0] m28_38;
   assign m28_38 =10'b0;

   // m28_39 = W*in
   wire signed [9:0] m28_39;
   assign m28_39 =10'b0;

   // m28_40 = W*in
   wire signed [9:0] m28_40;
   assign m28_40 =10'b0;

   // m28_41 = W*in
   wire signed [9:0] m28_41;
   assign m28_41 =10'b0;

   // m28_42 = W*in
   wire signed [9:0] m28_42;
   assign m28_42 =10'b0;

   // m28_43 = W*in
   wire signed [9:0] m28_43;
   assign m28_43 =10'b0;

   // m28_44 = W*in
   wire signed [9:0] m28_44;
   assign m28_44 =10'b0;

   // m28_45 = W*in
   wire signed [9:0] m28_45;
   assign m28_45 =10'b0;

   // m28_46 = W*in
   wire signed [9:0] m28_46;
   assign m28_46 =10'b0;

   // m28_47 = W*in
   wire signed [9:0] m28_47;
   assign m28_47 =10'b0;

   // m28_48 = W*in
   wire signed [9:0] m28_48;
   assign m28_48 =10'b0;

   // m28_49 = W*in
   wire signed [9:0] m28_49;
   assign m28_49 =10'b0;

   // m28_50 = W*in
   wire signed [9:0] m28_50;
   assign m28_50 =10'b0;

   // m28_51 = W*in
   wire signed [9:0] m28_51;
   assign m28_51 =10'b0;

   // m28_52 = W*in
   wire signed [9:0] m28_52;
   assign m28_52 =10'b0;

   // m28_53 = W*in
   wire signed [9:0] m28_53;
   assign m28_53 =10'b0;

   // m28_54 = W*in
   wire signed [9:0] m28_54;
   assign m28_54 =10'b0;

   // m28_55 = W*in
   wire signed [9:0] m28_55;
   assign m28_55 =10'b0;

   // m28_56 = W*in
   wire signed [9:0] m28_56;
   assign m28_56 =10'b0;

   // m28_57 = W*in
   wire signed [9:0] m28_57;
   assign m28_57 =10'b0;

   // m28_58 = W*in
   wire signed [9:0] m28_58;
   assign m28_58 =10'b0;

   // m28_59 = W*in
   wire signed [9:0] m28_59;
   assign m28_59 =10'b0;

   // m28_60 = W*in
   wire signed [9:0] m28_60;
   assign m28_60 =10'b0;

   // m28_61 = W*in
   wire signed [9:0] m28_61;
   assign m28_61 =10'b0;

   // m28_62 = W*in
   wire signed [9:0] m28_62;
   assign m28_62 =10'b0;

   // m28_63 = W*in
   wire signed [9:0] m28_63;
   assign m28_63 =10'b0;

   // m28_64 = W*in
   wire signed [9:0] m28_64;
   assign m28_64 ={ {5{neg28[5]}} , neg28[5:1] };

   // m28_65 = W*in
   wire signed [9:0] m28_65;
   assign m28_65 =10'b0;

   // m28_66 = W*in
   wire signed [9:0] m28_66;
   assign m28_66 =10'b0;

   // m28_67 = W*in
   wire signed [9:0] m28_67;
   assign m28_67 =10'b0;

   // m28_68 = W*in
   wire signed [9:0] m28_68;
   assign m28_68 =10'b0;

   // m28_69 = W*in
   wire signed [9:0] m28_69;
   assign m28_69 =10'b0;

   // m28_70 = W*in
   wire signed [9:0] m28_70;
   assign m28_70 =10'b0;

   // m28_71 = W*in
   wire signed [9:0] m28_71;
   assign m28_71 =10'b0;

   // m28_72 = W*in
   wire signed [9:0] m28_72;
   assign m28_72 =10'b0;

   // m28_73 = W*in
   wire signed [9:0] m28_73;
   assign m28_73 =10'b0;

   // m28_74 = W*in
   wire signed [9:0] m28_74;
   assign m28_74 =10'b0;

   // m28_75 = W*in
   wire signed [9:0] m28_75;
   assign m28_75 =10'b0;

   // m28_76 = W*in
   wire signed [9:0] m28_76;
   assign m28_76 =10'b0;

   // m28_77 = W*in
   wire signed [9:0] m28_77;
   assign m28_77 =10'b0;

   // m28_78 = W*in
   wire signed [9:0] m28_78;
   assign m28_78 =10'b0;

   // m28_79 = W*in
   wire signed [9:0] m28_79;
   assign m28_79 =10'b0;

   // m28_80 = W*in
   wire signed [9:0] m28_80;
   assign m28_80 =10'b0;

   // m28_81 = W*in
   wire signed [9:0] m28_81;
   assign m28_81 =10'b0;

   // m28_82 = W*in
   wire signed [9:0] m28_82;
   assign m28_82 =10'b0;

   // m28_83 = W*in
   wire signed [9:0] m28_83;
   assign m28_83 =10'b0;

   // m28_84 = W*in
   wire signed [9:0] m28_84;
   assign m28_84 =10'b0;

   // m28_85 = W*in
   wire signed [9:0] m28_85;
   assign m28_85 ={ {5{in28[5]}} , in28[5:1] };

   // m28_86 = W*in
   wire signed [9:0] m28_86;
   assign m28_86 =10'b0;

   // m28_87 = W*in
   wire signed [9:0] m28_87;
   assign m28_87 =10'b0;

   // m28_88 = W*in
   wire signed [9:0] m28_88;
   assign m28_88 =10'b0;

   // m28_89 = W*in
   wire signed [9:0] m28_89;
   assign m28_89 =10'b0;

   // m28_90 = W*in
   wire signed [9:0] m28_90;
   assign m28_90 =10'b0;

   // m28_91 = W*in
   wire signed [9:0] m28_91;
   assign m28_91 =10'b0;

   // m28_92 = W*in
   wire signed [9:0] m28_92;
   assign m28_92 =10'b0;

   // m28_93 = W*in
   wire signed [9:0] m28_93;
   assign m28_93 =10'b0;

   // m28_94 = W*in
   wire signed [9:0] m28_94;
   assign m28_94 =10'b0;

   // m28_95 = W*in
   wire signed [9:0] m28_95;
   assign m28_95 =10'b0;

   // m28_96 = W*in
   wire signed [9:0] m28_96;
   assign m28_96 =10'b0;

   // m28_97 = W*in
   wire signed [9:0] m28_97;
   assign m28_97 =10'b0;

   // m28_98 = W*in
   wire signed [9:0] m28_98;
   assign m28_98 =10'b0;

   // m28_99 = W*in
   wire signed [9:0] m28_99;
   assign m28_99 =10'b0;

   // m28_100 = W*in
   wire signed [9:0] m28_100;
   assign m28_100 =10'b0;

   // m28_101 = W*in
   wire signed [9:0] m28_101;
   assign m28_101 =10'b0;

   // m28_102 = W*in
   wire signed [9:0] m28_102;
   assign m28_102 =10'b0;

   // m28_103 = W*in
   wire signed [9:0] m28_103;
   assign m28_103 =10'b0;

   // m28_104 = W*in
   wire signed [9:0] m28_104;
   assign m28_104 =10'b0;

   // m28_105 = W*in
   wire signed [9:0] m28_105;
   assign m28_105 =10'b0;

   // m28_106 = W*in
   wire signed [9:0] m28_106;
   assign m28_106 =10'b0;

   // m28_107 = W*in
   wire signed [9:0] m28_107;
   assign m28_107 =10'b0;

   // m28_108 = W*in
   wire signed [9:0] m28_108;
   assign m28_108 =10'b0;

   // m28_109 = W*in
   wire signed [9:0] m28_109;
   assign m28_109 =10'b0;

   // m28_110 = W*in
   wire signed [9:0] m28_110;
   assign m28_110 =10'b0;

   // m28_111 = W*in
   wire signed [9:0] m28_111;
   assign m28_111 =10'b0;

   // m28_112 = W*in
   wire signed [9:0] m28_112;
   assign m28_112 =10'b0;

   // m28_113 = W*in
   wire signed [9:0] m28_113;
   assign m28_113 =10'b0;

   // m28_114 = W*in
   wire signed [9:0] m28_114;
   assign m28_114 =10'b0;

   // m28_115 = W*in
   wire signed [9:0] m28_115;
   assign m28_115 =10'b0;

   // m28_116 = W*in
   wire signed [9:0] m28_116;
   assign m28_116 =10'b0;

   // m28_117 = W*in
   wire signed [9:0] m28_117;
   assign m28_117 =10'b0;

   // m29_1 = W*in
   wire signed [9:0] m29_1;
   assign m29_1 =10'b0;

   // m29_2 = W*in
   wire signed [9:0] m29_2;
   assign m29_2 =10'b0;

   // m29_3 = W*in
   wire signed [9:0] m29_3;
   assign m29_3 =10'b0;

   // m29_4 = W*in
   wire signed [9:0] m29_4;
   assign m29_4 =10'b0;

   // m29_5 = W*in
   wire signed [9:0] m29_5;
   assign m29_5 =10'b0;

   // m29_6 = W*in
   wire signed [9:0] m29_6;
   assign m29_6 =10'b0;

   // m29_7 = W*in
   wire signed [9:0] m29_7;
   assign m29_7 =10'b0;

   // m29_8 = W*in
   wire signed [9:0] m29_8;
   assign m29_8 =10'b0;

   // m29_9 = W*in
   wire signed [9:0] m29_9;
   assign m29_9 =10'b0;

   // m29_10 = W*in
   wire signed [9:0] m29_10;
   assign m29_10 =10'b0;

   // m29_11 = W*in
   wire signed [9:0] m29_11;
   assign m29_11 =10'b0;

   // m29_12 = W*in
   wire signed [9:0] m29_12;
   assign m29_12 =10'b0;

   // m29_13 = W*in
   wire signed [9:0] m29_13;
   assign m29_13 =10'b0;

   // m29_14 = W*in
   wire signed [9:0] m29_14;
   assign m29_14 =10'b0;

   // m29_15 = W*in
   wire signed [9:0] m29_15;
   assign m29_15 =10'b0;

   // m29_16 = W*in
   wire signed [9:0] m29_16;
   assign m29_16 =10'b0;

   // m29_17 = W*in
   wire signed [9:0] m29_17;
   assign m29_17 =10'b0;

   // m29_18 = W*in
   wire signed [9:0] m29_18;
   assign m29_18 =10'b0;

   // m29_19 = W*in
   wire signed [9:0] m29_19;
   assign m29_19 =10'b0;

   // m29_20 = W*in
   wire signed [9:0] m29_20;
   assign m29_20 ={ {5{in29[5]}} , in29[5:1] };

   // m29_21 = W*in
   wire signed [9:0] m29_21;
   assign m29_21 =10'b0;

   // m29_22 = W*in
   wire signed [9:0] m29_22;
   assign m29_22 =10'b0;

   // m29_23 = W*in
   wire signed [9:0] m29_23;
   assign m29_23 =10'b0;

   // m29_24 = W*in
   wire signed [9:0] m29_24;
   assign m29_24 =10'b0;

   // m29_25 = W*in
   wire signed [9:0] m29_25;
   assign m29_25 ={ {4{neg29[5]}} , neg29[5:0] };

   // m29_26 = W*in
   wire signed [9:0] m29_26;
   assign m29_26 =10'b0;

   // m29_27 = W*in
   wire signed [9:0] m29_27;
   assign m29_27 =10'b0;

   // m29_28 = W*in
   wire signed [9:0] m29_28;
   assign m29_28 ={ {5{neg29[5]}} , neg29[5:1] };

   // m29_29 = W*in
   wire signed [9:0] m29_29;
   assign m29_29 ={ {5{neg29[5]}} , neg29[5:1] };

   // m29_30 = W*in
   wire signed [9:0] m29_30;
   assign m29_30 =10'b0;

   // m29_31 = W*in
   wire signed [9:0] m29_31;
   assign m29_31 =10'b0;

   // m29_32 = W*in
   wire signed [9:0] m29_32;
   assign m29_32 =10'b0;

   // m29_33 = W*in
   wire signed [9:0] m29_33;
   assign m29_33 =10'b0;

   // m29_34 = W*in
   wire signed [9:0] m29_34;
   assign m29_34 =10'b0;

   // m29_35 = W*in
   wire signed [9:0] m29_35;
   assign m29_35 =10'b0;

   // m29_36 = W*in
   wire signed [9:0] m29_36;
   assign m29_36 =10'b0;

   // m29_37 = W*in
   wire signed [9:0] m29_37;
   assign m29_37 =10'b0;

   // m29_38 = W*in
   wire signed [9:0] m29_38;
   assign m29_38 =10'b0;

   // m29_39 = W*in
   wire signed [9:0] m29_39;
   assign m29_39 =10'b0;

   // m29_40 = W*in
   wire signed [9:0] m29_40;
   assign m29_40 =10'b0;

   // m29_41 = W*in
   wire signed [9:0] m29_41;
   assign m29_41 =10'b0;

   // m29_42 = W*in
   wire signed [9:0] m29_42;
   assign m29_42 =10'b0;

   // m29_43 = W*in
   wire signed [9:0] m29_43;
   assign m29_43 =10'b0;

   // m29_44 = W*in
   wire signed [9:0] m29_44;
   assign m29_44 =10'b0;

   // m29_45 = W*in
   wire signed [9:0] m29_45;
   assign m29_45 =10'b0;

   // m29_46 = W*in
   wire signed [9:0] m29_46;
   assign m29_46 =10'b0;

   // m29_47 = W*in
   wire signed [9:0] m29_47;
   assign m29_47 =10'b0;

   // m29_48 = W*in
   wire signed [9:0] m29_48;
   assign m29_48 =10'b0;

   // m29_49 = W*in
   wire signed [9:0] m29_49;
   assign m29_49 =10'b0;

   // m29_50 = W*in
   wire signed [9:0] m29_50;
   assign m29_50 =10'b0;

   // m29_51 = W*in
   wire signed [9:0] m29_51;
   assign m29_51 =10'b0;

   // m29_52 = W*in
   wire signed [9:0] m29_52;
   assign m29_52 =10'b0;

   // m29_53 = W*in
   wire signed [9:0] m29_53;
   assign m29_53 =10'b0;

   // m29_54 = W*in
   wire signed [9:0] m29_54;
   assign m29_54 =10'b0;

   // m29_55 = W*in
   wire signed [9:0] m29_55;
   assign m29_55 =10'b0;

   // m29_56 = W*in
   wire signed [9:0] m29_56;
   assign m29_56 =10'b0;

   // m29_57 = W*in
   wire signed [9:0] m29_57;
   assign m29_57 =10'b0;

   // m29_58 = W*in
   wire signed [9:0] m29_58;
   assign m29_58 =10'b0;

   // m29_59 = W*in
   wire signed [9:0] m29_59;
   assign m29_59 ={ {4{neg29[5]}} , neg29[5:0] };

   // m29_60 = W*in
   wire signed [9:0] m29_60;
   assign m29_60 =10'b0;

   // m29_61 = W*in
   wire signed [9:0] m29_61;
   assign m29_61 =10'b0;

   // m29_62 = W*in
   wire signed [9:0] m29_62;
   assign m29_62 =10'b0;

   // m29_63 = W*in
   wire signed [9:0] m29_63;
   assign m29_63 =10'b0;

   // m29_64 = W*in
   wire signed [9:0] m29_64;
   assign m29_64 =10'b0;

   // m29_65 = W*in
   wire signed [9:0] m29_65;
   assign m29_65 =10'b0;

   // m29_66 = W*in
   wire signed [9:0] m29_66;
   assign m29_66 ={ {5{neg29[5]}} , neg29[5:1] };

   // m29_67 = W*in
   wire signed [9:0] m29_67;
   assign m29_67 =10'b0;

   // m29_68 = W*in
   wire signed [9:0] m29_68;
   assign m29_68 =10'b0;

   // m29_69 = W*in
   wire signed [9:0] m29_69;
   assign m29_69 ={ {5{in29[5]}} , in29[5:1] };

   // m29_70 = W*in
   wire signed [9:0] m29_70;
   assign m29_70 =10'b0;

   // m29_71 = W*in
   wire signed [9:0] m29_71;
   assign m29_71 =10'b0;

   // m29_72 = W*in
   wire signed [9:0] m29_72;
   assign m29_72 =10'b0;

   // m29_73 = W*in
   wire signed [9:0] m29_73;
   assign m29_73 =10'b0;

   // m29_74 = W*in
   wire signed [9:0] m29_74;
   assign m29_74 =10'b0;

   // m29_75 = W*in
   wire signed [9:0] m29_75;
   assign m29_75 =10'b0;

   // m29_76 = W*in
   wire signed [9:0] m29_76;
   assign m29_76 =10'b0;

   // m29_77 = W*in
   wire signed [9:0] m29_77;
   assign m29_77 =10'b0;

   // m29_78 = W*in
   wire signed [9:0] m29_78;
   assign m29_78 =10'b0;

   // m29_79 = W*in
   wire signed [9:0] m29_79;
   assign m29_79 =10'b0;

   // m29_80 = W*in
   wire signed [9:0] m29_80;
   assign m29_80 =10'b0;

   // m29_81 = W*in
   wire signed [9:0] m29_81;
   assign m29_81 =10'b0;

   // m29_82 = W*in
   wire signed [9:0] m29_82;
   assign m29_82 ={ {5{in29[5]}} , in29[5:1] };

   // m29_83 = W*in
   wire signed [9:0] m29_83;
   assign m29_83 =10'b0;

   // m29_84 = W*in
   wire signed [9:0] m29_84;
   assign m29_84 =10'b0;

   // m29_85 = W*in
   wire signed [9:0] m29_85;
   assign m29_85 =10'b0;

   // m29_86 = W*in
   wire signed [9:0] m29_86;
   assign m29_86 =10'b0;

   // m29_87 = W*in
   wire signed [9:0] m29_87;
   assign m29_87 =10'b0;

   // m29_88 = W*in
   wire signed [9:0] m29_88;
   assign m29_88 =10'b0;

   // m29_89 = W*in
   wire signed [9:0] m29_89;
   assign m29_89 =10'b0;

   // m29_90 = W*in
   wire signed [9:0] m29_90;
   assign m29_90 =10'b0;

   // m29_91 = W*in
   wire signed [9:0] m29_91;
   assign m29_91 =10'b0;

   // m29_92 = W*in
   wire signed [9:0] m29_92;
   assign m29_92 =10'b0;

   // m29_93 = W*in
   wire signed [9:0] m29_93;
   assign m29_93 =10'b0;

   // m29_94 = W*in
   wire signed [9:0] m29_94;
   assign m29_94 =10'b0;

   // m29_95 = W*in
   wire signed [9:0] m29_95;
   assign m29_95 =10'b0;

   // m29_96 = W*in
   wire signed [9:0] m29_96;
   assign m29_96 =10'b0;

   // m29_97 = W*in
   wire signed [9:0] m29_97;
   assign m29_97 =10'b0;

   // m29_98 = W*in
   wire signed [9:0] m29_98;
   assign m29_98 =10'b0;

   // m29_99 = W*in
   wire signed [9:0] m29_99;
   assign m29_99 =10'b0;

   // m29_100 = W*in
   wire signed [9:0] m29_100;
   assign m29_100 =10'b0;

   // m29_101 = W*in
   wire signed [9:0] m29_101;
   assign m29_101 =10'b0;

   // m29_102 = W*in
   wire signed [9:0] m29_102;
   assign m29_102 =10'b0;

   // m29_103 = W*in
   wire signed [9:0] m29_103;
   assign m29_103 =10'b0;

   // m29_104 = W*in
   wire signed [9:0] m29_104;
   assign m29_104 =10'b0;

   // m29_105 = W*in
   wire signed [9:0] m29_105;
   assign m29_105 =10'b0;

   // m29_106 = W*in
   wire signed [9:0] m29_106;
   assign m29_106 =10'b0;

   // m29_107 = W*in
   wire signed [9:0] m29_107;
   assign m29_107 =10'b0;

   // m29_108 = W*in
   wire signed [9:0] m29_108;
   assign m29_108 ={ {5{in29[5]}} , in29[5:1] };

   // m29_109 = W*in
   wire signed [9:0] m29_109;
   assign m29_109 ={ {5{in29[5]}} , in29[5:1] };

   // m29_110 = W*in
   wire signed [9:0] m29_110;
   assign m29_110 =10'b0;

   // m29_111 = W*in
   wire signed [9:0] m29_111;
   assign m29_111 =10'b0;

   // m29_112 = W*in
   wire signed [9:0] m29_112;
   assign m29_112 =10'b0;

   // m29_113 = W*in
   wire signed [9:0] m29_113;
   assign m29_113 =10'b0;

   // m29_114 = W*in
   wire signed [9:0] m29_114;
   assign m29_114 =10'b0;

   // m29_115 = W*in
   wire signed [9:0] m29_115;
   assign m29_115 =10'b0;

   // m29_116 = W*in
   wire signed [9:0] m29_116;
   assign m29_116 =10'b0;

   // m29_117 = W*in
   wire signed [9:0] m29_117;
   assign m29_117 =10'b0;

   // m30_1 = W*in
   wire signed [9:0] m30_1;
   assign m30_1 =10'b0;

   // m30_2 = W*in
   wire signed [9:0] m30_2;
   assign m30_2 =10'b0;

   // m30_3 = W*in
   wire signed [9:0] m30_3;
   assign m30_3 ={ {4{in30[5]}} , in30[5:0] };

   // m30_4 = W*in
   wire signed [9:0] m30_4;
   assign m30_4 =10'b0;

   // m30_5 = W*in
   wire signed [9:0] m30_5;
   assign m30_5 =10'b0;

   // m30_6 = W*in
   wire signed [9:0] m30_6;
   assign m30_6 =10'b0;

   // m30_7 = W*in
   wire signed [9:0] m30_7;
   assign m30_7 =10'b0;

   // m30_8 = W*in
   wire signed [9:0] m30_8;
   assign m30_8 =10'b0;

   // m30_9 = W*in
   wire signed [9:0] m30_9;
   assign m30_9 =10'b0;

   // m30_10 = W*in
   wire signed [9:0] m30_10;
   assign m30_10 =10'b0;

   // m30_11 = W*in
   wire signed [9:0] m30_11;
   assign m30_11 =10'b0;

   // m30_12 = W*in
   wire signed [9:0] m30_12;
   assign m30_12 =10'b0;

   // m30_13 = W*in
   wire signed [9:0] m30_13;
   assign m30_13 =10'b0;

   // m30_14 = W*in
   wire signed [9:0] m30_14;
   assign m30_14 =10'b0;

   // m30_15 = W*in
   wire signed [9:0] m30_15;
   assign m30_15 =10'b0;

   // m30_16 = W*in
   wire signed [9:0] m30_16;
   assign m30_16 =10'b0;

   // m30_17 = W*in
   wire signed [9:0] m30_17;
   assign m30_17 =10'b0;

   // m30_18 = W*in
   wire signed [9:0] m30_18;
   assign m30_18 =10'b0;

   // m30_19 = W*in
   wire signed [9:0] m30_19;
   assign m30_19 =10'b0;

   // m30_20 = W*in
   wire signed [9:0] m30_20;
   assign m30_20 =10'b0;

   // m30_21 = W*in
   wire signed [9:0] m30_21;
   assign m30_21 =10'b0;

   // m30_22 = W*in
   wire signed [9:0] m30_22;
   assign m30_22 ={ {5{in30[5]}} , in30[5:1] };

   // m30_23 = W*in
   wire signed [9:0] m30_23;
   assign m30_23 =10'b0;

   // m30_24 = W*in
   wire signed [9:0] m30_24;
   assign m30_24 =10'b0;

   // m30_25 = W*in
   wire signed [9:0] m30_25;
   assign m30_25 ={ {4{neg30[5]}} , neg30[5:0] };

   // m30_26 = W*in
   wire signed [9:0] m30_26;
   assign m30_26 =10'b0;

   // m30_27 = W*in
   wire signed [9:0] m30_27;
   assign m30_27 ={ {5{in30[5]}} , in30[5:1] };

   // m30_28 = W*in
   wire signed [9:0] m30_28;
   assign m30_28 ={ {5{neg30[5]}} , neg30[5:1] };

   // m30_29 = W*in
   wire signed [9:0] m30_29;
   assign m30_29 ={ {5{neg30[5]}} , neg30[5:1] };

   // m30_30 = W*in
   wire signed [9:0] m30_30;
   assign m30_30 =10'b0;

   // m30_31 = W*in
   wire signed [9:0] m30_31;
   assign m30_31 ={ {5{in30[5]}} , in30[5:1] };

   // m30_32 = W*in
   wire signed [9:0] m30_32;
   assign m30_32 =10'b0;

   // m30_33 = W*in
   wire signed [9:0] m30_33;
   assign m30_33 =10'b0;

   // m30_34 = W*in
   wire signed [9:0] m30_34;
   assign m30_34 =10'b0;

   // m30_35 = W*in
   wire signed [9:0] m30_35;
   assign m30_35 ={ {4{neg30[5]}} , neg30[5:0] };

   // m30_36 = W*in
   wire signed [9:0] m30_36;
   assign m30_36 ={ {5{neg30[5]}} , neg30[5:1] };

   // m30_37 = W*in
   wire signed [9:0] m30_37;
   assign m30_37 =10'b0;

   // m30_38 = W*in
   wire signed [9:0] m30_38;
   assign m30_38 =10'b0;

   // m30_39 = W*in
   wire signed [9:0] m30_39;
   assign m30_39 =10'b0;

   // m30_40 = W*in
   wire signed [9:0] m30_40;
   assign m30_40 =10'b0;

   // m30_41 = W*in
   wire signed [9:0] m30_41;
   assign m30_41 =10'b0;

   // m30_42 = W*in
   wire signed [9:0] m30_42;
   assign m30_42 =10'b0;

   // m30_43 = W*in
   wire signed [9:0] m30_43;
   assign m30_43 =10'b0;

   // m30_44 = W*in
   wire signed [9:0] m30_44;
   assign m30_44 =10'b0;

   // m30_45 = W*in
   wire signed [9:0] m30_45;
   assign m30_45 =10'b0;

   // m30_46 = W*in
   wire signed [9:0] m30_46;
   assign m30_46 =10'b0;

   // m30_47 = W*in
   wire signed [9:0] m30_47;
   assign m30_47 =10'b0;

   // m30_48 = W*in
   wire signed [9:0] m30_48;
   assign m30_48 =10'b0;

   // m30_49 = W*in
   wire signed [9:0] m30_49;
   assign m30_49 =10'b0;

   // m30_50 = W*in
   wire signed [9:0] m30_50;
   assign m30_50 =10'b0;

   // m30_51 = W*in
   wire signed [9:0] m30_51;
   assign m30_51 =10'b0;

   // m30_52 = W*in
   wire signed [9:0] m30_52;
   assign m30_52 =10'b0;

   // m30_53 = W*in
   wire signed [9:0] m30_53;
   assign m30_53 =10'b0;

   // m30_54 = W*in
   wire signed [9:0] m30_54;
   assign m30_54 =10'b0;

   // m30_55 = W*in
   wire signed [9:0] m30_55;
   assign m30_55 =10'b0;

   // m30_56 = W*in
   wire signed [9:0] m30_56;
   assign m30_56 =10'b0;

   // m30_57 = W*in
   wire signed [9:0] m30_57;
   assign m30_57 =10'b0;

   // m30_58 = W*in
   wire signed [9:0] m30_58;
   assign m30_58 =10'b0;

   // m30_59 = W*in
   wire signed [9:0] m30_59;
   assign m30_59 =10'b0;

   // m30_60 = W*in
   wire signed [9:0] m30_60;
   assign m30_60 =10'b0;

   // m30_61 = W*in
   wire signed [9:0] m30_61;
   assign m30_61 =10'b0;

   // m30_62 = W*in
   wire signed [9:0] m30_62;
   assign m30_62 =10'b0;

   // m30_63 = W*in
   wire signed [9:0] m30_63;
   assign m30_63 =10'b0;

   // m30_64 = W*in
   wire signed [9:0] m30_64;
   assign m30_64 =10'b0;

   // m30_65 = W*in
   wire signed [9:0] m30_65;
   assign m30_65 =10'b0;

   // m30_66 = W*in
   wire signed [9:0] m30_66;
   assign m30_66 ={ {5{neg30[5]}} , neg30[5:1] };

   // m30_67 = W*in
   wire signed [9:0] m30_67;
   assign m30_67 =10'b0;

   // m30_68 = W*in
   wire signed [9:0] m30_68;
   assign m30_68 =10'b0;

   // m30_69 = W*in
   wire signed [9:0] m30_69;
   assign m30_69 ={ {4{in30[5]}} , in30[5:0] };

   // m30_70 = W*in
   wire signed [9:0] m30_70;
   assign m30_70 ={ {5{neg30[5]}} , neg30[5:1] };

   // m30_71 = W*in
   wire signed [9:0] m30_71;
   assign m30_71 =10'b0;

   // m30_72 = W*in
   wire signed [9:0] m30_72;
   assign m30_72 ={ {4{neg30[5]}} , neg30[5:0] };

   // m30_73 = W*in
   wire signed [9:0] m30_73;
   assign m30_73 =10'b0;

   // m30_74 = W*in
   wire signed [9:0] m30_74;
   assign m30_74 =10'b0;

   // m30_75 = W*in
   wire signed [9:0] m30_75;
   assign m30_75 ={ {4{neg30[5]}} , neg30[5:0] };

   // m30_76 = W*in
   wire signed [9:0] m30_76;
   assign m30_76 ={ {4{in30[5]}} , in30[5:0] };

   // m30_77 = W*in
   wire signed [9:0] m30_77;
   assign m30_77 =10'b0;

   // m30_78 = W*in
   wire signed [9:0] m30_78;
   assign m30_78 =10'b0;

   // m30_79 = W*in
   wire signed [9:0] m30_79;
   assign m30_79 =10'b0;

   // m30_80 = W*in
   wire signed [9:0] m30_80;
   assign m30_80 ={ {4{in30[5]}} , in30[5:0] };

   // m30_81 = W*in
   wire signed [9:0] m30_81;
   assign m30_81 =10'b0;

   // m30_82 = W*in
   wire signed [9:0] m30_82;
   assign m30_82 ={ {4{in30[5]}} , in30[5:0] };

   // m30_83 = W*in
   wire signed [9:0] m30_83;
   assign m30_83 =10'b0;

   // m30_84 = W*in
   wire signed [9:0] m30_84;
   assign m30_84 =10'b0;

   // m30_85 = W*in
   wire signed [9:0] m30_85;
   assign m30_85 ={ {5{in30[5]}} , in30[5:1] };

   // m30_86 = W*in
   wire signed [9:0] m30_86;
   assign m30_86 =10'b0;

   // m30_87 = W*in
   wire signed [9:0] m30_87;
   assign m30_87 =10'b0;

   // m30_88 = W*in
   wire signed [9:0] m30_88;
   assign m30_88 =10'b0;

   // m30_89 = W*in
   wire signed [9:0] m30_89;
   assign m30_89 ={ {4{in30[5]}} , in30[5:0] };

   // m30_90 = W*in
   wire signed [9:0] m30_90;
   assign m30_90 =10'b0;

   // m30_91 = W*in
   wire signed [9:0] m30_91;
   assign m30_91 =10'b0;

   // m30_92 = W*in
   wire signed [9:0] m30_92;
   assign m30_92 =10'b0;

   // m30_93 = W*in
   wire signed [9:0] m30_93;
   assign m30_93 =10'b0;

   // m30_94 = W*in
   wire signed [9:0] m30_94;
   assign m30_94 ={ {4{neg30[5]}} , neg30[5:0] };

   // m30_95 = W*in
   wire signed [9:0] m30_95;
   assign m30_95 =10'b0;

   // m30_96 = W*in
   wire signed [9:0] m30_96;
   assign m30_96 =10'b0;

   // m30_97 = W*in
   wire signed [9:0] m30_97;
   assign m30_97 =10'b0;

   // m30_98 = W*in
   wire signed [9:0] m30_98;
   assign m30_98 ={ {4{in30[5]}} , in30[5:0] };

   // m30_99 = W*in
   wire signed [9:0] m30_99;
   assign m30_99 =10'b0;

   // m30_100 = W*in
   wire signed [9:0] m30_100;
   assign m30_100 =10'b0;

   // m30_101 = W*in
   wire signed [9:0] m30_101;
   assign m30_101 =10'b0;

   // m30_102 = W*in
   wire signed [9:0] m30_102;
   assign m30_102 =10'b0;

   // m30_103 = W*in
   wire signed [9:0] m30_103;
   assign m30_103 =10'b0;

   // m30_104 = W*in
   wire signed [9:0] m30_104;
   assign m30_104 =10'b0;

   // m30_105 = W*in
   wire signed [9:0] m30_105;
   assign m30_105 =10'b0;

   // m30_106 = W*in
   wire signed [9:0] m30_106;
   assign m30_106 =10'b0;

   // m30_107 = W*in
   wire signed [9:0] m30_107;
   assign m30_107 ={ {5{in30[5]}} , in30[5:1] };

   // m30_108 = W*in
   wire signed [9:0] m30_108;
   assign m30_108 =10'b0;

   // m30_109 = W*in
   wire signed [9:0] m30_109;
   assign m30_109 ={ {4{in30[5]}} , in30[5:0] };

   // m30_110 = W*in
   wire signed [9:0] m30_110;
   assign m30_110 =10'b0;

   // m30_111 = W*in
   wire signed [9:0] m30_111;
   assign m30_111 =10'b0;

   // m30_112 = W*in
   wire signed [9:0] m30_112;
   assign m30_112 =10'b0;

   // m30_113 = W*in
   wire signed [9:0] m30_113;
   assign m30_113 =10'b0;

   // m30_114 = W*in
   wire signed [9:0] m30_114;
   assign m30_114 =10'b0;

   // m30_115 = W*in
   wire signed [9:0] m30_115;
   assign m30_115 =10'b0;

   // m30_116 = W*in
   wire signed [9:0] m30_116;
   assign m30_116 =10'b0;

   // m30_117 = W*in
   wire signed [9:0] m30_117;
   assign m30_117 =10'b0;

   // m31_1 = W*in
   wire signed [9:0] m31_1;
   assign m31_1 =10'b0;

   // m31_2 = W*in
   wire signed [9:0] m31_2;
   assign m31_2 ={ {4{in31[5]}} , in31[5:0] };

   // m31_3 = W*in
   wire signed [9:0] m31_3;
   assign m31_3 =10'b0;

   // m31_4 = W*in
   wire signed [9:0] m31_4;
   assign m31_4 =10'b0;

   // m31_5 = W*in
   wire signed [9:0] m31_5;
   assign m31_5 =10'b0;

   // m31_6 = W*in
   wire signed [9:0] m31_6;
   assign m31_6 =10'b0;

   // m31_7 = W*in
   wire signed [9:0] m31_7;
   assign m31_7 =10'b0;

   // m31_8 = W*in
   wire signed [9:0] m31_8;
   assign m31_8 =10'b0;

   // m31_9 = W*in
   wire signed [9:0] m31_9;
   assign m31_9 =10'b0;

   // m31_10 = W*in
   wire signed [9:0] m31_10;
   assign m31_10 ={ {4{in31[5]}} , in31[5:0] };

   // m31_11 = W*in
   wire signed [9:0] m31_11;
   assign m31_11 =10'b0;

   // m31_12 = W*in
   wire signed [9:0] m31_12;
   assign m31_12 =10'b0;

   // m31_13 = W*in
   wire signed [9:0] m31_13;
   assign m31_13 =10'b0;

   // m31_14 = W*in
   wire signed [9:0] m31_14;
   assign m31_14 =10'b0;

   // m31_15 = W*in
   wire signed [9:0] m31_15;
   assign m31_15 =10'b0;

   // m31_16 = W*in
   wire signed [9:0] m31_16;
   assign m31_16 =10'b0;

   // m31_17 = W*in
   wire signed [9:0] m31_17;
   assign m31_17 ={ {5{in31[5]}} , in31[5:1] };

   // m31_18 = W*in
   wire signed [9:0] m31_18;
   assign m31_18 =10'b0;

   // m31_19 = W*in
   wire signed [9:0] m31_19;
   assign m31_19 =10'b0;

   // m31_20 = W*in
   wire signed [9:0] m31_20;
   assign m31_20 =10'b0;

   // m31_21 = W*in
   wire signed [9:0] m31_21;
   assign m31_21 =10'b0;

   // m31_22 = W*in
   wire signed [9:0] m31_22;
   assign m31_22 ={ {5{in31[5]}} , in31[5:1] };

   // m31_23 = W*in
   wire signed [9:0] m31_23;
   assign m31_23 =10'b0;

   // m31_24 = W*in
   wire signed [9:0] m31_24;
   assign m31_24 =10'b0;

   // m31_25 = W*in
   wire signed [9:0] m31_25;
   assign m31_25 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_26 = W*in
   wire signed [9:0] m31_26;
   assign m31_26 =10'b0;

   // m31_27 = W*in
   wire signed [9:0] m31_27;
   assign m31_27 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_28 = W*in
   wire signed [9:0] m31_28;
   assign m31_28 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_29 = W*in
   wire signed [9:0] m31_29;
   assign m31_29 ={ {4{in31[5]}} , in31[5:0] };

   // m31_30 = W*in
   wire signed [9:0] m31_30;
   assign m31_30 =10'b0;

   // m31_31 = W*in
   wire signed [9:0] m31_31;
   assign m31_31 ={ {5{in31[5]}} , in31[5:1] };

   // m31_32 = W*in
   wire signed [9:0] m31_32;
   assign m31_32 =10'b0;

   // m31_33 = W*in
   wire signed [9:0] m31_33;
   assign m31_33 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_34 = W*in
   wire signed [9:0] m31_34;
   assign m31_34 =10'b0;

   // m31_35 = W*in
   wire signed [9:0] m31_35;
   assign m31_35 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_36 = W*in
   wire signed [9:0] m31_36;
   assign m31_36 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_37 = W*in
   wire signed [9:0] m31_37;
   assign m31_37 =10'b0;

   // m31_38 = W*in
   wire signed [9:0] m31_38;
   assign m31_38 =10'b0;

   // m31_39 = W*in
   wire signed [9:0] m31_39;
   assign m31_39 =10'b0;

   // m31_40 = W*in
   wire signed [9:0] m31_40;
   assign m31_40 =10'b0;

   // m31_41 = W*in
   wire signed [9:0] m31_41;
   assign m31_41 =10'b0;

   // m31_42 = W*in
   wire signed [9:0] m31_42;
   assign m31_42 =10'b0;

   // m31_43 = W*in
   wire signed [9:0] m31_43;
   assign m31_43 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_44 = W*in
   wire signed [9:0] m31_44;
   assign m31_44 =10'b0;

   // m31_45 = W*in
   wire signed [9:0] m31_45;
   assign m31_45 =10'b0;

   // m31_46 = W*in
   wire signed [9:0] m31_46;
   assign m31_46 =10'b0;

   // m31_47 = W*in
   wire signed [9:0] m31_47;
   assign m31_47 =10'b0;

   // m31_48 = W*in
   wire signed [9:0] m31_48;
   assign m31_48 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_49 = W*in
   wire signed [9:0] m31_49;
   assign m31_49 =10'b0;

   // m31_50 = W*in
   wire signed [9:0] m31_50;
   assign m31_50 =10'b0;

   // m31_51 = W*in
   wire signed [9:0] m31_51;
   assign m31_51 =10'b0;

   // m31_52 = W*in
   wire signed [9:0] m31_52;
   assign m31_52 ={ {4{in31[5]}} , in31[5:0] };

   // m31_53 = W*in
   wire signed [9:0] m31_53;
   assign m31_53 ={ {4{in31[5]}} , in31[5:0] };

   // m31_54 = W*in
   wire signed [9:0] m31_54;
   assign m31_54 =10'b0;

   // m31_55 = W*in
   wire signed [9:0] m31_55;
   assign m31_55 =10'b0;

   // m31_56 = W*in
   wire signed [9:0] m31_56;
   assign m31_56 =10'b0;

   // m31_57 = W*in
   wire signed [9:0] m31_57;
   assign m31_57 =10'b0;

   // m31_58 = W*in
   wire signed [9:0] m31_58;
   assign m31_58 =10'b0;

   // m31_59 = W*in
   wire signed [9:0] m31_59;
   assign m31_59 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_60 = W*in
   wire signed [9:0] m31_60;
   assign m31_60 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_61 = W*in
   wire signed [9:0] m31_61;
   assign m31_61 =10'b0;

   // m31_62 = W*in
   wire signed [9:0] m31_62;
   assign m31_62 =10'b0;

   // m31_63 = W*in
   wire signed [9:0] m31_63;
   assign m31_63 =10'b0;

   // m31_64 = W*in
   wire signed [9:0] m31_64;
   assign m31_64 =10'b0;

   // m31_65 = W*in
   wire signed [9:0] m31_65;
   assign m31_65 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_66 = W*in
   wire signed [9:0] m31_66;
   assign m31_66 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_67 = W*in
   wire signed [9:0] m31_67;
   assign m31_67 =10'b0;

   // m31_68 = W*in
   wire signed [9:0] m31_68;
   assign m31_68 =10'b0;

   // m31_69 = W*in
   wire signed [9:0] m31_69;
   assign m31_69 ={ {5{in31[5]}} , in31[5:1] };

   // m31_70 = W*in
   wire signed [9:0] m31_70;
   assign m31_70 ={ {5{in31[5]}} , in31[5:1] };

   // m31_71 = W*in
   wire signed [9:0] m31_71;
   assign m31_71 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_72 = W*in
   wire signed [9:0] m31_72;
   assign m31_72 =10'b0;

   // m31_73 = W*in
   wire signed [9:0] m31_73;
   assign m31_73 =10'b0;

   // m31_74 = W*in
   wire signed [9:0] m31_74;
   assign m31_74 =10'b0;

   // m31_75 = W*in
   wire signed [9:0] m31_75;
   assign m31_75 ={ {5{neg31[5]}} , neg31[5:1] };

   // m31_76 = W*in
   wire signed [9:0] m31_76;
   assign m31_76 ={ {4{in31[5]}} , in31[5:0] };

   // m31_77 = W*in
   wire signed [9:0] m31_77;
   assign m31_77 ={ {4{in31[5]}} , in31[5:0] };

   // m31_78 = W*in
   wire signed [9:0] m31_78;
   assign m31_78 =10'b0;

   // m31_79 = W*in
   wire signed [9:0] m31_79;
   assign m31_79 =10'b0;

   // m31_80 = W*in
   wire signed [9:0] m31_80;
   assign m31_80 =10'b0;

   // m31_81 = W*in
   wire signed [9:0] m31_81;
   assign m31_81 =10'b0;

   // m31_82 = W*in
   wire signed [9:0] m31_82;
   assign m31_82 =10'b0;

   // m31_83 = W*in
   wire signed [9:0] m31_83;
   assign m31_83 =10'b0;

   // m31_84 = W*in
   wire signed [9:0] m31_84;
   assign m31_84 =10'b0;

   // m31_85 = W*in
   wire signed [9:0] m31_85;
   assign m31_85 ={ {4{in31[5]}} , in31[5:0] };

   // m31_86 = W*in
   wire signed [9:0] m31_86;
   assign m31_86 =10'b0;

   // m31_87 = W*in
   wire signed [9:0] m31_87;
   assign m31_87 =10'b0;

   // m31_88 = W*in
   wire signed [9:0] m31_88;
   assign m31_88 =10'b0;

   // m31_89 = W*in
   wire signed [9:0] m31_89;
   assign m31_89 =10'b0;

   // m31_90 = W*in
   wire signed [9:0] m31_90;
   assign m31_90 =10'b0;

   // m31_91 = W*in
   wire signed [9:0] m31_91;
   assign m31_91 =10'b0;

   // m31_92 = W*in
   wire signed [9:0] m31_92;
   assign m31_92 =10'b0;

   // m31_93 = W*in
   wire signed [9:0] m31_93;
   assign m31_93 =10'b0;

   // m31_94 = W*in
   wire signed [9:0] m31_94;
   assign m31_94 =10'b0;

   // m31_95 = W*in
   wire signed [9:0] m31_95;
   assign m31_95 =10'b0;

   // m31_96 = W*in
   wire signed [9:0] m31_96;
   assign m31_96 =10'b0;

   // m31_97 = W*in
   wire signed [9:0] m31_97;
   assign m31_97 =10'b0;

   // m31_98 = W*in
   wire signed [9:0] m31_98;
   assign m31_98 ={ {4{in31[5]}} , in31[5:0] };

   // m31_99 = W*in
   wire signed [9:0] m31_99;
   assign m31_99 =10'b0;

   // m31_100 = W*in
   wire signed [9:0] m31_100;
   assign m31_100 =10'b0;

   // m31_101 = W*in
   wire signed [9:0] m31_101;
   assign m31_101 =10'b0;

   // m31_102 = W*in
   wire signed [9:0] m31_102;
   assign m31_102 =10'b0;

   // m31_103 = W*in
   wire signed [9:0] m31_103;
   assign m31_103 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_104 = W*in
   wire signed [9:0] m31_104;
   assign m31_104 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_105 = W*in
   wire signed [9:0] m31_105;
   assign m31_105 =10'b0;

   // m31_106 = W*in
   wire signed [9:0] m31_106;
   assign m31_106 =10'b0;

   // m31_107 = W*in
   wire signed [9:0] m31_107;
   assign m31_107 =10'b0;

   // m31_108 = W*in
   wire signed [9:0] m31_108;
   assign m31_108 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_109 = W*in
   wire signed [9:0] m31_109;
   assign m31_109 ={ {4{neg31[5]}} , neg31[5:0] };

   // m31_110 = W*in
   wire signed [9:0] m31_110;
   assign m31_110 =10'b0;

   // m31_111 = W*in
   wire signed [9:0] m31_111;
   assign m31_111 =10'b0;

   // m31_112 = W*in
   wire signed [9:0] m31_112;
   assign m31_112 =10'b0;

   // m31_113 = W*in
   wire signed [9:0] m31_113;
   assign m31_113 =10'b0;

   // m31_114 = W*in
   wire signed [9:0] m31_114;
   assign m31_114 =10'b0;

   // m31_115 = W*in
   wire signed [9:0] m31_115;
   assign m31_115 =10'b0;

   // m31_116 = W*in
   wire signed [9:0] m31_116;
   assign m31_116 =10'b0;

   // m31_117 = W*in
   wire signed [9:0] m31_117;
   assign m31_117 ={ {4{neg31[5]}} , neg31[5:0] };

   // m32_1 = W*in
   wire signed [9:0] m32_1;
   assign m32_1 =10'b0;

   // m32_2 = W*in
   wire signed [9:0] m32_2;
   assign m32_2 ={ {4{in32[5]}} , in32[5:0] };

   // m32_3 = W*in
   wire signed [9:0] m32_3;
   assign m32_3 ={ {4{in32[5]}} , in32[5:0] };

   // m32_4 = W*in
   wire signed [9:0] m32_4;
   assign m32_4 =10'b0;

   // m32_5 = W*in
   wire signed [9:0] m32_5;
   assign m32_5 ={ {4{in32[5]}} , in32[5:0] };

   // m32_6 = W*in
   wire signed [9:0] m32_6;
   assign m32_6 =10'b0;

   // m32_7 = W*in
   wire signed [9:0] m32_7;
   assign m32_7 =10'b0;

   // m32_8 = W*in
   wire signed [9:0] m32_8;
   assign m32_8 ={ {4{in32[5]}} , in32[5:0] };

   // m32_9 = W*in
   wire signed [9:0] m32_9;
   assign m32_9 =10'b0;

   // m32_10 = W*in
   wire signed [9:0] m32_10;
   assign m32_10 =10'b0;

   // m32_11 = W*in
   wire signed [9:0] m32_11;
   assign m32_11 =10'b0;

   // m32_12 = W*in
   wire signed [9:0] m32_12;
   assign m32_12 =10'b0;

   // m32_13 = W*in
   wire signed [9:0] m32_13;
   assign m32_13 ={ {4{in32[5]}} , in32[5:0] };

   // m32_14 = W*in
   wire signed [9:0] m32_14;
   assign m32_14 =10'b0;

   // m32_15 = W*in
   wire signed [9:0] m32_15;
   assign m32_15 =10'b0;

   // m32_16 = W*in
   wire signed [9:0] m32_16;
   assign m32_16 =10'b0;

   // m32_17 = W*in
   wire signed [9:0] m32_17;
   assign m32_17 ={ {5{in32[5]}} , in32[5:1] };

   // m32_18 = W*in
   wire signed [9:0] m32_18;
   assign m32_18 =10'b0;

   // m32_19 = W*in
   wire signed [9:0] m32_19;
   assign m32_19 ={ {5{in32[5]}} , in32[5:1] };

   // m32_20 = W*in
   wire signed [9:0] m32_20;
   assign m32_20 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_21 = W*in
   wire signed [9:0] m32_21;
   assign m32_21 =10'b0;

   // m32_22 = W*in
   wire signed [9:0] m32_22;
   assign m32_22 =10'b0;

   // m32_23 = W*in
   wire signed [9:0] m32_23;
   assign m32_23 =10'b0;

   // m32_24 = W*in
   wire signed [9:0] m32_24;
   assign m32_24 =10'b0;

   // m32_25 = W*in
   wire signed [9:0] m32_25;
   assign m32_25 =10'b0;

   // m32_26 = W*in
   wire signed [9:0] m32_26;
   assign m32_26 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_27 = W*in
   wire signed [9:0] m32_27;
   assign m32_27 =10'b0;

   // m32_28 = W*in
   wire signed [9:0] m32_28;
   assign m32_28 =10'b0;

   // m32_29 = W*in
   wire signed [9:0] m32_29;
   assign m32_29 ={ {4{in32[5]}} , in32[5:0] };

   // m32_30 = W*in
   wire signed [9:0] m32_30;
   assign m32_30 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_31 = W*in
   wire signed [9:0] m32_31;
   assign m32_31 ={ {4{in32[5]}} , in32[5:0] };

   // m32_32 = W*in
   wire signed [9:0] m32_32;
   assign m32_32 =10'b0;

   // m32_33 = W*in
   wire signed [9:0] m32_33;
   assign m32_33 =10'b0;

   // m32_34 = W*in
   wire signed [9:0] m32_34;
   assign m32_34 =10'b0;

   // m32_35 = W*in
   wire signed [9:0] m32_35;
   assign m32_35 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_36 = W*in
   wire signed [9:0] m32_36;
   assign m32_36 =10'b0;

   // m32_37 = W*in
   wire signed [9:0] m32_37;
   assign m32_37 =10'b0;

   // m32_38 = W*in
   wire signed [9:0] m32_38;
   assign m32_38 =10'b0;

   // m32_39 = W*in
   wire signed [9:0] m32_39;
   assign m32_39 =10'b0;

   // m32_40 = W*in
   wire signed [9:0] m32_40;
   assign m32_40 =10'b0;

   // m32_41 = W*in
   wire signed [9:0] m32_41;
   assign m32_41 =10'b0;

   // m32_42 = W*in
   wire signed [9:0] m32_42;
   assign m32_42 =10'b0;

   // m32_43 = W*in
   wire signed [9:0] m32_43;
   assign m32_43 =10'b0;

   // m32_44 = W*in
   wire signed [9:0] m32_44;
   assign m32_44 =10'b0;

   // m32_45 = W*in
   wire signed [9:0] m32_45;
   assign m32_45 =10'b0;

   // m32_46 = W*in
   wire signed [9:0] m32_46;
   assign m32_46 =10'b0;

   // m32_47 = W*in
   wire signed [9:0] m32_47;
   assign m32_47 =10'b0;

   // m32_48 = W*in
   wire signed [9:0] m32_48;
   assign m32_48 =10'b0;

   // m32_49 = W*in
   wire signed [9:0] m32_49;
   assign m32_49 =10'b0;

   // m32_50 = W*in
   wire signed [9:0] m32_50;
   assign m32_50 =10'b0;

   // m32_51 = W*in
   wire signed [9:0] m32_51;
   assign m32_51 ={ {4{in32[5]}} , in32[5:0] };

   // m32_52 = W*in
   wire signed [9:0] m32_52;
   assign m32_52 ={ {4{in32[5]}} , in32[5:0] };

   // m32_53 = W*in
   wire signed [9:0] m32_53;
   assign m32_53 ={ {4{in32[5]}} , in32[5:0] };

   // m32_54 = W*in
   wire signed [9:0] m32_54;
   assign m32_54 =10'b0;

   // m32_55 = W*in
   wire signed [9:0] m32_55;
   assign m32_55 =10'b0;

   // m32_56 = W*in
   wire signed [9:0] m32_56;
   assign m32_56 =10'b0;

   // m32_57 = W*in
   wire signed [9:0] m32_57;
   assign m32_57 =10'b0;

   // m32_58 = W*in
   wire signed [9:0] m32_58;
   assign m32_58 =10'b0;

   // m32_59 = W*in
   wire signed [9:0] m32_59;
   assign m32_59 =10'b0;

   // m32_60 = W*in
   wire signed [9:0] m32_60;
   assign m32_60 =10'b0;

   // m32_61 = W*in
   wire signed [9:0] m32_61;
   assign m32_61 =10'b0;

   // m32_62 = W*in
   wire signed [9:0] m32_62;
   assign m32_62 =10'b0;

   // m32_63 = W*in
   wire signed [9:0] m32_63;
   assign m32_63 =10'b0;

   // m32_64 = W*in
   wire signed [9:0] m32_64;
   assign m32_64 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_65 = W*in
   wire signed [9:0] m32_65;
   assign m32_65 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_66 = W*in
   wire signed [9:0] m32_66;
   assign m32_66 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_67 = W*in
   wire signed [9:0] m32_67;
   assign m32_67 ={ {4{in32[5]}} , in32[5:0] };

   // m32_68 = W*in
   wire signed [9:0] m32_68;
   assign m32_68 =10'b0;

   // m32_69 = W*in
   wire signed [9:0] m32_69;
   assign m32_69 =10'b0;

   // m32_70 = W*in
   wire signed [9:0] m32_70;
   assign m32_70 =10'b0;

   // m32_71 = W*in
   wire signed [9:0] m32_71;
   assign m32_71 =10'b0;

   // m32_72 = W*in
   wire signed [9:0] m32_72;
   assign m32_72 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_73 = W*in
   wire signed [9:0] m32_73;
   assign m32_73 ={ {4{in32[5]}} , in32[5:0] };

   // m32_74 = W*in
   wire signed [9:0] m32_74;
   assign m32_74 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_75 = W*in
   wire signed [9:0] m32_75;
   assign m32_75 =10'b0;

   // m32_76 = W*in
   wire signed [9:0] m32_76;
   assign m32_76 =10'b0;

   // m32_77 = W*in
   wire signed [9:0] m32_77;
   assign m32_77 =10'b0;

   // m32_78 = W*in
   wire signed [9:0] m32_78;
   assign m32_78 =10'b0;

   // m32_79 = W*in
   wire signed [9:0] m32_79;
   assign m32_79 =10'b0;

   // m32_80 = W*in
   wire signed [9:0] m32_80;
   assign m32_80 ={ {4{in32[5]}} , in32[5:0] };

   // m32_81 = W*in
   wire signed [9:0] m32_81;
   assign m32_81 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_82 = W*in
   wire signed [9:0] m32_82;
   assign m32_82 =10'b0;

   // m32_83 = W*in
   wire signed [9:0] m32_83;
   assign m32_83 =10'b0;

   // m32_84 = W*in
   wire signed [9:0] m32_84;
   assign m32_84 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_85 = W*in
   wire signed [9:0] m32_85;
   assign m32_85 =10'b0;

   // m32_86 = W*in
   wire signed [9:0] m32_86;
   assign m32_86 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_87 = W*in
   wire signed [9:0] m32_87;
   assign m32_87 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_88 = W*in
   wire signed [9:0] m32_88;
   assign m32_88 =10'b0;

   // m32_89 = W*in
   wire signed [9:0] m32_89;
   assign m32_89 =10'b0;

   // m32_90 = W*in
   wire signed [9:0] m32_90;
   assign m32_90 =10'b0;

   // m32_91 = W*in
   wire signed [9:0] m32_91;
   assign m32_91 =10'b0;

   // m32_92 = W*in
   wire signed [9:0] m32_92;
   assign m32_92 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_93 = W*in
   wire signed [9:0] m32_93;
   assign m32_93 =10'b0;

   // m32_94 = W*in
   wire signed [9:0] m32_94;
   assign m32_94 =10'b0;

   // m32_95 = W*in
   wire signed [9:0] m32_95;
   assign m32_95 =10'b0;

   // m32_96 = W*in
   wire signed [9:0] m32_96;
   assign m32_96 =10'b0;

   // m32_97 = W*in
   wire signed [9:0] m32_97;
   assign m32_97 =10'b0;

   // m32_98 = W*in
   wire signed [9:0] m32_98;
   assign m32_98 ={ {4{in32[5]}} , in32[5:0] };

   // m32_99 = W*in
   wire signed [9:0] m32_99;
   assign m32_99 =10'b0;

   // m32_100 = W*in
   wire signed [9:0] m32_100;
   assign m32_100 =10'b0;

   // m32_101 = W*in
   wire signed [9:0] m32_101;
   assign m32_101 =10'b0;

   // m32_102 = W*in
   wire signed [9:0] m32_102;
   assign m32_102 =10'b0;

   // m32_103 = W*in
   wire signed [9:0] m32_103;
   assign m32_103 =10'b0;

   // m32_104 = W*in
   wire signed [9:0] m32_104;
   assign m32_104 =10'b0;

   // m32_105 = W*in
   wire signed [9:0] m32_105;
   assign m32_105 ={ {4{in32[5]}} , in32[5:0] };

   // m32_106 = W*in
   wire signed [9:0] m32_106;
   assign m32_106 =10'b0;

   // m32_107 = W*in
   wire signed [9:0] m32_107;
   assign m32_107 ={ {4{in32[5]}} , in32[5:0] };

   // m32_108 = W*in
   wire signed [9:0] m32_108;
   assign m32_108 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_109 = W*in
   wire signed [9:0] m32_109;
   assign m32_109 =10'b0;

   // m32_110 = W*in
   wire signed [9:0] m32_110;
   assign m32_110 ={ {4{neg32[5]}} , neg32[5:0] };

   // m32_111 = W*in
   wire signed [9:0] m32_111;
   assign m32_111 =10'b0;

   // m32_112 = W*in
   wire signed [9:0] m32_112;
   assign m32_112 =10'b0;

   // m32_113 = W*in
   wire signed [9:0] m32_113;
   assign m32_113 =10'b0;

   // m32_114 = W*in
   wire signed [9:0] m32_114;
   assign m32_114 =10'b0;

   // m32_115 = W*in
   wire signed [9:0] m32_115;
   assign m32_115 =10'b0;

   // m32_116 = W*in
   wire signed [9:0] m32_116;
   assign m32_116 ={ {5{neg32[5]}} , neg32[5:1] };

   // m32_117 = W*in
   wire signed [9:0] m32_117;
   assign m32_117 =10'b0;

   // m33_1 = W*in
   wire signed [9:0] m33_1;
   assign m33_1 =10'b0;

   // m33_2 = W*in
   wire signed [9:0] m33_2;
   assign m33_2 =10'b0;

   // m33_3 = W*in
   wire signed [9:0] m33_3;
   assign m33_3 =10'b0;

   // m33_4 = W*in
   wire signed [9:0] m33_4;
   assign m33_4 =10'b0;

   // m33_5 = W*in
   wire signed [9:0] m33_5;
   assign m33_5 =10'b0;

   // m33_6 = W*in
   wire signed [9:0] m33_6;
   assign m33_6 =10'b0;

   // m33_7 = W*in
   wire signed [9:0] m33_7;
   assign m33_7 =10'b0;

   // m33_8 = W*in
   wire signed [9:0] m33_8;
   assign m33_8 =10'b0;

   // m33_9 = W*in
   wire signed [9:0] m33_9;
   assign m33_9 =10'b0;

   // m33_10 = W*in
   wire signed [9:0] m33_10;
   assign m33_10 =10'b0;

   // m33_11 = W*in
   wire signed [9:0] m33_11;
   assign m33_11 =10'b0;

   // m33_12 = W*in
   wire signed [9:0] m33_12;
   assign m33_12 =10'b0;

   // m33_13 = W*in
   wire signed [9:0] m33_13;
   assign m33_13 =10'b0;

   // m33_14 = W*in
   wire signed [9:0] m33_14;
   assign m33_14 =10'b0;

   // m33_15 = W*in
   wire signed [9:0] m33_15;
   assign m33_15 =10'b0;

   // m33_16 = W*in
   wire signed [9:0] m33_16;
   assign m33_16 =10'b0;

   // m33_17 = W*in
   wire signed [9:0] m33_17;
   assign m33_17 =10'b0;

   // m33_18 = W*in
   wire signed [9:0] m33_18;
   assign m33_18 =10'b0;

   // m33_19 = W*in
   wire signed [9:0] m33_19;
   assign m33_19 =10'b0;

   // m33_20 = W*in
   wire signed [9:0] m33_20;
   assign m33_20 =10'b0;

   // m33_21 = W*in
   wire signed [9:0] m33_21;
   assign m33_21 =10'b0;

   // m33_22 = W*in
   wire signed [9:0] m33_22;
   assign m33_22 =10'b0;

   // m33_23 = W*in
   wire signed [9:0] m33_23;
   assign m33_23 =10'b0;

   // m33_24 = W*in
   wire signed [9:0] m33_24;
   assign m33_24 =10'b0;

   // m33_25 = W*in
   wire signed [9:0] m33_25;
   assign m33_25 =10'b0;

   // m33_26 = W*in
   wire signed [9:0] m33_26;
   assign m33_26 =10'b0;

   // m33_27 = W*in
   wire signed [9:0] m33_27;
   assign m33_27 ={ {5{in33[5]}} , in33[5:1] };

   // m33_28 = W*in
   wire signed [9:0] m33_28;
   assign m33_28 =10'b0;

   // m33_29 = W*in
   wire signed [9:0] m33_29;
   assign m33_29 ={ {5{neg33[5]}} , neg33[5:1] };

   // m33_30 = W*in
   wire signed [9:0] m33_30;
   assign m33_30 =10'b0;

   // m33_31 = W*in
   wire signed [9:0] m33_31;
   assign m33_31 =10'b0;

   // m33_32 = W*in
   wire signed [9:0] m33_32;
   assign m33_32 =10'b0;

   // m33_33 = W*in
   wire signed [9:0] m33_33;
   assign m33_33 =10'b0;

   // m33_34 = W*in
   wire signed [9:0] m33_34;
   assign m33_34 =10'b0;

   // m33_35 = W*in
   wire signed [9:0] m33_35;
   assign m33_35 =10'b0;

   // m33_36 = W*in
   wire signed [9:0] m33_36;
   assign m33_36 ={ {5{in33[5]}} , in33[5:1] };

   // m33_37 = W*in
   wire signed [9:0] m33_37;
   assign m33_37 =10'b0;

   // m33_38 = W*in
   wire signed [9:0] m33_38;
   assign m33_38 =10'b0;

   // m33_39 = W*in
   wire signed [9:0] m33_39;
   assign m33_39 =10'b0;

   // m33_40 = W*in
   wire signed [9:0] m33_40;
   assign m33_40 =10'b0;

   // m33_41 = W*in
   wire signed [9:0] m33_41;
   assign m33_41 =10'b0;

   // m33_42 = W*in
   wire signed [9:0] m33_42;
   assign m33_42 =10'b0;

   // m33_43 = W*in
   wire signed [9:0] m33_43;
   assign m33_43 =10'b0;

   // m33_44 = W*in
   wire signed [9:0] m33_44;
   assign m33_44 =10'b0;

   // m33_45 = W*in
   wire signed [9:0] m33_45;
   assign m33_45 =10'b0;

   // m33_46 = W*in
   wire signed [9:0] m33_46;
   assign m33_46 =10'b0;

   // m33_47 = W*in
   wire signed [9:0] m33_47;
   assign m33_47 =10'b0;

   // m33_48 = W*in
   wire signed [9:0] m33_48;
   assign m33_48 =10'b0;

   // m33_49 = W*in
   wire signed [9:0] m33_49;
   assign m33_49 =10'b0;

   // m33_50 = W*in
   wire signed [9:0] m33_50;
   assign m33_50 =10'b0;

   // m33_51 = W*in
   wire signed [9:0] m33_51;
   assign m33_51 =10'b0;

   // m33_52 = W*in
   wire signed [9:0] m33_52;
   assign m33_52 =10'b0;

   // m33_53 = W*in
   wire signed [9:0] m33_53;
   assign m33_53 =10'b0;

   // m33_54 = W*in
   wire signed [9:0] m33_54;
   assign m33_54 =10'b0;

   // m33_55 = W*in
   wire signed [9:0] m33_55;
   assign m33_55 =10'b0;

   // m33_56 = W*in
   wire signed [9:0] m33_56;
   assign m33_56 =10'b0;

   // m33_57 = W*in
   wire signed [9:0] m33_57;
   assign m33_57 =10'b0;

   // m33_58 = W*in
   wire signed [9:0] m33_58;
   assign m33_58 =10'b0;

   // m33_59 = W*in
   wire signed [9:0] m33_59;
   assign m33_59 =10'b0;

   // m33_60 = W*in
   wire signed [9:0] m33_60;
   assign m33_60 =10'b0;

   // m33_61 = W*in
   wire signed [9:0] m33_61;
   assign m33_61 =10'b0;

   // m33_62 = W*in
   wire signed [9:0] m33_62;
   assign m33_62 =10'b0;

   // m33_63 = W*in
   wire signed [9:0] m33_63;
   assign m33_63 =10'b0;

   // m33_64 = W*in
   wire signed [9:0] m33_64;
   assign m33_64 =10'b0;

   // m33_65 = W*in
   wire signed [9:0] m33_65;
   assign m33_65 =10'b0;

   // m33_66 = W*in
   wire signed [9:0] m33_66;
   assign m33_66 =10'b0;

   // m33_67 = W*in
   wire signed [9:0] m33_67;
   assign m33_67 =10'b0;

   // m33_68 = W*in
   wire signed [9:0] m33_68;
   assign m33_68 =10'b0;

   // m33_69 = W*in
   wire signed [9:0] m33_69;
   assign m33_69 =10'b0;

   // m33_70 = W*in
   wire signed [9:0] m33_70;
   assign m33_70 =10'b0;

   // m33_71 = W*in
   wire signed [9:0] m33_71;
   assign m33_71 =10'b0;

   // m33_72 = W*in
   wire signed [9:0] m33_72;
   assign m33_72 =10'b0;

   // m33_73 = W*in
   wire signed [9:0] m33_73;
   assign m33_73 =10'b0;

   // m33_74 = W*in
   wire signed [9:0] m33_74;
   assign m33_74 =10'b0;

   // m33_75 = W*in
   wire signed [9:0] m33_75;
   assign m33_75 =10'b0;

   // m33_76 = W*in
   wire signed [9:0] m33_76;
   assign m33_76 =10'b0;

   // m33_77 = W*in
   wire signed [9:0] m33_77;
   assign m33_77 =10'b0;

   // m33_78 = W*in
   wire signed [9:0] m33_78;
   assign m33_78 =10'b0;

   // m33_79 = W*in
   wire signed [9:0] m33_79;
   assign m33_79 =10'b0;

   // m33_80 = W*in
   wire signed [9:0] m33_80;
   assign m33_80 =10'b0;

   // m33_81 = W*in
   wire signed [9:0] m33_81;
   assign m33_81 =10'b0;

   // m33_82 = W*in
   wire signed [9:0] m33_82;
   assign m33_82 =10'b0;

   // m33_83 = W*in
   wire signed [9:0] m33_83;
   assign m33_83 =10'b0;

   // m33_84 = W*in
   wire signed [9:0] m33_84;
   assign m33_84 =10'b0;

   // m33_85 = W*in
   wire signed [9:0] m33_85;
   assign m33_85 =10'b0;

   // m33_86 = W*in
   wire signed [9:0] m33_86;
   assign m33_86 =10'b0;

   // m33_87 = W*in
   wire signed [9:0] m33_87;
   assign m33_87 =10'b0;

   // m33_88 = W*in
   wire signed [9:0] m33_88;
   assign m33_88 =10'b0;

   // m33_89 = W*in
   wire signed [9:0] m33_89;
   assign m33_89 =10'b0;

   // m33_90 = W*in
   wire signed [9:0] m33_90;
   assign m33_90 =10'b0;

   // m33_91 = W*in
   wire signed [9:0] m33_91;
   assign m33_91 =10'b0;

   // m33_92 = W*in
   wire signed [9:0] m33_92;
   assign m33_92 =10'b0;

   // m33_93 = W*in
   wire signed [9:0] m33_93;
   assign m33_93 =10'b0;

   // m33_94 = W*in
   wire signed [9:0] m33_94;
   assign m33_94 =10'b0;

   // m33_95 = W*in
   wire signed [9:0] m33_95;
   assign m33_95 =10'b0;

   // m33_96 = W*in
   wire signed [9:0] m33_96;
   assign m33_96 =10'b0;

   // m33_97 = W*in
   wire signed [9:0] m33_97;
   assign m33_97 =10'b0;

   // m33_98 = W*in
   wire signed [9:0] m33_98;
   assign m33_98 =10'b0;

   // m33_99 = W*in
   wire signed [9:0] m33_99;
   assign m33_99 =10'b0;

   // m33_100 = W*in
   wire signed [9:0] m33_100;
   assign m33_100 =10'b0;

   // m33_101 = W*in
   wire signed [9:0] m33_101;
   assign m33_101 =10'b0;

   // m33_102 = W*in
   wire signed [9:0] m33_102;
   assign m33_102 =10'b0;

   // m33_103 = W*in
   wire signed [9:0] m33_103;
   assign m33_103 =10'b0;

   // m33_104 = W*in
   wire signed [9:0] m33_104;
   assign m33_104 =10'b0;

   // m33_105 = W*in
   wire signed [9:0] m33_105;
   assign m33_105 =10'b0;

   // m33_106 = W*in
   wire signed [9:0] m33_106;
   assign m33_106 =10'b0;

   // m33_107 = W*in
   wire signed [9:0] m33_107;
   assign m33_107 =10'b0;

   // m33_108 = W*in
   wire signed [9:0] m33_108;
   assign m33_108 =10'b0;

   // m33_109 = W*in
   wire signed [9:0] m33_109;
   assign m33_109 =10'b0;

   // m33_110 = W*in
   wire signed [9:0] m33_110;
   assign m33_110 =10'b0;

   // m33_111 = W*in
   wire signed [9:0] m33_111;
   assign m33_111 =10'b0;

   // m33_112 = W*in
   wire signed [9:0] m33_112;
   assign m33_112 =10'b0;

   // m33_113 = W*in
   wire signed [9:0] m33_113;
   assign m33_113 =10'b0;

   // m33_114 = W*in
   wire signed [9:0] m33_114;
   assign m33_114 =10'b0;

   // m33_115 = W*in
   wire signed [9:0] m33_115;
   assign m33_115 =10'b0;

   // m33_116 = W*in
   wire signed [9:0] m33_116;
   assign m33_116 =10'b0;

   // m33_117 = W*in
   wire signed [9:0] m33_117;
   assign m33_117 =10'b0;

   // m34_1 = W*in
   wire signed [9:0] m34_1;
   assign m34_1 =10'b0;

   // m34_2 = W*in
   wire signed [9:0] m34_2;
   assign m34_2 =10'b0;

   // m34_3 = W*in
   wire signed [9:0] m34_3;
   assign m34_3 =10'b0;

   // m34_4 = W*in
   wire signed [9:0] m34_4;
   assign m34_4 =10'b0;

   // m34_5 = W*in
   wire signed [9:0] m34_5;
   assign m34_5 =10'b0;

   // m34_6 = W*in
   wire signed [9:0] m34_6;
   assign m34_6 =10'b0;

   // m34_7 = W*in
   wire signed [9:0] m34_7;
   assign m34_7 =10'b0;

   // m34_8 = W*in
   wire signed [9:0] m34_8;
   assign m34_8 ={ {4{in34[5]}} , in34[5:0] };

   // m34_9 = W*in
   wire signed [9:0] m34_9;
   assign m34_9 =10'b0;

   // m34_10 = W*in
   wire signed [9:0] m34_10;
   assign m34_10 ={ {4{neg34[5]}} , neg34[5:0] };

   // m34_11 = W*in
   wire signed [9:0] m34_11;
   assign m34_11 =10'b0;

   // m34_12 = W*in
   wire signed [9:0] m34_12;
   assign m34_12 =10'b0;

   // m34_13 = W*in
   wire signed [9:0] m34_13;
   assign m34_13 =10'b0;

   // m34_14 = W*in
   wire signed [9:0] m34_14;
   assign m34_14 =10'b0;

   // m34_15 = W*in
   wire signed [9:0] m34_15;
   assign m34_15 =10'b0;

   // m34_16 = W*in
   wire signed [9:0] m34_16;
   assign m34_16 =10'b0;

   // m34_17 = W*in
   wire signed [9:0] m34_17;
   assign m34_17 =10'b0;

   // m34_18 = W*in
   wire signed [9:0] m34_18;
   assign m34_18 =10'b0;

   // m34_19 = W*in
   wire signed [9:0] m34_19;
   assign m34_19 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_20 = W*in
   wire signed [9:0] m34_20;
   assign m34_20 ={ {5{in34[5]}} , in34[5:1] };

   // m34_21 = W*in
   wire signed [9:0] m34_21;
   assign m34_21 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_22 = W*in
   wire signed [9:0] m34_22;
   assign m34_22 =10'b0;

   // m34_23 = W*in
   wire signed [9:0] m34_23;
   assign m34_23 =10'b0;

   // m34_24 = W*in
   wire signed [9:0] m34_24;
   assign m34_24 =10'b0;

   // m34_25 = W*in
   wire signed [9:0] m34_25;
   assign m34_25 =10'b0;

   // m34_26 = W*in
   wire signed [9:0] m34_26;
   assign m34_26 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_27 = W*in
   wire signed [9:0] m34_27;
   assign m34_27 ={ {5{in34[5]}} , in34[5:1] };

   // m34_28 = W*in
   wire signed [9:0] m34_28;
   assign m34_28 =10'b0;

   // m34_29 = W*in
   wire signed [9:0] m34_29;
   assign m34_29 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_30 = W*in
   wire signed [9:0] m34_30;
   assign m34_30 =10'b0;

   // m34_31 = W*in
   wire signed [9:0] m34_31;
   assign m34_31 ={ {4{in34[5]}} , in34[5:0] };

   // m34_32 = W*in
   wire signed [9:0] m34_32;
   assign m34_32 =10'b0;

   // m34_33 = W*in
   wire signed [9:0] m34_33;
   assign m34_33 =10'b0;

   // m34_34 = W*in
   wire signed [9:0] m34_34;
   assign m34_34 ={ {4{in34[5]}} , in34[5:0] };

   // m34_35 = W*in
   wire signed [9:0] m34_35;
   assign m34_35 =10'b0;

   // m34_36 = W*in
   wire signed [9:0] m34_36;
   assign m34_36 =10'b0;

   // m34_37 = W*in
   wire signed [9:0] m34_37;
   assign m34_37 =10'b0;

   // m34_38 = W*in
   wire signed [9:0] m34_38;
   assign m34_38 =10'b0;

   // m34_39 = W*in
   wire signed [9:0] m34_39;
   assign m34_39 =10'b0;

   // m34_40 = W*in
   wire signed [9:0] m34_40;
   assign m34_40 =10'b0;

   // m34_41 = W*in
   wire signed [9:0] m34_41;
   assign m34_41 =10'b0;

   // m34_42 = W*in
   wire signed [9:0] m34_42;
   assign m34_42 =10'b0;

   // m34_43 = W*in
   wire signed [9:0] m34_43;
   assign m34_43 =10'b0;

   // m34_44 = W*in
   wire signed [9:0] m34_44;
   assign m34_44 =10'b0;

   // m34_45 = W*in
   wire signed [9:0] m34_45;
   assign m34_45 =10'b0;

   // m34_46 = W*in
   wire signed [9:0] m34_46;
   assign m34_46 =10'b0;

   // m34_47 = W*in
   wire signed [9:0] m34_47;
   assign m34_47 =10'b0;

   // m34_48 = W*in
   wire signed [9:0] m34_48;
   assign m34_48 =10'b0;

   // m34_49 = W*in
   wire signed [9:0] m34_49;
   assign m34_49 =10'b0;

   // m34_50 = W*in
   wire signed [9:0] m34_50;
   assign m34_50 =10'b0;

   // m34_51 = W*in
   wire signed [9:0] m34_51;
   assign m34_51 =10'b0;

   // m34_52 = W*in
   wire signed [9:0] m34_52;
   assign m34_52 ={ {4{in34[5]}} , in34[5:0] };

   // m34_53 = W*in
   wire signed [9:0] m34_53;
   assign m34_53 =10'b0;

   // m34_54 = W*in
   wire signed [9:0] m34_54;
   assign m34_54 =10'b0;

   // m34_55 = W*in
   wire signed [9:0] m34_55;
   assign m34_55 =10'b0;

   // m34_56 = W*in
   wire signed [9:0] m34_56;
   assign m34_56 =10'b0;

   // m34_57 = W*in
   wire signed [9:0] m34_57;
   assign m34_57 =10'b0;

   // m34_58 = W*in
   wire signed [9:0] m34_58;
   assign m34_58 =10'b0;

   // m34_59 = W*in
   wire signed [9:0] m34_59;
   assign m34_59 =10'b0;

   // m34_60 = W*in
   wire signed [9:0] m34_60;
   assign m34_60 =10'b0;

   // m34_61 = W*in
   wire signed [9:0] m34_61;
   assign m34_61 =10'b0;

   // m34_62 = W*in
   wire signed [9:0] m34_62;
   assign m34_62 =10'b0;

   // m34_63 = W*in
   wire signed [9:0] m34_63;
   assign m34_63 =10'b0;

   // m34_64 = W*in
   wire signed [9:0] m34_64;
   assign m34_64 ={ {5{in34[5]}} , in34[5:1] };

   // m34_65 = W*in
   wire signed [9:0] m34_65;
   assign m34_65 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_66 = W*in
   wire signed [9:0] m34_66;
   assign m34_66 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_67 = W*in
   wire signed [9:0] m34_67;
   assign m34_67 =10'b0;

   // m34_68 = W*in
   wire signed [9:0] m34_68;
   assign m34_68 =10'b0;

   // m34_69 = W*in
   wire signed [9:0] m34_69;
   assign m34_69 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_70 = W*in
   wire signed [9:0] m34_70;
   assign m34_70 =10'b0;

   // m34_71 = W*in
   wire signed [9:0] m34_71;
   assign m34_71 =10'b0;

   // m34_72 = W*in
   wire signed [9:0] m34_72;
   assign m34_72 ={ {5{neg34[5]}} , neg34[5:1] };

   // m34_73 = W*in
   wire signed [9:0] m34_73;
   assign m34_73 ={ {5{in34[5]}} , in34[5:1] };

   // m34_74 = W*in
   wire signed [9:0] m34_74;
   assign m34_74 =10'b0;

   // m34_75 = W*in
   wire signed [9:0] m34_75;
   assign m34_75 =10'b0;

   // m34_76 = W*in
   wire signed [9:0] m34_76;
   assign m34_76 =10'b0;

   // m34_77 = W*in
   wire signed [9:0] m34_77;
   assign m34_77 =10'b0;

   // m34_78 = W*in
   wire signed [9:0] m34_78;
   assign m34_78 =10'b0;

   // m34_79 = W*in
   wire signed [9:0] m34_79;
   assign m34_79 =10'b0;

   // m34_80 = W*in
   wire signed [9:0] m34_80;
   assign m34_80 =10'b0;

   // m34_81 = W*in
   wire signed [9:0] m34_81;
   assign m34_81 =10'b0;

   // m34_82 = W*in
   wire signed [9:0] m34_82;
   assign m34_82 =10'b0;

   // m34_83 = W*in
   wire signed [9:0] m34_83;
   assign m34_83 =10'b0;

   // m34_84 = W*in
   wire signed [9:0] m34_84;
   assign m34_84 ={ {4{neg34[5]}} , neg34[5:0] };

   // m34_85 = W*in
   wire signed [9:0] m34_85;
   assign m34_85 =10'b0;

   // m34_86 = W*in
   wire signed [9:0] m34_86;
   assign m34_86 =10'b0;

   // m34_87 = W*in
   wire signed [9:0] m34_87;
   assign m34_87 =10'b0;

   // m34_88 = W*in
   wire signed [9:0] m34_88;
   assign m34_88 =10'b0;

   // m34_89 = W*in
   wire signed [9:0] m34_89;
   assign m34_89 =10'b0;

   // m34_90 = W*in
   wire signed [9:0] m34_90;
   assign m34_90 =10'b0;

   // m34_91 = W*in
   wire signed [9:0] m34_91;
   assign m34_91 =10'b0;

   // m34_92 = W*in
   wire signed [9:0] m34_92;
   assign m34_92 =10'b0;

   // m34_93 = W*in
   wire signed [9:0] m34_93;
   assign m34_93 =10'b0;

   // m34_94 = W*in
   wire signed [9:0] m34_94;
   assign m34_94 =10'b0;

   // m34_95 = W*in
   wire signed [9:0] m34_95;
   assign m34_95 =10'b0;

   // m34_96 = W*in
   wire signed [9:0] m34_96;
   assign m34_96 =10'b0;

   // m34_97 = W*in
   wire signed [9:0] m34_97;
   assign m34_97 =10'b0;

   // m34_98 = W*in
   wire signed [9:0] m34_98;
   assign m34_98 ={ {4{in34[5]}} , in34[5:0] };

   // m34_99 = W*in
   wire signed [9:0] m34_99;
   assign m34_99 =10'b0;

   // m34_100 = W*in
   wire signed [9:0] m34_100;
   assign m34_100 =10'b0;

   // m34_101 = W*in
   wire signed [9:0] m34_101;
   assign m34_101 =10'b0;

   // m34_102 = W*in
   wire signed [9:0] m34_102;
   assign m34_102 =10'b0;

   // m34_103 = W*in
   wire signed [9:0] m34_103;
   assign m34_103 =10'b0;

   // m34_104 = W*in
   wire signed [9:0] m34_104;
   assign m34_104 =10'b0;

   // m34_105 = W*in
   wire signed [9:0] m34_105;
   assign m34_105 =10'b0;

   // m34_106 = W*in
   wire signed [9:0] m34_106;
   assign m34_106 =10'b0;

   // m34_107 = W*in
   wire signed [9:0] m34_107;
   assign m34_107 =10'b0;

   // m34_108 = W*in
   wire signed [9:0] m34_108;
   assign m34_108 =10'b0;

   // m34_109 = W*in
   wire signed [9:0] m34_109;
   assign m34_109 =10'b0;

   // m34_110 = W*in
   wire signed [9:0] m34_110;
   assign m34_110 =10'b0;

   // m34_111 = W*in
   wire signed [9:0] m34_111;
   assign m34_111 =10'b0;

   // m34_112 = W*in
   wire signed [9:0] m34_112;
   assign m34_112 =10'b0;

   // m34_113 = W*in
   wire signed [9:0] m34_113;
   assign m34_113 =10'b0;

   // m34_114 = W*in
   wire signed [9:0] m34_114;
   assign m34_114 =10'b0;

   // m34_115 = W*in
   wire signed [9:0] m34_115;
   assign m34_115 =10'b0;

   // m34_116 = W*in
   wire signed [9:0] m34_116;
   assign m34_116 =10'b0;

   // m34_117 = W*in
   wire signed [9:0] m34_117;
   assign m34_117 =10'b0;

   // m35_1 = W*in
   wire signed [9:0] m35_1;
   assign m35_1 =10'b0;

   // m35_2 = W*in
   wire signed [9:0] m35_2;
   assign m35_2 =10'b0;

   // m35_3 = W*in
   wire signed [9:0] m35_3;
   assign m35_3 =10'b0;

   // m35_4 = W*in
   wire signed [9:0] m35_4;
   assign m35_4 =10'b0;

   // m35_5 = W*in
   wire signed [9:0] m35_5;
   assign m35_5 =10'b0;

   // m35_6 = W*in
   wire signed [9:0] m35_6;
   assign m35_6 =10'b0;

   // m35_7 = W*in
   wire signed [9:0] m35_7;
   assign m35_7 =10'b0;

   // m35_8 = W*in
   wire signed [9:0] m35_8;
   assign m35_8 =10'b0;

   // m35_9 = W*in
   wire signed [9:0] m35_9;
   assign m35_9 =10'b0;

   // m35_10 = W*in
   wire signed [9:0] m35_10;
   assign m35_10 =10'b0;

   // m35_11 = W*in
   wire signed [9:0] m35_11;
   assign m35_11 =10'b0;

   // m35_12 = W*in
   wire signed [9:0] m35_12;
   assign m35_12 =10'b0;

   // m35_13 = W*in
   wire signed [9:0] m35_13;
   assign m35_13 =10'b0;

   // m35_14 = W*in
   wire signed [9:0] m35_14;
   assign m35_14 =10'b0;

   // m35_15 = W*in
   wire signed [9:0] m35_15;
   assign m35_15 =10'b0;

   // m35_16 = W*in
   wire signed [9:0] m35_16;
   assign m35_16 =10'b0;

   // m35_17 = W*in
   wire signed [9:0] m35_17;
   assign m35_17 =10'b0;

   // m35_18 = W*in
   wire signed [9:0] m35_18;
   assign m35_18 =10'b0;

   // m35_19 = W*in
   wire signed [9:0] m35_19;
   assign m35_19 =10'b0;

   // m35_20 = W*in
   wire signed [9:0] m35_20;
   assign m35_20 =10'b0;

   // m35_21 = W*in
   wire signed [9:0] m35_21;
   assign m35_21 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_22 = W*in
   wire signed [9:0] m35_22;
   assign m35_22 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_23 = W*in
   wire signed [9:0] m35_23;
   assign m35_23 =10'b0;

   // m35_24 = W*in
   wire signed [9:0] m35_24;
   assign m35_24 =10'b0;

   // m35_25 = W*in
   wire signed [9:0] m35_25;
   assign m35_25 =10'b0;

   // m35_26 = W*in
   wire signed [9:0] m35_26;
   assign m35_26 =10'b0;

   // m35_27 = W*in
   wire signed [9:0] m35_27;
   assign m35_27 =10'b0;

   // m35_28 = W*in
   wire signed [9:0] m35_28;
   assign m35_28 =10'b0;

   // m35_29 = W*in
   wire signed [9:0] m35_29;
   assign m35_29 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_30 = W*in
   wire signed [9:0] m35_30;
   assign m35_30 =10'b0;

   // m35_31 = W*in
   wire signed [9:0] m35_31;
   assign m35_31 =10'b0;

   // m35_32 = W*in
   wire signed [9:0] m35_32;
   assign m35_32 =10'b0;

   // m35_33 = W*in
   wire signed [9:0] m35_33;
   assign m35_33 =10'b0;

   // m35_34 = W*in
   wire signed [9:0] m35_34;
   assign m35_34 =10'b0;

   // m35_35 = W*in
   wire signed [9:0] m35_35;
   assign m35_35 =10'b0;

   // m35_36 = W*in
   wire signed [9:0] m35_36;
   assign m35_36 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_37 = W*in
   wire signed [9:0] m35_37;
   assign m35_37 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_38 = W*in
   wire signed [9:0] m35_38;
   assign m35_38 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_39 = W*in
   wire signed [9:0] m35_39;
   assign m35_39 =10'b0;

   // m35_40 = W*in
   wire signed [9:0] m35_40;
   assign m35_40 =10'b0;

   // m35_41 = W*in
   wire signed [9:0] m35_41;
   assign m35_41 =10'b0;

   // m35_42 = W*in
   wire signed [9:0] m35_42;
   assign m35_42 ={ {4{in35[5]}} , in35[5:0] };

   // m35_43 = W*in
   wire signed [9:0] m35_43;
   assign m35_43 =10'b0;

   // m35_44 = W*in
   wire signed [9:0] m35_44;
   assign m35_44 =10'b0;

   // m35_45 = W*in
   wire signed [9:0] m35_45;
   assign m35_45 =10'b0;

   // m35_46 = W*in
   wire signed [9:0] m35_46;
   assign m35_46 =10'b0;

   // m35_47 = W*in
   wire signed [9:0] m35_47;
   assign m35_47 =10'b0;

   // m35_48 = W*in
   wire signed [9:0] m35_48;
   assign m35_48 =10'b0;

   // m35_49 = W*in
   wire signed [9:0] m35_49;
   assign m35_49 =10'b0;

   // m35_50 = W*in
   wire signed [9:0] m35_50;
   assign m35_50 =10'b0;

   // m35_51 = W*in
   wire signed [9:0] m35_51;
   assign m35_51 =10'b0;

   // m35_52 = W*in
   wire signed [9:0] m35_52;
   assign m35_52 =10'b0;

   // m35_53 = W*in
   wire signed [9:0] m35_53;
   assign m35_53 =10'b0;

   // m35_54 = W*in
   wire signed [9:0] m35_54;
   assign m35_54 =10'b0;

   // m35_55 = W*in
   wire signed [9:0] m35_55;
   assign m35_55 =10'b0;

   // m35_56 = W*in
   wire signed [9:0] m35_56;
   assign m35_56 =10'b0;

   // m35_57 = W*in
   wire signed [9:0] m35_57;
   assign m35_57 =10'b0;

   // m35_58 = W*in
   wire signed [9:0] m35_58;
   assign m35_58 =10'b0;

   // m35_59 = W*in
   wire signed [9:0] m35_59;
   assign m35_59 =10'b0;

   // m35_60 = W*in
   wire signed [9:0] m35_60;
   assign m35_60 =10'b0;

   // m35_61 = W*in
   wire signed [9:0] m35_61;
   assign m35_61 =10'b0;

   // m35_62 = W*in
   wire signed [9:0] m35_62;
   assign m35_62 =10'b0;

   // m35_63 = W*in
   wire signed [9:0] m35_63;
   assign m35_63 =10'b0;

   // m35_64 = W*in
   wire signed [9:0] m35_64;
   assign m35_64 ={ {4{in35[5]}} , in35[5:0] };

   // m35_65 = W*in
   wire signed [9:0] m35_65;
   assign m35_65 ={ {4{in35[5]}} , in35[5:0] };

   // m35_66 = W*in
   wire signed [9:0] m35_66;
   assign m35_66 =10'b0;

   // m35_67 = W*in
   wire signed [9:0] m35_67;
   assign m35_67 =10'b0;

   // m35_68 = W*in
   wire signed [9:0] m35_68;
   assign m35_68 =10'b0;

   // m35_69 = W*in
   wire signed [9:0] m35_69;
   assign m35_69 =10'b0;

   // m35_70 = W*in
   wire signed [9:0] m35_70;
   assign m35_70 =10'b0;

   // m35_71 = W*in
   wire signed [9:0] m35_71;
   assign m35_71 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_72 = W*in
   wire signed [9:0] m35_72;
   assign m35_72 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_73 = W*in
   wire signed [9:0] m35_73;
   assign m35_73 =10'b0;

   // m35_74 = W*in
   wire signed [9:0] m35_74;
   assign m35_74 =10'b0;

   // m35_75 = W*in
   wire signed [9:0] m35_75;
   assign m35_75 ={ {4{in35[5]}} , in35[5:0] };

   // m35_76 = W*in
   wire signed [9:0] m35_76;
   assign m35_76 =10'b0;

   // m35_77 = W*in
   wire signed [9:0] m35_77;
   assign m35_77 =10'b0;

   // m35_78 = W*in
   wire signed [9:0] m35_78;
   assign m35_78 =10'b0;

   // m35_79 = W*in
   wire signed [9:0] m35_79;
   assign m35_79 =10'b0;

   // m35_80 = W*in
   wire signed [9:0] m35_80;
   assign m35_80 =10'b0;

   // m35_81 = W*in
   wire signed [9:0] m35_81;
   assign m35_81 ={ {5{in35[5]}} , in35[5:1] };

   // m35_82 = W*in
   wire signed [9:0] m35_82;
   assign m35_82 =10'b0;

   // m35_83 = W*in
   wire signed [9:0] m35_83;
   assign m35_83 =10'b0;

   // m35_84 = W*in
   wire signed [9:0] m35_84;
   assign m35_84 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_85 = W*in
   wire signed [9:0] m35_85;
   assign m35_85 ={ {5{neg35[5]}} , neg35[5:1] };

   // m35_86 = W*in
   wire signed [9:0] m35_86;
   assign m35_86 =10'b0;

   // m35_87 = W*in
   wire signed [9:0] m35_87;
   assign m35_87 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_88 = W*in
   wire signed [9:0] m35_88;
   assign m35_88 =10'b0;

   // m35_89 = W*in
   wire signed [9:0] m35_89;
   assign m35_89 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_90 = W*in
   wire signed [9:0] m35_90;
   assign m35_90 =10'b0;

   // m35_91 = W*in
   wire signed [9:0] m35_91;
   assign m35_91 =10'b0;

   // m35_92 = W*in
   wire signed [9:0] m35_92;
   assign m35_92 =10'b0;

   // m35_93 = W*in
   wire signed [9:0] m35_93;
   assign m35_93 =10'b0;

   // m35_94 = W*in
   wire signed [9:0] m35_94;
   assign m35_94 ={ {4{in35[5]}} , in35[5:0] };

   // m35_95 = W*in
   wire signed [9:0] m35_95;
   assign m35_95 =10'b0;

   // m35_96 = W*in
   wire signed [9:0] m35_96;
   assign m35_96 =10'b0;

   // m35_97 = W*in
   wire signed [9:0] m35_97;
   assign m35_97 =10'b0;

   // m35_98 = W*in
   wire signed [9:0] m35_98;
   assign m35_98 =10'b0;

   // m35_99 = W*in
   wire signed [9:0] m35_99;
   assign m35_99 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_100 = W*in
   wire signed [9:0] m35_100;
   assign m35_100 ={ {4{in35[5]}} , in35[5:0] };

   // m35_101 = W*in
   wire signed [9:0] m35_101;
   assign m35_101 =10'b0;

   // m35_102 = W*in
   wire signed [9:0] m35_102;
   assign m35_102 =10'b0;

   // m35_103 = W*in
   wire signed [9:0] m35_103;
   assign m35_103 =10'b0;

   // m35_104 = W*in
   wire signed [9:0] m35_104;
   assign m35_104 =10'b0;

   // m35_105 = W*in
   wire signed [9:0] m35_105;
   assign m35_105 =10'b0;

   // m35_106 = W*in
   wire signed [9:0] m35_106;
   assign m35_106 =10'b0;

   // m35_107 = W*in
   wire signed [9:0] m35_107;
   assign m35_107 =10'b0;

   // m35_108 = W*in
   wire signed [9:0] m35_108;
   assign m35_108 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_109 = W*in
   wire signed [9:0] m35_109;
   assign m35_109 ={ {4{neg35[5]}} , neg35[5:0] };

   // m35_110 = W*in
   wire signed [9:0] m35_110;
   assign m35_110 ={ {4{in35[5]}} , in35[5:0] };

   // m35_111 = W*in
   wire signed [9:0] m35_111;
   assign m35_111 =10'b0;

   // m35_112 = W*in
   wire signed [9:0] m35_112;
   assign m35_112 =10'b0;

   // m35_113 = W*in
   wire signed [9:0] m35_113;
   assign m35_113 =10'b0;

   // m35_114 = W*in
   wire signed [9:0] m35_114;
   assign m35_114 =10'b0;

   // m35_115 = W*in
   wire signed [9:0] m35_115;
   assign m35_115 =10'b0;

   // m35_116 = W*in
   wire signed [9:0] m35_116;
   assign m35_116 =10'b0;

   // m35_117 = W*in
   wire signed [9:0] m35_117;
   assign m35_117 =10'b0;

   // m36_1 = W*in
   wire signed [9:0] m36_1;
   assign m36_1 ={ {4{in36[5]}} , in36[5:0] };

   // m36_2 = W*in
   wire signed [9:0] m36_2;
   assign m36_2 =10'b0;

   // m36_3 = W*in
   wire signed [9:0] m36_3;
   assign m36_3 =10'b0;

   // m36_4 = W*in
   wire signed [9:0] m36_4;
   assign m36_4 =10'b0;

   // m36_5 = W*in
   wire signed [9:0] m36_5;
   assign m36_5 =10'b0;

   // m36_6 = W*in
   wire signed [9:0] m36_6;
   assign m36_6 =10'b0;

   // m36_7 = W*in
   wire signed [9:0] m36_7;
   assign m36_7 =10'b0;

   // m36_8 = W*in
   wire signed [9:0] m36_8;
   assign m36_8 =10'b0;

   // m36_9 = W*in
   wire signed [9:0] m36_9;
   assign m36_9 =10'b0;

   // m36_10 = W*in
   wire signed [9:0] m36_10;
   assign m36_10 =10'b0;

   // m36_11 = W*in
   wire signed [9:0] m36_11;
   assign m36_11 =10'b0;

   // m36_12 = W*in
   wire signed [9:0] m36_12;
   assign m36_12 =10'b0;

   // m36_13 = W*in
   wire signed [9:0] m36_13;
   assign m36_13 =10'b0;

   // m36_14 = W*in
   wire signed [9:0] m36_14;
   assign m36_14 =10'b0;

   // m36_15 = W*in
   wire signed [9:0] m36_15;
   assign m36_15 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_16 = W*in
   wire signed [9:0] m36_16;
   assign m36_16 ={ {4{in36[5]}} , in36[5:0] };

   // m36_17 = W*in
   wire signed [9:0] m36_17;
   assign m36_17 ={ {5{in36[5]}} , in36[5:1] };

   // m36_18 = W*in
   wire signed [9:0] m36_18;
   assign m36_18 =10'b0;

   // m36_19 = W*in
   wire signed [9:0] m36_19;
   assign m36_19 =10'b0;

   // m36_20 = W*in
   wire signed [9:0] m36_20;
   assign m36_20 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_21 = W*in
   wire signed [9:0] m36_21;
   assign m36_21 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_22 = W*in
   wire signed [9:0] m36_22;
   assign m36_22 =10'b0;

   // m36_23 = W*in
   wire signed [9:0] m36_23;
   assign m36_23 =10'b0;

   // m36_24 = W*in
   wire signed [9:0] m36_24;
   assign m36_24 =10'b0;

   // m36_25 = W*in
   wire signed [9:0] m36_25;
   assign m36_25 ={ {4{in36[5]}} , in36[5:0] };

   // m36_26 = W*in
   wire signed [9:0] m36_26;
   assign m36_26 =10'b0;

   // m36_27 = W*in
   wire signed [9:0] m36_27;
   assign m36_27 =10'b0;

   // m36_28 = W*in
   wire signed [9:0] m36_28;
   assign m36_28 ={ {5{in36[5]}} , in36[5:1] };

   // m36_29 = W*in
   wire signed [9:0] m36_29;
   assign m36_29 =10'b0;

   // m36_30 = W*in
   wire signed [9:0] m36_30;
   assign m36_30 =10'b0;

   // m36_31 = W*in
   wire signed [9:0] m36_31;
   assign m36_31 =10'b0;

   // m36_32 = W*in
   wire signed [9:0] m36_32;
   assign m36_32 =10'b0;

   // m36_33 = W*in
   wire signed [9:0] m36_33;
   assign m36_33 ={ {4{in36[5]}} , in36[5:0] };

   // m36_34 = W*in
   wire signed [9:0] m36_34;
   assign m36_34 =10'b0;

   // m36_35 = W*in
   wire signed [9:0] m36_35;
   assign m36_35 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_36 = W*in
   wire signed [9:0] m36_36;
   assign m36_36 ={ {5{in36[5]}} , in36[5:1] };

   // m36_37 = W*in
   wire signed [9:0] m36_37;
   assign m36_37 =10'b0;

   // m36_38 = W*in
   wire signed [9:0] m36_38;
   assign m36_38 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_39 = W*in
   wire signed [9:0] m36_39;
   assign m36_39 =10'b0;

   // m36_40 = W*in
   wire signed [9:0] m36_40;
   assign m36_40 =10'b0;

   // m36_41 = W*in
   wire signed [9:0] m36_41;
   assign m36_41 =10'b0;

   // m36_42 = W*in
   wire signed [9:0] m36_42;
   assign m36_42 =10'b0;

   // m36_43 = W*in
   wire signed [9:0] m36_43;
   assign m36_43 =10'b0;

   // m36_44 = W*in
   wire signed [9:0] m36_44;
   assign m36_44 =10'b0;

   // m36_45 = W*in
   wire signed [9:0] m36_45;
   assign m36_45 ={ {4{in36[5]}} , in36[5:0] };

   // m36_46 = W*in
   wire signed [9:0] m36_46;
   assign m36_46 =10'b0;

   // m36_47 = W*in
   wire signed [9:0] m36_47;
   assign m36_47 =10'b0;

   // m36_48 = W*in
   wire signed [9:0] m36_48;
   assign m36_48 =10'b0;

   // m36_49 = W*in
   wire signed [9:0] m36_49;
   assign m36_49 =10'b0;

   // m36_50 = W*in
   wire signed [9:0] m36_50;
   assign m36_50 =10'b0;

   // m36_51 = W*in
   wire signed [9:0] m36_51;
   assign m36_51 =10'b0;

   // m36_52 = W*in
   wire signed [9:0] m36_52;
   assign m36_52 =10'b0;

   // m36_53 = W*in
   wire signed [9:0] m36_53;
   assign m36_53 =10'b0;

   // m36_54 = W*in
   wire signed [9:0] m36_54;
   assign m36_54 =10'b0;

   // m36_55 = W*in
   wire signed [9:0] m36_55;
   assign m36_55 =10'b0;

   // m36_56 = W*in
   wire signed [9:0] m36_56;
   assign m36_56 ={ {4{in36[5]}} , in36[5:0] };

   // m36_57 = W*in
   wire signed [9:0] m36_57;
   assign m36_57 =10'b0;

   // m36_58 = W*in
   wire signed [9:0] m36_58;
   assign m36_58 =10'b0;

   // m36_59 = W*in
   wire signed [9:0] m36_59;
   assign m36_59 =10'b0;

   // m36_60 = W*in
   wire signed [9:0] m36_60;
   assign m36_60 =10'b0;

   // m36_61 = W*in
   wire signed [9:0] m36_61;
   assign m36_61 =10'b0;

   // m36_62 = W*in
   wire signed [9:0] m36_62;
   assign m36_62 =10'b0;

   // m36_63 = W*in
   wire signed [9:0] m36_63;
   assign m36_63 =10'b0;

   // m36_64 = W*in
   wire signed [9:0] m36_64;
   assign m36_64 =10'b0;

   // m36_65 = W*in
   wire signed [9:0] m36_65;
   assign m36_65 =10'b0;

   // m36_66 = W*in
   wire signed [9:0] m36_66;
   assign m36_66 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_67 = W*in
   wire signed [9:0] m36_67;
   assign m36_67 =10'b0;

   // m36_68 = W*in
   wire signed [9:0] m36_68;
   assign m36_68 =10'b0;

   // m36_69 = W*in
   wire signed [9:0] m36_69;
   assign m36_69 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_70 = W*in
   wire signed [9:0] m36_70;
   assign m36_70 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_71 = W*in
   wire signed [9:0] m36_71;
   assign m36_71 =10'b0;

   // m36_72 = W*in
   wire signed [9:0] m36_72;
   assign m36_72 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_73 = W*in
   wire signed [9:0] m36_73;
   assign m36_73 =10'b0;

   // m36_74 = W*in
   wire signed [9:0] m36_74;
   assign m36_74 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_75 = W*in
   wire signed [9:0] m36_75;
   assign m36_75 =10'b0;

   // m36_76 = W*in
   wire signed [9:0] m36_76;
   assign m36_76 =10'b0;

   // m36_77 = W*in
   wire signed [9:0] m36_77;
   assign m36_77 =10'b0;

   // m36_78 = W*in
   wire signed [9:0] m36_78;
   assign m36_78 =10'b0;

   // m36_79 = W*in
   wire signed [9:0] m36_79;
   assign m36_79 =10'b0;

   // m36_80 = W*in
   wire signed [9:0] m36_80;
   assign m36_80 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_81 = W*in
   wire signed [9:0] m36_81;
   assign m36_81 ={ {5{in36[5]}} , in36[5:1] };

   // m36_82 = W*in
   wire signed [9:0] m36_82;
   assign m36_82 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_83 = W*in
   wire signed [9:0] m36_83;
   assign m36_83 =10'b0;

   // m36_84 = W*in
   wire signed [9:0] m36_84;
   assign m36_84 =10'b0;

   // m36_85 = W*in
   wire signed [9:0] m36_85;
   assign m36_85 =10'b0;

   // m36_86 = W*in
   wire signed [9:0] m36_86;
   assign m36_86 =10'b0;

   // m36_87 = W*in
   wire signed [9:0] m36_87;
   assign m36_87 =10'b0;

   // m36_88 = W*in
   wire signed [9:0] m36_88;
   assign m36_88 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_89 = W*in
   wire signed [9:0] m36_89;
   assign m36_89 =10'b0;

   // m36_90 = W*in
   wire signed [9:0] m36_90;
   assign m36_90 =10'b0;

   // m36_91 = W*in
   wire signed [9:0] m36_91;
   assign m36_91 =10'b0;

   // m36_92 = W*in
   wire signed [9:0] m36_92;
   assign m36_92 =10'b0;

   // m36_93 = W*in
   wire signed [9:0] m36_93;
   assign m36_93 =10'b0;

   // m36_94 = W*in
   wire signed [9:0] m36_94;
   assign m36_94 =10'b0;

   // m36_95 = W*in
   wire signed [9:0] m36_95;
   assign m36_95 =10'b0;

   // m36_96 = W*in
   wire signed [9:0] m36_96;
   assign m36_96 =10'b0;

   // m36_97 = W*in
   wire signed [9:0] m36_97;
   assign m36_97 =10'b0;

   // m36_98 = W*in
   wire signed [9:0] m36_98;
   assign m36_98 =10'b0;

   // m36_99 = W*in
   wire signed [9:0] m36_99;
   assign m36_99 =10'b0;

   // m36_100 = W*in
   wire signed [9:0] m36_100;
   assign m36_100 =10'b0;

   // m36_101 = W*in
   wire signed [9:0] m36_101;
   assign m36_101 =10'b0;

   // m36_102 = W*in
   wire signed [9:0] m36_102;
   assign m36_102 =10'b0;

   // m36_103 = W*in
   wire signed [9:0] m36_103;
   assign m36_103 =10'b0;

   // m36_104 = W*in
   wire signed [9:0] m36_104;
   assign m36_104 =10'b0;

   // m36_105 = W*in
   wire signed [9:0] m36_105;
   assign m36_105 =10'b0;

   // m36_106 = W*in
   wire signed [9:0] m36_106;
   assign m36_106 =10'b0;

   // m36_107 = W*in
   wire signed [9:0] m36_107;
   assign m36_107 =10'b0;

   // m36_108 = W*in
   wire signed [9:0] m36_108;
   assign m36_108 ={ {5{neg36[5]}} , neg36[5:1] };

   // m36_109 = W*in
   wire signed [9:0] m36_109;
   assign m36_109 ={ {4{neg36[5]}} , neg36[5:0] };

   // m36_110 = W*in
   wire signed [9:0] m36_110;
   assign m36_110 =10'b0;

   // m36_111 = W*in
   wire signed [9:0] m36_111;
   assign m36_111 =10'b0;

   // m36_112 = W*in
   wire signed [9:0] m36_112;
   assign m36_112 =10'b0;

   // m36_113 = W*in
   wire signed [9:0] m36_113;
   assign m36_113 =10'b0;

   // m36_114 = W*in
   wire signed [9:0] m36_114;
   assign m36_114 =10'b0;

   // m36_115 = W*in
   wire signed [9:0] m36_115;
   assign m36_115 =10'b0;

   // m36_116 = W*in
   wire signed [9:0] m36_116;
   assign m36_116 =10'b0;

   // m36_117 = W*in
   wire signed [9:0] m36_117;
   assign m36_117 =10'b0;

   // m37_1 = W*in
   wire signed [9:0] m37_1;
   assign m37_1 =10'b0;

   // m37_2 = W*in
   wire signed [9:0] m37_2;
   assign m37_2 =10'b0;

   // m37_3 = W*in
   wire signed [9:0] m37_3;
   assign m37_3 =10'b0;

   // m37_4 = W*in
   wire signed [9:0] m37_4;
   assign m37_4 =10'b0;

   // m37_5 = W*in
   wire signed [9:0] m37_5;
   assign m37_5 =10'b0;

   // m37_6 = W*in
   wire signed [9:0] m37_6;
   assign m37_6 =10'b0;

   // m37_7 = W*in
   wire signed [9:0] m37_7;
   assign m37_7 =10'b0;

   // m37_8 = W*in
   wire signed [9:0] m37_8;
   assign m37_8 =10'b0;

   // m37_9 = W*in
   wire signed [9:0] m37_9;
   assign m37_9 =10'b0;

   // m37_10 = W*in
   wire signed [9:0] m37_10;
   assign m37_10 =10'b0;

   // m37_11 = W*in
   wire signed [9:0] m37_11;
   assign m37_11 =10'b0;

   // m37_12 = W*in
   wire signed [9:0] m37_12;
   assign m37_12 =10'b0;

   // m37_13 = W*in
   wire signed [9:0] m37_13;
   assign m37_13 =10'b0;

   // m37_14 = W*in
   wire signed [9:0] m37_14;
   assign m37_14 =10'b0;

   // m37_15 = W*in
   wire signed [9:0] m37_15;
   assign m37_15 =10'b0;

   // m37_16 = W*in
   wire signed [9:0] m37_16;
   assign m37_16 =10'b0;

   // m37_17 = W*in
   wire signed [9:0] m37_17;
   assign m37_17 =10'b0;

   // m37_18 = W*in
   wire signed [9:0] m37_18;
   assign m37_18 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_19 = W*in
   wire signed [9:0] m37_19;
   assign m37_19 =10'b0;

   // m37_20 = W*in
   wire signed [9:0] m37_20;
   assign m37_20 ={ {5{in37[5]}} , in37[5:1] };

   // m37_21 = W*in
   wire signed [9:0] m37_21;
   assign m37_21 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_22 = W*in
   wire signed [9:0] m37_22;
   assign m37_22 =10'b0;

   // m37_23 = W*in
   wire signed [9:0] m37_23;
   assign m37_23 =10'b0;

   // m37_24 = W*in
   wire signed [9:0] m37_24;
   assign m37_24 =10'b0;

   // m37_25 = W*in
   wire signed [9:0] m37_25;
   assign m37_25 =10'b0;

   // m37_26 = W*in
   wire signed [9:0] m37_26;
   assign m37_26 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_27 = W*in
   wire signed [9:0] m37_27;
   assign m37_27 =10'b0;

   // m37_28 = W*in
   wire signed [9:0] m37_28;
   assign m37_28 =10'b0;

   // m37_29 = W*in
   wire signed [9:0] m37_29;
   assign m37_29 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_30 = W*in
   wire signed [9:0] m37_30;
   assign m37_30 =10'b0;

   // m37_31 = W*in
   wire signed [9:0] m37_31;
   assign m37_31 ={ {5{in37[5]}} , in37[5:1] };

   // m37_32 = W*in
   wire signed [9:0] m37_32;
   assign m37_32 =10'b0;

   // m37_33 = W*in
   wire signed [9:0] m37_33;
   assign m37_33 =10'b0;

   // m37_34 = W*in
   wire signed [9:0] m37_34;
   assign m37_34 =10'b0;

   // m37_35 = W*in
   wire signed [9:0] m37_35;
   assign m37_35 =10'b0;

   // m37_36 = W*in
   wire signed [9:0] m37_36;
   assign m37_36 ={ {5{in37[5]}} , in37[5:1] };

   // m37_37 = W*in
   wire signed [9:0] m37_37;
   assign m37_37 =10'b0;

   // m37_38 = W*in
   wire signed [9:0] m37_38;
   assign m37_38 =10'b0;

   // m37_39 = W*in
   wire signed [9:0] m37_39;
   assign m37_39 =10'b0;

   // m37_40 = W*in
   wire signed [9:0] m37_40;
   assign m37_40 =10'b0;

   // m37_41 = W*in
   wire signed [9:0] m37_41;
   assign m37_41 =10'b0;

   // m37_42 = W*in
   wire signed [9:0] m37_42;
   assign m37_42 =10'b0;

   // m37_43 = W*in
   wire signed [9:0] m37_43;
   assign m37_43 =10'b0;

   // m37_44 = W*in
   wire signed [9:0] m37_44;
   assign m37_44 =10'b0;

   // m37_45 = W*in
   wire signed [9:0] m37_45;
   assign m37_45 =10'b0;

   // m37_46 = W*in
   wire signed [9:0] m37_46;
   assign m37_46 =10'b0;

   // m37_47 = W*in
   wire signed [9:0] m37_47;
   assign m37_47 =10'b0;

   // m37_48 = W*in
   wire signed [9:0] m37_48;
   assign m37_48 =10'b0;

   // m37_49 = W*in
   wire signed [9:0] m37_49;
   assign m37_49 =10'b0;

   // m37_50 = W*in
   wire signed [9:0] m37_50;
   assign m37_50 =10'b0;

   // m37_51 = W*in
   wire signed [9:0] m37_51;
   assign m37_51 =10'b0;

   // m37_52 = W*in
   wire signed [9:0] m37_52;
   assign m37_52 =10'b0;

   // m37_53 = W*in
   wire signed [9:0] m37_53;
   assign m37_53 =10'b0;

   // m37_54 = W*in
   wire signed [9:0] m37_54;
   assign m37_54 =10'b0;

   // m37_55 = W*in
   wire signed [9:0] m37_55;
   assign m37_55 =10'b0;

   // m37_56 = W*in
   wire signed [9:0] m37_56;
   assign m37_56 =10'b0;

   // m37_57 = W*in
   wire signed [9:0] m37_57;
   assign m37_57 =10'b0;

   // m37_58 = W*in
   wire signed [9:0] m37_58;
   assign m37_58 =10'b0;

   // m37_59 = W*in
   wire signed [9:0] m37_59;
   assign m37_59 =10'b0;

   // m37_60 = W*in
   wire signed [9:0] m37_60;
   assign m37_60 =10'b0;

   // m37_61 = W*in
   wire signed [9:0] m37_61;
   assign m37_61 =10'b0;

   // m37_62 = W*in
   wire signed [9:0] m37_62;
   assign m37_62 =10'b0;

   // m37_63 = W*in
   wire signed [9:0] m37_63;
   assign m37_63 =10'b0;

   // m37_64 = W*in
   wire signed [9:0] m37_64;
   assign m37_64 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_65 = W*in
   wire signed [9:0] m37_65;
   assign m37_65 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_66 = W*in
   wire signed [9:0] m37_66;
   assign m37_66 ={ {4{neg37[5]}} , neg37[5:0] };

   // m37_67 = W*in
   wire signed [9:0] m37_67;
   assign m37_67 =10'b0;

   // m37_68 = W*in
   wire signed [9:0] m37_68;
   assign m37_68 =10'b0;

   // m37_69 = W*in
   wire signed [9:0] m37_69;
   assign m37_69 =10'b0;

   // m37_70 = W*in
   wire signed [9:0] m37_70;
   assign m37_70 =10'b0;

   // m37_71 = W*in
   wire signed [9:0] m37_71;
   assign m37_71 =10'b0;

   // m37_72 = W*in
   wire signed [9:0] m37_72;
   assign m37_72 ={ {5{neg37[5]}} , neg37[5:1] };

   // m37_73 = W*in
   wire signed [9:0] m37_73;
   assign m37_73 =10'b0;

   // m37_74 = W*in
   wire signed [9:0] m37_74;
   assign m37_74 =10'b0;

   // m37_75 = W*in
   wire signed [9:0] m37_75;
   assign m37_75 =10'b0;

   // m37_76 = W*in
   wire signed [9:0] m37_76;
   assign m37_76 =10'b0;

   // m37_77 = W*in
   wire signed [9:0] m37_77;
   assign m37_77 =10'b0;

   // m37_78 = W*in
   wire signed [9:0] m37_78;
   assign m37_78 =10'b0;

   // m37_79 = W*in
   wire signed [9:0] m37_79;
   assign m37_79 =10'b0;

   // m37_80 = W*in
   wire signed [9:0] m37_80;
   assign m37_80 =10'b0;

   // m37_81 = W*in
   wire signed [9:0] m37_81;
   assign m37_81 =10'b0;

   // m37_82 = W*in
   wire signed [9:0] m37_82;
   assign m37_82 =10'b0;

   // m37_83 = W*in
   wire signed [9:0] m37_83;
   assign m37_83 =10'b0;

   // m37_84 = W*in
   wire signed [9:0] m37_84;
   assign m37_84 =10'b0;

   // m37_85 = W*in
   wire signed [9:0] m37_85;
   assign m37_85 =10'b0;

   // m37_86 = W*in
   wire signed [9:0] m37_86;
   assign m37_86 =10'b0;

   // m37_87 = W*in
   wire signed [9:0] m37_87;
   assign m37_87 =10'b0;

   // m37_88 = W*in
   wire signed [9:0] m37_88;
   assign m37_88 =10'b0;

   // m37_89 = W*in
   wire signed [9:0] m37_89;
   assign m37_89 =10'b0;

   // m37_90 = W*in
   wire signed [9:0] m37_90;
   assign m37_90 =10'b0;

   // m37_91 = W*in
   wire signed [9:0] m37_91;
   assign m37_91 =10'b0;

   // m37_92 = W*in
   wire signed [9:0] m37_92;
   assign m37_92 =10'b0;

   // m37_93 = W*in
   wire signed [9:0] m37_93;
   assign m37_93 =10'b0;

   // m37_94 = W*in
   wire signed [9:0] m37_94;
   assign m37_94 =10'b0;

   // m37_95 = W*in
   wire signed [9:0] m37_95;
   assign m37_95 =10'b0;

   // m37_96 = W*in
   wire signed [9:0] m37_96;
   assign m37_96 =10'b0;

   // m37_97 = W*in
   wire signed [9:0] m37_97;
   assign m37_97 =10'b0;

   // m37_98 = W*in
   wire signed [9:0] m37_98;
   assign m37_98 =10'b0;

   // m37_99 = W*in
   wire signed [9:0] m37_99;
   assign m37_99 =10'b0;

   // m37_100 = W*in
   wire signed [9:0] m37_100;
   assign m37_100 ={ {4{neg37[5]}} , neg37[5:0] };

   // m37_101 = W*in
   wire signed [9:0] m37_101;
   assign m37_101 =10'b0;

   // m37_102 = W*in
   wire signed [9:0] m37_102;
   assign m37_102 =10'b0;

   // m37_103 = W*in
   wire signed [9:0] m37_103;
   assign m37_103 =10'b0;

   // m37_104 = W*in
   wire signed [9:0] m37_104;
   assign m37_104 =10'b0;

   // m37_105 = W*in
   wire signed [9:0] m37_105;
   assign m37_105 =10'b0;

   // m37_106 = W*in
   wire signed [9:0] m37_106;
   assign m37_106 =10'b0;

   // m37_107 = W*in
   wire signed [9:0] m37_107;
   assign m37_107 =10'b0;

   // m37_108 = W*in
   wire signed [9:0] m37_108;
   assign m37_108 =10'b0;

   // m37_109 = W*in
   wire signed [9:0] m37_109;
   assign m37_109 =10'b0;

   // m37_110 = W*in
   wire signed [9:0] m37_110;
   assign m37_110 =10'b0;

   // m37_111 = W*in
   wire signed [9:0] m37_111;
   assign m37_111 =10'b0;

   // m37_112 = W*in
   wire signed [9:0] m37_112;
   assign m37_112 =10'b0;

   // m37_113 = W*in
   wire signed [9:0] m37_113;
   assign m37_113 =10'b0;

   // m37_114 = W*in
   wire signed [9:0] m37_114;
   assign m37_114 =10'b0;

   // m37_115 = W*in
   wire signed [9:0] m37_115;
   assign m37_115 =10'b0;

   // m37_116 = W*in
   wire signed [9:0] m37_116;
   assign m37_116 ={ {4{in37[5]}} , in37[5:0] };

   // m37_117 = W*in
   wire signed [9:0] m37_117;
   assign m37_117 =10'b0;

   // m38_1 = W*in
   wire signed [9:0] m38_1;
   assign m38_1 =10'b0;

   // m38_2 = W*in
   wire signed [9:0] m38_2;
   assign m38_2 =10'b0;

   // m38_3 = W*in
   wire signed [9:0] m38_3;
   assign m38_3 =10'b0;

   // m38_4 = W*in
   wire signed [9:0] m38_4;
   assign m38_4 =10'b0;

   // m38_5 = W*in
   wire signed [9:0] m38_5;
   assign m38_5 =10'b0;

   // m38_6 = W*in
   wire signed [9:0] m38_6;
   assign m38_6 =10'b0;

   // m38_7 = W*in
   wire signed [9:0] m38_7;
   assign m38_7 =10'b0;

   // m38_8 = W*in
   wire signed [9:0] m38_8;
   assign m38_8 =10'b0;

   // m38_9 = W*in
   wire signed [9:0] m38_9;
   assign m38_9 =10'b0;

   // m38_10 = W*in
   wire signed [9:0] m38_10;
   assign m38_10 =10'b0;

   // m38_11 = W*in
   wire signed [9:0] m38_11;
   assign m38_11 =10'b0;

   // m38_12 = W*in
   wire signed [9:0] m38_12;
   assign m38_12 =10'b0;

   // m38_13 = W*in
   wire signed [9:0] m38_13;
   assign m38_13 =10'b0;

   // m38_14 = W*in
   wire signed [9:0] m38_14;
   assign m38_14 =10'b0;

   // m38_15 = W*in
   wire signed [9:0] m38_15;
   assign m38_15 =10'b0;

   // m38_16 = W*in
   wire signed [9:0] m38_16;
   assign m38_16 =10'b0;

   // m38_17 = W*in
   wire signed [9:0] m38_17;
   assign m38_17 =10'b0;

   // m38_18 = W*in
   wire signed [9:0] m38_18;
   assign m38_18 =10'b0;

   // m38_19 = W*in
   wire signed [9:0] m38_19;
   assign m38_19 =10'b0;

   // m38_20 = W*in
   wire signed [9:0] m38_20;
   assign m38_20 ={ {5{in38[5]}} , in38[5:1] };

   // m38_21 = W*in
   wire signed [9:0] m38_21;
   assign m38_21 =10'b0;

   // m38_22 = W*in
   wire signed [9:0] m38_22;
   assign m38_22 =10'b0;

   // m38_23 = W*in
   wire signed [9:0] m38_23;
   assign m38_23 =10'b0;

   // m38_24 = W*in
   wire signed [9:0] m38_24;
   assign m38_24 =10'b0;

   // m38_25 = W*in
   wire signed [9:0] m38_25;
   assign m38_25 =10'b0;

   // m38_26 = W*in
   wire signed [9:0] m38_26;
   assign m38_26 ={ {5{neg38[5]}} , neg38[5:1] };

   // m38_27 = W*in
   wire signed [9:0] m38_27;
   assign m38_27 =10'b0;

   // m38_28 = W*in
   wire signed [9:0] m38_28;
   assign m38_28 =10'b0;

   // m38_29 = W*in
   wire signed [9:0] m38_29;
   assign m38_29 ={ {5{neg38[5]}} , neg38[5:1] };

   // m38_30 = W*in
   wire signed [9:0] m38_30;
   assign m38_30 =10'b0;

   // m38_31 = W*in
   wire signed [9:0] m38_31;
   assign m38_31 ={ {5{in38[5]}} , in38[5:1] };

   // m38_32 = W*in
   wire signed [9:0] m38_32;
   assign m38_32 =10'b0;

   // m38_33 = W*in
   wire signed [9:0] m38_33;
   assign m38_33 =10'b0;

   // m38_34 = W*in
   wire signed [9:0] m38_34;
   assign m38_34 =10'b0;

   // m38_35 = W*in
   wire signed [9:0] m38_35;
   assign m38_35 =10'b0;

   // m38_36 = W*in
   wire signed [9:0] m38_36;
   assign m38_36 =10'b0;

   // m38_37 = W*in
   wire signed [9:0] m38_37;
   assign m38_37 =10'b0;

   // m38_38 = W*in
   wire signed [9:0] m38_38;
   assign m38_38 =10'b0;

   // m38_39 = W*in
   wire signed [9:0] m38_39;
   assign m38_39 =10'b0;

   // m38_40 = W*in
   wire signed [9:0] m38_40;
   assign m38_40 =10'b0;

   // m38_41 = W*in
   wire signed [9:0] m38_41;
   assign m38_41 =10'b0;

   // m38_42 = W*in
   wire signed [9:0] m38_42;
   assign m38_42 =10'b0;

   // m38_43 = W*in
   wire signed [9:0] m38_43;
   assign m38_43 =10'b0;

   // m38_44 = W*in
   wire signed [9:0] m38_44;
   assign m38_44 =10'b0;

   // m38_45 = W*in
   wire signed [9:0] m38_45;
   assign m38_45 =10'b0;

   // m38_46 = W*in
   wire signed [9:0] m38_46;
   assign m38_46 =10'b0;

   // m38_47 = W*in
   wire signed [9:0] m38_47;
   assign m38_47 =10'b0;

   // m38_48 = W*in
   wire signed [9:0] m38_48;
   assign m38_48 =10'b0;

   // m38_49 = W*in
   wire signed [9:0] m38_49;
   assign m38_49 =10'b0;

   // m38_50 = W*in
   wire signed [9:0] m38_50;
   assign m38_50 =10'b0;

   // m38_51 = W*in
   wire signed [9:0] m38_51;
   assign m38_51 =10'b0;

   // m38_52 = W*in
   wire signed [9:0] m38_52;
   assign m38_52 =10'b0;

   // m38_53 = W*in
   wire signed [9:0] m38_53;
   assign m38_53 =10'b0;

   // m38_54 = W*in
   wire signed [9:0] m38_54;
   assign m38_54 =10'b0;

   // m38_55 = W*in
   wire signed [9:0] m38_55;
   assign m38_55 =10'b0;

   // m38_56 = W*in
   wire signed [9:0] m38_56;
   assign m38_56 =10'b0;

   // m38_57 = W*in
   wire signed [9:0] m38_57;
   assign m38_57 =10'b0;

   // m38_58 = W*in
   wire signed [9:0] m38_58;
   assign m38_58 =10'b0;

   // m38_59 = W*in
   wire signed [9:0] m38_59;
   assign m38_59 =10'b0;

   // m38_60 = W*in
   wire signed [9:0] m38_60;
   assign m38_60 =10'b0;

   // m38_61 = W*in
   wire signed [9:0] m38_61;
   assign m38_61 =10'b0;

   // m38_62 = W*in
   wire signed [9:0] m38_62;
   assign m38_62 =10'b0;

   // m38_63 = W*in
   wire signed [9:0] m38_63;
   assign m38_63 =10'b0;

   // m38_64 = W*in
   wire signed [9:0] m38_64;
   assign m38_64 =10'b0;

   // m38_65 = W*in
   wire signed [9:0] m38_65;
   assign m38_65 =10'b0;

   // m38_66 = W*in
   wire signed [9:0] m38_66;
   assign m38_66 ={ {5{neg38[5]}} , neg38[5:1] };

   // m38_67 = W*in
   wire signed [9:0] m38_67;
   assign m38_67 =10'b0;

   // m38_68 = W*in
   wire signed [9:0] m38_68;
   assign m38_68 =10'b0;

   // m38_69 = W*in
   wire signed [9:0] m38_69;
   assign m38_69 =10'b0;

   // m38_70 = W*in
   wire signed [9:0] m38_70;
   assign m38_70 =10'b0;

   // m38_71 = W*in
   wire signed [9:0] m38_71;
   assign m38_71 =10'b0;

   // m38_72 = W*in
   wire signed [9:0] m38_72;
   assign m38_72 =10'b0;

   // m38_73 = W*in
   wire signed [9:0] m38_73;
   assign m38_73 =10'b0;

   // m38_74 = W*in
   wire signed [9:0] m38_74;
   assign m38_74 =10'b0;

   // m38_75 = W*in
   wire signed [9:0] m38_75;
   assign m38_75 =10'b0;

   // m38_76 = W*in
   wire signed [9:0] m38_76;
   assign m38_76 =10'b0;

   // m38_77 = W*in
   wire signed [9:0] m38_77;
   assign m38_77 =10'b0;

   // m38_78 = W*in
   wire signed [9:0] m38_78;
   assign m38_78 =10'b0;

   // m38_79 = W*in
   wire signed [9:0] m38_79;
   assign m38_79 =10'b0;

   // m38_80 = W*in
   wire signed [9:0] m38_80;
   assign m38_80 =10'b0;

   // m38_81 = W*in
   wire signed [9:0] m38_81;
   assign m38_81 =10'b0;

   // m38_82 = W*in
   wire signed [9:0] m38_82;
   assign m38_82 =10'b0;

   // m38_83 = W*in
   wire signed [9:0] m38_83;
   assign m38_83 =10'b0;

   // m38_84 = W*in
   wire signed [9:0] m38_84;
   assign m38_84 =10'b0;

   // m38_85 = W*in
   wire signed [9:0] m38_85;
   assign m38_85 =10'b0;

   // m38_86 = W*in
   wire signed [9:0] m38_86;
   assign m38_86 =10'b0;

   // m38_87 = W*in
   wire signed [9:0] m38_87;
   assign m38_87 =10'b0;

   // m38_88 = W*in
   wire signed [9:0] m38_88;
   assign m38_88 =10'b0;

   // m38_89 = W*in
   wire signed [9:0] m38_89;
   assign m38_89 =10'b0;

   // m38_90 = W*in
   wire signed [9:0] m38_90;
   assign m38_90 =10'b0;

   // m38_91 = W*in
   wire signed [9:0] m38_91;
   assign m38_91 =10'b0;

   // m38_92 = W*in
   wire signed [9:0] m38_92;
   assign m38_92 =10'b0;

   // m38_93 = W*in
   wire signed [9:0] m38_93;
   assign m38_93 =10'b0;

   // m38_94 = W*in
   wire signed [9:0] m38_94;
   assign m38_94 =10'b0;

   // m38_95 = W*in
   wire signed [9:0] m38_95;
   assign m38_95 =10'b0;

   // m38_96 = W*in
   wire signed [9:0] m38_96;
   assign m38_96 =10'b0;

   // m38_97 = W*in
   wire signed [9:0] m38_97;
   assign m38_97 =10'b0;

   // m38_98 = W*in
   wire signed [9:0] m38_98;
   assign m38_98 =10'b0;

   // m38_99 = W*in
   wire signed [9:0] m38_99;
   assign m38_99 =10'b0;

   // m38_100 = W*in
   wire signed [9:0] m38_100;
   assign m38_100 =10'b0;

   // m38_101 = W*in
   wire signed [9:0] m38_101;
   assign m38_101 =10'b0;

   // m38_102 = W*in
   wire signed [9:0] m38_102;
   assign m38_102 =10'b0;

   // m38_103 = W*in
   wire signed [9:0] m38_103;
   assign m38_103 =10'b0;

   // m38_104 = W*in
   wire signed [9:0] m38_104;
   assign m38_104 =10'b0;

   // m38_105 = W*in
   wire signed [9:0] m38_105;
   assign m38_105 =10'b0;

   // m38_106 = W*in
   wire signed [9:0] m38_106;
   assign m38_106 =10'b0;

   // m38_107 = W*in
   wire signed [9:0] m38_107;
   assign m38_107 =10'b0;

   // m38_108 = W*in
   wire signed [9:0] m38_108;
   assign m38_108 =10'b0;

   // m38_109 = W*in
   wire signed [9:0] m38_109;
   assign m38_109 ={ {5{in38[5]}} , in38[5:1] };

   // m38_110 = W*in
   wire signed [9:0] m38_110;
   assign m38_110 =10'b0;

   // m38_111 = W*in
   wire signed [9:0] m38_111;
   assign m38_111 =10'b0;

   // m38_112 = W*in
   wire signed [9:0] m38_112;
   assign m38_112 =10'b0;

   // m38_113 = W*in
   wire signed [9:0] m38_113;
   assign m38_113 =10'b0;

   // m38_114 = W*in
   wire signed [9:0] m38_114;
   assign m38_114 =10'b0;

   // m38_115 = W*in
   wire signed [9:0] m38_115;
   assign m38_115 =10'b0;

   // m38_116 = W*in
   wire signed [9:0] m38_116;
   assign m38_116 =10'b0;

   // m38_117 = W*in
   wire signed [9:0] m38_117;
   assign m38_117 =10'b0;

   // m39_1 = W*in
   wire signed [9:0] m39_1;
   assign m39_1 =10'b0;

   // m39_2 = W*in
   wire signed [9:0] m39_2;
   assign m39_2 =10'b0;

   // m39_3 = W*in
   wire signed [9:0] m39_3;
   assign m39_3 =10'b0;

   // m39_4 = W*in
   wire signed [9:0] m39_4;
   assign m39_4 =10'b0;

   // m39_5 = W*in
   wire signed [9:0] m39_5;
   assign m39_5 =10'b0;

   // m39_6 = W*in
   wire signed [9:0] m39_6;
   assign m39_6 =10'b0;

   // m39_7 = W*in
   wire signed [9:0] m39_7;
   assign m39_7 =10'b0;

   // m39_8 = W*in
   wire signed [9:0] m39_8;
   assign m39_8 =10'b0;

   // m39_9 = W*in
   wire signed [9:0] m39_9;
   assign m39_9 =10'b0;

   // m39_10 = W*in
   wire signed [9:0] m39_10;
   assign m39_10 =10'b0;

   // m39_11 = W*in
   wire signed [9:0] m39_11;
   assign m39_11 =10'b0;

   // m39_12 = W*in
   wire signed [9:0] m39_12;
   assign m39_12 =10'b0;

   // m39_13 = W*in
   wire signed [9:0] m39_13;
   assign m39_13 =10'b0;

   // m39_14 = W*in
   wire signed [9:0] m39_14;
   assign m39_14 =10'b0;

   // m39_15 = W*in
   wire signed [9:0] m39_15;
   assign m39_15 =10'b0;

   // m39_16 = W*in
   wire signed [9:0] m39_16;
   assign m39_16 =10'b0;

   // m39_17 = W*in
   wire signed [9:0] m39_17;
   assign m39_17 =10'b0;

   // m39_18 = W*in
   wire signed [9:0] m39_18;
   assign m39_18 ={ {5{in39[5]}} , in39[5:1] };

   // m39_19 = W*in
   wire signed [9:0] m39_19;
   assign m39_19 =10'b0;

   // m39_20 = W*in
   wire signed [9:0] m39_20;
   assign m39_20 =10'b0;

   // m39_21 = W*in
   wire signed [9:0] m39_21;
   assign m39_21 =10'b0;

   // m39_22 = W*in
   wire signed [9:0] m39_22;
   assign m39_22 ={ {5{in39[5]}} , in39[5:1] };

   // m39_23 = W*in
   wire signed [9:0] m39_23;
   assign m39_23 =10'b0;

   // m39_24 = W*in
   wire signed [9:0] m39_24;
   assign m39_24 =10'b0;

   // m39_25 = W*in
   wire signed [9:0] m39_25;
   assign m39_25 =10'b0;

   // m39_26 = W*in
   wire signed [9:0] m39_26;
   assign m39_26 ={ {5{in39[5]}} , in39[5:1] };

   // m39_27 = W*in
   wire signed [9:0] m39_27;
   assign m39_27 ={ {5{in39[5]}} , in39[5:1] };

   // m39_28 = W*in
   wire signed [9:0] m39_28;
   assign m39_28 ={ {5{in39[5]}} , in39[5:1] };

   // m39_29 = W*in
   wire signed [9:0] m39_29;
   assign m39_29 ={ {5{neg39[5]}} , neg39[5:1] };

   // m39_30 = W*in
   wire signed [9:0] m39_30;
   assign m39_30 =10'b0;

   // m39_31 = W*in
   wire signed [9:0] m39_31;
   assign m39_31 =10'b0;

   // m39_32 = W*in
   wire signed [9:0] m39_32;
   assign m39_32 =10'b0;

   // m39_33 = W*in
   wire signed [9:0] m39_33;
   assign m39_33 =10'b0;

   // m39_34 = W*in
   wire signed [9:0] m39_34;
   assign m39_34 =10'b0;

   // m39_35 = W*in
   wire signed [9:0] m39_35;
   assign m39_35 =10'b0;

   // m39_36 = W*in
   wire signed [9:0] m39_36;
   assign m39_36 =10'b0;

   // m39_37 = W*in
   wire signed [9:0] m39_37;
   assign m39_37 =10'b0;

   // m39_38 = W*in
   wire signed [9:0] m39_38;
   assign m39_38 =10'b0;

   // m39_39 = W*in
   wire signed [9:0] m39_39;
   assign m39_39 =10'b0;

   // m39_40 = W*in
   wire signed [9:0] m39_40;
   assign m39_40 =10'b0;

   // m39_41 = W*in
   wire signed [9:0] m39_41;
   assign m39_41 =10'b0;

   // m39_42 = W*in
   wire signed [9:0] m39_42;
   assign m39_42 ={ {4{in39[5]}} , in39[5:0] };

   // m39_43 = W*in
   wire signed [9:0] m39_43;
   assign m39_43 =10'b0;

   // m39_44 = W*in
   wire signed [9:0] m39_44;
   assign m39_44 =10'b0;

   // m39_45 = W*in
   wire signed [9:0] m39_45;
   assign m39_45 =10'b0;

   // m39_46 = W*in
   wire signed [9:0] m39_46;
   assign m39_46 =10'b0;

   // m39_47 = W*in
   wire signed [9:0] m39_47;
   assign m39_47 =10'b0;

   // m39_48 = W*in
   wire signed [9:0] m39_48;
   assign m39_48 =10'b0;

   // m39_49 = W*in
   wire signed [9:0] m39_49;
   assign m39_49 =10'b0;

   // m39_50 = W*in
   wire signed [9:0] m39_50;
   assign m39_50 =10'b0;

   // m39_51 = W*in
   wire signed [9:0] m39_51;
   assign m39_51 =10'b0;

   // m39_52 = W*in
   wire signed [9:0] m39_52;
   assign m39_52 =10'b0;

   // m39_53 = W*in
   wire signed [9:0] m39_53;
   assign m39_53 =10'b0;

   // m39_54 = W*in
   wire signed [9:0] m39_54;
   assign m39_54 =10'b0;

   // m39_55 = W*in
   wire signed [9:0] m39_55;
   assign m39_55 =10'b0;

   // m39_56 = W*in
   wire signed [9:0] m39_56;
   assign m39_56 =10'b0;

   // m39_57 = W*in
   wire signed [9:0] m39_57;
   assign m39_57 =10'b0;

   // m39_58 = W*in
   wire signed [9:0] m39_58;
   assign m39_58 =10'b0;

   // m39_59 = W*in
   wire signed [9:0] m39_59;
   assign m39_59 =10'b0;

   // m39_60 = W*in
   wire signed [9:0] m39_60;
   assign m39_60 =10'b0;

   // m39_61 = W*in
   wire signed [9:0] m39_61;
   assign m39_61 =10'b0;

   // m39_62 = W*in
   wire signed [9:0] m39_62;
   assign m39_62 =10'b0;

   // m39_63 = W*in
   wire signed [9:0] m39_63;
   assign m39_63 =10'b0;

   // m39_64 = W*in
   wire signed [9:0] m39_64;
   assign m39_64 =10'b0;

   // m39_65 = W*in
   wire signed [9:0] m39_65;
   assign m39_65 =10'b0;

   // m39_66 = W*in
   wire signed [9:0] m39_66;
   assign m39_66 =10'b0;

   // m39_67 = W*in
   wire signed [9:0] m39_67;
   assign m39_67 =10'b0;

   // m39_68 = W*in
   wire signed [9:0] m39_68;
   assign m39_68 =10'b0;

   // m39_69 = W*in
   wire signed [9:0] m39_69;
   assign m39_69 ={ {4{neg39[5]}} , neg39[5:0] };

   // m39_70 = W*in
   wire signed [9:0] m39_70;
   assign m39_70 =10'b0;

   // m39_71 = W*in
   wire signed [9:0] m39_71;
   assign m39_71 =10'b0;

   // m39_72 = W*in
   wire signed [9:0] m39_72;
   assign m39_72 =10'b0;

   // m39_73 = W*in
   wire signed [9:0] m39_73;
   assign m39_73 =10'b0;

   // m39_74 = W*in
   wire signed [9:0] m39_74;
   assign m39_74 =10'b0;

   // m39_75 = W*in
   wire signed [9:0] m39_75;
   assign m39_75 =10'b0;

   // m39_76 = W*in
   wire signed [9:0] m39_76;
   assign m39_76 =10'b0;

   // m39_77 = W*in
   wire signed [9:0] m39_77;
   assign m39_77 =10'b0;

   // m39_78 = W*in
   wire signed [9:0] m39_78;
   assign m39_78 =10'b0;

   // m39_79 = W*in
   wire signed [9:0] m39_79;
   assign m39_79 =10'b0;

   // m39_80 = W*in
   wire signed [9:0] m39_80;
   assign m39_80 =10'b0;

   // m39_81 = W*in
   wire signed [9:0] m39_81;
   assign m39_81 ={ {5{in39[5]}} , in39[5:1] };

   // m39_82 = W*in
   wire signed [9:0] m39_82;
   assign m39_82 =10'b0;

   // m39_83 = W*in
   wire signed [9:0] m39_83;
   assign m39_83 =10'b0;

   // m39_84 = W*in
   wire signed [9:0] m39_84;
   assign m39_84 =10'b0;

   // m39_85 = W*in
   wire signed [9:0] m39_85;
   assign m39_85 ={ {5{neg39[5]}} , neg39[5:1] };

   // m39_86 = W*in
   wire signed [9:0] m39_86;
   assign m39_86 =10'b0;

   // m39_87 = W*in
   wire signed [9:0] m39_87;
   assign m39_87 =10'b0;

   // m39_88 = W*in
   wire signed [9:0] m39_88;
   assign m39_88 =10'b0;

   // m39_89 = W*in
   wire signed [9:0] m39_89;
   assign m39_89 =10'b0;

   // m39_90 = W*in
   wire signed [9:0] m39_90;
   assign m39_90 =10'b0;

   // m39_91 = W*in
   wire signed [9:0] m39_91;
   assign m39_91 =10'b0;

   // m39_92 = W*in
   wire signed [9:0] m39_92;
   assign m39_92 =10'b0;

   // m39_93 = W*in
   wire signed [9:0] m39_93;
   assign m39_93 ={ {4{neg39[5]}} , neg39[5:0] };

   // m39_94 = W*in
   wire signed [9:0] m39_94;
   assign m39_94 =10'b0;

   // m39_95 = W*in
   wire signed [9:0] m39_95;
   assign m39_95 =10'b0;

   // m39_96 = W*in
   wire signed [9:0] m39_96;
   assign m39_96 =10'b0;

   // m39_97 = W*in
   wire signed [9:0] m39_97;
   assign m39_97 =10'b0;

   // m39_98 = W*in
   wire signed [9:0] m39_98;
   assign m39_98 =10'b0;

   // m39_99 = W*in
   wire signed [9:0] m39_99;
   assign m39_99 =10'b0;

   // m39_100 = W*in
   wire signed [9:0] m39_100;
   assign m39_100 =10'b0;

   // m39_101 = W*in
   wire signed [9:0] m39_101;
   assign m39_101 =10'b0;

   // m39_102 = W*in
   wire signed [9:0] m39_102;
   assign m39_102 =10'b0;

   // m39_103 = W*in
   wire signed [9:0] m39_103;
   assign m39_103 =10'b0;

   // m39_104 = W*in
   wire signed [9:0] m39_104;
   assign m39_104 =10'b0;

   // m39_105 = W*in
   wire signed [9:0] m39_105;
   assign m39_105 =10'b0;

   // m39_106 = W*in
   wire signed [9:0] m39_106;
   assign m39_106 =10'b0;

   // m39_107 = W*in
   wire signed [9:0] m39_107;
   assign m39_107 =10'b0;

   // m39_108 = W*in
   wire signed [9:0] m39_108;
   assign m39_108 =10'b0;

   // m39_109 = W*in
   wire signed [9:0] m39_109;
   assign m39_109 ={ {5{neg39[5]}} , neg39[5:1] };

   // m39_110 = W*in
   wire signed [9:0] m39_110;
   assign m39_110 =10'b0;

   // m39_111 = W*in
   wire signed [9:0] m39_111;
   assign m39_111 =10'b0;

   // m39_112 = W*in
   wire signed [9:0] m39_112;
   assign m39_112 =10'b0;

   // m39_113 = W*in
   wire signed [9:0] m39_113;
   assign m39_113 =10'b0;

   // m39_114 = W*in
   wire signed [9:0] m39_114;
   assign m39_114 =10'b0;

   // m39_115 = W*in
   wire signed [9:0] m39_115;
   assign m39_115 =10'b0;

   // m39_116 = W*in
   wire signed [9:0] m39_116;
   assign m39_116 =10'b0;

   // m39_117 = W*in
   wire signed [9:0] m39_117;
   assign m39_117 =10'b0;

   // m40_1 = W*in
   wire signed [9:0] m40_1;
   assign m40_1 =10'b0;

   // m40_2 = W*in
   wire signed [9:0] m40_2;
   assign m40_2 =10'b0;

   // m40_3 = W*in
   wire signed [9:0] m40_3;
   assign m40_3 =10'b0;

   // m40_4 = W*in
   wire signed [9:0] m40_4;
   assign m40_4 =10'b0;

   // m40_5 = W*in
   wire signed [9:0] m40_5;
   assign m40_5 =10'b0;

   // m40_6 = W*in
   wire signed [9:0] m40_6;
   assign m40_6 =10'b0;

   // m40_7 = W*in
   wire signed [9:0] m40_7;
   assign m40_7 =10'b0;

   // m40_8 = W*in
   wire signed [9:0] m40_8;
   assign m40_8 =10'b0;

   // m40_9 = W*in
   wire signed [9:0] m40_9;
   assign m40_9 =10'b0;

   // m40_10 = W*in
   wire signed [9:0] m40_10;
   assign m40_10 =10'b0;

   // m40_11 = W*in
   wire signed [9:0] m40_11;
   assign m40_11 =10'b0;

   // m40_12 = W*in
   wire signed [9:0] m40_12;
   assign m40_12 =10'b0;

   // m40_13 = W*in
   wire signed [9:0] m40_13;
   assign m40_13 =10'b0;

   // m40_14 = W*in
   wire signed [9:0] m40_14;
   assign m40_14 =10'b0;

   // m40_15 = W*in
   wire signed [9:0] m40_15;
   assign m40_15 =10'b0;

   // m40_16 = W*in
   wire signed [9:0] m40_16;
   assign m40_16 =10'b0;

   // m40_17 = W*in
   wire signed [9:0] m40_17;
   assign m40_17 =10'b0;

   // m40_18 = W*in
   wire signed [9:0] m40_18;
   assign m40_18 =10'b0;

   // m40_19 = W*in
   wire signed [9:0] m40_19;
   assign m40_19 =10'b0;

   // m40_20 = W*in
   wire signed [9:0] m40_20;
   assign m40_20 ={ {5{neg40[5]}} , neg40[5:1] };

   // m40_21 = W*in
   wire signed [9:0] m40_21;
   assign m40_21 =10'b0;

   // m40_22 = W*in
   wire signed [9:0] m40_22;
   assign m40_22 =10'b0;

   // m40_23 = W*in
   wire signed [9:0] m40_23;
   assign m40_23 =10'b0;

   // m40_24 = W*in
   wire signed [9:0] m40_24;
   assign m40_24 =10'b0;

   // m40_25 = W*in
   wire signed [9:0] m40_25;
   assign m40_25 =10'b0;

   // m40_26 = W*in
   wire signed [9:0] m40_26;
   assign m40_26 ={ {4{in40[5]}} , in40[5:0] };

   // m40_27 = W*in
   wire signed [9:0] m40_27;
   assign m40_27 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_28 = W*in
   wire signed [9:0] m40_28;
   assign m40_28 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_29 = W*in
   wire signed [9:0] m40_29;
   assign m40_29 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_30 = W*in
   wire signed [9:0] m40_30;
   assign m40_30 =10'b0;

   // m40_31 = W*in
   wire signed [9:0] m40_31;
   assign m40_31 =10'b0;

   // m40_32 = W*in
   wire signed [9:0] m40_32;
   assign m40_32 =10'b0;

   // m40_33 = W*in
   wire signed [9:0] m40_33;
   assign m40_33 =10'b0;

   // m40_34 = W*in
   wire signed [9:0] m40_34;
   assign m40_34 =10'b0;

   // m40_35 = W*in
   wire signed [9:0] m40_35;
   assign m40_35 ={ {5{neg40[5]}} , neg40[5:1] };

   // m40_36 = W*in
   wire signed [9:0] m40_36;
   assign m40_36 =10'b0;

   // m40_37 = W*in
   wire signed [9:0] m40_37;
   assign m40_37 =10'b0;

   // m40_38 = W*in
   wire signed [9:0] m40_38;
   assign m40_38 =10'b0;

   // m40_39 = W*in
   wire signed [9:0] m40_39;
   assign m40_39 =10'b0;

   // m40_40 = W*in
   wire signed [9:0] m40_40;
   assign m40_40 =10'b0;

   // m40_41 = W*in
   wire signed [9:0] m40_41;
   assign m40_41 =10'b0;

   // m40_42 = W*in
   wire signed [9:0] m40_42;
   assign m40_42 ={ {4{in40[5]}} , in40[5:0] };

   // m40_43 = W*in
   wire signed [9:0] m40_43;
   assign m40_43 =10'b0;

   // m40_44 = W*in
   wire signed [9:0] m40_44;
   assign m40_44 =10'b0;

   // m40_45 = W*in
   wire signed [9:0] m40_45;
   assign m40_45 =10'b0;

   // m40_46 = W*in
   wire signed [9:0] m40_46;
   assign m40_46 =10'b0;

   // m40_47 = W*in
   wire signed [9:0] m40_47;
   assign m40_47 =10'b0;

   // m40_48 = W*in
   wire signed [9:0] m40_48;
   assign m40_48 =10'b0;

   // m40_49 = W*in
   wire signed [9:0] m40_49;
   assign m40_49 =10'b0;

   // m40_50 = W*in
   wire signed [9:0] m40_50;
   assign m40_50 =10'b0;

   // m40_51 = W*in
   wire signed [9:0] m40_51;
   assign m40_51 =10'b0;

   // m40_52 = W*in
   wire signed [9:0] m40_52;
   assign m40_52 =10'b0;

   // m40_53 = W*in
   wire signed [9:0] m40_53;
   assign m40_53 =10'b0;

   // m40_54 = W*in
   wire signed [9:0] m40_54;
   assign m40_54 =10'b0;

   // m40_55 = W*in
   wire signed [9:0] m40_55;
   assign m40_55 =10'b0;

   // m40_56 = W*in
   wire signed [9:0] m40_56;
   assign m40_56 =10'b0;

   // m40_57 = W*in
   wire signed [9:0] m40_57;
   assign m40_57 =10'b0;

   // m40_58 = W*in
   wire signed [9:0] m40_58;
   assign m40_58 =10'b0;

   // m40_59 = W*in
   wire signed [9:0] m40_59;
   assign m40_59 =10'b0;

   // m40_60 = W*in
   wire signed [9:0] m40_60;
   assign m40_60 =10'b0;

   // m40_61 = W*in
   wire signed [9:0] m40_61;
   assign m40_61 =10'b0;

   // m40_62 = W*in
   wire signed [9:0] m40_62;
   assign m40_62 =10'b0;

   // m40_63 = W*in
   wire signed [9:0] m40_63;
   assign m40_63 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_64 = W*in
   wire signed [9:0] m40_64;
   assign m40_64 ={ {5{in40[5]}} , in40[5:1] };

   // m40_65 = W*in
   wire signed [9:0] m40_65;
   assign m40_65 =10'b0;

   // m40_66 = W*in
   wire signed [9:0] m40_66;
   assign m40_66 ={ {5{in40[5]}} , in40[5:1] };

   // m40_67 = W*in
   wire signed [9:0] m40_67;
   assign m40_67 =10'b0;

   // m40_68 = W*in
   wire signed [9:0] m40_68;
   assign m40_68 =10'b0;

   // m40_69 = W*in
   wire signed [9:0] m40_69;
   assign m40_69 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_70 = W*in
   wire signed [9:0] m40_70;
   assign m40_70 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_71 = W*in
   wire signed [9:0] m40_71;
   assign m40_71 =10'b0;

   // m40_72 = W*in
   wire signed [9:0] m40_72;
   assign m40_72 ={ {5{neg40[5]}} , neg40[5:1] };

   // m40_73 = W*in
   wire signed [9:0] m40_73;
   assign m40_73 =10'b0;

   // m40_74 = W*in
   wire signed [9:0] m40_74;
   assign m40_74 =10'b0;

   // m40_75 = W*in
   wire signed [9:0] m40_75;
   assign m40_75 ={ {4{in40[5]}} , in40[5:0] };

   // m40_76 = W*in
   wire signed [9:0] m40_76;
   assign m40_76 =10'b0;

   // m40_77 = W*in
   wire signed [9:0] m40_77;
   assign m40_77 ={ {4{in40[5]}} , in40[5:0] };

   // m40_78 = W*in
   wire signed [9:0] m40_78;
   assign m40_78 =10'b0;

   // m40_79 = W*in
   wire signed [9:0] m40_79;
   assign m40_79 =10'b0;

   // m40_80 = W*in
   wire signed [9:0] m40_80;
   assign m40_80 =10'b0;

   // m40_81 = W*in
   wire signed [9:0] m40_81;
   assign m40_81 ={ {5{in40[5]}} , in40[5:1] };

   // m40_82 = W*in
   wire signed [9:0] m40_82;
   assign m40_82 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_83 = W*in
   wire signed [9:0] m40_83;
   assign m40_83 =10'b0;

   // m40_84 = W*in
   wire signed [9:0] m40_84;
   assign m40_84 =10'b0;

   // m40_85 = W*in
   wire signed [9:0] m40_85;
   assign m40_85 =10'b0;

   // m40_86 = W*in
   wire signed [9:0] m40_86;
   assign m40_86 =10'b0;

   // m40_87 = W*in
   wire signed [9:0] m40_87;
   assign m40_87 =10'b0;

   // m40_88 = W*in
   wire signed [9:0] m40_88;
   assign m40_88 =10'b0;

   // m40_89 = W*in
   wire signed [9:0] m40_89;
   assign m40_89 =10'b0;

   // m40_90 = W*in
   wire signed [9:0] m40_90;
   assign m40_90 =10'b0;

   // m40_91 = W*in
   wire signed [9:0] m40_91;
   assign m40_91 =10'b0;

   // m40_92 = W*in
   wire signed [9:0] m40_92;
   assign m40_92 =10'b0;

   // m40_93 = W*in
   wire signed [9:0] m40_93;
   assign m40_93 =10'b0;

   // m40_94 = W*in
   wire signed [9:0] m40_94;
   assign m40_94 ={ {4{in40[5]}} , in40[5:0] };

   // m40_95 = W*in
   wire signed [9:0] m40_95;
   assign m40_95 ={ {4{neg40[5]}} , neg40[5:0] };

   // m40_96 = W*in
   wire signed [9:0] m40_96;
   assign m40_96 =10'b0;

   // m40_97 = W*in
   wire signed [9:0] m40_97;
   assign m40_97 =10'b0;

   // m40_98 = W*in
   wire signed [9:0] m40_98;
   assign m40_98 =10'b0;

   // m40_99 = W*in
   wire signed [9:0] m40_99;
   assign m40_99 =10'b0;

   // m40_100 = W*in
   wire signed [9:0] m40_100;
   assign m40_100 ={ {4{in40[5]}} , in40[5:0] };

   // m40_101 = W*in
   wire signed [9:0] m40_101;
   assign m40_101 =10'b0;

   // m40_102 = W*in
   wire signed [9:0] m40_102;
   assign m40_102 =10'b0;

   // m40_103 = W*in
   wire signed [9:0] m40_103;
   assign m40_103 =10'b0;

   // m40_104 = W*in
   wire signed [9:0] m40_104;
   assign m40_104 =10'b0;

   // m40_105 = W*in
   wire signed [9:0] m40_105;
   assign m40_105 =10'b0;

   // m40_106 = W*in
   wire signed [9:0] m40_106;
   assign m40_106 =10'b0;

   // m40_107 = W*in
   wire signed [9:0] m40_107;
   assign m40_107 =10'b0;

   // m40_108 = W*in
   wire signed [9:0] m40_108;
   assign m40_108 =10'b0;

   // m40_109 = W*in
   wire signed [9:0] m40_109;
   assign m40_109 ={ {5{neg40[5]}} , neg40[5:1] };

   // m40_110 = W*in
   wire signed [9:0] m40_110;
   assign m40_110 =10'b0;

   // m40_111 = W*in
   wire signed [9:0] m40_111;
   assign m40_111 =10'b0;

   // m40_112 = W*in
   wire signed [9:0] m40_112;
   assign m40_112 =10'b0;

   // m40_113 = W*in
   wire signed [9:0] m40_113;
   assign m40_113 =10'b0;

   // m40_114 = W*in
   wire signed [9:0] m40_114;
   assign m40_114 =10'b0;

   // m40_115 = W*in
   wire signed [9:0] m40_115;
   assign m40_115 =10'b0;

   // m40_116 = W*in
   wire signed [9:0] m40_116;
   assign m40_116 =10'b0;

   // m40_117 = W*in
   wire signed [9:0] m40_117;
   assign m40_117 ={ {4{neg40[5]}} , neg40[5:0] };

   // m41_1 = W*in
   wire signed [9:0] m41_1;
   assign m41_1 ={ {4{in41[5]}} , in41[5:0] };

   // m41_2 = W*in
   wire signed [9:0] m41_2;
   assign m41_2 ={ {4{in41[5]}} , in41[5:0] };

   // m41_3 = W*in
   wire signed [9:0] m41_3;
   assign m41_3 =10'b0;

   // m41_4 = W*in
   wire signed [9:0] m41_4;
   assign m41_4 =10'b0;

   // m41_5 = W*in
   wire signed [9:0] m41_5;
   assign m41_5 =10'b0;

   // m41_6 = W*in
   wire signed [9:0] m41_6;
   assign m41_6 =10'b0;

   // m41_7 = W*in
   wire signed [9:0] m41_7;
   assign m41_7 =10'b0;

   // m41_8 = W*in
   wire signed [9:0] m41_8;
   assign m41_8 ={ {4{in41[5]}} , in41[5:0] };

   // m41_9 = W*in
   wire signed [9:0] m41_9;
   assign m41_9 =10'b0;

   // m41_10 = W*in
   wire signed [9:0] m41_10;
   assign m41_10 =10'b0;

   // m41_11 = W*in
   wire signed [9:0] m41_11;
   assign m41_11 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_12 = W*in
   wire signed [9:0] m41_12;
   assign m41_12 =10'b0;

   // m41_13 = W*in
   wire signed [9:0] m41_13;
   assign m41_13 =10'b0;

   // m41_14 = W*in
   wire signed [9:0] m41_14;
   assign m41_14 =10'b0;

   // m41_15 = W*in
   wire signed [9:0] m41_15;
   assign m41_15 ={ {4{in41[5]}} , in41[5:0] };

   // m41_16 = W*in
   wire signed [9:0] m41_16;
   assign m41_16 =10'b0;

   // m41_17 = W*in
   wire signed [9:0] m41_17;
   assign m41_17 =10'b0;

   // m41_18 = W*in
   wire signed [9:0] m41_18;
   assign m41_18 =10'b0;

   // m41_19 = W*in
   wire signed [9:0] m41_19;
   assign m41_19 =10'b0;

   // m41_20 = W*in
   wire signed [9:0] m41_20;
   assign m41_20 =10'b0;

   // m41_21 = W*in
   wire signed [9:0] m41_21;
   assign m41_21 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_22 = W*in
   wire signed [9:0] m41_22;
   assign m41_22 =10'b0;

   // m41_23 = W*in
   wire signed [9:0] m41_23;
   assign m41_23 =10'b0;

   // m41_24 = W*in
   wire signed [9:0] m41_24;
   assign m41_24 =10'b0;

   // m41_25 = W*in
   wire signed [9:0] m41_25;
   assign m41_25 ={ {4{in41[5]}} , in41[5:0] };

   // m41_26 = W*in
   wire signed [9:0] m41_26;
   assign m41_26 ={ {5{in41[5]}} , in41[5:1] };

   // m41_27 = W*in
   wire signed [9:0] m41_27;
   assign m41_27 ={ {5{neg41[5]}} , neg41[5:1] };

   // m41_28 = W*in
   wire signed [9:0] m41_28;
   assign m41_28 =10'b0;

   // m41_29 = W*in
   wire signed [9:0] m41_29;
   assign m41_29 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_30 = W*in
   wire signed [9:0] m41_30;
   assign m41_30 =10'b0;

   // m41_31 = W*in
   wire signed [9:0] m41_31;
   assign m41_31 =10'b0;

   // m41_32 = W*in
   wire signed [9:0] m41_32;
   assign m41_32 =10'b0;

   // m41_33 = W*in
   wire signed [9:0] m41_33;
   assign m41_33 ={ {4{in41[5]}} , in41[5:0] };

   // m41_34 = W*in
   wire signed [9:0] m41_34;
   assign m41_34 =10'b0;

   // m41_35 = W*in
   wire signed [9:0] m41_35;
   assign m41_35 =10'b0;

   // m41_36 = W*in
   wire signed [9:0] m41_36;
   assign m41_36 ={ {4{in41[5]}} , in41[5:0] };

   // m41_37 = W*in
   wire signed [9:0] m41_37;
   assign m41_37 =10'b0;

   // m41_38 = W*in
   wire signed [9:0] m41_38;
   assign m41_38 =10'b0;

   // m41_39 = W*in
   wire signed [9:0] m41_39;
   assign m41_39 =10'b0;

   // m41_40 = W*in
   wire signed [9:0] m41_40;
   assign m41_40 =10'b0;

   // m41_41 = W*in
   wire signed [9:0] m41_41;
   assign m41_41 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_42 = W*in
   wire signed [9:0] m41_42;
   assign m41_42 =10'b0;

   // m41_43 = W*in
   wire signed [9:0] m41_43;
   assign m41_43 =10'b0;

   // m41_44 = W*in
   wire signed [9:0] m41_44;
   assign m41_44 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_45 = W*in
   wire signed [9:0] m41_45;
   assign m41_45 ={ {4{in41[5]}} , in41[5:0] };

   // m41_46 = W*in
   wire signed [9:0] m41_46;
   assign m41_46 =10'b0;

   // m41_47 = W*in
   wire signed [9:0] m41_47;
   assign m41_47 =10'b0;

   // m41_48 = W*in
   wire signed [9:0] m41_48;
   assign m41_48 =10'b0;

   // m41_49 = W*in
   wire signed [9:0] m41_49;
   assign m41_49 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_50 = W*in
   wire signed [9:0] m41_50;
   assign m41_50 =10'b0;

   // m41_51 = W*in
   wire signed [9:0] m41_51;
   assign m41_51 ={ {4{in41[5]}} , in41[5:0] };

   // m41_52 = W*in
   wire signed [9:0] m41_52;
   assign m41_52 =10'b0;

   // m41_53 = W*in
   wire signed [9:0] m41_53;
   assign m41_53 =10'b0;

   // m41_54 = W*in
   wire signed [9:0] m41_54;
   assign m41_54 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_55 = W*in
   wire signed [9:0] m41_55;
   assign m41_55 =10'b0;

   // m41_56 = W*in
   wire signed [9:0] m41_56;
   assign m41_56 ={ {4{in41[5]}} , in41[5:0] };

   // m41_57 = W*in
   wire signed [9:0] m41_57;
   assign m41_57 =10'b0;

   // m41_58 = W*in
   wire signed [9:0] m41_58;
   assign m41_58 =10'b0;

   // m41_59 = W*in
   wire signed [9:0] m41_59;
   assign m41_59 =10'b0;

   // m41_60 = W*in
   wire signed [9:0] m41_60;
   assign m41_60 =10'b0;

   // m41_61 = W*in
   wire signed [9:0] m41_61;
   assign m41_61 =10'b0;

   // m41_62 = W*in
   wire signed [9:0] m41_62;
   assign m41_62 =10'b0;

   // m41_63 = W*in
   wire signed [9:0] m41_63;
   assign m41_63 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_64 = W*in
   wire signed [9:0] m41_64;
   assign m41_64 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_65 = W*in
   wire signed [9:0] m41_65;
   assign m41_65 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_66 = W*in
   wire signed [9:0] m41_66;
   assign m41_66 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_67 = W*in
   wire signed [9:0] m41_67;
   assign m41_67 =10'b0;

   // m41_68 = W*in
   wire signed [9:0] m41_68;
   assign m41_68 ={ {4{in41[5]}} , in41[5:0] };

   // m41_69 = W*in
   wire signed [9:0] m41_69;
   assign m41_69 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_70 = W*in
   wire signed [9:0] m41_70;
   assign m41_70 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_71 = W*in
   wire signed [9:0] m41_71;
   assign m41_71 =10'b0;

   // m41_72 = W*in
   wire signed [9:0] m41_72;
   assign m41_72 =10'b0;

   // m41_73 = W*in
   wire signed [9:0] m41_73;
   assign m41_73 ={ {4{in41[5]}} , in41[5:0] };

   // m41_74 = W*in
   wire signed [9:0] m41_74;
   assign m41_74 =10'b0;

   // m41_75 = W*in
   wire signed [9:0] m41_75;
   assign m41_75 ={ {5{in41[5]}} , in41[5:1] };

   // m41_76 = W*in
   wire signed [9:0] m41_76;
   assign m41_76 =10'b0;

   // m41_77 = W*in
   wire signed [9:0] m41_77;
   assign m41_77 =10'b0;

   // m41_78 = W*in
   wire signed [9:0] m41_78;
   assign m41_78 ={ {4{in41[5]}} , in41[5:0] };

   // m41_79 = W*in
   wire signed [9:0] m41_79;
   assign m41_79 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_80 = W*in
   wire signed [9:0] m41_80;
   assign m41_80 =10'b0;

   // m41_81 = W*in
   wire signed [9:0] m41_81;
   assign m41_81 =10'b0;

   // m41_82 = W*in
   wire signed [9:0] m41_82;
   assign m41_82 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_83 = W*in
   wire signed [9:0] m41_83;
   assign m41_83 =10'b0;

   // m41_84 = W*in
   wire signed [9:0] m41_84;
   assign m41_84 =10'b0;

   // m41_85 = W*in
   wire signed [9:0] m41_85;
   assign m41_85 =10'b0;

   // m41_86 = W*in
   wire signed [9:0] m41_86;
   assign m41_86 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_87 = W*in
   wire signed [9:0] m41_87;
   assign m41_87 =10'b0;

   // m41_88 = W*in
   wire signed [9:0] m41_88;
   assign m41_88 =10'b0;

   // m41_89 = W*in
   wire signed [9:0] m41_89;
   assign m41_89 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_90 = W*in
   wire signed [9:0] m41_90;
   assign m41_90 ={ {4{in41[5]}} , in41[5:0] };

   // m41_91 = W*in
   wire signed [9:0] m41_91;
   assign m41_91 =10'b0;

   // m41_92 = W*in
   wire signed [9:0] m41_92;
   assign m41_92 =10'b0;

   // m41_93 = W*in
   wire signed [9:0] m41_93;
   assign m41_93 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_94 = W*in
   wire signed [9:0] m41_94;
   assign m41_94 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_95 = W*in
   wire signed [9:0] m41_95;
   assign m41_95 =10'b0;

   // m41_96 = W*in
   wire signed [9:0] m41_96;
   assign m41_96 =10'b0;

   // m41_97 = W*in
   wire signed [9:0] m41_97;
   assign m41_97 =10'b0;

   // m41_98 = W*in
   wire signed [9:0] m41_98;
   assign m41_98 =10'b0;

   // m41_99 = W*in
   wire signed [9:0] m41_99;
   assign m41_99 =10'b0;

   // m41_100 = W*in
   wire signed [9:0] m41_100;
   assign m41_100 =10'b0;

   // m41_101 = W*in
   wire signed [9:0] m41_101;
   assign m41_101 =10'b0;

   // m41_102 = W*in
   wire signed [9:0] m41_102;
   assign m41_102 ={ {4{in41[5]}} , in41[5:0] };

   // m41_103 = W*in
   wire signed [9:0] m41_103;
   assign m41_103 =10'b0;

   // m41_104 = W*in
   wire signed [9:0] m41_104;
   assign m41_104 =10'b0;

   // m41_105 = W*in
   wire signed [9:0] m41_105;
   assign m41_105 =10'b0;

   // m41_106 = W*in
   wire signed [9:0] m41_106;
   assign m41_106 =10'b0;

   // m41_107 = W*in
   wire signed [9:0] m41_107;
   assign m41_107 ={ {4{in41[5]}} , in41[5:0] };

   // m41_108 = W*in
   wire signed [9:0] m41_108;
   assign m41_108 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_109 = W*in
   wire signed [9:0] m41_109;
   assign m41_109 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_110 = W*in
   wire signed [9:0] m41_110;
   assign m41_110 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_111 = W*in
   wire signed [9:0] m41_111;
   assign m41_111 ={ {3{in41[5]}} , in41 , {1{1'b0}} };

   // m41_112 = W*in
   wire signed [9:0] m41_112;
   assign m41_112 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_113 = W*in
   wire signed [9:0] m41_113;
   assign m41_113 ={ {4{in41[5]}} , in41[5:0] };

   // m41_114 = W*in
   wire signed [9:0] m41_114;
   assign m41_114 =10'b0;

   // m41_115 = W*in
   wire signed [9:0] m41_115;
   assign m41_115 =10'b0;

   // m41_116 = W*in
   wire signed [9:0] m41_116;
   assign m41_116 ={ {4{neg41[5]}} , neg41[5:0] };

   // m41_117 = W*in
   wire signed [9:0] m41_117;
   assign m41_117 =10'b0;

   // m42_1 = W*in
   wire signed [9:0] m42_1;
   assign m42_1 =10'b0;

   // m42_2 = W*in
   wire signed [9:0] m42_2;
   assign m42_2 =10'b0;

   // m42_3 = W*in
   wire signed [9:0] m42_3;
   assign m42_3 =10'b0;

   // m42_4 = W*in
   wire signed [9:0] m42_4;
   assign m42_4 =10'b0;

   // m42_5 = W*in
   wire signed [9:0] m42_5;
   assign m42_5 ={ {4{in42[5]}} , in42[5:0] };

   // m42_6 = W*in
   wire signed [9:0] m42_6;
   assign m42_6 =10'b0;

   // m42_7 = W*in
   wire signed [9:0] m42_7;
   assign m42_7 =10'b0;

   // m42_8 = W*in
   wire signed [9:0] m42_8;
   assign m42_8 =10'b0;

   // m42_9 = W*in
   wire signed [9:0] m42_9;
   assign m42_9 =10'b0;

   // m42_10 = W*in
   wire signed [9:0] m42_10;
   assign m42_10 =10'b0;

   // m42_11 = W*in
   wire signed [9:0] m42_11;
   assign m42_11 =10'b0;

   // m42_12 = W*in
   wire signed [9:0] m42_12;
   assign m42_12 =10'b0;

   // m42_13 = W*in
   wire signed [9:0] m42_13;
   assign m42_13 =10'b0;

   // m42_14 = W*in
   wire signed [9:0] m42_14;
   assign m42_14 =10'b0;

   // m42_15 = W*in
   wire signed [9:0] m42_15;
   assign m42_15 ={ {4{in42[5]}} , in42[5:0] };

   // m42_16 = W*in
   wire signed [9:0] m42_16;
   assign m42_16 =10'b0;

   // m42_17 = W*in
   wire signed [9:0] m42_17;
   assign m42_17 =10'b0;

   // m42_18 = W*in
   wire signed [9:0] m42_18;
   assign m42_18 =10'b0;

   // m42_19 = W*in
   wire signed [9:0] m42_19;
   assign m42_19 =10'b0;

   // m42_20 = W*in
   wire signed [9:0] m42_20;
   assign m42_20 =10'b0;

   // m42_21 = W*in
   wire signed [9:0] m42_21;
   assign m42_21 =10'b0;

   // m42_22 = W*in
   wire signed [9:0] m42_22;
   assign m42_22 ={ {5{neg42[5]}} , neg42[5:1] };

   // m42_23 = W*in
   wire signed [9:0] m42_23;
   assign m42_23 =10'b0;

   // m42_24 = W*in
   wire signed [9:0] m42_24;
   assign m42_24 =10'b0;

   // m42_25 = W*in
   wire signed [9:0] m42_25;
   assign m42_25 =10'b0;

   // m42_26 = W*in
   wire signed [9:0] m42_26;
   assign m42_26 =10'b0;

   // m42_27 = W*in
   wire signed [9:0] m42_27;
   assign m42_27 =10'b0;

   // m42_28 = W*in
   wire signed [9:0] m42_28;
   assign m42_28 ={ {4{in42[5]}} , in42[5:0] };

   // m42_29 = W*in
   wire signed [9:0] m42_29;
   assign m42_29 =10'b0;

   // m42_30 = W*in
   wire signed [9:0] m42_30;
   assign m42_30 =10'b0;

   // m42_31 = W*in
   wire signed [9:0] m42_31;
   assign m42_31 =10'b0;

   // m42_32 = W*in
   wire signed [9:0] m42_32;
   assign m42_32 =10'b0;

   // m42_33 = W*in
   wire signed [9:0] m42_33;
   assign m42_33 =10'b0;

   // m42_34 = W*in
   wire signed [9:0] m42_34;
   assign m42_34 =10'b0;

   // m42_35 = W*in
   wire signed [9:0] m42_35;
   assign m42_35 =10'b0;

   // m42_36 = W*in
   wire signed [9:0] m42_36;
   assign m42_36 =10'b0;

   // m42_37 = W*in
   wire signed [9:0] m42_37;
   assign m42_37 =10'b0;

   // m42_38 = W*in
   wire signed [9:0] m42_38;
   assign m42_38 =10'b0;

   // m42_39 = W*in
   wire signed [9:0] m42_39;
   assign m42_39 =10'b0;

   // m42_40 = W*in
   wire signed [9:0] m42_40;
   assign m42_40 =10'b0;

   // m42_41 = W*in
   wire signed [9:0] m42_41;
   assign m42_41 =10'b0;

   // m42_42 = W*in
   wire signed [9:0] m42_42;
   assign m42_42 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_43 = W*in
   wire signed [9:0] m42_43;
   assign m42_43 ={ {4{in42[5]}} , in42[5:0] };

   // m42_44 = W*in
   wire signed [9:0] m42_44;
   assign m42_44 =10'b0;

   // m42_45 = W*in
   wire signed [9:0] m42_45;
   assign m42_45 =10'b0;

   // m42_46 = W*in
   wire signed [9:0] m42_46;
   assign m42_46 =10'b0;

   // m42_47 = W*in
   wire signed [9:0] m42_47;
   assign m42_47 =10'b0;

   // m42_48 = W*in
   wire signed [9:0] m42_48;
   assign m42_48 ={ {4{in42[5]}} , in42[5:0] };

   // m42_49 = W*in
   wire signed [9:0] m42_49;
   assign m42_49 =10'b0;

   // m42_50 = W*in
   wire signed [9:0] m42_50;
   assign m42_50 =10'b0;

   // m42_51 = W*in
   wire signed [9:0] m42_51;
   assign m42_51 ={ {4{in42[5]}} , in42[5:0] };

   // m42_52 = W*in
   wire signed [9:0] m42_52;
   assign m42_52 =10'b0;

   // m42_53 = W*in
   wire signed [9:0] m42_53;
   assign m42_53 =10'b0;

   // m42_54 = W*in
   wire signed [9:0] m42_54;
   assign m42_54 =10'b0;

   // m42_55 = W*in
   wire signed [9:0] m42_55;
   assign m42_55 =10'b0;

   // m42_56 = W*in
   wire signed [9:0] m42_56;
   assign m42_56 =10'b0;

   // m42_57 = W*in
   wire signed [9:0] m42_57;
   assign m42_57 =10'b0;

   // m42_58 = W*in
   wire signed [9:0] m42_58;
   assign m42_58 =10'b0;

   // m42_59 = W*in
   wire signed [9:0] m42_59;
   assign m42_59 ={ {4{in42[5]}} , in42[5:0] };

   // m42_60 = W*in
   wire signed [9:0] m42_60;
   assign m42_60 =10'b0;

   // m42_61 = W*in
   wire signed [9:0] m42_61;
   assign m42_61 =10'b0;

   // m42_62 = W*in
   wire signed [9:0] m42_62;
   assign m42_62 =10'b0;

   // m42_63 = W*in
   wire signed [9:0] m42_63;
   assign m42_63 =10'b0;

   // m42_64 = W*in
   wire signed [9:0] m42_64;
   assign m42_64 ={ {3{neg42[5]}} , neg42 , {1{1'b0}} };

   // m42_65 = W*in
   wire signed [9:0] m42_65;
   assign m42_65 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_66 = W*in
   wire signed [9:0] m42_66;
   assign m42_66 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_67 = W*in
   wire signed [9:0] m42_67;
   assign m42_67 =10'b0;

   // m42_68 = W*in
   wire signed [9:0] m42_68;
   assign m42_68 ={ {4{in42[5]}} , in42[5:0] };

   // m42_69 = W*in
   wire signed [9:0] m42_69;
   assign m42_69 =10'b0;

   // m42_70 = W*in
   wire signed [9:0] m42_70;
   assign m42_70 ={ {4{in42[5]}} , in42[5:0] };

   // m42_71 = W*in
   wire signed [9:0] m42_71;
   assign m42_71 ={ {4{in42[5]}} , in42[5:0] };

   // m42_72 = W*in
   wire signed [9:0] m42_72;
   assign m42_72 ={ {4{in42[5]}} , in42[5:0] };

   // m42_73 = W*in
   wire signed [9:0] m42_73;
   assign m42_73 =10'b0;

   // m42_74 = W*in
   wire signed [9:0] m42_74;
   assign m42_74 =10'b0;

   // m42_75 = W*in
   wire signed [9:0] m42_75;
   assign m42_75 =10'b0;

   // m42_76 = W*in
   wire signed [9:0] m42_76;
   assign m42_76 =10'b0;

   // m42_77 = W*in
   wire signed [9:0] m42_77;
   assign m42_77 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_78 = W*in
   wire signed [9:0] m42_78;
   assign m42_78 =10'b0;

   // m42_79 = W*in
   wire signed [9:0] m42_79;
   assign m42_79 =10'b0;

   // m42_80 = W*in
   wire signed [9:0] m42_80;
   assign m42_80 =10'b0;

   // m42_81 = W*in
   wire signed [9:0] m42_81;
   assign m42_81 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_82 = W*in
   wire signed [9:0] m42_82;
   assign m42_82 ={ {5{neg42[5]}} , neg42[5:1] };

   // m42_83 = W*in
   wire signed [9:0] m42_83;
   assign m42_83 =10'b0;

   // m42_84 = W*in
   wire signed [9:0] m42_84;
   assign m42_84 =10'b0;

   // m42_85 = W*in
   wire signed [9:0] m42_85;
   assign m42_85 ={ {5{neg42[5]}} , neg42[5:1] };

   // m42_86 = W*in
   wire signed [9:0] m42_86;
   assign m42_86 =10'b0;

   // m42_87 = W*in
   wire signed [9:0] m42_87;
   assign m42_87 =10'b0;

   // m42_88 = W*in
   wire signed [9:0] m42_88;
   assign m42_88 ={ {4{in42[5]}} , in42[5:0] };

   // m42_89 = W*in
   wire signed [9:0] m42_89;
   assign m42_89 =10'b0;

   // m42_90 = W*in
   wire signed [9:0] m42_90;
   assign m42_90 ={ {4{in42[5]}} , in42[5:0] };

   // m42_91 = W*in
   wire signed [9:0] m42_91;
   assign m42_91 =10'b0;

   // m42_92 = W*in
   wire signed [9:0] m42_92;
   assign m42_92 ={ {4{in42[5]}} , in42[5:0] };

   // m42_93 = W*in
   wire signed [9:0] m42_93;
   assign m42_93 =10'b0;

   // m42_94 = W*in
   wire signed [9:0] m42_94;
   assign m42_94 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_95 = W*in
   wire signed [9:0] m42_95;
   assign m42_95 =10'b0;

   // m42_96 = W*in
   wire signed [9:0] m42_96;
   assign m42_96 =10'b0;

   // m42_97 = W*in
   wire signed [9:0] m42_97;
   assign m42_97 =10'b0;

   // m42_98 = W*in
   wire signed [9:0] m42_98;
   assign m42_98 =10'b0;

   // m42_99 = W*in
   wire signed [9:0] m42_99;
   assign m42_99 =10'b0;

   // m42_100 = W*in
   wire signed [9:0] m42_100;
   assign m42_100 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_101 = W*in
   wire signed [9:0] m42_101;
   assign m42_101 =10'b0;

   // m42_102 = W*in
   wire signed [9:0] m42_102;
   assign m42_102 =10'b0;

   // m42_103 = W*in
   wire signed [9:0] m42_103;
   assign m42_103 =10'b0;

   // m42_104 = W*in
   wire signed [9:0] m42_104;
   assign m42_104 =10'b0;

   // m42_105 = W*in
   wire signed [9:0] m42_105;
   assign m42_105 =10'b0;

   // m42_106 = W*in
   wire signed [9:0] m42_106;
   assign m42_106 =10'b0;

   // m42_107 = W*in
   wire signed [9:0] m42_107;
   assign m42_107 =10'b0;

   // m42_108 = W*in
   wire signed [9:0] m42_108;
   assign m42_108 ={ {5{neg42[5]}} , neg42[5:1] };

   // m42_109 = W*in
   wire signed [9:0] m42_109;
   assign m42_109 ={ {5{neg42[5]}} , neg42[5:1] };

   // m42_110 = W*in
   wire signed [9:0] m42_110;
   assign m42_110 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_111 = W*in
   wire signed [9:0] m42_111;
   assign m42_111 ={ {4{in42[5]}} , in42[5:0] };

   // m42_112 = W*in
   wire signed [9:0] m42_112;
   assign m42_112 ={ {4{neg42[5]}} , neg42[5:0] };

   // m42_113 = W*in
   wire signed [9:0] m42_113;
   assign m42_113 =10'b0;

   // m42_114 = W*in
   wire signed [9:0] m42_114;
   assign m42_114 =10'b0;

   // m42_115 = W*in
   wire signed [9:0] m42_115;
   assign m42_115 ={ {5{neg42[5]}} , neg42[5:1] };

   // m42_116 = W*in
   wire signed [9:0] m42_116;
   assign m42_116 =10'b0;

   // m42_117 = W*in
   wire signed [9:0] m42_117;
   assign m42_117 =10'b0;

   // m43_1 = W*in
   wire signed [9:0] m43_1;
   assign m43_1 =10'b0;

   // m43_2 = W*in
   wire signed [9:0] m43_2;
   assign m43_2 =10'b0;

   // m43_3 = W*in
   wire signed [9:0] m43_3;
   assign m43_3 =10'b0;

   // m43_4 = W*in
   wire signed [9:0] m43_4;
   assign m43_4 =10'b0;

   // m43_5 = W*in
   wire signed [9:0] m43_5;
   assign m43_5 =10'b0;

   // m43_6 = W*in
   wire signed [9:0] m43_6;
   assign m43_6 =10'b0;

   // m43_7 = W*in
   wire signed [9:0] m43_7;
   assign m43_7 =10'b0;

   // m43_8 = W*in
   wire signed [9:0] m43_8;
   assign m43_8 =10'b0;

   // m43_9 = W*in
   wire signed [9:0] m43_9;
   assign m43_9 =10'b0;

   // m43_10 = W*in
   wire signed [9:0] m43_10;
   assign m43_10 =10'b0;

   // m43_11 = W*in
   wire signed [9:0] m43_11;
   assign m43_11 =10'b0;

   // m43_12 = W*in
   wire signed [9:0] m43_12;
   assign m43_12 =10'b0;

   // m43_13 = W*in
   wire signed [9:0] m43_13;
   assign m43_13 =10'b0;

   // m43_14 = W*in
   wire signed [9:0] m43_14;
   assign m43_14 =10'b0;

   // m43_15 = W*in
   wire signed [9:0] m43_15;
   assign m43_15 =10'b0;

   // m43_16 = W*in
   wire signed [9:0] m43_16;
   assign m43_16 =10'b0;

   // m43_17 = W*in
   wire signed [9:0] m43_17;
   assign m43_17 =10'b0;

   // m43_18 = W*in
   wire signed [9:0] m43_18;
   assign m43_18 =10'b0;

   // m43_19 = W*in
   wire signed [9:0] m43_19;
   assign m43_19 =10'b0;

   // m43_20 = W*in
   wire signed [9:0] m43_20;
   assign m43_20 ={ {5{neg43[5]}} , neg43[5:1] };

   // m43_21 = W*in
   wire signed [9:0] m43_21;
   assign m43_21 =10'b0;

   // m43_22 = W*in
   wire signed [9:0] m43_22;
   assign m43_22 =10'b0;

   // m43_23 = W*in
   wire signed [9:0] m43_23;
   assign m43_23 =10'b0;

   // m43_24 = W*in
   wire signed [9:0] m43_24;
   assign m43_24 =10'b0;

   // m43_25 = W*in
   wire signed [9:0] m43_25;
   assign m43_25 =10'b0;

   // m43_26 = W*in
   wire signed [9:0] m43_26;
   assign m43_26 ={ {5{in43[5]}} , in43[5:1] };

   // m43_27 = W*in
   wire signed [9:0] m43_27;
   assign m43_27 =10'b0;

   // m43_28 = W*in
   wire signed [9:0] m43_28;
   assign m43_28 =10'b0;

   // m43_29 = W*in
   wire signed [9:0] m43_29;
   assign m43_29 =10'b0;

   // m43_30 = W*in
   wire signed [9:0] m43_30;
   assign m43_30 =10'b0;

   // m43_31 = W*in
   wire signed [9:0] m43_31;
   assign m43_31 =10'b0;

   // m43_32 = W*in
   wire signed [9:0] m43_32;
   assign m43_32 =10'b0;

   // m43_33 = W*in
   wire signed [9:0] m43_33;
   assign m43_33 =10'b0;

   // m43_34 = W*in
   wire signed [9:0] m43_34;
   assign m43_34 =10'b0;

   // m43_35 = W*in
   wire signed [9:0] m43_35;
   assign m43_35 =10'b0;

   // m43_36 = W*in
   wire signed [9:0] m43_36;
   assign m43_36 =10'b0;

   // m43_37 = W*in
   wire signed [9:0] m43_37;
   assign m43_37 =10'b0;

   // m43_38 = W*in
   wire signed [9:0] m43_38;
   assign m43_38 =10'b0;

   // m43_39 = W*in
   wire signed [9:0] m43_39;
   assign m43_39 =10'b0;

   // m43_40 = W*in
   wire signed [9:0] m43_40;
   assign m43_40 =10'b0;

   // m43_41 = W*in
   wire signed [9:0] m43_41;
   assign m43_41 =10'b0;

   // m43_42 = W*in
   wire signed [9:0] m43_42;
   assign m43_42 =10'b0;

   // m43_43 = W*in
   wire signed [9:0] m43_43;
   assign m43_43 =10'b0;

   // m43_44 = W*in
   wire signed [9:0] m43_44;
   assign m43_44 =10'b0;

   // m43_45 = W*in
   wire signed [9:0] m43_45;
   assign m43_45 =10'b0;

   // m43_46 = W*in
   wire signed [9:0] m43_46;
   assign m43_46 =10'b0;

   // m43_47 = W*in
   wire signed [9:0] m43_47;
   assign m43_47 =10'b0;

   // m43_48 = W*in
   wire signed [9:0] m43_48;
   assign m43_48 =10'b0;

   // m43_49 = W*in
   wire signed [9:0] m43_49;
   assign m43_49 =10'b0;

   // m43_50 = W*in
   wire signed [9:0] m43_50;
   assign m43_50 =10'b0;

   // m43_51 = W*in
   wire signed [9:0] m43_51;
   assign m43_51 =10'b0;

   // m43_52 = W*in
   wire signed [9:0] m43_52;
   assign m43_52 =10'b0;

   // m43_53 = W*in
   wire signed [9:0] m43_53;
   assign m43_53 =10'b0;

   // m43_54 = W*in
   wire signed [9:0] m43_54;
   assign m43_54 =10'b0;

   // m43_55 = W*in
   wire signed [9:0] m43_55;
   assign m43_55 =10'b0;

   // m43_56 = W*in
   wire signed [9:0] m43_56;
   assign m43_56 =10'b0;

   // m43_57 = W*in
   wire signed [9:0] m43_57;
   assign m43_57 =10'b0;

   // m43_58 = W*in
   wire signed [9:0] m43_58;
   assign m43_58 =10'b0;

   // m43_59 = W*in
   wire signed [9:0] m43_59;
   assign m43_59 =10'b0;

   // m43_60 = W*in
   wire signed [9:0] m43_60;
   assign m43_60 =10'b0;

   // m43_61 = W*in
   wire signed [9:0] m43_61;
   assign m43_61 =10'b0;

   // m43_62 = W*in
   wire signed [9:0] m43_62;
   assign m43_62 =10'b0;

   // m43_63 = W*in
   wire signed [9:0] m43_63;
   assign m43_63 =10'b0;

   // m43_64 = W*in
   wire signed [9:0] m43_64;
   assign m43_64 ={ {5{neg43[5]}} , neg43[5:1] };

   // m43_65 = W*in
   wire signed [9:0] m43_65;
   assign m43_65 ={ {5{neg43[5]}} , neg43[5:1] };

   // m43_66 = W*in
   wire signed [9:0] m43_66;
   assign m43_66 ={ {5{neg43[5]}} , neg43[5:1] };

   // m43_67 = W*in
   wire signed [9:0] m43_67;
   assign m43_67 =10'b0;

   // m43_68 = W*in
   wire signed [9:0] m43_68;
   assign m43_68 =10'b0;

   // m43_69 = W*in
   wire signed [9:0] m43_69;
   assign m43_69 =10'b0;

   // m43_70 = W*in
   wire signed [9:0] m43_70;
   assign m43_70 =10'b0;

   // m43_71 = W*in
   wire signed [9:0] m43_71;
   assign m43_71 =10'b0;

   // m43_72 = W*in
   wire signed [9:0] m43_72;
   assign m43_72 ={ {5{in43[5]}} , in43[5:1] };

   // m43_73 = W*in
   wire signed [9:0] m43_73;
   assign m43_73 =10'b0;

   // m43_74 = W*in
   wire signed [9:0] m43_74;
   assign m43_74 =10'b0;

   // m43_75 = W*in
   wire signed [9:0] m43_75;
   assign m43_75 =10'b0;

   // m43_76 = W*in
   wire signed [9:0] m43_76;
   assign m43_76 =10'b0;

   // m43_77 = W*in
   wire signed [9:0] m43_77;
   assign m43_77 =10'b0;

   // m43_78 = W*in
   wire signed [9:0] m43_78;
   assign m43_78 ={ {4{in43[5]}} , in43[5:0] };

   // m43_79 = W*in
   wire signed [9:0] m43_79;
   assign m43_79 =10'b0;

   // m43_80 = W*in
   wire signed [9:0] m43_80;
   assign m43_80 =10'b0;

   // m43_81 = W*in
   wire signed [9:0] m43_81;
   assign m43_81 ={ {5{neg43[5]}} , neg43[5:1] };

   // m43_82 = W*in
   wire signed [9:0] m43_82;
   assign m43_82 =10'b0;

   // m43_83 = W*in
   wire signed [9:0] m43_83;
   assign m43_83 =10'b0;

   // m43_84 = W*in
   wire signed [9:0] m43_84;
   assign m43_84 =10'b0;

   // m43_85 = W*in
   wire signed [9:0] m43_85;
   assign m43_85 =10'b0;

   // m43_86 = W*in
   wire signed [9:0] m43_86;
   assign m43_86 =10'b0;

   // m43_87 = W*in
   wire signed [9:0] m43_87;
   assign m43_87 =10'b0;

   // m43_88 = W*in
   wire signed [9:0] m43_88;
   assign m43_88 =10'b0;

   // m43_89 = W*in
   wire signed [9:0] m43_89;
   assign m43_89 =10'b0;

   // m43_90 = W*in
   wire signed [9:0] m43_90;
   assign m43_90 =10'b0;

   // m43_91 = W*in
   wire signed [9:0] m43_91;
   assign m43_91 =10'b0;

   // m43_92 = W*in
   wire signed [9:0] m43_92;
   assign m43_92 =10'b0;

   // m43_93 = W*in
   wire signed [9:0] m43_93;
   assign m43_93 =10'b0;

   // m43_94 = W*in
   wire signed [9:0] m43_94;
   assign m43_94 =10'b0;

   // m43_95 = W*in
   wire signed [9:0] m43_95;
   assign m43_95 =10'b0;

   // m43_96 = W*in
   wire signed [9:0] m43_96;
   assign m43_96 =10'b0;

   // m43_97 = W*in
   wire signed [9:0] m43_97;
   assign m43_97 =10'b0;

   // m43_98 = W*in
   wire signed [9:0] m43_98;
   assign m43_98 =10'b0;

   // m43_99 = W*in
   wire signed [9:0] m43_99;
   assign m43_99 =10'b0;

   // m43_100 = W*in
   wire signed [9:0] m43_100;
   assign m43_100 =10'b0;

   // m43_101 = W*in
   wire signed [9:0] m43_101;
   assign m43_101 =10'b0;

   // m43_102 = W*in
   wire signed [9:0] m43_102;
   assign m43_102 =10'b0;

   // m43_103 = W*in
   wire signed [9:0] m43_103;
   assign m43_103 =10'b0;

   // m43_104 = W*in
   wire signed [9:0] m43_104;
   assign m43_104 =10'b0;

   // m43_105 = W*in
   wire signed [9:0] m43_105;
   assign m43_105 =10'b0;

   // m43_106 = W*in
   wire signed [9:0] m43_106;
   assign m43_106 =10'b0;

   // m43_107 = W*in
   wire signed [9:0] m43_107;
   assign m43_107 =10'b0;

   // m43_108 = W*in
   wire signed [9:0] m43_108;
   assign m43_108 ={ {5{neg43[5]}} , neg43[5:1] };

   // m43_109 = W*in
   wire signed [9:0] m43_109;
   assign m43_109 =10'b0;

   // m43_110 = W*in
   wire signed [9:0] m43_110;
   assign m43_110 =10'b0;

   // m43_111 = W*in
   wire signed [9:0] m43_111;
   assign m43_111 =10'b0;

   // m43_112 = W*in
   wire signed [9:0] m43_112;
   assign m43_112 =10'b0;

   // m43_113 = W*in
   wire signed [9:0] m43_113;
   assign m43_113 =10'b0;

   // m43_114 = W*in
   wire signed [9:0] m43_114;
   assign m43_114 =10'b0;

   // m43_115 = W*in
   wire signed [9:0] m43_115;
   assign m43_115 =10'b0;

   // m43_116 = W*in
   wire signed [9:0] m43_116;
   assign m43_116 =10'b0;

   // m43_117 = W*in
   wire signed [9:0] m43_117;
   assign m43_117 =10'b0;

   // m44_1 = W*in
   wire signed [9:0] m44_1;
   assign m44_1 =10'b0;

   // m44_2 = W*in
   wire signed [9:0] m44_2;
   assign m44_2 =10'b0;

   // m44_3 = W*in
   wire signed [9:0] m44_3;
   assign m44_3 =10'b0;

   // m44_4 = W*in
   wire signed [9:0] m44_4;
   assign m44_4 =10'b0;

   // m44_5 = W*in
   wire signed [9:0] m44_5;
   assign m44_5 =10'b0;

   // m44_6 = W*in
   wire signed [9:0] m44_6;
   assign m44_6 =10'b0;

   // m44_7 = W*in
   wire signed [9:0] m44_7;
   assign m44_7 =10'b0;

   // m44_8 = W*in
   wire signed [9:0] m44_8;
   assign m44_8 =10'b0;

   // m44_9 = W*in
   wire signed [9:0] m44_9;
   assign m44_9 =10'b0;

   // m44_10 = W*in
   wire signed [9:0] m44_10;
   assign m44_10 =10'b0;

   // m44_11 = W*in
   wire signed [9:0] m44_11;
   assign m44_11 =10'b0;

   // m44_12 = W*in
   wire signed [9:0] m44_12;
   assign m44_12 =10'b0;

   // m44_13 = W*in
   wire signed [9:0] m44_13;
   assign m44_13 =10'b0;

   // m44_14 = W*in
   wire signed [9:0] m44_14;
   assign m44_14 =10'b0;

   // m44_15 = W*in
   wire signed [9:0] m44_15;
   assign m44_15 =10'b0;

   // m44_16 = W*in
   wire signed [9:0] m44_16;
   assign m44_16 =10'b0;

   // m44_17 = W*in
   wire signed [9:0] m44_17;
   assign m44_17 =10'b0;

   // m44_18 = W*in
   wire signed [9:0] m44_18;
   assign m44_18 =10'b0;

   // m44_19 = W*in
   wire signed [9:0] m44_19;
   assign m44_19 ={ {5{in44[5]}} , in44[5:1] };

   // m44_20 = W*in
   wire signed [9:0] m44_20;
   assign m44_20 =10'b0;

   // m44_21 = W*in
   wire signed [9:0] m44_21;
   assign m44_21 =10'b0;

   // m44_22 = W*in
   wire signed [9:0] m44_22;
   assign m44_22 =10'b0;

   // m44_23 = W*in
   wire signed [9:0] m44_23;
   assign m44_23 =10'b0;

   // m44_24 = W*in
   wire signed [9:0] m44_24;
   assign m44_24 =10'b0;

   // m44_25 = W*in
   wire signed [9:0] m44_25;
   assign m44_25 =10'b0;

   // m44_26 = W*in
   wire signed [9:0] m44_26;
   assign m44_26 =10'b0;

   // m44_27 = W*in
   wire signed [9:0] m44_27;
   assign m44_27 =10'b0;

   // m44_28 = W*in
   wire signed [9:0] m44_28;
   assign m44_28 =10'b0;

   // m44_29 = W*in
   wire signed [9:0] m44_29;
   assign m44_29 ={ {5{in44[5]}} , in44[5:1] };

   // m44_30 = W*in
   wire signed [9:0] m44_30;
   assign m44_30 =10'b0;

   // m44_31 = W*in
   wire signed [9:0] m44_31;
   assign m44_31 =10'b0;

   // m44_32 = W*in
   wire signed [9:0] m44_32;
   assign m44_32 =10'b0;

   // m44_33 = W*in
   wire signed [9:0] m44_33;
   assign m44_33 =10'b0;

   // m44_34 = W*in
   wire signed [9:0] m44_34;
   assign m44_34 =10'b0;

   // m44_35 = W*in
   wire signed [9:0] m44_35;
   assign m44_35 ={ {5{neg44[5]}} , neg44[5:1] };

   // m44_36 = W*in
   wire signed [9:0] m44_36;
   assign m44_36 =10'b0;

   // m44_37 = W*in
   wire signed [9:0] m44_37;
   assign m44_37 =10'b0;

   // m44_38 = W*in
   wire signed [9:0] m44_38;
   assign m44_38 =10'b0;

   // m44_39 = W*in
   wire signed [9:0] m44_39;
   assign m44_39 =10'b0;

   // m44_40 = W*in
   wire signed [9:0] m44_40;
   assign m44_40 =10'b0;

   // m44_41 = W*in
   wire signed [9:0] m44_41;
   assign m44_41 =10'b0;

   // m44_42 = W*in
   wire signed [9:0] m44_42;
   assign m44_42 =10'b0;

   // m44_43 = W*in
   wire signed [9:0] m44_43;
   assign m44_43 =10'b0;

   // m44_44 = W*in
   wire signed [9:0] m44_44;
   assign m44_44 =10'b0;

   // m44_45 = W*in
   wire signed [9:0] m44_45;
   assign m44_45 =10'b0;

   // m44_46 = W*in
   wire signed [9:0] m44_46;
   assign m44_46 =10'b0;

   // m44_47 = W*in
   wire signed [9:0] m44_47;
   assign m44_47 =10'b0;

   // m44_48 = W*in
   wire signed [9:0] m44_48;
   assign m44_48 =10'b0;

   // m44_49 = W*in
   wire signed [9:0] m44_49;
   assign m44_49 =10'b0;

   // m44_50 = W*in
   wire signed [9:0] m44_50;
   assign m44_50 =10'b0;

   // m44_51 = W*in
   wire signed [9:0] m44_51;
   assign m44_51 =10'b0;

   // m44_52 = W*in
   wire signed [9:0] m44_52;
   assign m44_52 =10'b0;

   // m44_53 = W*in
   wire signed [9:0] m44_53;
   assign m44_53 =10'b0;

   // m44_54 = W*in
   wire signed [9:0] m44_54;
   assign m44_54 =10'b0;

   // m44_55 = W*in
   wire signed [9:0] m44_55;
   assign m44_55 =10'b0;

   // m44_56 = W*in
   wire signed [9:0] m44_56;
   assign m44_56 =10'b0;

   // m44_57 = W*in
   wire signed [9:0] m44_57;
   assign m44_57 =10'b0;

   // m44_58 = W*in
   wire signed [9:0] m44_58;
   assign m44_58 =10'b0;

   // m44_59 = W*in
   wire signed [9:0] m44_59;
   assign m44_59 =10'b0;

   // m44_60 = W*in
   wire signed [9:0] m44_60;
   assign m44_60 =10'b0;

   // m44_61 = W*in
   wire signed [9:0] m44_61;
   assign m44_61 =10'b0;

   // m44_62 = W*in
   wire signed [9:0] m44_62;
   assign m44_62 =10'b0;

   // m44_63 = W*in
   wire signed [9:0] m44_63;
   assign m44_63 =10'b0;

   // m44_64 = W*in
   wire signed [9:0] m44_64;
   assign m44_64 =10'b0;

   // m44_65 = W*in
   wire signed [9:0] m44_65;
   assign m44_65 =10'b0;

   // m44_66 = W*in
   wire signed [9:0] m44_66;
   assign m44_66 =10'b0;

   // m44_67 = W*in
   wire signed [9:0] m44_67;
   assign m44_67 =10'b0;

   // m44_68 = W*in
   wire signed [9:0] m44_68;
   assign m44_68 =10'b0;

   // m44_69 = W*in
   wire signed [9:0] m44_69;
   assign m44_69 =10'b0;

   // m44_70 = W*in
   wire signed [9:0] m44_70;
   assign m44_70 =10'b0;

   // m44_71 = W*in
   wire signed [9:0] m44_71;
   assign m44_71 =10'b0;

   // m44_72 = W*in
   wire signed [9:0] m44_72;
   assign m44_72 ={ {5{neg44[5]}} , neg44[5:1] };

   // m44_73 = W*in
   wire signed [9:0] m44_73;
   assign m44_73 =10'b0;

   // m44_74 = W*in
   wire signed [9:0] m44_74;
   assign m44_74 =10'b0;

   // m44_75 = W*in
   wire signed [9:0] m44_75;
   assign m44_75 =10'b0;

   // m44_76 = W*in
   wire signed [9:0] m44_76;
   assign m44_76 =10'b0;

   // m44_77 = W*in
   wire signed [9:0] m44_77;
   assign m44_77 =10'b0;

   // m44_78 = W*in
   wire signed [9:0] m44_78;
   assign m44_78 =10'b0;

   // m44_79 = W*in
   wire signed [9:0] m44_79;
   assign m44_79 =10'b0;

   // m44_80 = W*in
   wire signed [9:0] m44_80;
   assign m44_80 =10'b0;

   // m44_81 = W*in
   wire signed [9:0] m44_81;
   assign m44_81 =10'b0;

   // m44_82 = W*in
   wire signed [9:0] m44_82;
   assign m44_82 =10'b0;

   // m44_83 = W*in
   wire signed [9:0] m44_83;
   assign m44_83 =10'b0;

   // m44_84 = W*in
   wire signed [9:0] m44_84;
   assign m44_84 =10'b0;

   // m44_85 = W*in
   wire signed [9:0] m44_85;
   assign m44_85 ={ {5{in44[5]}} , in44[5:1] };

   // m44_86 = W*in
   wire signed [9:0] m44_86;
   assign m44_86 =10'b0;

   // m44_87 = W*in
   wire signed [9:0] m44_87;
   assign m44_87 =10'b0;

   // m44_88 = W*in
   wire signed [9:0] m44_88;
   assign m44_88 =10'b0;

   // m44_89 = W*in
   wire signed [9:0] m44_89;
   assign m44_89 =10'b0;

   // m44_90 = W*in
   wire signed [9:0] m44_90;
   assign m44_90 =10'b0;

   // m44_91 = W*in
   wire signed [9:0] m44_91;
   assign m44_91 =10'b0;

   // m44_92 = W*in
   wire signed [9:0] m44_92;
   assign m44_92 =10'b0;

   // m44_93 = W*in
   wire signed [9:0] m44_93;
   assign m44_93 =10'b0;

   // m44_94 = W*in
   wire signed [9:0] m44_94;
   assign m44_94 =10'b0;

   // m44_95 = W*in
   wire signed [9:0] m44_95;
   assign m44_95 =10'b0;

   // m44_96 = W*in
   wire signed [9:0] m44_96;
   assign m44_96 =10'b0;

   // m44_97 = W*in
   wire signed [9:0] m44_97;
   assign m44_97 =10'b0;

   // m44_98 = W*in
   wire signed [9:0] m44_98;
   assign m44_98 =10'b0;

   // m44_99 = W*in
   wire signed [9:0] m44_99;
   assign m44_99 =10'b0;

   // m44_100 = W*in
   wire signed [9:0] m44_100;
   assign m44_100 =10'b0;

   // m44_101 = W*in
   wire signed [9:0] m44_101;
   assign m44_101 =10'b0;

   // m44_102 = W*in
   wire signed [9:0] m44_102;
   assign m44_102 =10'b0;

   // m44_103 = W*in
   wire signed [9:0] m44_103;
   assign m44_103 =10'b0;

   // m44_104 = W*in
   wire signed [9:0] m44_104;
   assign m44_104 =10'b0;

   // m44_105 = W*in
   wire signed [9:0] m44_105;
   assign m44_105 =10'b0;

   // m44_106 = W*in
   wire signed [9:0] m44_106;
   assign m44_106 =10'b0;

   // m44_107 = W*in
   wire signed [9:0] m44_107;
   assign m44_107 =10'b0;

   // m44_108 = W*in
   wire signed [9:0] m44_108;
   assign m44_108 =10'b0;

   // m44_109 = W*in
   wire signed [9:0] m44_109;
   assign m44_109 =10'b0;

   // m44_110 = W*in
   wire signed [9:0] m44_110;
   assign m44_110 =10'b0;

   // m44_111 = W*in
   wire signed [9:0] m44_111;
   assign m44_111 =10'b0;

   // m44_112 = W*in
   wire signed [9:0] m44_112;
   assign m44_112 =10'b0;

   // m44_113 = W*in
   wire signed [9:0] m44_113;
   assign m44_113 =10'b0;

   // m44_114 = W*in
   wire signed [9:0] m44_114;
   assign m44_114 =10'b0;

   // m44_115 = W*in
   wire signed [9:0] m44_115;
   assign m44_115 =10'b0;

   // m44_116 = W*in
   wire signed [9:0] m44_116;
   assign m44_116 =10'b0;

   // m44_117 = W*in
   wire signed [9:0] m44_117;
   assign m44_117 =10'b0;

   // m45_1 = W*in
   wire signed [9:0] m45_1;
   assign m45_1 =10'b0;

   // m45_2 = W*in
   wire signed [9:0] m45_2;
   assign m45_2 ={ {4{in45[5]}} , in45[5:0] };

   // m45_3 = W*in
   wire signed [9:0] m45_3;
   assign m45_3 =10'b0;

   // m45_4 = W*in
   wire signed [9:0] m45_4;
   assign m45_4 =10'b0;

   // m45_5 = W*in
   wire signed [9:0] m45_5;
   assign m45_5 =10'b0;

   // m45_6 = W*in
   wire signed [9:0] m45_6;
   assign m45_6 =10'b0;

   // m45_7 = W*in
   wire signed [9:0] m45_7;
   assign m45_7 ={ {4{in45[5]}} , in45[5:0] };

   // m45_8 = W*in
   wire signed [9:0] m45_8;
   assign m45_8 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_9 = W*in
   wire signed [9:0] m45_9;
   assign m45_9 =10'b0;

   // m45_10 = W*in
   wire signed [9:0] m45_10;
   assign m45_10 =10'b0;

   // m45_11 = W*in
   wire signed [9:0] m45_11;
   assign m45_11 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_12 = W*in
   wire signed [9:0] m45_12;
   assign m45_12 =10'b0;

   // m45_13 = W*in
   wire signed [9:0] m45_13;
   assign m45_13 =10'b0;

   // m45_14 = W*in
   wire signed [9:0] m45_14;
   assign m45_14 =10'b0;

   // m45_15 = W*in
   wire signed [9:0] m45_15;
   assign m45_15 ={ {4{in45[5]}} , in45[5:0] };

   // m45_16 = W*in
   wire signed [9:0] m45_16;
   assign m45_16 =10'b0;

   // m45_17 = W*in
   wire signed [9:0] m45_17;
   assign m45_17 =10'b0;

   // m45_18 = W*in
   wire signed [9:0] m45_18;
   assign m45_18 =10'b0;

   // m45_19 = W*in
   wire signed [9:0] m45_19;
   assign m45_19 ={ {5{in45[5]}} , in45[5:1] };

   // m45_20 = W*in
   wire signed [9:0] m45_20;
   assign m45_20 ={ {5{in45[5]}} , in45[5:1] };

   // m45_21 = W*in
   wire signed [9:0] m45_21;
   assign m45_21 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_22 = W*in
   wire signed [9:0] m45_22;
   assign m45_22 =10'b0;

   // m45_23 = W*in
   wire signed [9:0] m45_23;
   assign m45_23 =10'b0;

   // m45_24 = W*in
   wire signed [9:0] m45_24;
   assign m45_24 =10'b0;

   // m45_25 = W*in
   wire signed [9:0] m45_25;
   assign m45_25 =10'b0;

   // m45_26 = W*in
   wire signed [9:0] m45_26;
   assign m45_26 =10'b0;

   // m45_27 = W*in
   wire signed [9:0] m45_27;
   assign m45_27 =10'b0;

   // m45_28 = W*in
   wire signed [9:0] m45_28;
   assign m45_28 =10'b0;

   // m45_29 = W*in
   wire signed [9:0] m45_29;
   assign m45_29 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_30 = W*in
   wire signed [9:0] m45_30;
   assign m45_30 =10'b0;

   // m45_31 = W*in
   wire signed [9:0] m45_31;
   assign m45_31 ={ {5{in45[5]}} , in45[5:1] };

   // m45_32 = W*in
   wire signed [9:0] m45_32;
   assign m45_32 =10'b0;

   // m45_33 = W*in
   wire signed [9:0] m45_33;
   assign m45_33 =10'b0;

   // m45_34 = W*in
   wire signed [9:0] m45_34;
   assign m45_34 =10'b0;

   // m45_35 = W*in
   wire signed [9:0] m45_35;
   assign m45_35 =10'b0;

   // m45_36 = W*in
   wire signed [9:0] m45_36;
   assign m45_36 =10'b0;

   // m45_37 = W*in
   wire signed [9:0] m45_37;
   assign m45_37 =10'b0;

   // m45_38 = W*in
   wire signed [9:0] m45_38;
   assign m45_38 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_39 = W*in
   wire signed [9:0] m45_39;
   assign m45_39 =10'b0;

   // m45_40 = W*in
   wire signed [9:0] m45_40;
   assign m45_40 =10'b0;

   // m45_41 = W*in
   wire signed [9:0] m45_41;
   assign m45_41 =10'b0;

   // m45_42 = W*in
   wire signed [9:0] m45_42;
   assign m45_42 =10'b0;

   // m45_43 = W*in
   wire signed [9:0] m45_43;
   assign m45_43 =10'b0;

   // m45_44 = W*in
   wire signed [9:0] m45_44;
   assign m45_44 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_45 = W*in
   wire signed [9:0] m45_45;
   assign m45_45 =10'b0;

   // m45_46 = W*in
   wire signed [9:0] m45_46;
   assign m45_46 =10'b0;

   // m45_47 = W*in
   wire signed [9:0] m45_47;
   assign m45_47 =10'b0;

   // m45_48 = W*in
   wire signed [9:0] m45_48;
   assign m45_48 =10'b0;

   // m45_49 = W*in
   wire signed [9:0] m45_49;
   assign m45_49 =10'b0;

   // m45_50 = W*in
   wire signed [9:0] m45_50;
   assign m45_50 ={ {4{in45[5]}} , in45[5:0] };

   // m45_51 = W*in
   wire signed [9:0] m45_51;
   assign m45_51 ={ {4{in45[5]}} , in45[5:0] };

   // m45_52 = W*in
   wire signed [9:0] m45_52;
   assign m45_52 =10'b0;

   // m45_53 = W*in
   wire signed [9:0] m45_53;
   assign m45_53 =10'b0;

   // m45_54 = W*in
   wire signed [9:0] m45_54;
   assign m45_54 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_55 = W*in
   wire signed [9:0] m45_55;
   assign m45_55 =10'b0;

   // m45_56 = W*in
   wire signed [9:0] m45_56;
   assign m45_56 =10'b0;

   // m45_57 = W*in
   wire signed [9:0] m45_57;
   assign m45_57 =10'b0;

   // m45_58 = W*in
   wire signed [9:0] m45_58;
   assign m45_58 =10'b0;

   // m45_59 = W*in
   wire signed [9:0] m45_59;
   assign m45_59 =10'b0;

   // m45_60 = W*in
   wire signed [9:0] m45_60;
   assign m45_60 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_61 = W*in
   wire signed [9:0] m45_61;
   assign m45_61 =10'b0;

   // m45_62 = W*in
   wire signed [9:0] m45_62;
   assign m45_62 =10'b0;

   // m45_63 = W*in
   wire signed [9:0] m45_63;
   assign m45_63 =10'b0;

   // m45_64 = W*in
   wire signed [9:0] m45_64;
   assign m45_64 =10'b0;

   // m45_65 = W*in
   wire signed [9:0] m45_65;
   assign m45_65 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_66 = W*in
   wire signed [9:0] m45_66;
   assign m45_66 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_67 = W*in
   wire signed [9:0] m45_67;
   assign m45_67 =10'b0;

   // m45_68 = W*in
   wire signed [9:0] m45_68;
   assign m45_68 ={ {3{in45[5]}} , in45 , {1{1'b0}} };

   // m45_69 = W*in
   wire signed [9:0] m45_69;
   assign m45_69 =10'b0;

   // m45_70 = W*in
   wire signed [9:0] m45_70;
   assign m45_70 =10'b0;

   // m45_71 = W*in
   wire signed [9:0] m45_71;
   assign m45_71 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_72 = W*in
   wire signed [9:0] m45_72;
   assign m45_72 =10'b0;

   // m45_73 = W*in
   wire signed [9:0] m45_73;
   assign m45_73 ={ {4{in45[5]}} , in45[5:0] };

   // m45_74 = W*in
   wire signed [9:0] m45_74;
   assign m45_74 =10'b0;

   // m45_75 = W*in
   wire signed [9:0] m45_75;
   assign m45_75 =10'b0;

   // m45_76 = W*in
   wire signed [9:0] m45_76;
   assign m45_76 =10'b0;

   // m45_77 = W*in
   wire signed [9:0] m45_77;
   assign m45_77 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_78 = W*in
   wire signed [9:0] m45_78;
   assign m45_78 =10'b0;

   // m45_79 = W*in
   wire signed [9:0] m45_79;
   assign m45_79 =10'b0;

   // m45_80 = W*in
   wire signed [9:0] m45_80;
   assign m45_80 =10'b0;

   // m45_81 = W*in
   wire signed [9:0] m45_81;
   assign m45_81 =10'b0;

   // m45_82 = W*in
   wire signed [9:0] m45_82;
   assign m45_82 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_83 = W*in
   wire signed [9:0] m45_83;
   assign m45_83 =10'b0;

   // m45_84 = W*in
   wire signed [9:0] m45_84;
   assign m45_84 =10'b0;

   // m45_85 = W*in
   wire signed [9:0] m45_85;
   assign m45_85 =10'b0;

   // m45_86 = W*in
   wire signed [9:0] m45_86;
   assign m45_86 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_87 = W*in
   wire signed [9:0] m45_87;
   assign m45_87 =10'b0;

   // m45_88 = W*in
   wire signed [9:0] m45_88;
   assign m45_88 ={ {4{in45[5]}} , in45[5:0] };

   // m45_89 = W*in
   wire signed [9:0] m45_89;
   assign m45_89 =10'b0;

   // m45_90 = W*in
   wire signed [9:0] m45_90;
   assign m45_90 ={ {4{in45[5]}} , in45[5:0] };

   // m45_91 = W*in
   wire signed [9:0] m45_91;
   assign m45_91 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_92 = W*in
   wire signed [9:0] m45_92;
   assign m45_92 =10'b0;

   // m45_93 = W*in
   wire signed [9:0] m45_93;
   assign m45_93 =10'b0;

   // m45_94 = W*in
   wire signed [9:0] m45_94;
   assign m45_94 =10'b0;

   // m45_95 = W*in
   wire signed [9:0] m45_95;
   assign m45_95 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_96 = W*in
   wire signed [9:0] m45_96;
   assign m45_96 =10'b0;

   // m45_97 = W*in
   wire signed [9:0] m45_97;
   assign m45_97 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_98 = W*in
   wire signed [9:0] m45_98;
   assign m45_98 =10'b0;

   // m45_99 = W*in
   wire signed [9:0] m45_99;
   assign m45_99 =10'b0;

   // m45_100 = W*in
   wire signed [9:0] m45_100;
   assign m45_100 =10'b0;

   // m45_101 = W*in
   wire signed [9:0] m45_101;
   assign m45_101 =10'b0;

   // m45_102 = W*in
   wire signed [9:0] m45_102;
   assign m45_102 =10'b0;

   // m45_103 = W*in
   wire signed [9:0] m45_103;
   assign m45_103 =10'b0;

   // m45_104 = W*in
   wire signed [9:0] m45_104;
   assign m45_104 =10'b0;

   // m45_105 = W*in
   wire signed [9:0] m45_105;
   assign m45_105 ={ {4{in45[5]}} , in45[5:0] };

   // m45_106 = W*in
   wire signed [9:0] m45_106;
   assign m45_106 =10'b0;

   // m45_107 = W*in
   wire signed [9:0] m45_107;
   assign m45_107 ={ {4{in45[5]}} , in45[5:0] };

   // m45_108 = W*in
   wire signed [9:0] m45_108;
   assign m45_108 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_109 = W*in
   wire signed [9:0] m45_109;
   assign m45_109 ={ {5{neg45[5]}} , neg45[5:1] };

   // m45_110 = W*in
   wire signed [9:0] m45_110;
   assign m45_110 ={ {4{neg45[5]}} , neg45[5:0] };

   // m45_111 = W*in
   wire signed [9:0] m45_111;
   assign m45_111 =10'b0;

   // m45_112 = W*in
   wire signed [9:0] m45_112;
   assign m45_112 =10'b0;

   // m45_113 = W*in
   wire signed [9:0] m45_113;
   assign m45_113 ={ {4{in45[5]}} , in45[5:0] };

   // m45_114 = W*in
   wire signed [9:0] m45_114;
   assign m45_114 =10'b0;

   // m45_115 = W*in
   wire signed [9:0] m45_115;
   assign m45_115 =10'b0;

   // m45_116 = W*in
   wire signed [9:0] m45_116;
   assign m45_116 =10'b0;

   // m45_117 = W*in
   wire signed [9:0] m45_117;
   assign m45_117 =10'b0;

   // m46_1 = W*in
   wire signed [9:0] m46_1;
   assign m46_1 =10'b0;

   // m46_2 = W*in
   wire signed [9:0] m46_2;
   assign m46_2 ={ {4{in46[5]}} , in46[5:0] };

   // m46_3 = W*in
   wire signed [9:0] m46_3;
   assign m46_3 =10'b0;

   // m46_4 = W*in
   wire signed [9:0] m46_4;
   assign m46_4 =10'b0;

   // m46_5 = W*in
   wire signed [9:0] m46_5;
   assign m46_5 ={ {4{in46[5]}} , in46[5:0] };

   // m46_6 = W*in
   wire signed [9:0] m46_6;
   assign m46_6 =10'b0;

   // m46_7 = W*in
   wire signed [9:0] m46_7;
   assign m46_7 =10'b0;

   // m46_8 = W*in
   wire signed [9:0] m46_8;
   assign m46_8 =10'b0;

   // m46_9 = W*in
   wire signed [9:0] m46_9;
   assign m46_9 =10'b0;

   // m46_10 = W*in
   wire signed [9:0] m46_10;
   assign m46_10 =10'b0;

   // m46_11 = W*in
   wire signed [9:0] m46_11;
   assign m46_11 =10'b0;

   // m46_12 = W*in
   wire signed [9:0] m46_12;
   assign m46_12 =10'b0;

   // m46_13 = W*in
   wire signed [9:0] m46_13;
   assign m46_13 =10'b0;

   // m46_14 = W*in
   wire signed [9:0] m46_14;
   assign m46_14 =10'b0;

   // m46_15 = W*in
   wire signed [9:0] m46_15;
   assign m46_15 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_16 = W*in
   wire signed [9:0] m46_16;
   assign m46_16 =10'b0;

   // m46_17 = W*in
   wire signed [9:0] m46_17;
   assign m46_17 =10'b0;

   // m46_18 = W*in
   wire signed [9:0] m46_18;
   assign m46_18 ={ {5{in46[5]}} , in46[5:1] };

   // m46_19 = W*in
   wire signed [9:0] m46_19;
   assign m46_19 =10'b0;

   // m46_20 = W*in
   wire signed [9:0] m46_20;
   assign m46_20 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_21 = W*in
   wire signed [9:0] m46_21;
   assign m46_21 =10'b0;

   // m46_22 = W*in
   wire signed [9:0] m46_22;
   assign m46_22 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_23 = W*in
   wire signed [9:0] m46_23;
   assign m46_23 =10'b0;

   // m46_24 = W*in
   wire signed [9:0] m46_24;
   assign m46_24 =10'b0;

   // m46_25 = W*in
   wire signed [9:0] m46_25;
   assign m46_25 =10'b0;

   // m46_26 = W*in
   wire signed [9:0] m46_26;
   assign m46_26 ={ {5{in46[5]}} , in46[5:1] };

   // m46_27 = W*in
   wire signed [9:0] m46_27;
   assign m46_27 =10'b0;

   // m46_28 = W*in
   wire signed [9:0] m46_28;
   assign m46_28 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_29 = W*in
   wire signed [9:0] m46_29;
   assign m46_29 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_30 = W*in
   wire signed [9:0] m46_30;
   assign m46_30 =10'b0;

   // m46_31 = W*in
   wire signed [9:0] m46_31;
   assign m46_31 ={ {5{in46[5]}} , in46[5:1] };

   // m46_32 = W*in
   wire signed [9:0] m46_32;
   assign m46_32 =10'b0;

   // m46_33 = W*in
   wire signed [9:0] m46_33;
   assign m46_33 =10'b0;

   // m46_34 = W*in
   wire signed [9:0] m46_34;
   assign m46_34 =10'b0;

   // m46_35 = W*in
   wire signed [9:0] m46_35;
   assign m46_35 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_36 = W*in
   wire signed [9:0] m46_36;
   assign m46_36 =10'b0;

   // m46_37 = W*in
   wire signed [9:0] m46_37;
   assign m46_37 =10'b0;

   // m46_38 = W*in
   wire signed [9:0] m46_38;
   assign m46_38 =10'b0;

   // m46_39 = W*in
   wire signed [9:0] m46_39;
   assign m46_39 =10'b0;

   // m46_40 = W*in
   wire signed [9:0] m46_40;
   assign m46_40 =10'b0;

   // m46_41 = W*in
   wire signed [9:0] m46_41;
   assign m46_41 =10'b0;

   // m46_42 = W*in
   wire signed [9:0] m46_42;
   assign m46_42 =10'b0;

   // m46_43 = W*in
   wire signed [9:0] m46_43;
   assign m46_43 =10'b0;

   // m46_44 = W*in
   wire signed [9:0] m46_44;
   assign m46_44 =10'b0;

   // m46_45 = W*in
   wire signed [9:0] m46_45;
   assign m46_45 =10'b0;

   // m46_46 = W*in
   wire signed [9:0] m46_46;
   assign m46_46 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_47 = W*in
   wire signed [9:0] m46_47;
   assign m46_47 =10'b0;

   // m46_48 = W*in
   wire signed [9:0] m46_48;
   assign m46_48 ={ {4{in46[5]}} , in46[5:0] };

   // m46_49 = W*in
   wire signed [9:0] m46_49;
   assign m46_49 =10'b0;

   // m46_50 = W*in
   wire signed [9:0] m46_50;
   assign m46_50 ={ {4{in46[5]}} , in46[5:0] };

   // m46_51 = W*in
   wire signed [9:0] m46_51;
   assign m46_51 ={ {4{in46[5]}} , in46[5:0] };

   // m46_52 = W*in
   wire signed [9:0] m46_52;
   assign m46_52 =10'b0;

   // m46_53 = W*in
   wire signed [9:0] m46_53;
   assign m46_53 =10'b0;

   // m46_54 = W*in
   wire signed [9:0] m46_54;
   assign m46_54 =10'b0;

   // m46_55 = W*in
   wire signed [9:0] m46_55;
   assign m46_55 =10'b0;

   // m46_56 = W*in
   wire signed [9:0] m46_56;
   assign m46_56 =10'b0;

   // m46_57 = W*in
   wire signed [9:0] m46_57;
   assign m46_57 =10'b0;

   // m46_58 = W*in
   wire signed [9:0] m46_58;
   assign m46_58 =10'b0;

   // m46_59 = W*in
   wire signed [9:0] m46_59;
   assign m46_59 =10'b0;

   // m46_60 = W*in
   wire signed [9:0] m46_60;
   assign m46_60 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_61 = W*in
   wire signed [9:0] m46_61;
   assign m46_61 =10'b0;

   // m46_62 = W*in
   wire signed [9:0] m46_62;
   assign m46_62 =10'b0;

   // m46_63 = W*in
   wire signed [9:0] m46_63;
   assign m46_63 =10'b0;

   // m46_64 = W*in
   wire signed [9:0] m46_64;
   assign m46_64 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_65 = W*in
   wire signed [9:0] m46_65;
   assign m46_65 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_66 = W*in
   wire signed [9:0] m46_66;
   assign m46_66 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_67 = W*in
   wire signed [9:0] m46_67;
   assign m46_67 =10'b0;

   // m46_68 = W*in
   wire signed [9:0] m46_68;
   assign m46_68 ={ {4{in46[5]}} , in46[5:0] };

   // m46_69 = W*in
   wire signed [9:0] m46_69;
   assign m46_69 ={ {5{in46[5]}} , in46[5:1] };

   // m46_70 = W*in
   wire signed [9:0] m46_70;
   assign m46_70 ={ {5{in46[5]}} , in46[5:1] };

   // m46_71 = W*in
   wire signed [9:0] m46_71;
   assign m46_71 =10'b0;

   // m46_72 = W*in
   wire signed [9:0] m46_72;
   assign m46_72 ={ {5{in46[5]}} , in46[5:1] };

   // m46_73 = W*in
   wire signed [9:0] m46_73;
   assign m46_73 =10'b0;

   // m46_74 = W*in
   wire signed [9:0] m46_74;
   assign m46_74 =10'b0;

   // m46_75 = W*in
   wire signed [9:0] m46_75;
   assign m46_75 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_76 = W*in
   wire signed [9:0] m46_76;
   assign m46_76 ={ {4{in46[5]}} , in46[5:0] };

   // m46_77 = W*in
   wire signed [9:0] m46_77;
   assign m46_77 =10'b0;

   // m46_78 = W*in
   wire signed [9:0] m46_78;
   assign m46_78 =10'b0;

   // m46_79 = W*in
   wire signed [9:0] m46_79;
   assign m46_79 =10'b0;

   // m46_80 = W*in
   wire signed [9:0] m46_80;
   assign m46_80 =10'b0;

   // m46_81 = W*in
   wire signed [9:0] m46_81;
   assign m46_81 ={ {5{neg46[5]}} , neg46[5:1] };

   // m46_82 = W*in
   wire signed [9:0] m46_82;
   assign m46_82 ={ {5{in46[5]}} , in46[5:1] };

   // m46_83 = W*in
   wire signed [9:0] m46_83;
   assign m46_83 =10'b0;

   // m46_84 = W*in
   wire signed [9:0] m46_84;
   assign m46_84 =10'b0;

   // m46_85 = W*in
   wire signed [9:0] m46_85;
   assign m46_85 =10'b0;

   // m46_86 = W*in
   wire signed [9:0] m46_86;
   assign m46_86 =10'b0;

   // m46_87 = W*in
   wire signed [9:0] m46_87;
   assign m46_87 =10'b0;

   // m46_88 = W*in
   wire signed [9:0] m46_88;
   assign m46_88 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_89 = W*in
   wire signed [9:0] m46_89;
   assign m46_89 =10'b0;

   // m46_90 = W*in
   wire signed [9:0] m46_90;
   assign m46_90 =10'b0;

   // m46_91 = W*in
   wire signed [9:0] m46_91;
   assign m46_91 =10'b0;

   // m46_92 = W*in
   wire signed [9:0] m46_92;
   assign m46_92 ={ {3{in46[5]}} , in46 , {1{1'b0}} };

   // m46_93 = W*in
   wire signed [9:0] m46_93;
   assign m46_93 =10'b0;

   // m46_94 = W*in
   wire signed [9:0] m46_94;
   assign m46_94 =10'b0;

   // m46_95 = W*in
   wire signed [9:0] m46_95;
   assign m46_95 =10'b0;

   // m46_96 = W*in
   wire signed [9:0] m46_96;
   assign m46_96 =10'b0;

   // m46_97 = W*in
   wire signed [9:0] m46_97;
   assign m46_97 =10'b0;

   // m46_98 = W*in
   wire signed [9:0] m46_98;
   assign m46_98 =10'b0;

   // m46_99 = W*in
   wire signed [9:0] m46_99;
   assign m46_99 =10'b0;

   // m46_100 = W*in
   wire signed [9:0] m46_100;
   assign m46_100 =10'b0;

   // m46_101 = W*in
   wire signed [9:0] m46_101;
   assign m46_101 =10'b0;

   // m46_102 = W*in
   wire signed [9:0] m46_102;
   assign m46_102 =10'b0;

   // m46_103 = W*in
   wire signed [9:0] m46_103;
   assign m46_103 =10'b0;

   // m46_104 = W*in
   wire signed [9:0] m46_104;
   assign m46_104 =10'b0;

   // m46_105 = W*in
   wire signed [9:0] m46_105;
   assign m46_105 =10'b0;

   // m46_106 = W*in
   wire signed [9:0] m46_106;
   assign m46_106 =10'b0;

   // m46_107 = W*in
   wire signed [9:0] m46_107;
   assign m46_107 =10'b0;

   // m46_108 = W*in
   wire signed [9:0] m46_108;
   assign m46_108 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_109 = W*in
   wire signed [9:0] m46_109;
   assign m46_109 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_110 = W*in
   wire signed [9:0] m46_110;
   assign m46_110 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_111 = W*in
   wire signed [9:0] m46_111;
   assign m46_111 =10'b0;

   // m46_112 = W*in
   wire signed [9:0] m46_112;
   assign m46_112 =10'b0;

   // m46_113 = W*in
   wire signed [9:0] m46_113;
   assign m46_113 =10'b0;

   // m46_114 = W*in
   wire signed [9:0] m46_114;
   assign m46_114 ={ {4{neg46[5]}} , neg46[5:0] };

   // m46_115 = W*in
   wire signed [9:0] m46_115;
   assign m46_115 =10'b0;

   // m46_116 = W*in
   wire signed [9:0] m46_116;
   assign m46_116 =10'b0;

   // m46_117 = W*in
   wire signed [9:0] m46_117;
   assign m46_117 ={ {4{neg46[5]}} , neg46[5:0] };

   // m47_1 = W*in
   wire signed [9:0] m47_1;
   assign m47_1 ={ {4{in47[5]}} , in47[5:0] };

   // m47_2 = W*in
   wire signed [9:0] m47_2;
   assign m47_2 =10'b0;

   // m47_3 = W*in
   wire signed [9:0] m47_3;
   assign m47_3 =10'b0;

   // m47_4 = W*in
   wire signed [9:0] m47_4;
   assign m47_4 =10'b0;

   // m47_5 = W*in
   wire signed [9:0] m47_5;
   assign m47_5 =10'b0;

   // m47_6 = W*in
   wire signed [9:0] m47_6;
   assign m47_6 =10'b0;

   // m47_7 = W*in
   wire signed [9:0] m47_7;
   assign m47_7 =10'b0;

   // m47_8 = W*in
   wire signed [9:0] m47_8;
   assign m47_8 =10'b0;

   // m47_9 = W*in
   wire signed [9:0] m47_9;
   assign m47_9 =10'b0;

   // m47_10 = W*in
   wire signed [9:0] m47_10;
   assign m47_10 =10'b0;

   // m47_11 = W*in
   wire signed [9:0] m47_11;
   assign m47_11 =10'b0;

   // m47_12 = W*in
   wire signed [9:0] m47_12;
   assign m47_12 =10'b0;

   // m47_13 = W*in
   wire signed [9:0] m47_13;
   assign m47_13 =10'b0;

   // m47_14 = W*in
   wire signed [9:0] m47_14;
   assign m47_14 =10'b0;

   // m47_15 = W*in
   wire signed [9:0] m47_15;
   assign m47_15 =10'b0;

   // m47_16 = W*in
   wire signed [9:0] m47_16;
   assign m47_16 =10'b0;

   // m47_17 = W*in
   wire signed [9:0] m47_17;
   assign m47_17 =10'b0;

   // m47_18 = W*in
   wire signed [9:0] m47_18;
   assign m47_18 ={ {5{neg47[5]}} , neg47[5:1] };

   // m47_19 = W*in
   wire signed [9:0] m47_19;
   assign m47_19 =10'b0;

   // m47_20 = W*in
   wire signed [9:0] m47_20;
   assign m47_20 =10'b0;

   // m47_21 = W*in
   wire signed [9:0] m47_21;
   assign m47_21 =10'b0;

   // m47_22 = W*in
   wire signed [9:0] m47_22;
   assign m47_22 =10'b0;

   // m47_23 = W*in
   wire signed [9:0] m47_23;
   assign m47_23 =10'b0;

   // m47_24 = W*in
   wire signed [9:0] m47_24;
   assign m47_24 =10'b0;

   // m47_25 = W*in
   wire signed [9:0] m47_25;
   assign m47_25 =10'b0;

   // m47_26 = W*in
   wire signed [9:0] m47_26;
   assign m47_26 ={ {5{neg47[5]}} , neg47[5:1] };

   // m47_27 = W*in
   wire signed [9:0] m47_27;
   assign m47_27 =10'b0;

   // m47_28 = W*in
   wire signed [9:0] m47_28;
   assign m47_28 ={ {5{in47[5]}} , in47[5:1] };

   // m47_29 = W*in
   wire signed [9:0] m47_29;
   assign m47_29 =10'b0;

   // m47_30 = W*in
   wire signed [9:0] m47_30;
   assign m47_30 =10'b0;

   // m47_31 = W*in
   wire signed [9:0] m47_31;
   assign m47_31 ={ {5{in47[5]}} , in47[5:1] };

   // m47_32 = W*in
   wire signed [9:0] m47_32;
   assign m47_32 =10'b0;

   // m47_33 = W*in
   wire signed [9:0] m47_33;
   assign m47_33 =10'b0;

   // m47_34 = W*in
   wire signed [9:0] m47_34;
   assign m47_34 =10'b0;

   // m47_35 = W*in
   wire signed [9:0] m47_35;
   assign m47_35 =10'b0;

   // m47_36 = W*in
   wire signed [9:0] m47_36;
   assign m47_36 ={ {5{in47[5]}} , in47[5:1] };

   // m47_37 = W*in
   wire signed [9:0] m47_37;
   assign m47_37 =10'b0;

   // m47_38 = W*in
   wire signed [9:0] m47_38;
   assign m47_38 ={ {4{neg47[5]}} , neg47[5:0] };

   // m47_39 = W*in
   wire signed [9:0] m47_39;
   assign m47_39 =10'b0;

   // m47_40 = W*in
   wire signed [9:0] m47_40;
   assign m47_40 =10'b0;

   // m47_41 = W*in
   wire signed [9:0] m47_41;
   assign m47_41 =10'b0;

   // m47_42 = W*in
   wire signed [9:0] m47_42;
   assign m47_42 =10'b0;

   // m47_43 = W*in
   wire signed [9:0] m47_43;
   assign m47_43 =10'b0;

   // m47_44 = W*in
   wire signed [9:0] m47_44;
   assign m47_44 =10'b0;

   // m47_45 = W*in
   wire signed [9:0] m47_45;
   assign m47_45 ={ {4{in47[5]}} , in47[5:0] };

   // m47_46 = W*in
   wire signed [9:0] m47_46;
   assign m47_46 =10'b0;

   // m47_47 = W*in
   wire signed [9:0] m47_47;
   assign m47_47 =10'b0;

   // m47_48 = W*in
   wire signed [9:0] m47_48;
   assign m47_48 =10'b0;

   // m47_49 = W*in
   wire signed [9:0] m47_49;
   assign m47_49 =10'b0;

   // m47_50 = W*in
   wire signed [9:0] m47_50;
   assign m47_50 =10'b0;

   // m47_51 = W*in
   wire signed [9:0] m47_51;
   assign m47_51 ={ {4{in47[5]}} , in47[5:0] };

   // m47_52 = W*in
   wire signed [9:0] m47_52;
   assign m47_52 =10'b0;

   // m47_53 = W*in
   wire signed [9:0] m47_53;
   assign m47_53 =10'b0;

   // m47_54 = W*in
   wire signed [9:0] m47_54;
   assign m47_54 =10'b0;

   // m47_55 = W*in
   wire signed [9:0] m47_55;
   assign m47_55 =10'b0;

   // m47_56 = W*in
   wire signed [9:0] m47_56;
   assign m47_56 =10'b0;

   // m47_57 = W*in
   wire signed [9:0] m47_57;
   assign m47_57 =10'b0;

   // m47_58 = W*in
   wire signed [9:0] m47_58;
   assign m47_58 =10'b0;

   // m47_59 = W*in
   wire signed [9:0] m47_59;
   assign m47_59 =10'b0;

   // m47_60 = W*in
   wire signed [9:0] m47_60;
   assign m47_60 =10'b0;

   // m47_61 = W*in
   wire signed [9:0] m47_61;
   assign m47_61 =10'b0;

   // m47_62 = W*in
   wire signed [9:0] m47_62;
   assign m47_62 =10'b0;

   // m47_63 = W*in
   wire signed [9:0] m47_63;
   assign m47_63 =10'b0;

   // m47_64 = W*in
   wire signed [9:0] m47_64;
   assign m47_64 =10'b0;

   // m47_65 = W*in
   wire signed [9:0] m47_65;
   assign m47_65 =10'b0;

   // m47_66 = W*in
   wire signed [9:0] m47_66;
   assign m47_66 =10'b0;

   // m47_67 = W*in
   wire signed [9:0] m47_67;
   assign m47_67 =10'b0;

   // m47_68 = W*in
   wire signed [9:0] m47_68;
   assign m47_68 =10'b0;

   // m47_69 = W*in
   wire signed [9:0] m47_69;
   assign m47_69 ={ {5{neg47[5]}} , neg47[5:1] };

   // m47_70 = W*in
   wire signed [9:0] m47_70;
   assign m47_70 ={ {5{neg47[5]}} , neg47[5:1] };

   // m47_71 = W*in
   wire signed [9:0] m47_71;
   assign m47_71 ={ {5{neg47[5]}} , neg47[5:1] };

   // m47_72 = W*in
   wire signed [9:0] m47_72;
   assign m47_72 ={ {4{neg47[5]}} , neg47[5:0] };

   // m47_73 = W*in
   wire signed [9:0] m47_73;
   assign m47_73 ={ {5{in47[5]}} , in47[5:1] };

   // m47_74 = W*in
   wire signed [9:0] m47_74;
   assign m47_74 ={ {4{neg47[5]}} , neg47[5:0] };

   // m47_75 = W*in
   wire signed [9:0] m47_75;
   assign m47_75 =10'b0;

   // m47_76 = W*in
   wire signed [9:0] m47_76;
   assign m47_76 =10'b0;

   // m47_77 = W*in
   wire signed [9:0] m47_77;
   assign m47_77 =10'b0;

   // m47_78 = W*in
   wire signed [9:0] m47_78;
   assign m47_78 =10'b0;

   // m47_79 = W*in
   wire signed [9:0] m47_79;
   assign m47_79 =10'b0;

   // m47_80 = W*in
   wire signed [9:0] m47_80;
   assign m47_80 =10'b0;

   // m47_81 = W*in
   wire signed [9:0] m47_81;
   assign m47_81 =10'b0;

   // m47_82 = W*in
   wire signed [9:0] m47_82;
   assign m47_82 =10'b0;

   // m47_83 = W*in
   wire signed [9:0] m47_83;
   assign m47_83 =10'b0;

   // m47_84 = W*in
   wire signed [9:0] m47_84;
   assign m47_84 =10'b0;

   // m47_85 = W*in
   wire signed [9:0] m47_85;
   assign m47_85 =10'b0;

   // m47_86 = W*in
   wire signed [9:0] m47_86;
   assign m47_86 =10'b0;

   // m47_87 = W*in
   wire signed [9:0] m47_87;
   assign m47_87 =10'b0;

   // m47_88 = W*in
   wire signed [9:0] m47_88;
   assign m47_88 =10'b0;

   // m47_89 = W*in
   wire signed [9:0] m47_89;
   assign m47_89 =10'b0;

   // m47_90 = W*in
   wire signed [9:0] m47_90;
   assign m47_90 =10'b0;

   // m47_91 = W*in
   wire signed [9:0] m47_91;
   assign m47_91 =10'b0;

   // m47_92 = W*in
   wire signed [9:0] m47_92;
   assign m47_92 =10'b0;

   // m47_93 = W*in
   wire signed [9:0] m47_93;
   assign m47_93 =10'b0;

   // m47_94 = W*in
   wire signed [9:0] m47_94;
   assign m47_94 =10'b0;

   // m47_95 = W*in
   wire signed [9:0] m47_95;
   assign m47_95 =10'b0;

   // m47_96 = W*in
   wire signed [9:0] m47_96;
   assign m47_96 =10'b0;

   // m47_97 = W*in
   wire signed [9:0] m47_97;
   assign m47_97 =10'b0;

   // m47_98 = W*in
   wire signed [9:0] m47_98;
   assign m47_98 =10'b0;

   // m47_99 = W*in
   wire signed [9:0] m47_99;
   assign m47_99 ={ {4{neg47[5]}} , neg47[5:0] };

   // m47_100 = W*in
   wire signed [9:0] m47_100;
   assign m47_100 =10'b0;

   // m47_101 = W*in
   wire signed [9:0] m47_101;
   assign m47_101 =10'b0;

   // m47_102 = W*in
   wire signed [9:0] m47_102;
   assign m47_102 ={ {4{in47[5]}} , in47[5:0] };

   // m47_103 = W*in
   wire signed [9:0] m47_103;
   assign m47_103 =10'b0;

   // m47_104 = W*in
   wire signed [9:0] m47_104;
   assign m47_104 =10'b0;

   // m47_105 = W*in
   wire signed [9:0] m47_105;
   assign m47_105 =10'b0;

   // m47_106 = W*in
   wire signed [9:0] m47_106;
   assign m47_106 =10'b0;

   // m47_107 = W*in
   wire signed [9:0] m47_107;
   assign m47_107 =10'b0;

   // m47_108 = W*in
   wire signed [9:0] m47_108;
   assign m47_108 =10'b0;

   // m47_109 = W*in
   wire signed [9:0] m47_109;
   assign m47_109 =10'b0;

   // m47_110 = W*in
   wire signed [9:0] m47_110;
   assign m47_110 =10'b0;

   // m47_111 = W*in
   wire signed [9:0] m47_111;
   assign m47_111 =10'b0;

   // m47_112 = W*in
   wire signed [9:0] m47_112;
   assign m47_112 =10'b0;

   // m47_113 = W*in
   wire signed [9:0] m47_113;
   assign m47_113 =10'b0;

   // m47_114 = W*in
   wire signed [9:0] m47_114;
   assign m47_114 =10'b0;

   // m47_115 = W*in
   wire signed [9:0] m47_115;
   assign m47_115 =10'b0;

   // m47_116 = W*in
   wire signed [9:0] m47_116;
   assign m47_116 =10'b0;

   // m47_117 = W*in
   wire signed [9:0] m47_117;
   assign m47_117 =10'b0;

   // m48_1 = W*in
   wire signed [9:0] m48_1;
   assign m48_1 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_2 = W*in
   wire signed [9:0] m48_2;
   assign m48_2 ={ {4{in48[5]}} , in48[5:0] };

   // m48_3 = W*in
   wire signed [9:0] m48_3;
   assign m48_3 ={ {4{in48[5]}} , in48[5:0] };

   // m48_4 = W*in
   wire signed [9:0] m48_4;
   assign m48_4 =10'b0;

   // m48_5 = W*in
   wire signed [9:0] m48_5;
   assign m48_5 =10'b0;

   // m48_6 = W*in
   wire signed [9:0] m48_6;
   assign m48_6 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_7 = W*in
   wire signed [9:0] m48_7;
   assign m48_7 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_8 = W*in
   wire signed [9:0] m48_8;
   assign m48_8 =10'b0;

   // m48_9 = W*in
   wire signed [9:0] m48_9;
   assign m48_9 =10'b0;

   // m48_10 = W*in
   wire signed [9:0] m48_10;
   assign m48_10 =10'b0;

   // m48_11 = W*in
   wire signed [9:0] m48_11;
   assign m48_11 =10'b0;

   // m48_12 = W*in
   wire signed [9:0] m48_12;
   assign m48_12 =10'b0;

   // m48_13 = W*in
   wire signed [9:0] m48_13;
   assign m48_13 ={ {4{in48[5]}} , in48[5:0] };

   // m48_14 = W*in
   wire signed [9:0] m48_14;
   assign m48_14 =10'b0;

   // m48_15 = W*in
   wire signed [9:0] m48_15;
   assign m48_15 =10'b0;

   // m48_16 = W*in
   wire signed [9:0] m48_16;
   assign m48_16 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_17 = W*in
   wire signed [9:0] m48_17;
   assign m48_17 =10'b0;

   // m48_18 = W*in
   wire signed [9:0] m48_18;
   assign m48_18 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_19 = W*in
   wire signed [9:0] m48_19;
   assign m48_19 ={ {5{neg48[5]}} , neg48[5:1] };

   // m48_20 = W*in
   wire signed [9:0] m48_20;
   assign m48_20 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_21 = W*in
   wire signed [9:0] m48_21;
   assign m48_21 =10'b0;

   // m48_22 = W*in
   wire signed [9:0] m48_22;
   assign m48_22 =10'b0;

   // m48_23 = W*in
   wire signed [9:0] m48_23;
   assign m48_23 ={ {4{in48[5]}} , in48[5:0] };

   // m48_24 = W*in
   wire signed [9:0] m48_24;
   assign m48_24 =10'b0;

   // m48_25 = W*in
   wire signed [9:0] m48_25;
   assign m48_25 ={ {4{in48[5]}} , in48[5:0] };

   // m48_26 = W*in
   wire signed [9:0] m48_26;
   assign m48_26 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_27 = W*in
   wire signed [9:0] m48_27;
   assign m48_27 ={ {5{in48[5]}} , in48[5:1] };

   // m48_28 = W*in
   wire signed [9:0] m48_28;
   assign m48_28 ={ {4{in48[5]}} , in48[5:0] };

   // m48_29 = W*in
   wire signed [9:0] m48_29;
   assign m48_29 ={ {5{in48[5]}} , in48[5:1] };

   // m48_30 = W*in
   wire signed [9:0] m48_30;
   assign m48_30 ={ {5{neg48[5]}} , neg48[5:1] };

   // m48_31 = W*in
   wire signed [9:0] m48_31;
   assign m48_31 ={ {4{in48[5]}} , in48[5:0] };

   // m48_32 = W*in
   wire signed [9:0] m48_32;
   assign m48_32 =10'b0;

   // m48_33 = W*in
   wire signed [9:0] m48_33;
   assign m48_33 ={ {4{in48[5]}} , in48[5:0] };

   // m48_34 = W*in
   wire signed [9:0] m48_34;
   assign m48_34 =10'b0;

   // m48_35 = W*in
   wire signed [9:0] m48_35;
   assign m48_35 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_36 = W*in
   wire signed [9:0] m48_36;
   assign m48_36 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_37 = W*in
   wire signed [9:0] m48_37;
   assign m48_37 =10'b0;

   // m48_38 = W*in
   wire signed [9:0] m48_38;
   assign m48_38 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_39 = W*in
   wire signed [9:0] m48_39;
   assign m48_39 =10'b0;

   // m48_40 = W*in
   wire signed [9:0] m48_40;
   assign m48_40 =10'b0;

   // m48_41 = W*in
   wire signed [9:0] m48_41;
   assign m48_41 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_42 = W*in
   wire signed [9:0] m48_42;
   assign m48_42 =10'b0;

   // m48_43 = W*in
   wire signed [9:0] m48_43;
   assign m48_43 ={ {4{in48[5]}} , in48[5:0] };

   // m48_44 = W*in
   wire signed [9:0] m48_44;
   assign m48_44 =10'b0;

   // m48_45 = W*in
   wire signed [9:0] m48_45;
   assign m48_45 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_46 = W*in
   wire signed [9:0] m48_46;
   assign m48_46 =10'b0;

   // m48_47 = W*in
   wire signed [9:0] m48_47;
   assign m48_47 =10'b0;

   // m48_48 = W*in
   wire signed [9:0] m48_48;
   assign m48_48 =10'b0;

   // m48_49 = W*in
   wire signed [9:0] m48_49;
   assign m48_49 =10'b0;

   // m48_50 = W*in
   wire signed [9:0] m48_50;
   assign m48_50 =10'b0;

   // m48_51 = W*in
   wire signed [9:0] m48_51;
   assign m48_51 ={ {4{in48[5]}} , in48[5:0] };

   // m48_52 = W*in
   wire signed [9:0] m48_52;
   assign m48_52 =10'b0;

   // m48_53 = W*in
   wire signed [9:0] m48_53;
   assign m48_53 ={ {4{in48[5]}} , in48[5:0] };

   // m48_54 = W*in
   wire signed [9:0] m48_54;
   assign m48_54 =10'b0;

   // m48_55 = W*in
   wire signed [9:0] m48_55;
   assign m48_55 =10'b0;

   // m48_56 = W*in
   wire signed [9:0] m48_56;
   assign m48_56 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_57 = W*in
   wire signed [9:0] m48_57;
   assign m48_57 =10'b0;

   // m48_58 = W*in
   wire signed [9:0] m48_58;
   assign m48_58 =10'b0;

   // m48_59 = W*in
   wire signed [9:0] m48_59;
   assign m48_59 ={ {4{in48[5]}} , in48[5:0] };

   // m48_60 = W*in
   wire signed [9:0] m48_60;
   assign m48_60 =10'b0;

   // m48_61 = W*in
   wire signed [9:0] m48_61;
   assign m48_61 =10'b0;

   // m48_62 = W*in
   wire signed [9:0] m48_62;
   assign m48_62 =10'b0;

   // m48_63 = W*in
   wire signed [9:0] m48_63;
   assign m48_63 =10'b0;

   // m48_64 = W*in
   wire signed [9:0] m48_64;
   assign m48_64 ={ {5{neg48[5]}} , neg48[5:1] };

   // m48_65 = W*in
   wire signed [9:0] m48_65;
   assign m48_65 =10'b0;

   // m48_66 = W*in
   wire signed [9:0] m48_66;
   assign m48_66 =10'b0;

   // m48_67 = W*in
   wire signed [9:0] m48_67;
   assign m48_67 =10'b0;

   // m48_68 = W*in
   wire signed [9:0] m48_68;
   assign m48_68 =10'b0;

   // m48_69 = W*in
   wire signed [9:0] m48_69;
   assign m48_69 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_70 = W*in
   wire signed [9:0] m48_70;
   assign m48_70 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_71 = W*in
   wire signed [9:0] m48_71;
   assign m48_71 ={ {5{neg48[5]}} , neg48[5:1] };

   // m48_72 = W*in
   wire signed [9:0] m48_72;
   assign m48_72 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_73 = W*in
   wire signed [9:0] m48_73;
   assign m48_73 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_74 = W*in
   wire signed [9:0] m48_74;
   assign m48_74 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_75 = W*in
   wire signed [9:0] m48_75;
   assign m48_75 ={ {5{neg48[5]}} , neg48[5:1] };

   // m48_76 = W*in
   wire signed [9:0] m48_76;
   assign m48_76 =10'b0;

   // m48_77 = W*in
   wire signed [9:0] m48_77;
   assign m48_77 ={ {4{in48[5]}} , in48[5:0] };

   // m48_78 = W*in
   wire signed [9:0] m48_78;
   assign m48_78 =10'b0;

   // m48_79 = W*in
   wire signed [9:0] m48_79;
   assign m48_79 =10'b0;

   // m48_80 = W*in
   wire signed [9:0] m48_80;
   assign m48_80 =10'b0;

   // m48_81 = W*in
   wire signed [9:0] m48_81;
   assign m48_81 =10'b0;

   // m48_82 = W*in
   wire signed [9:0] m48_82;
   assign m48_82 =10'b0;

   // m48_83 = W*in
   wire signed [9:0] m48_83;
   assign m48_83 =10'b0;

   // m48_84 = W*in
   wire signed [9:0] m48_84;
   assign m48_84 =10'b0;

   // m48_85 = W*in
   wire signed [9:0] m48_85;
   assign m48_85 =10'b0;

   // m48_86 = W*in
   wire signed [9:0] m48_86;
   assign m48_86 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_87 = W*in
   wire signed [9:0] m48_87;
   assign m48_87 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_88 = W*in
   wire signed [9:0] m48_88;
   assign m48_88 =10'b0;

   // m48_89 = W*in
   wire signed [9:0] m48_89;
   assign m48_89 =10'b0;

   // m48_90 = W*in
   wire signed [9:0] m48_90;
   assign m48_90 =10'b0;

   // m48_91 = W*in
   wire signed [9:0] m48_91;
   assign m48_91 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_92 = W*in
   wire signed [9:0] m48_92;
   assign m48_92 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_93 = W*in
   wire signed [9:0] m48_93;
   assign m48_93 =10'b0;

   // m48_94 = W*in
   wire signed [9:0] m48_94;
   assign m48_94 ={ {5{neg48[5]}} , neg48[5:1] };

   // m48_95 = W*in
   wire signed [9:0] m48_95;
   assign m48_95 ={ {4{in48[5]}} , in48[5:0] };

   // m48_96 = W*in
   wire signed [9:0] m48_96;
   assign m48_96 =10'b0;

   // m48_97 = W*in
   wire signed [9:0] m48_97;
   assign m48_97 =10'b0;

   // m48_98 = W*in
   wire signed [9:0] m48_98;
   assign m48_98 ={ {3{in48[5]}} , in48 , {1{1'b0}} };

   // m48_99 = W*in
   wire signed [9:0] m48_99;
   assign m48_99 ={ {3{neg48[5]}} , neg48 , {1{1'b0}} };

   // m48_100 = W*in
   wire signed [9:0] m48_100;
   assign m48_100 =10'b0;

   // m48_101 = W*in
   wire signed [9:0] m48_101;
   assign m48_101 =10'b0;

   // m48_102 = W*in
   wire signed [9:0] m48_102;
   assign m48_102 ={ {4{in48[5]}} , in48[5:0] };

   // m48_103 = W*in
   wire signed [9:0] m48_103;
   assign m48_103 =10'b0;

   // m48_104 = W*in
   wire signed [9:0] m48_104;
   assign m48_104 =10'b0;

   // m48_105 = W*in
   wire signed [9:0] m48_105;
   assign m48_105 ={ {4{in48[5]}} , in48[5:0] };

   // m48_106 = W*in
   wire signed [9:0] m48_106;
   assign m48_106 ={ {4{in48[5]}} , in48[5:0] };

   // m48_107 = W*in
   wire signed [9:0] m48_107;
   assign m48_107 =10'b0;

   // m48_108 = W*in
   wire signed [9:0] m48_108;
   assign m48_108 ={ {4{neg48[5]}} , neg48[5:0] };

   // m48_109 = W*in
   wire signed [9:0] m48_109;
   assign m48_109 =10'b0;

   // m48_110 = W*in
   wire signed [9:0] m48_110;
   assign m48_110 =10'b0;

   // m48_111 = W*in
   wire signed [9:0] m48_111;
   assign m48_111 =10'b0;

   // m48_112 = W*in
   wire signed [9:0] m48_112;
   assign m48_112 =10'b0;

   // m48_113 = W*in
   wire signed [9:0] m48_113;
   assign m48_113 =10'b0;

   // m48_114 = W*in
   wire signed [9:0] m48_114;
   assign m48_114 =10'b0;

   // m48_115 = W*in
   wire signed [9:0] m48_115;
   assign m48_115 =10'b0;

   // m48_116 = W*in
   wire signed [9:0] m48_116;
   assign m48_116 =10'b0;

   // m48_117 = W*in
   wire signed [9:0] m48_117;
   assign m48_117 =10'b0;

   // m49_1 = W*in
   wire signed [9:0] m49_1;
   assign m49_1 ={ {4{in49[5]}} , in49[5:0] };

   // m49_2 = W*in
   wire signed [9:0] m49_2;
   assign m49_2 ={ {4{in49[5]}} , in49[5:0] };

   // m49_3 = W*in
   wire signed [9:0] m49_3;
   assign m49_3 =10'b0;

   // m49_4 = W*in
   wire signed [9:0] m49_4;
   assign m49_4 ={ {4{in49[5]}} , in49[5:0] };

   // m49_5 = W*in
   wire signed [9:0] m49_5;
   assign m49_5 =10'b0;

   // m49_6 = W*in
   wire signed [9:0] m49_6;
   assign m49_6 ={ {4{in49[5]}} , in49[5:0] };

   // m49_7 = W*in
   wire signed [9:0] m49_7;
   assign m49_7 =10'b0;

   // m49_8 = W*in
   wire signed [9:0] m49_8;
   assign m49_8 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_9 = W*in
   wire signed [9:0] m49_9;
   assign m49_9 =10'b0;

   // m49_10 = W*in
   wire signed [9:0] m49_10;
   assign m49_10 =10'b0;

   // m49_11 = W*in
   wire signed [9:0] m49_11;
   assign m49_11 ={ {4{in49[5]}} , in49[5:0] };

   // m49_12 = W*in
   wire signed [9:0] m49_12;
   assign m49_12 =10'b0;

   // m49_13 = W*in
   wire signed [9:0] m49_13;
   assign m49_13 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_14 = W*in
   wire signed [9:0] m49_14;
   assign m49_14 =10'b0;

   // m49_15 = W*in
   wire signed [9:0] m49_15;
   assign m49_15 =10'b0;

   // m49_16 = W*in
   wire signed [9:0] m49_16;
   assign m49_16 ={ {4{in49[5]}} , in49[5:0] };

   // m49_17 = W*in
   wire signed [9:0] m49_17;
   assign m49_17 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_18 = W*in
   wire signed [9:0] m49_18;
   assign m49_18 =10'b0;

   // m49_19 = W*in
   wire signed [9:0] m49_19;
   assign m49_19 =10'b0;

   // m49_20 = W*in
   wire signed [9:0] m49_20;
   assign m49_20 =10'b0;

   // m49_21 = W*in
   wire signed [9:0] m49_21;
   assign m49_21 =10'b0;

   // m49_22 = W*in
   wire signed [9:0] m49_22;
   assign m49_22 ={ {4{in49[5]}} , in49[5:0] };

   // m49_23 = W*in
   wire signed [9:0] m49_23;
   assign m49_23 =10'b0;

   // m49_24 = W*in
   wire signed [9:0] m49_24;
   assign m49_24 =10'b0;

   // m49_25 = W*in
   wire signed [9:0] m49_25;
   assign m49_25 =10'b0;

   // m49_26 = W*in
   wire signed [9:0] m49_26;
   assign m49_26 =10'b0;

   // m49_27 = W*in
   wire signed [9:0] m49_27;
   assign m49_27 ={ {4{in49[5]}} , in49[5:0] };

   // m49_28 = W*in
   wire signed [9:0] m49_28;
   assign m49_28 =10'b0;

   // m49_29 = W*in
   wire signed [9:0] m49_29;
   assign m49_29 ={ {5{neg49[5]}} , neg49[5:1] };

   // m49_30 = W*in
   wire signed [9:0] m49_30;
   assign m49_30 ={ {5{neg49[5]}} , neg49[5:1] };

   // m49_31 = W*in
   wire signed [9:0] m49_31;
   assign m49_31 ={ {5{neg49[5]}} , neg49[5:1] };

   // m49_32 = W*in
   wire signed [9:0] m49_32;
   assign m49_32 =10'b0;

   // m49_33 = W*in
   wire signed [9:0] m49_33;
   assign m49_33 ={ {4{in49[5]}} , in49[5:0] };

   // m49_34 = W*in
   wire signed [9:0] m49_34;
   assign m49_34 =10'b0;

   // m49_35 = W*in
   wire signed [9:0] m49_35;
   assign m49_35 =10'b0;

   // m49_36 = W*in
   wire signed [9:0] m49_36;
   assign m49_36 ={ {4{in49[5]}} , in49[5:0] };

   // m49_37 = W*in
   wire signed [9:0] m49_37;
   assign m49_37 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_38 = W*in
   wire signed [9:0] m49_38;
   assign m49_38 =10'b0;

   // m49_39 = W*in
   wire signed [9:0] m49_39;
   assign m49_39 =10'b0;

   // m49_40 = W*in
   wire signed [9:0] m49_40;
   assign m49_40 =10'b0;

   // m49_41 = W*in
   wire signed [9:0] m49_41;
   assign m49_41 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_42 = W*in
   wire signed [9:0] m49_42;
   assign m49_42 =10'b0;

   // m49_43 = W*in
   wire signed [9:0] m49_43;
   assign m49_43 ={ {4{in49[5]}} , in49[5:0] };

   // m49_44 = W*in
   wire signed [9:0] m49_44;
   assign m49_44 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_45 = W*in
   wire signed [9:0] m49_45;
   assign m49_45 =10'b0;

   // m49_46 = W*in
   wire signed [9:0] m49_46;
   assign m49_46 ={ {4{in49[5]}} , in49[5:0] };

   // m49_47 = W*in
   wire signed [9:0] m49_47;
   assign m49_47 =10'b0;

   // m49_48 = W*in
   wire signed [9:0] m49_48;
   assign m49_48 =10'b0;

   // m49_49 = W*in
   wire signed [9:0] m49_49;
   assign m49_49 ={ {3{in49[5]}} , in49 , {1{1'b0}} };

   // m49_50 = W*in
   wire signed [9:0] m49_50;
   assign m49_50 =10'b0;

   // m49_51 = W*in
   wire signed [9:0] m49_51;
   assign m49_51 =10'b0;

   // m49_52 = W*in
   wire signed [9:0] m49_52;
   assign m49_52 =10'b0;

   // m49_53 = W*in
   wire signed [9:0] m49_53;
   assign m49_53 =10'b0;

   // m49_54 = W*in
   wire signed [9:0] m49_54;
   assign m49_54 =10'b0;

   // m49_55 = W*in
   wire signed [9:0] m49_55;
   assign m49_55 =10'b0;

   // m49_56 = W*in
   wire signed [9:0] m49_56;
   assign m49_56 ={ {4{in49[5]}} , in49[5:0] };

   // m49_57 = W*in
   wire signed [9:0] m49_57;
   assign m49_57 =10'b0;

   // m49_58 = W*in
   wire signed [9:0] m49_58;
   assign m49_58 ={ {4{in49[5]}} , in49[5:0] };

   // m49_59 = W*in
   wire signed [9:0] m49_59;
   assign m49_59 ={ {5{in49[5]}} , in49[5:1] };

   // m49_60 = W*in
   wire signed [9:0] m49_60;
   assign m49_60 =10'b0;

   // m49_61 = W*in
   wire signed [9:0] m49_61;
   assign m49_61 ={ {4{in49[5]}} , in49[5:0] };

   // m49_62 = W*in
   wire signed [9:0] m49_62;
   assign m49_62 ={ {4{in49[5]}} , in49[5:0] };

   // m49_63 = W*in
   wire signed [9:0] m49_63;
   assign m49_63 =10'b0;

   // m49_64 = W*in
   wire signed [9:0] m49_64;
   assign m49_64 =10'b0;

   // m49_65 = W*in
   wire signed [9:0] m49_65;
   assign m49_65 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_66 = W*in
   wire signed [9:0] m49_66;
   assign m49_66 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_67 = W*in
   wire signed [9:0] m49_67;
   assign m49_67 =10'b0;

   // m49_68 = W*in
   wire signed [9:0] m49_68;
   assign m49_68 =10'b0;

   // m49_69 = W*in
   wire signed [9:0] m49_69;
   assign m49_69 =10'b0;

   // m49_70 = W*in
   wire signed [9:0] m49_70;
   assign m49_70 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_71 = W*in
   wire signed [9:0] m49_71;
   assign m49_71 ={ {4{in49[5]}} , in49[5:0] };

   // m49_72 = W*in
   wire signed [9:0] m49_72;
   assign m49_72 ={ {4{in49[5]}} , in49[5:0] };

   // m49_73 = W*in
   wire signed [9:0] m49_73;
   assign m49_73 ={ {4{in49[5]}} , in49[5:0] };

   // m49_74 = W*in
   wire signed [9:0] m49_74;
   assign m49_74 =10'b0;

   // m49_75 = W*in
   wire signed [9:0] m49_75;
   assign m49_75 ={ {4{in49[5]}} , in49[5:0] };

   // m49_76 = W*in
   wire signed [9:0] m49_76;
   assign m49_76 =10'b0;

   // m49_77 = W*in
   wire signed [9:0] m49_77;
   assign m49_77 ={ {4{in49[5]}} , in49[5:0] };

   // m49_78 = W*in
   wire signed [9:0] m49_78;
   assign m49_78 =10'b0;

   // m49_79 = W*in
   wire signed [9:0] m49_79;
   assign m49_79 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_80 = W*in
   wire signed [9:0] m49_80;
   assign m49_80 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_81 = W*in
   wire signed [9:0] m49_81;
   assign m49_81 ={ {5{in49[5]}} , in49[5:1] };

   // m49_82 = W*in
   wire signed [9:0] m49_82;
   assign m49_82 =10'b0;

   // m49_83 = W*in
   wire signed [9:0] m49_83;
   assign m49_83 =10'b0;

   // m49_84 = W*in
   wire signed [9:0] m49_84;
   assign m49_84 =10'b0;

   // m49_85 = W*in
   wire signed [9:0] m49_85;
   assign m49_85 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_86 = W*in
   wire signed [9:0] m49_86;
   assign m49_86 =10'b0;

   // m49_87 = W*in
   wire signed [9:0] m49_87;
   assign m49_87 =10'b0;

   // m49_88 = W*in
   wire signed [9:0] m49_88;
   assign m49_88 =10'b0;

   // m49_89 = W*in
   wire signed [9:0] m49_89;
   assign m49_89 =10'b0;

   // m49_90 = W*in
   wire signed [9:0] m49_90;
   assign m49_90 =10'b0;

   // m49_91 = W*in
   wire signed [9:0] m49_91;
   assign m49_91 =10'b0;

   // m49_92 = W*in
   wire signed [9:0] m49_92;
   assign m49_92 =10'b0;

   // m49_93 = W*in
   wire signed [9:0] m49_93;
   assign m49_93 =10'b0;

   // m49_94 = W*in
   wire signed [9:0] m49_94;
   assign m49_94 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_95 = W*in
   wire signed [9:0] m49_95;
   assign m49_95 ={ {4{in49[5]}} , in49[5:0] };

   // m49_96 = W*in
   wire signed [9:0] m49_96;
   assign m49_96 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_97 = W*in
   wire signed [9:0] m49_97;
   assign m49_97 =10'b0;

   // m49_98 = W*in
   wire signed [9:0] m49_98;
   assign m49_98 =10'b0;

   // m49_99 = W*in
   wire signed [9:0] m49_99;
   assign m49_99 =10'b0;

   // m49_100 = W*in
   wire signed [9:0] m49_100;
   assign m49_100 =10'b0;

   // m49_101 = W*in
   wire signed [9:0] m49_101;
   assign m49_101 ={ {4{in49[5]}} , in49[5:0] };

   // m49_102 = W*in
   wire signed [9:0] m49_102;
   assign m49_102 =10'b0;

   // m49_103 = W*in
   wire signed [9:0] m49_103;
   assign m49_103 =10'b0;

   // m49_104 = W*in
   wire signed [9:0] m49_104;
   assign m49_104 =10'b0;

   // m49_105 = W*in
   wire signed [9:0] m49_105;
   assign m49_105 =10'b0;

   // m49_106 = W*in
   wire signed [9:0] m49_106;
   assign m49_106 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_107 = W*in
   wire signed [9:0] m49_107;
   assign m49_107 ={ {4{in49[5]}} , in49[5:0] };

   // m49_108 = W*in
   wire signed [9:0] m49_108;
   assign m49_108 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_109 = W*in
   wire signed [9:0] m49_109;
   assign m49_109 ={ {4{neg49[5]}} , neg49[5:0] };

   // m49_110 = W*in
   wire signed [9:0] m49_110;
   assign m49_110 =10'b0;

   // m49_111 = W*in
   wire signed [9:0] m49_111;
   assign m49_111 =10'b0;

   // m49_112 = W*in
   wire signed [9:0] m49_112;
   assign m49_112 =10'b0;

   // m49_113 = W*in
   wire signed [9:0] m49_113;
   assign m49_113 =10'b0;

   // m49_114 = W*in
   wire signed [9:0] m49_114;
   assign m49_114 =10'b0;

   // m49_115 = W*in
   wire signed [9:0] m49_115;
   assign m49_115 =10'b0;

   // m49_116 = W*in
   wire signed [9:0] m49_116;
   assign m49_116 ={ {3{neg49[5]}} , neg49 , {1{1'b0}} };

   // m49_117 = W*in
   wire signed [9:0] m49_117;
   assign m49_117 =10'b0;

   // m50_1 = W*in
   wire signed [9:0] m50_1;
   assign m50_1 =10'b0;

   // m50_2 = W*in
   wire signed [9:0] m50_2;
   assign m50_2 =10'b0;

   // m50_3 = W*in
   wire signed [9:0] m50_3;
   assign m50_3 =10'b0;

   // m50_4 = W*in
   wire signed [9:0] m50_4;
   assign m50_4 =10'b0;

   // m50_5 = W*in
   wire signed [9:0] m50_5;
   assign m50_5 ={ {4{in50[5]}} , in50[5:0] };

   // m50_6 = W*in
   wire signed [9:0] m50_6;
   assign m50_6 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_7 = W*in
   wire signed [9:0] m50_7;
   assign m50_7 =10'b0;

   // m50_8 = W*in
   wire signed [9:0] m50_8;
   assign m50_8 =10'b0;

   // m50_9 = W*in
   wire signed [9:0] m50_9;
   assign m50_9 =10'b0;

   // m50_10 = W*in
   wire signed [9:0] m50_10;
   assign m50_10 =10'b0;

   // m50_11 = W*in
   wire signed [9:0] m50_11;
   assign m50_11 ={ {4{in50[5]}} , in50[5:0] };

   // m50_12 = W*in
   wire signed [9:0] m50_12;
   assign m50_12 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_13 = W*in
   wire signed [9:0] m50_13;
   assign m50_13 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_14 = W*in
   wire signed [9:0] m50_14;
   assign m50_14 =10'b0;

   // m50_15 = W*in
   wire signed [9:0] m50_15;
   assign m50_15 =10'b0;

   // m50_16 = W*in
   wire signed [9:0] m50_16;
   assign m50_16 =10'b0;

   // m50_17 = W*in
   wire signed [9:0] m50_17;
   assign m50_17 ={ {5{in50[5]}} , in50[5:1] };

   // m50_18 = W*in
   wire signed [9:0] m50_18;
   assign m50_18 =10'b0;

   // m50_19 = W*in
   wire signed [9:0] m50_19;
   assign m50_19 ={ {4{in50[5]}} , in50[5:0] };

   // m50_20 = W*in
   wire signed [9:0] m50_20;
   assign m50_20 ={ {5{in50[5]}} , in50[5:1] };

   // m50_21 = W*in
   wire signed [9:0] m50_21;
   assign m50_21 =10'b0;

   // m50_22 = W*in
   wire signed [9:0] m50_22;
   assign m50_22 ={ {4{in50[5]}} , in50[5:0] };

   // m50_23 = W*in
   wire signed [9:0] m50_23;
   assign m50_23 =10'b0;

   // m50_24 = W*in
   wire signed [9:0] m50_24;
   assign m50_24 ={ {5{in50[5]}} , in50[5:1] };

   // m50_25 = W*in
   wire signed [9:0] m50_25;
   assign m50_25 ={ {4{in50[5]}} , in50[5:0] };

   // m50_26 = W*in
   wire signed [9:0] m50_26;
   assign m50_26 =10'b0;

   // m50_27 = W*in
   wire signed [9:0] m50_27;
   assign m50_27 ={ {5{in50[5]}} , in50[5:1] };

   // m50_28 = W*in
   wire signed [9:0] m50_28;
   assign m50_28 ={ {4{in50[5]}} , in50[5:0] };

   // m50_29 = W*in
   wire signed [9:0] m50_29;
   assign m50_29 =10'b0;

   // m50_30 = W*in
   wire signed [9:0] m50_30;
   assign m50_30 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_31 = W*in
   wire signed [9:0] m50_31;
   assign m50_31 =10'b0;

   // m50_32 = W*in
   wire signed [9:0] m50_32;
   assign m50_32 =10'b0;

   // m50_33 = W*in
   wire signed [9:0] m50_33;
   assign m50_33 =10'b0;

   // m50_34 = W*in
   wire signed [9:0] m50_34;
   assign m50_34 ={ {4{in50[5]}} , in50[5:0] };

   // m50_35 = W*in
   wire signed [9:0] m50_35;
   assign m50_35 =10'b0;

   // m50_36 = W*in
   wire signed [9:0] m50_36;
   assign m50_36 =10'b0;

   // m50_37 = W*in
   wire signed [9:0] m50_37;
   assign m50_37 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_38 = W*in
   wire signed [9:0] m50_38;
   assign m50_38 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_39 = W*in
   wire signed [9:0] m50_39;
   assign m50_39 =10'b0;

   // m50_40 = W*in
   wire signed [9:0] m50_40;
   assign m50_40 =10'b0;

   // m50_41 = W*in
   wire signed [9:0] m50_41;
   assign m50_41 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_42 = W*in
   wire signed [9:0] m50_42;
   assign m50_42 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_43 = W*in
   wire signed [9:0] m50_43;
   assign m50_43 ={ {4{in50[5]}} , in50[5:0] };

   // m50_44 = W*in
   wire signed [9:0] m50_44;
   assign m50_44 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_45 = W*in
   wire signed [9:0] m50_45;
   assign m50_45 =10'b0;

   // m50_46 = W*in
   wire signed [9:0] m50_46;
   assign m50_46 =10'b0;

   // m50_47 = W*in
   wire signed [9:0] m50_47;
   assign m50_47 ={ {4{in50[5]}} , in50[5:0] };

   // m50_48 = W*in
   wire signed [9:0] m50_48;
   assign m50_48 =10'b0;

   // m50_49 = W*in
   wire signed [9:0] m50_49;
   assign m50_49 ={ {4{in50[5]}} , in50[5:0] };

   // m50_50 = W*in
   wire signed [9:0] m50_50;
   assign m50_50 =10'b0;

   // m50_51 = W*in
   wire signed [9:0] m50_51;
   assign m50_51 =10'b0;

   // m50_52 = W*in
   wire signed [9:0] m50_52;
   assign m50_52 =10'b0;

   // m50_53 = W*in
   wire signed [9:0] m50_53;
   assign m50_53 ={ {5{in50[5]}} , in50[5:1] };

   // m50_54 = W*in
   wire signed [9:0] m50_54;
   assign m50_54 ={ {4{in50[5]}} , in50[5:0] };

   // m50_55 = W*in
   wire signed [9:0] m50_55;
   assign m50_55 =10'b0;

   // m50_56 = W*in
   wire signed [9:0] m50_56;
   assign m50_56 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_57 = W*in
   wire signed [9:0] m50_57;
   assign m50_57 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_58 = W*in
   wire signed [9:0] m50_58;
   assign m50_58 =10'b0;

   // m50_59 = W*in
   wire signed [9:0] m50_59;
   assign m50_59 ={ {4{in50[5]}} , in50[5:0] };

   // m50_60 = W*in
   wire signed [9:0] m50_60;
   assign m50_60 =10'b0;

   // m50_61 = W*in
   wire signed [9:0] m50_61;
   assign m50_61 =10'b0;

   // m50_62 = W*in
   wire signed [9:0] m50_62;
   assign m50_62 =10'b0;

   // m50_63 = W*in
   wire signed [9:0] m50_63;
   assign m50_63 =10'b0;

   // m50_64 = W*in
   wire signed [9:0] m50_64;
   assign m50_64 =10'b0;

   // m50_65 = W*in
   wire signed [9:0] m50_65;
   assign m50_65 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_66 = W*in
   wire signed [9:0] m50_66;
   assign m50_66 ={ {5{in50[5]}} , in50[5:1] };

   // m50_67 = W*in
   wire signed [9:0] m50_67;
   assign m50_67 ={ {4{in50[5]}} , in50[5:0] };

   // m50_68 = W*in
   wire signed [9:0] m50_68;
   assign m50_68 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_69 = W*in
   wire signed [9:0] m50_69;
   assign m50_69 =10'b0;

   // m50_70 = W*in
   wire signed [9:0] m50_70;
   assign m50_70 ={ {4{in50[5]}} , in50[5:0] };

   // m50_71 = W*in
   wire signed [9:0] m50_71;
   assign m50_71 =10'b0;

   // m50_72 = W*in
   wire signed [9:0] m50_72;
   assign m50_72 =10'b0;

   // m50_73 = W*in
   wire signed [9:0] m50_73;
   assign m50_73 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_74 = W*in
   wire signed [9:0] m50_74;
   assign m50_74 ={ {5{in50[5]}} , in50[5:1] };

   // m50_75 = W*in
   wire signed [9:0] m50_75;
   assign m50_75 =10'b0;

   // m50_76 = W*in
   wire signed [9:0] m50_76;
   assign m50_76 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_77 = W*in
   wire signed [9:0] m50_77;
   assign m50_77 =10'b0;

   // m50_78 = W*in
   wire signed [9:0] m50_78;
   assign m50_78 =10'b0;

   // m50_79 = W*in
   wire signed [9:0] m50_79;
   assign m50_79 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_80 = W*in
   wire signed [9:0] m50_80;
   assign m50_80 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_81 = W*in
   wire signed [9:0] m50_81;
   assign m50_81 =10'b0;

   // m50_82 = W*in
   wire signed [9:0] m50_82;
   assign m50_82 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_83 = W*in
   wire signed [9:0] m50_83;
   assign m50_83 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_84 = W*in
   wire signed [9:0] m50_84;
   assign m50_84 =10'b0;

   // m50_85 = W*in
   wire signed [9:0] m50_85;
   assign m50_85 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_86 = W*in
   wire signed [9:0] m50_86;
   assign m50_86 =10'b0;

   // m50_87 = W*in
   wire signed [9:0] m50_87;
   assign m50_87 ={ {4{in50[5]}} , in50[5:0] };

   // m50_88 = W*in
   wire signed [9:0] m50_88;
   assign m50_88 ={ {4{in50[5]}} , in50[5:0] };

   // m50_89 = W*in
   wire signed [9:0] m50_89;
   assign m50_89 =10'b0;

   // m50_90 = W*in
   wire signed [9:0] m50_90;
   assign m50_90 =10'b0;

   // m50_91 = W*in
   wire signed [9:0] m50_91;
   assign m50_91 ={ {3{in50[5]}} , in50 , {1{1'b0}} };

   // m50_92 = W*in
   wire signed [9:0] m50_92;
   assign m50_92 =10'b0;

   // m50_93 = W*in
   wire signed [9:0] m50_93;
   assign m50_93 =10'b0;

   // m50_94 = W*in
   wire signed [9:0] m50_94;
   assign m50_94 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_95 = W*in
   wire signed [9:0] m50_95;
   assign m50_95 =10'b0;

   // m50_96 = W*in
   wire signed [9:0] m50_96;
   assign m50_96 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_97 = W*in
   wire signed [9:0] m50_97;
   assign m50_97 ={ {4{in50[5]}} , in50[5:0] };

   // m50_98 = W*in
   wire signed [9:0] m50_98;
   assign m50_98 =10'b0;

   // m50_99 = W*in
   wire signed [9:0] m50_99;
   assign m50_99 =10'b0;

   // m50_100 = W*in
   wire signed [9:0] m50_100;
   assign m50_100 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_101 = W*in
   wire signed [9:0] m50_101;
   assign m50_101 =10'b0;

   // m50_102 = W*in
   wire signed [9:0] m50_102;
   assign m50_102 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_103 = W*in
   wire signed [9:0] m50_103;
   assign m50_103 =10'b0;

   // m50_104 = W*in
   wire signed [9:0] m50_104;
   assign m50_104 =10'b0;

   // m50_105 = W*in
   wire signed [9:0] m50_105;
   assign m50_105 =10'b0;

   // m50_106 = W*in
   wire signed [9:0] m50_106;
   assign m50_106 =10'b0;

   // m50_107 = W*in
   wire signed [9:0] m50_107;
   assign m50_107 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_108 = W*in
   wire signed [9:0] m50_108;
   assign m50_108 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_109 = W*in
   wire signed [9:0] m50_109;
   assign m50_109 ={ {4{neg50[5]}} , neg50[5:0] };

   // m50_110 = W*in
   wire signed [9:0] m50_110;
   assign m50_110 ={ {4{in50[5]}} , in50[5:0] };

   // m50_111 = W*in
   wire signed [9:0] m50_111;
   assign m50_111 =10'b0;

   // m50_112 = W*in
   wire signed [9:0] m50_112;
   assign m50_112 ={ {5{neg50[5]}} , neg50[5:1] };

   // m50_113 = W*in
   wire signed [9:0] m50_113;
   assign m50_113 =10'b0;

   // m50_114 = W*in
   wire signed [9:0] m50_114;
   assign m50_114 ={ {4{in50[5]}} , in50[5:0] };

   // m50_115 = W*in
   wire signed [9:0] m50_115;
   assign m50_115 =10'b0;

   // m50_116 = W*in
   wire signed [9:0] m50_116;
   assign m50_116 ={ {3{neg50[5]}} , neg50 , {1{1'b0}} };

   // m50_117 = W*in
   wire signed [9:0] m50_117;
   assign m50_117 =10'b0;

   // m51_1 = W*in
   wire signed [9:0] m51_1;
   assign m51_1 =10'b0;

   // m51_2 = W*in
   wire signed [9:0] m51_2;
   assign m51_2 =10'b0;

   // m51_3 = W*in
   wire signed [9:0] m51_3;
   assign m51_3 =10'b0;

   // m51_4 = W*in
   wire signed [9:0] m51_4;
   assign m51_4 =10'b0;

   // m51_5 = W*in
   wire signed [9:0] m51_5;
   assign m51_5 =10'b0;

   // m51_6 = W*in
   wire signed [9:0] m51_6;
   assign m51_6 ={ {4{in51[5]}} , in51[5:0] };

   // m51_7 = W*in
   wire signed [9:0] m51_7;
   assign m51_7 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_8 = W*in
   wire signed [9:0] m51_8;
   assign m51_8 =10'b0;

   // m51_9 = W*in
   wire signed [9:0] m51_9;
   assign m51_9 =10'b0;

   // m51_10 = W*in
   wire signed [9:0] m51_10;
   assign m51_10 =10'b0;

   // m51_11 = W*in
   wire signed [9:0] m51_11;
   assign m51_11 =10'b0;

   // m51_12 = W*in
   wire signed [9:0] m51_12;
   assign m51_12 =10'b0;

   // m51_13 = W*in
   wire signed [9:0] m51_13;
   assign m51_13 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_14 = W*in
   wire signed [9:0] m51_14;
   assign m51_14 =10'b0;

   // m51_15 = W*in
   wire signed [9:0] m51_15;
   assign m51_15 =10'b0;

   // m51_16 = W*in
   wire signed [9:0] m51_16;
   assign m51_16 =10'b0;

   // m51_17 = W*in
   wire signed [9:0] m51_17;
   assign m51_17 =10'b0;

   // m51_18 = W*in
   wire signed [9:0] m51_18;
   assign m51_18 =10'b0;

   // m51_19 = W*in
   wire signed [9:0] m51_19;
   assign m51_19 ={ {4{in51[5]}} , in51[5:0] };

   // m51_20 = W*in
   wire signed [9:0] m51_20;
   assign m51_20 =10'b0;

   // m51_21 = W*in
   wire signed [9:0] m51_21;
   assign m51_21 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_22 = W*in
   wire signed [9:0] m51_22;
   assign m51_22 ={ {4{in51[5]}} , in51[5:0] };

   // m51_23 = W*in
   wire signed [9:0] m51_23;
   assign m51_23 =10'b0;

   // m51_24 = W*in
   wire signed [9:0] m51_24;
   assign m51_24 ={ {4{in51[5]}} , in51[5:0] };

   // m51_25 = W*in
   wire signed [9:0] m51_25;
   assign m51_25 =10'b0;

   // m51_26 = W*in
   wire signed [9:0] m51_26;
   assign m51_26 ={ {5{in51[5]}} , in51[5:1] };

   // m51_27 = W*in
   wire signed [9:0] m51_27;
   assign m51_27 =10'b0;

   // m51_28 = W*in
   wire signed [9:0] m51_28;
   assign m51_28 =10'b0;

   // m51_29 = W*in
   wire signed [9:0] m51_29;
   assign m51_29 =10'b0;

   // m51_30 = W*in
   wire signed [9:0] m51_30;
   assign m51_30 =10'b0;

   // m51_31 = W*in
   wire signed [9:0] m51_31;
   assign m51_31 =10'b0;

   // m51_32 = W*in
   wire signed [9:0] m51_32;
   assign m51_32 =10'b0;

   // m51_33 = W*in
   wire signed [9:0] m51_33;
   assign m51_33 =10'b0;

   // m51_34 = W*in
   wire signed [9:0] m51_34;
   assign m51_34 ={ {4{in51[5]}} , in51[5:0] };

   // m51_35 = W*in
   wire signed [9:0] m51_35;
   assign m51_35 ={ {4{in51[5]}} , in51[5:0] };

   // m51_36 = W*in
   wire signed [9:0] m51_36;
   assign m51_36 =10'b0;

   // m51_37 = W*in
   wire signed [9:0] m51_37;
   assign m51_37 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_38 = W*in
   wire signed [9:0] m51_38;
   assign m51_38 ={ {4{in51[5]}} , in51[5:0] };

   // m51_39 = W*in
   wire signed [9:0] m51_39;
   assign m51_39 ={ {5{in51[5]}} , in51[5:1] };

   // m51_40 = W*in
   wire signed [9:0] m51_40;
   assign m51_40 =10'b0;

   // m51_41 = W*in
   wire signed [9:0] m51_41;
   assign m51_41 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_42 = W*in
   wire signed [9:0] m51_42;
   assign m51_42 =10'b0;

   // m51_43 = W*in
   wire signed [9:0] m51_43;
   assign m51_43 =10'b0;

   // m51_44 = W*in
   wire signed [9:0] m51_44;
   assign m51_44 ={ {4{in51[5]}} , in51[5:0] };

   // m51_45 = W*in
   wire signed [9:0] m51_45;
   assign m51_45 =10'b0;

   // m51_46 = W*in
   wire signed [9:0] m51_46;
   assign m51_46 =10'b0;

   // m51_47 = W*in
   wire signed [9:0] m51_47;
   assign m51_47 =10'b0;

   // m51_48 = W*in
   wire signed [9:0] m51_48;
   assign m51_48 =10'b0;

   // m51_49 = W*in
   wire signed [9:0] m51_49;
   assign m51_49 =10'b0;

   // m51_50 = W*in
   wire signed [9:0] m51_50;
   assign m51_50 =10'b0;

   // m51_51 = W*in
   wire signed [9:0] m51_51;
   assign m51_51 =10'b0;

   // m51_52 = W*in
   wire signed [9:0] m51_52;
   assign m51_52 =10'b0;

   // m51_53 = W*in
   wire signed [9:0] m51_53;
   assign m51_53 ={ {4{in51[5]}} , in51[5:0] };

   // m51_54 = W*in
   wire signed [9:0] m51_54;
   assign m51_54 ={ {4{in51[5]}} , in51[5:0] };

   // m51_55 = W*in
   wire signed [9:0] m51_55;
   assign m51_55 =10'b0;

   // m51_56 = W*in
   wire signed [9:0] m51_56;
   assign m51_56 =10'b0;

   // m51_57 = W*in
   wire signed [9:0] m51_57;
   assign m51_57 =10'b0;

   // m51_58 = W*in
   wire signed [9:0] m51_58;
   assign m51_58 =10'b0;

   // m51_59 = W*in
   wire signed [9:0] m51_59;
   assign m51_59 =10'b0;

   // m51_60 = W*in
   wire signed [9:0] m51_60;
   assign m51_60 =10'b0;

   // m51_61 = W*in
   wire signed [9:0] m51_61;
   assign m51_61 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_62 = W*in
   wire signed [9:0] m51_62;
   assign m51_62 =10'b0;

   // m51_63 = W*in
   wire signed [9:0] m51_63;
   assign m51_63 =10'b0;

   // m51_64 = W*in
   wire signed [9:0] m51_64;
   assign m51_64 =10'b0;

   // m51_65 = W*in
   wire signed [9:0] m51_65;
   assign m51_65 ={ {5{neg51[5]}} , neg51[5:1] };

   // m51_66 = W*in
   wire signed [9:0] m51_66;
   assign m51_66 =10'b0;

   // m51_67 = W*in
   wire signed [9:0] m51_67;
   assign m51_67 =10'b0;

   // m51_68 = W*in
   wire signed [9:0] m51_68;
   assign m51_68 =10'b0;

   // m51_69 = W*in
   wire signed [9:0] m51_69;
   assign m51_69 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_70 = W*in
   wire signed [9:0] m51_70;
   assign m51_70 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_71 = W*in
   wire signed [9:0] m51_71;
   assign m51_71 =10'b0;

   // m51_72 = W*in
   wire signed [9:0] m51_72;
   assign m51_72 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_73 = W*in
   wire signed [9:0] m51_73;
   assign m51_73 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_74 = W*in
   wire signed [9:0] m51_74;
   assign m51_74 =10'b0;

   // m51_75 = W*in
   wire signed [9:0] m51_75;
   assign m51_75 ={ {4{in51[5]}} , in51[5:0] };

   // m51_76 = W*in
   wire signed [9:0] m51_76;
   assign m51_76 ={ {4{in51[5]}} , in51[5:0] };

   // m51_77 = W*in
   wire signed [9:0] m51_77;
   assign m51_77 =10'b0;

   // m51_78 = W*in
   wire signed [9:0] m51_78;
   assign m51_78 =10'b0;

   // m51_79 = W*in
   wire signed [9:0] m51_79;
   assign m51_79 =10'b0;

   // m51_80 = W*in
   wire signed [9:0] m51_80;
   assign m51_80 =10'b0;

   // m51_81 = W*in
   wire signed [9:0] m51_81;
   assign m51_81 =10'b0;

   // m51_82 = W*in
   wire signed [9:0] m51_82;
   assign m51_82 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_83 = W*in
   wire signed [9:0] m51_83;
   assign m51_83 =10'b0;

   // m51_84 = W*in
   wire signed [9:0] m51_84;
   assign m51_84 =10'b0;

   // m51_85 = W*in
   wire signed [9:0] m51_85;
   assign m51_85 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_86 = W*in
   wire signed [9:0] m51_86;
   assign m51_86 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_87 = W*in
   wire signed [9:0] m51_87;
   assign m51_87 =10'b0;

   // m51_88 = W*in
   wire signed [9:0] m51_88;
   assign m51_88 =10'b0;

   // m51_89 = W*in
   wire signed [9:0] m51_89;
   assign m51_89 =10'b0;

   // m51_90 = W*in
   wire signed [9:0] m51_90;
   assign m51_90 =10'b0;

   // m51_91 = W*in
   wire signed [9:0] m51_91;
   assign m51_91 ={ {4{in51[5]}} , in51[5:0] };

   // m51_92 = W*in
   wire signed [9:0] m51_92;
   assign m51_92 =10'b0;

   // m51_93 = W*in
   wire signed [9:0] m51_93;
   assign m51_93 =10'b0;

   // m51_94 = W*in
   wire signed [9:0] m51_94;
   assign m51_94 =10'b0;

   // m51_95 = W*in
   wire signed [9:0] m51_95;
   assign m51_95 ={ {4{in51[5]}} , in51[5:0] };

   // m51_96 = W*in
   wire signed [9:0] m51_96;
   assign m51_96 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_97 = W*in
   wire signed [9:0] m51_97;
   assign m51_97 =10'b0;

   // m51_98 = W*in
   wire signed [9:0] m51_98;
   assign m51_98 =10'b0;

   // m51_99 = W*in
   wire signed [9:0] m51_99;
   assign m51_99 =10'b0;

   // m51_100 = W*in
   wire signed [9:0] m51_100;
   assign m51_100 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_101 = W*in
   wire signed [9:0] m51_101;
   assign m51_101 =10'b0;

   // m51_102 = W*in
   wire signed [9:0] m51_102;
   assign m51_102 =10'b0;

   // m51_103 = W*in
   wire signed [9:0] m51_103;
   assign m51_103 =10'b0;

   // m51_104 = W*in
   wire signed [9:0] m51_104;
   assign m51_104 =10'b0;

   // m51_105 = W*in
   wire signed [9:0] m51_105;
   assign m51_105 =10'b0;

   // m51_106 = W*in
   wire signed [9:0] m51_106;
   assign m51_106 =10'b0;

   // m51_107 = W*in
   wire signed [9:0] m51_107;
   assign m51_107 =10'b0;

   // m51_108 = W*in
   wire signed [9:0] m51_108;
   assign m51_108 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_109 = W*in
   wire signed [9:0] m51_109;
   assign m51_109 =10'b0;

   // m51_110 = W*in
   wire signed [9:0] m51_110;
   assign m51_110 ={ {4{in51[5]}} , in51[5:0] };

   // m51_111 = W*in
   wire signed [9:0] m51_111;
   assign m51_111 =10'b0;

   // m51_112 = W*in
   wire signed [9:0] m51_112;
   assign m51_112 =10'b0;

   // m51_113 = W*in
   wire signed [9:0] m51_113;
   assign m51_113 =10'b0;

   // m51_114 = W*in
   wire signed [9:0] m51_114;
   assign m51_114 =10'b0;

   // m51_115 = W*in
   wire signed [9:0] m51_115;
   assign m51_115 =10'b0;

   // m51_116 = W*in
   wire signed [9:0] m51_116;
   assign m51_116 ={ {4{neg51[5]}} , neg51[5:0] };

   // m51_117 = W*in
   wire signed [9:0] m51_117;
   assign m51_117 =10'b0;

   // m52_1 = W*in
   wire signed [9:0] m52_1;
   assign m52_1 =10'b0;

   // m52_2 = W*in
   wire signed [9:0] m52_2;
   assign m52_2 =10'b0;

   // m52_3 = W*in
   wire signed [9:0] m52_3;
   assign m52_3 =10'b0;

   // m52_4 = W*in
   wire signed [9:0] m52_4;
   assign m52_4 =10'b0;

   // m52_5 = W*in
   wire signed [9:0] m52_5;
   assign m52_5 =10'b0;

   // m52_6 = W*in
   wire signed [9:0] m52_6;
   assign m52_6 =10'b0;

   // m52_7 = W*in
   wire signed [9:0] m52_7;
   assign m52_7 =10'b0;

   // m52_8 = W*in
   wire signed [9:0] m52_8;
   assign m52_8 =10'b0;

   // m52_9 = W*in
   wire signed [9:0] m52_9;
   assign m52_9 =10'b0;

   // m52_10 = W*in
   wire signed [9:0] m52_10;
   assign m52_10 =10'b0;

   // m52_11 = W*in
   wire signed [9:0] m52_11;
   assign m52_11 =10'b0;

   // m52_12 = W*in
   wire signed [9:0] m52_12;
   assign m52_12 =10'b0;

   // m52_13 = W*in
   wire signed [9:0] m52_13;
   assign m52_13 =10'b0;

   // m52_14 = W*in
   wire signed [9:0] m52_14;
   assign m52_14 =10'b0;

   // m52_15 = W*in
   wire signed [9:0] m52_15;
   assign m52_15 =10'b0;

   // m52_16 = W*in
   wire signed [9:0] m52_16;
   assign m52_16 =10'b0;

   // m52_17 = W*in
   wire signed [9:0] m52_17;
   assign m52_17 =10'b0;

   // m52_18 = W*in
   wire signed [9:0] m52_18;
   assign m52_18 =10'b0;

   // m52_19 = W*in
   wire signed [9:0] m52_19;
   assign m52_19 =10'b0;

   // m52_20 = W*in
   wire signed [9:0] m52_20;
   assign m52_20 =10'b0;

   // m52_21 = W*in
   wire signed [9:0] m52_21;
   assign m52_21 ={ {5{neg52[5]}} , neg52[5:1] };

   // m52_22 = W*in
   wire signed [9:0] m52_22;
   assign m52_22 =10'b0;

   // m52_23 = W*in
   wire signed [9:0] m52_23;
   assign m52_23 =10'b0;

   // m52_24 = W*in
   wire signed [9:0] m52_24;
   assign m52_24 =10'b0;

   // m52_25 = W*in
   wire signed [9:0] m52_25;
   assign m52_25 ={ {4{in52[5]}} , in52[5:0] };

   // m52_26 = W*in
   wire signed [9:0] m52_26;
   assign m52_26 =10'b0;

   // m52_27 = W*in
   wire signed [9:0] m52_27;
   assign m52_27 =10'b0;

   // m52_28 = W*in
   wire signed [9:0] m52_28;
   assign m52_28 ={ {5{in52[5]}} , in52[5:1] };

   // m52_29 = W*in
   wire signed [9:0] m52_29;
   assign m52_29 =10'b0;

   // m52_30 = W*in
   wire signed [9:0] m52_30;
   assign m52_30 =10'b0;

   // m52_31 = W*in
   wire signed [9:0] m52_31;
   assign m52_31 ={ {5{in52[5]}} , in52[5:1] };

   // m52_32 = W*in
   wire signed [9:0] m52_32;
   assign m52_32 =10'b0;

   // m52_33 = W*in
   wire signed [9:0] m52_33;
   assign m52_33 =10'b0;

   // m52_34 = W*in
   wire signed [9:0] m52_34;
   assign m52_34 =10'b0;

   // m52_35 = W*in
   wire signed [9:0] m52_35;
   assign m52_35 =10'b0;

   // m52_36 = W*in
   wire signed [9:0] m52_36;
   assign m52_36 ={ {5{in52[5]}} , in52[5:1] };

   // m52_37 = W*in
   wire signed [9:0] m52_37;
   assign m52_37 =10'b0;

   // m52_38 = W*in
   wire signed [9:0] m52_38;
   assign m52_38 =10'b0;

   // m52_39 = W*in
   wire signed [9:0] m52_39;
   assign m52_39 =10'b0;

   // m52_40 = W*in
   wire signed [9:0] m52_40;
   assign m52_40 =10'b0;

   // m52_41 = W*in
   wire signed [9:0] m52_41;
   assign m52_41 =10'b0;

   // m52_42 = W*in
   wire signed [9:0] m52_42;
   assign m52_42 =10'b0;

   // m52_43 = W*in
   wire signed [9:0] m52_43;
   assign m52_43 =10'b0;

   // m52_44 = W*in
   wire signed [9:0] m52_44;
   assign m52_44 =10'b0;

   // m52_45 = W*in
   wire signed [9:0] m52_45;
   assign m52_45 =10'b0;

   // m52_46 = W*in
   wire signed [9:0] m52_46;
   assign m52_46 =10'b0;

   // m52_47 = W*in
   wire signed [9:0] m52_47;
   assign m52_47 =10'b0;

   // m52_48 = W*in
   wire signed [9:0] m52_48;
   assign m52_48 =10'b0;

   // m52_49 = W*in
   wire signed [9:0] m52_49;
   assign m52_49 =10'b0;

   // m52_50 = W*in
   wire signed [9:0] m52_50;
   assign m52_50 =10'b0;

   // m52_51 = W*in
   wire signed [9:0] m52_51;
   assign m52_51 =10'b0;

   // m52_52 = W*in
   wire signed [9:0] m52_52;
   assign m52_52 =10'b0;

   // m52_53 = W*in
   wire signed [9:0] m52_53;
   assign m52_53 =10'b0;

   // m52_54 = W*in
   wire signed [9:0] m52_54;
   assign m52_54 =10'b0;

   // m52_55 = W*in
   wire signed [9:0] m52_55;
   assign m52_55 =10'b0;

   // m52_56 = W*in
   wire signed [9:0] m52_56;
   assign m52_56 =10'b0;

   // m52_57 = W*in
   wire signed [9:0] m52_57;
   assign m52_57 =10'b0;

   // m52_58 = W*in
   wire signed [9:0] m52_58;
   assign m52_58 =10'b0;

   // m52_59 = W*in
   wire signed [9:0] m52_59;
   assign m52_59 ={ {4{in52[5]}} , in52[5:0] };

   // m52_60 = W*in
   wire signed [9:0] m52_60;
   assign m52_60 =10'b0;

   // m52_61 = W*in
   wire signed [9:0] m52_61;
   assign m52_61 =10'b0;

   // m52_62 = W*in
   wire signed [9:0] m52_62;
   assign m52_62 =10'b0;

   // m52_63 = W*in
   wire signed [9:0] m52_63;
   assign m52_63 =10'b0;

   // m52_64 = W*in
   wire signed [9:0] m52_64;
   assign m52_64 =10'b0;

   // m52_65 = W*in
   wire signed [9:0] m52_65;
   assign m52_65 =10'b0;

   // m52_66 = W*in
   wire signed [9:0] m52_66;
   assign m52_66 =10'b0;

   // m52_67 = W*in
   wire signed [9:0] m52_67;
   assign m52_67 =10'b0;

   // m52_68 = W*in
   wire signed [9:0] m52_68;
   assign m52_68 =10'b0;

   // m52_69 = W*in
   wire signed [9:0] m52_69;
   assign m52_69 ={ {5{neg52[5]}} , neg52[5:1] };

   // m52_70 = W*in
   wire signed [9:0] m52_70;
   assign m52_70 ={ {4{neg52[5]}} , neg52[5:0] };

   // m52_71 = W*in
   wire signed [9:0] m52_71;
   assign m52_71 =10'b0;

   // m52_72 = W*in
   wire signed [9:0] m52_72;
   assign m52_72 ={ {5{neg52[5]}} , neg52[5:1] };

   // m52_73 = W*in
   wire signed [9:0] m52_73;
   assign m52_73 ={ {5{in52[5]}} , in52[5:1] };

   // m52_74 = W*in
   wire signed [9:0] m52_74;
   assign m52_74 =10'b0;

   // m52_75 = W*in
   wire signed [9:0] m52_75;
   assign m52_75 =10'b0;

   // m52_76 = W*in
   wire signed [9:0] m52_76;
   assign m52_76 =10'b0;

   // m52_77 = W*in
   wire signed [9:0] m52_77;
   assign m52_77 =10'b0;

   // m52_78 = W*in
   wire signed [9:0] m52_78;
   assign m52_78 =10'b0;

   // m52_79 = W*in
   wire signed [9:0] m52_79;
   assign m52_79 =10'b0;

   // m52_80 = W*in
   wire signed [9:0] m52_80;
   assign m52_80 =10'b0;

   // m52_81 = W*in
   wire signed [9:0] m52_81;
   assign m52_81 =10'b0;

   // m52_82 = W*in
   wire signed [9:0] m52_82;
   assign m52_82 =10'b0;

   // m52_83 = W*in
   wire signed [9:0] m52_83;
   assign m52_83 =10'b0;

   // m52_84 = W*in
   wire signed [9:0] m52_84;
   assign m52_84 =10'b0;

   // m52_85 = W*in
   wire signed [9:0] m52_85;
   assign m52_85 =10'b0;

   // m52_86 = W*in
   wire signed [9:0] m52_86;
   assign m52_86 =10'b0;

   // m52_87 = W*in
   wire signed [9:0] m52_87;
   assign m52_87 =10'b0;

   // m52_88 = W*in
   wire signed [9:0] m52_88;
   assign m52_88 =10'b0;

   // m52_89 = W*in
   wire signed [9:0] m52_89;
   assign m52_89 =10'b0;

   // m52_90 = W*in
   wire signed [9:0] m52_90;
   assign m52_90 =10'b0;

   // m52_91 = W*in
   wire signed [9:0] m52_91;
   assign m52_91 =10'b0;

   // m52_92 = W*in
   wire signed [9:0] m52_92;
   assign m52_92 =10'b0;

   // m52_93 = W*in
   wire signed [9:0] m52_93;
   assign m52_93 =10'b0;

   // m52_94 = W*in
   wire signed [9:0] m52_94;
   assign m52_94 =10'b0;

   // m52_95 = W*in
   wire signed [9:0] m52_95;
   assign m52_95 =10'b0;

   // m52_96 = W*in
   wire signed [9:0] m52_96;
   assign m52_96 =10'b0;

   // m52_97 = W*in
   wire signed [9:0] m52_97;
   assign m52_97 =10'b0;

   // m52_98 = W*in
   wire signed [9:0] m52_98;
   assign m52_98 =10'b0;

   // m52_99 = W*in
   wire signed [9:0] m52_99;
   assign m52_99 ={ {4{neg52[5]}} , neg52[5:0] };

   // m52_100 = W*in
   wire signed [9:0] m52_100;
   assign m52_100 =10'b0;

   // m52_101 = W*in
   wire signed [9:0] m52_101;
   assign m52_101 =10'b0;

   // m52_102 = W*in
   wire signed [9:0] m52_102;
   assign m52_102 =10'b0;

   // m52_103 = W*in
   wire signed [9:0] m52_103;
   assign m52_103 =10'b0;

   // m52_104 = W*in
   wire signed [9:0] m52_104;
   assign m52_104 =10'b0;

   // m52_105 = W*in
   wire signed [9:0] m52_105;
   assign m52_105 =10'b0;

   // m52_106 = W*in
   wire signed [9:0] m52_106;
   assign m52_106 =10'b0;

   // m52_107 = W*in
   wire signed [9:0] m52_107;
   assign m52_107 =10'b0;

   // m52_108 = W*in
   wire signed [9:0] m52_108;
   assign m52_108 =10'b0;

   // m52_109 = W*in
   wire signed [9:0] m52_109;
   assign m52_109 =10'b0;

   // m52_110 = W*in
   wire signed [9:0] m52_110;
   assign m52_110 =10'b0;

   // m52_111 = W*in
   wire signed [9:0] m52_111;
   assign m52_111 =10'b0;

   // m52_112 = W*in
   wire signed [9:0] m52_112;
   assign m52_112 =10'b0;

   // m52_113 = W*in
   wire signed [9:0] m52_113;
   assign m52_113 =10'b0;

   // m52_114 = W*in
   wire signed [9:0] m52_114;
   assign m52_114 =10'b0;

   // m52_115 = W*in
   wire signed [9:0] m52_115;
   assign m52_115 =10'b0;

   // m52_116 = W*in
   wire signed [9:0] m52_116;
   assign m52_116 =10'b0;

   // m52_117 = W*in
   wire signed [9:0] m52_117;
   assign m52_117 =10'b0;

   // m53_1 = W*in
   wire signed [9:0] m53_1;
   assign m53_1 =10'b0;

   // m53_2 = W*in
   wire signed [9:0] m53_2;
   assign m53_2 =10'b0;

   // m53_3 = W*in
   wire signed [9:0] m53_3;
   assign m53_3 =10'b0;

   // m53_4 = W*in
   wire signed [9:0] m53_4;
   assign m53_4 =10'b0;

   // m53_5 = W*in
   wire signed [9:0] m53_5;
   assign m53_5 =10'b0;

   // m53_6 = W*in
   wire signed [9:0] m53_6;
   assign m53_6 =10'b0;

   // m53_7 = W*in
   wire signed [9:0] m53_7;
   assign m53_7 =10'b0;

   // m53_8 = W*in
   wire signed [9:0] m53_8;
   assign m53_8 =10'b0;

   // m53_9 = W*in
   wire signed [9:0] m53_9;
   assign m53_9 =10'b0;

   // m53_10 = W*in
   wire signed [9:0] m53_10;
   assign m53_10 =10'b0;

   // m53_11 = W*in
   wire signed [9:0] m53_11;
   assign m53_11 =10'b0;

   // m53_12 = W*in
   wire signed [9:0] m53_12;
   assign m53_12 =10'b0;

   // m53_13 = W*in
   wire signed [9:0] m53_13;
   assign m53_13 ={ {4{in53[5]}} , in53[5:0] };

   // m53_14 = W*in
   wire signed [9:0] m53_14;
   assign m53_14 =10'b0;

   // m53_15 = W*in
   wire signed [9:0] m53_15;
   assign m53_15 =10'b0;

   // m53_16 = W*in
   wire signed [9:0] m53_16;
   assign m53_16 =10'b0;

   // m53_17 = W*in
   wire signed [9:0] m53_17;
   assign m53_17 =10'b0;

   // m53_18 = W*in
   wire signed [9:0] m53_18;
   assign m53_18 =10'b0;

   // m53_19 = W*in
   wire signed [9:0] m53_19;
   assign m53_19 =10'b0;

   // m53_20 = W*in
   wire signed [9:0] m53_20;
   assign m53_20 =10'b0;

   // m53_21 = W*in
   wire signed [9:0] m53_21;
   assign m53_21 ={ {5{neg53[5]}} , neg53[5:1] };

   // m53_22 = W*in
   wire signed [9:0] m53_22;
   assign m53_22 =10'b0;

   // m53_23 = W*in
   wire signed [9:0] m53_23;
   assign m53_23 =10'b0;

   // m53_24 = W*in
   wire signed [9:0] m53_24;
   assign m53_24 =10'b0;

   // m53_25 = W*in
   wire signed [9:0] m53_25;
   assign m53_25 =10'b0;

   // m53_26 = W*in
   wire signed [9:0] m53_26;
   assign m53_26 =10'b0;

   // m53_27 = W*in
   wire signed [9:0] m53_27;
   assign m53_27 =10'b0;

   // m53_28 = W*in
   wire signed [9:0] m53_28;
   assign m53_28 =10'b0;

   // m53_29 = W*in
   wire signed [9:0] m53_29;
   assign m53_29 ={ {5{in53[5]}} , in53[5:1] };

   // m53_30 = W*in
   wire signed [9:0] m53_30;
   assign m53_30 =10'b0;

   // m53_31 = W*in
   wire signed [9:0] m53_31;
   assign m53_31 =10'b0;

   // m53_32 = W*in
   wire signed [9:0] m53_32;
   assign m53_32 =10'b0;

   // m53_33 = W*in
   wire signed [9:0] m53_33;
   assign m53_33 =10'b0;

   // m53_34 = W*in
   wire signed [9:0] m53_34;
   assign m53_34 =10'b0;

   // m53_35 = W*in
   wire signed [9:0] m53_35;
   assign m53_35 ={ {4{neg53[5]}} , neg53[5:0] };

   // m53_36 = W*in
   wire signed [9:0] m53_36;
   assign m53_36 =10'b0;

   // m53_37 = W*in
   wire signed [9:0] m53_37;
   assign m53_37 =10'b0;

   // m53_38 = W*in
   wire signed [9:0] m53_38;
   assign m53_38 =10'b0;

   // m53_39 = W*in
   wire signed [9:0] m53_39;
   assign m53_39 =10'b0;

   // m53_40 = W*in
   wire signed [9:0] m53_40;
   assign m53_40 =10'b0;

   // m53_41 = W*in
   wire signed [9:0] m53_41;
   assign m53_41 =10'b0;

   // m53_42 = W*in
   wire signed [9:0] m53_42;
   assign m53_42 =10'b0;

   // m53_43 = W*in
   wire signed [9:0] m53_43;
   assign m53_43 =10'b0;

   // m53_44 = W*in
   wire signed [9:0] m53_44;
   assign m53_44 =10'b0;

   // m53_45 = W*in
   wire signed [9:0] m53_45;
   assign m53_45 =10'b0;

   // m53_46 = W*in
   wire signed [9:0] m53_46;
   assign m53_46 =10'b0;

   // m53_47 = W*in
   wire signed [9:0] m53_47;
   assign m53_47 =10'b0;

   // m53_48 = W*in
   wire signed [9:0] m53_48;
   assign m53_48 =10'b0;

   // m53_49 = W*in
   wire signed [9:0] m53_49;
   assign m53_49 =10'b0;

   // m53_50 = W*in
   wire signed [9:0] m53_50;
   assign m53_50 =10'b0;

   // m53_51 = W*in
   wire signed [9:0] m53_51;
   assign m53_51 =10'b0;

   // m53_52 = W*in
   wire signed [9:0] m53_52;
   assign m53_52 =10'b0;

   // m53_53 = W*in
   wire signed [9:0] m53_53;
   assign m53_53 =10'b0;

   // m53_54 = W*in
   wire signed [9:0] m53_54;
   assign m53_54 =10'b0;

   // m53_55 = W*in
   wire signed [9:0] m53_55;
   assign m53_55 =10'b0;

   // m53_56 = W*in
   wire signed [9:0] m53_56;
   assign m53_56 =10'b0;

   // m53_57 = W*in
   wire signed [9:0] m53_57;
   assign m53_57 =10'b0;

   // m53_58 = W*in
   wire signed [9:0] m53_58;
   assign m53_58 =10'b0;

   // m53_59 = W*in
   wire signed [9:0] m53_59;
   assign m53_59 =10'b0;

   // m53_60 = W*in
   wire signed [9:0] m53_60;
   assign m53_60 =10'b0;

   // m53_61 = W*in
   wire signed [9:0] m53_61;
   assign m53_61 =10'b0;

   // m53_62 = W*in
   wire signed [9:0] m53_62;
   assign m53_62 =10'b0;

   // m53_63 = W*in
   wire signed [9:0] m53_63;
   assign m53_63 =10'b0;

   // m53_64 = W*in
   wire signed [9:0] m53_64;
   assign m53_64 =10'b0;

   // m53_65 = W*in
   wire signed [9:0] m53_65;
   assign m53_65 =10'b0;

   // m53_66 = W*in
   wire signed [9:0] m53_66;
   assign m53_66 =10'b0;

   // m53_67 = W*in
   wire signed [9:0] m53_67;
   assign m53_67 =10'b0;

   // m53_68 = W*in
   wire signed [9:0] m53_68;
   assign m53_68 =10'b0;

   // m53_69 = W*in
   wire signed [9:0] m53_69;
   assign m53_69 ={ {4{neg53[5]}} , neg53[5:0] };

   // m53_70 = W*in
   wire signed [9:0] m53_70;
   assign m53_70 =10'b0;

   // m53_71 = W*in
   wire signed [9:0] m53_71;
   assign m53_71 =10'b0;

   // m53_72 = W*in
   wire signed [9:0] m53_72;
   assign m53_72 ={ {5{neg53[5]}} , neg53[5:1] };

   // m53_73 = W*in
   wire signed [9:0] m53_73;
   assign m53_73 =10'b0;

   // m53_74 = W*in
   wire signed [9:0] m53_74;
   assign m53_74 ={ {5{neg53[5]}} , neg53[5:1] };

   // m53_75 = W*in
   wire signed [9:0] m53_75;
   assign m53_75 =10'b0;

   // m53_76 = W*in
   wire signed [9:0] m53_76;
   assign m53_76 =10'b0;

   // m53_77 = W*in
   wire signed [9:0] m53_77;
   assign m53_77 =10'b0;

   // m53_78 = W*in
   wire signed [9:0] m53_78;
   assign m53_78 =10'b0;

   // m53_79 = W*in
   wire signed [9:0] m53_79;
   assign m53_79 =10'b0;

   // m53_80 = W*in
   wire signed [9:0] m53_80;
   assign m53_80 =10'b0;

   // m53_81 = W*in
   wire signed [9:0] m53_81;
   assign m53_81 =10'b0;

   // m53_82 = W*in
   wire signed [9:0] m53_82;
   assign m53_82 ={ {5{neg53[5]}} , neg53[5:1] };

   // m53_83 = W*in
   wire signed [9:0] m53_83;
   assign m53_83 =10'b0;

   // m53_84 = W*in
   wire signed [9:0] m53_84;
   assign m53_84 =10'b0;

   // m53_85 = W*in
   wire signed [9:0] m53_85;
   assign m53_85 =10'b0;

   // m53_86 = W*in
   wire signed [9:0] m53_86;
   assign m53_86 =10'b0;

   // m53_87 = W*in
   wire signed [9:0] m53_87;
   assign m53_87 =10'b0;

   // m53_88 = W*in
   wire signed [9:0] m53_88;
   assign m53_88 =10'b0;

   // m53_89 = W*in
   wire signed [9:0] m53_89;
   assign m53_89 =10'b0;

   // m53_90 = W*in
   wire signed [9:0] m53_90;
   assign m53_90 =10'b0;

   // m53_91 = W*in
   wire signed [9:0] m53_91;
   assign m53_91 ={ {4{neg53[5]}} , neg53[5:0] };

   // m53_92 = W*in
   wire signed [9:0] m53_92;
   assign m53_92 =10'b0;

   // m53_93 = W*in
   wire signed [9:0] m53_93;
   assign m53_93 =10'b0;

   // m53_94 = W*in
   wire signed [9:0] m53_94;
   assign m53_94 =10'b0;

   // m53_95 = W*in
   wire signed [9:0] m53_95;
   assign m53_95 =10'b0;

   // m53_96 = W*in
   wire signed [9:0] m53_96;
   assign m53_96 =10'b0;

   // m53_97 = W*in
   wire signed [9:0] m53_97;
   assign m53_97 =10'b0;

   // m53_98 = W*in
   wire signed [9:0] m53_98;
   assign m53_98 =10'b0;

   // m53_99 = W*in
   wire signed [9:0] m53_99;
   assign m53_99 =10'b0;

   // m53_100 = W*in
   wire signed [9:0] m53_100;
   assign m53_100 =10'b0;

   // m53_101 = W*in
   wire signed [9:0] m53_101;
   assign m53_101 =10'b0;

   // m53_102 = W*in
   wire signed [9:0] m53_102;
   assign m53_102 =10'b0;

   // m53_103 = W*in
   wire signed [9:0] m53_103;
   assign m53_103 =10'b0;

   // m53_104 = W*in
   wire signed [9:0] m53_104;
   assign m53_104 =10'b0;

   // m53_105 = W*in
   wire signed [9:0] m53_105;
   assign m53_105 =10'b0;

   // m53_106 = W*in
   wire signed [9:0] m53_106;
   assign m53_106 =10'b0;

   // m53_107 = W*in
   wire signed [9:0] m53_107;
   assign m53_107 =10'b0;

   // m53_108 = W*in
   wire signed [9:0] m53_108;
   assign m53_108 =10'b0;

   // m53_109 = W*in
   wire signed [9:0] m53_109;
   assign m53_109 =10'b0;

   // m53_110 = W*in
   wire signed [9:0] m53_110;
   assign m53_110 =10'b0;

   // m53_111 = W*in
   wire signed [9:0] m53_111;
   assign m53_111 =10'b0;

   // m53_112 = W*in
   wire signed [9:0] m53_112;
   assign m53_112 =10'b0;

   // m53_113 = W*in
   wire signed [9:0] m53_113;
   assign m53_113 =10'b0;

   // m53_114 = W*in
   wire signed [9:0] m53_114;
   assign m53_114 =10'b0;

   // m53_115 = W*in
   wire signed [9:0] m53_115;
   assign m53_115 =10'b0;

   // m53_116 = W*in
   wire signed [9:0] m53_116;
   assign m53_116 =10'b0;

   // m53_117 = W*in
   wire signed [9:0] m53_117;
   assign m53_117 =10'b0;

   // m54_1 = W*in
   wire signed [9:0] m54_1;
   assign m54_1 =10'b0;

   // m54_2 = W*in
   wire signed [9:0] m54_2;
   assign m54_2 =10'b0;

   // m54_3 = W*in
   wire signed [9:0] m54_3;
   assign m54_3 =10'b0;

   // m54_4 = W*in
   wire signed [9:0] m54_4;
   assign m54_4 =10'b0;

   // m54_5 = W*in
   wire signed [9:0] m54_5;
   assign m54_5 =10'b0;

   // m54_6 = W*in
   wire signed [9:0] m54_6;
   assign m54_6 =10'b0;

   // m54_7 = W*in
   wire signed [9:0] m54_7;
   assign m54_7 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_8 = W*in
   wire signed [9:0] m54_8;
   assign m54_8 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_9 = W*in
   wire signed [9:0] m54_9;
   assign m54_9 =10'b0;

   // m54_10 = W*in
   wire signed [9:0] m54_10;
   assign m54_10 =10'b0;

   // m54_11 = W*in
   wire signed [9:0] m54_11;
   assign m54_11 ={ {4{in54[5]}} , in54[5:0] };

   // m54_12 = W*in
   wire signed [9:0] m54_12;
   assign m54_12 =10'b0;

   // m54_13 = W*in
   wire signed [9:0] m54_13;
   assign m54_13 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_14 = W*in
   wire signed [9:0] m54_14;
   assign m54_14 =10'b0;

   // m54_15 = W*in
   wire signed [9:0] m54_15;
   assign m54_15 =10'b0;

   // m54_16 = W*in
   wire signed [9:0] m54_16;
   assign m54_16 =10'b0;

   // m54_17 = W*in
   wire signed [9:0] m54_17;
   assign m54_17 ={ {5{neg54[5]}} , neg54[5:1] };

   // m54_18 = W*in
   wire signed [9:0] m54_18;
   assign m54_18 =10'b0;

   // m54_19 = W*in
   wire signed [9:0] m54_19;
   assign m54_19 ={ {5{neg54[5]}} , neg54[5:1] };

   // m54_20 = W*in
   wire signed [9:0] m54_20;
   assign m54_20 =10'b0;

   // m54_21 = W*in
   wire signed [9:0] m54_21;
   assign m54_21 =10'b0;

   // m54_22 = W*in
   wire signed [9:0] m54_22;
   assign m54_22 =10'b0;

   // m54_23 = W*in
   wire signed [9:0] m54_23;
   assign m54_23 =10'b0;

   // m54_24 = W*in
   wire signed [9:0] m54_24;
   assign m54_24 ={ {4{in54[5]}} , in54[5:0] };

   // m54_25 = W*in
   wire signed [9:0] m54_25;
   assign m54_25 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_26 = W*in
   wire signed [9:0] m54_26;
   assign m54_26 ={ {4{in54[5]}} , in54[5:0] };

   // m54_27 = W*in
   wire signed [9:0] m54_27;
   assign m54_27 =10'b0;

   // m54_28 = W*in
   wire signed [9:0] m54_28;
   assign m54_28 =10'b0;

   // m54_29 = W*in
   wire signed [9:0] m54_29;
   assign m54_29 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_30 = W*in
   wire signed [9:0] m54_30;
   assign m54_30 ={ {5{neg54[5]}} , neg54[5:1] };

   // m54_31 = W*in
   wire signed [9:0] m54_31;
   assign m54_31 ={ {5{neg54[5]}} , neg54[5:1] };

   // m54_32 = W*in
   wire signed [9:0] m54_32;
   assign m54_32 =10'b0;

   // m54_33 = W*in
   wire signed [9:0] m54_33;
   assign m54_33 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_34 = W*in
   wire signed [9:0] m54_34;
   assign m54_34 =10'b0;

   // m54_35 = W*in
   wire signed [9:0] m54_35;
   assign m54_35 =10'b0;

   // m54_36 = W*in
   wire signed [9:0] m54_36;
   assign m54_36 ={ {5{neg54[5]}} , neg54[5:1] };

   // m54_37 = W*in
   wire signed [9:0] m54_37;
   assign m54_37 =10'b0;

   // m54_38 = W*in
   wire signed [9:0] m54_38;
   assign m54_38 =10'b0;

   // m54_39 = W*in
   wire signed [9:0] m54_39;
   assign m54_39 =10'b0;

   // m54_40 = W*in
   wire signed [9:0] m54_40;
   assign m54_40 =10'b0;

   // m54_41 = W*in
   wire signed [9:0] m54_41;
   assign m54_41 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_42 = W*in
   wire signed [9:0] m54_42;
   assign m54_42 =10'b0;

   // m54_43 = W*in
   wire signed [9:0] m54_43;
   assign m54_43 =10'b0;

   // m54_44 = W*in
   wire signed [9:0] m54_44;
   assign m54_44 =10'b0;

   // m54_45 = W*in
   wire signed [9:0] m54_45;
   assign m54_45 =10'b0;

   // m54_46 = W*in
   wire signed [9:0] m54_46;
   assign m54_46 =10'b0;

   // m54_47 = W*in
   wire signed [9:0] m54_47;
   assign m54_47 =10'b0;

   // m54_48 = W*in
   wire signed [9:0] m54_48;
   assign m54_48 ={ {4{in54[5]}} , in54[5:0] };

   // m54_49 = W*in
   wire signed [9:0] m54_49;
   assign m54_49 =10'b0;

   // m54_50 = W*in
   wire signed [9:0] m54_50;
   assign m54_50 =10'b0;

   // m54_51 = W*in
   wire signed [9:0] m54_51;
   assign m54_51 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_52 = W*in
   wire signed [9:0] m54_52;
   assign m54_52 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_53 = W*in
   wire signed [9:0] m54_53;
   assign m54_53 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_54 = W*in
   wire signed [9:0] m54_54;
   assign m54_54 =10'b0;

   // m54_55 = W*in
   wire signed [9:0] m54_55;
   assign m54_55 =10'b0;

   // m54_56 = W*in
   wire signed [9:0] m54_56;
   assign m54_56 =10'b0;

   // m54_57 = W*in
   wire signed [9:0] m54_57;
   assign m54_57 =10'b0;

   // m54_58 = W*in
   wire signed [9:0] m54_58;
   assign m54_58 =10'b0;

   // m54_59 = W*in
   wire signed [9:0] m54_59;
   assign m54_59 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_60 = W*in
   wire signed [9:0] m54_60;
   assign m54_60 ={ {4{in54[5]}} , in54[5:0] };

   // m54_61 = W*in
   wire signed [9:0] m54_61;
   assign m54_61 =10'b0;

   // m54_62 = W*in
   wire signed [9:0] m54_62;
   assign m54_62 =10'b0;

   // m54_63 = W*in
   wire signed [9:0] m54_63;
   assign m54_63 =10'b0;

   // m54_64 = W*in
   wire signed [9:0] m54_64;
   assign m54_64 =10'b0;

   // m54_65 = W*in
   wire signed [9:0] m54_65;
   assign m54_65 =10'b0;

   // m54_66 = W*in
   wire signed [9:0] m54_66;
   assign m54_66 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_67 = W*in
   wire signed [9:0] m54_67;
   assign m54_67 =10'b0;

   // m54_68 = W*in
   wire signed [9:0] m54_68;
   assign m54_68 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_69 = W*in
   wire signed [9:0] m54_69;
   assign m54_69 =10'b0;

   // m54_70 = W*in
   wire signed [9:0] m54_70;
   assign m54_70 =10'b0;

   // m54_71 = W*in
   wire signed [9:0] m54_71;
   assign m54_71 ={ {4{in54[5]}} , in54[5:0] };

   // m54_72 = W*in
   wire signed [9:0] m54_72;
   assign m54_72 ={ {4{in54[5]}} , in54[5:0] };

   // m54_73 = W*in
   wire signed [9:0] m54_73;
   assign m54_73 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_74 = W*in
   wire signed [9:0] m54_74;
   assign m54_74 ={ {5{in54[5]}} , in54[5:1] };

   // m54_75 = W*in
   wire signed [9:0] m54_75;
   assign m54_75 ={ {5{neg54[5]}} , neg54[5:1] };

   // m54_76 = W*in
   wire signed [9:0] m54_76;
   assign m54_76 ={ {4{in54[5]}} , in54[5:0] };

   // m54_77 = W*in
   wire signed [9:0] m54_77;
   assign m54_77 ={ {4{in54[5]}} , in54[5:0] };

   // m54_78 = W*in
   wire signed [9:0] m54_78;
   assign m54_78 =10'b0;

   // m54_79 = W*in
   wire signed [9:0] m54_79;
   assign m54_79 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_80 = W*in
   wire signed [9:0] m54_80;
   assign m54_80 =10'b0;

   // m54_81 = W*in
   wire signed [9:0] m54_81;
   assign m54_81 =10'b0;

   // m54_82 = W*in
   wire signed [9:0] m54_82;
   assign m54_82 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_83 = W*in
   wire signed [9:0] m54_83;
   assign m54_83 ={ {4{in54[5]}} , in54[5:0] };

   // m54_84 = W*in
   wire signed [9:0] m54_84;
   assign m54_84 =10'b0;

   // m54_85 = W*in
   wire signed [9:0] m54_85;
   assign m54_85 =10'b0;

   // m54_86 = W*in
   wire signed [9:0] m54_86;
   assign m54_86 =10'b0;

   // m54_87 = W*in
   wire signed [9:0] m54_87;
   assign m54_87 ={ {4{in54[5]}} , in54[5:0] };

   // m54_88 = W*in
   wire signed [9:0] m54_88;
   assign m54_88 =10'b0;

   // m54_89 = W*in
   wire signed [9:0] m54_89;
   assign m54_89 =10'b0;

   // m54_90 = W*in
   wire signed [9:0] m54_90;
   assign m54_90 =10'b0;

   // m54_91 = W*in
   wire signed [9:0] m54_91;
   assign m54_91 =10'b0;

   // m54_92 = W*in
   wire signed [9:0] m54_92;
   assign m54_92 =10'b0;

   // m54_93 = W*in
   wire signed [9:0] m54_93;
   assign m54_93 =10'b0;

   // m54_94 = W*in
   wire signed [9:0] m54_94;
   assign m54_94 =10'b0;

   // m54_95 = W*in
   wire signed [9:0] m54_95;
   assign m54_95 =10'b0;

   // m54_96 = W*in
   wire signed [9:0] m54_96;
   assign m54_96 =10'b0;

   // m54_97 = W*in
   wire signed [9:0] m54_97;
   assign m54_97 =10'b0;

   // m54_98 = W*in
   wire signed [9:0] m54_98;
   assign m54_98 =10'b0;

   // m54_99 = W*in
   wire signed [9:0] m54_99;
   assign m54_99 ={ {4{in54[5]}} , in54[5:0] };

   // m54_100 = W*in
   wire signed [9:0] m54_100;
   assign m54_100 =10'b0;

   // m54_101 = W*in
   wire signed [9:0] m54_101;
   assign m54_101 =10'b0;

   // m54_102 = W*in
   wire signed [9:0] m54_102;
   assign m54_102 =10'b0;

   // m54_103 = W*in
   wire signed [9:0] m54_103;
   assign m54_103 =10'b0;

   // m54_104 = W*in
   wire signed [9:0] m54_104;
   assign m54_104 =10'b0;

   // m54_105 = W*in
   wire signed [9:0] m54_105;
   assign m54_105 =10'b0;

   // m54_106 = W*in
   wire signed [9:0] m54_106;
   assign m54_106 =10'b0;

   // m54_107 = W*in
   wire signed [9:0] m54_107;
   assign m54_107 =10'b0;

   // m54_108 = W*in
   wire signed [9:0] m54_108;
   assign m54_108 =10'b0;

   // m54_109 = W*in
   wire signed [9:0] m54_109;
   assign m54_109 =10'b0;

   // m54_110 = W*in
   wire signed [9:0] m54_110;
   assign m54_110 ={ {4{in54[5]}} , in54[5:0] };

   // m54_111 = W*in
   wire signed [9:0] m54_111;
   assign m54_111 =10'b0;

   // m54_112 = W*in
   wire signed [9:0] m54_112;
   assign m54_112 ={ {4{in54[5]}} , in54[5:0] };

   // m54_113 = W*in
   wire signed [9:0] m54_113;
   assign m54_113 =10'b0;

   // m54_114 = W*in
   wire signed [9:0] m54_114;
   assign m54_114 =10'b0;

   // m54_115 = W*in
   wire signed [9:0] m54_115;
   assign m54_115 =10'b0;

   // m54_116 = W*in
   wire signed [9:0] m54_116;
   assign m54_116 ={ {4{neg54[5]}} , neg54[5:0] };

   // m54_117 = W*in
   wire signed [9:0] m54_117;
   assign m54_117 =10'b0;

   // m55_1 = W*in
   wire signed [9:0] m55_1;
   assign m55_1 =10'b0;

   // m55_2 = W*in
   wire signed [9:0] m55_2;
   assign m55_2 =10'b0;

   // m55_3 = W*in
   wire signed [9:0] m55_3;
   assign m55_3 =10'b0;

   // m55_4 = W*in
   wire signed [9:0] m55_4;
   assign m55_4 =10'b0;

   // m55_5 = W*in
   wire signed [9:0] m55_5;
   assign m55_5 =10'b0;

   // m55_6 = W*in
   wire signed [9:0] m55_6;
   assign m55_6 =10'b0;

   // m55_7 = W*in
   wire signed [9:0] m55_7;
   assign m55_7 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_8 = W*in
   wire signed [9:0] m55_8;
   assign m55_8 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_9 = W*in
   wire signed [9:0] m55_9;
   assign m55_9 =10'b0;

   // m55_10 = W*in
   wire signed [9:0] m55_10;
   assign m55_10 =10'b0;

   // m55_11 = W*in
   wire signed [9:0] m55_11;
   assign m55_11 =10'b0;

   // m55_12 = W*in
   wire signed [9:0] m55_12;
   assign m55_12 =10'b0;

   // m55_13 = W*in
   wire signed [9:0] m55_13;
   assign m55_13 =10'b0;

   // m55_14 = W*in
   wire signed [9:0] m55_14;
   assign m55_14 =10'b0;

   // m55_15 = W*in
   wire signed [9:0] m55_15;
   assign m55_15 =10'b0;

   // m55_16 = W*in
   wire signed [9:0] m55_16;
   assign m55_16 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_17 = W*in
   wire signed [9:0] m55_17;
   assign m55_17 ={ {5{neg55[5]}} , neg55[5:1] };

   // m55_18 = W*in
   wire signed [9:0] m55_18;
   assign m55_18 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_19 = W*in
   wire signed [9:0] m55_19;
   assign m55_19 =10'b0;

   // m55_20 = W*in
   wire signed [9:0] m55_20;
   assign m55_20 ={ {5{in55[5]}} , in55[5:1] };

   // m55_21 = W*in
   wire signed [9:0] m55_21;
   assign m55_21 ={ {5{neg55[5]}} , neg55[5:1] };

   // m55_22 = W*in
   wire signed [9:0] m55_22;
   assign m55_22 =10'b0;

   // m55_23 = W*in
   wire signed [9:0] m55_23;
   assign m55_23 ={ {4{in55[5]}} , in55[5:0] };

   // m55_24 = W*in
   wire signed [9:0] m55_24;
   assign m55_24 =10'b0;

   // m55_25 = W*in
   wire signed [9:0] m55_25;
   assign m55_25 ={ {4{in55[5]}} , in55[5:0] };

   // m55_26 = W*in
   wire signed [9:0] m55_26;
   assign m55_26 =10'b0;

   // m55_27 = W*in
   wire signed [9:0] m55_27;
   assign m55_27 ={ {4{in55[5]}} , in55[5:0] };

   // m55_28 = W*in
   wire signed [9:0] m55_28;
   assign m55_28 ={ {4{in55[5]}} , in55[5:0] };

   // m55_29 = W*in
   wire signed [9:0] m55_29;
   assign m55_29 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_30 = W*in
   wire signed [9:0] m55_30;
   assign m55_30 =10'b0;

   // m55_31 = W*in
   wire signed [9:0] m55_31;
   assign m55_31 =10'b0;

   // m55_32 = W*in
   wire signed [9:0] m55_32;
   assign m55_32 =10'b0;

   // m55_33 = W*in
   wire signed [9:0] m55_33;
   assign m55_33 =10'b0;

   // m55_34 = W*in
   wire signed [9:0] m55_34;
   assign m55_34 =10'b0;

   // m55_35 = W*in
   wire signed [9:0] m55_35;
   assign m55_35 ={ {5{in55[5]}} , in55[5:1] };

   // m55_36 = W*in
   wire signed [9:0] m55_36;
   assign m55_36 =10'b0;

   // m55_37 = W*in
   wire signed [9:0] m55_37;
   assign m55_37 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_38 = W*in
   wire signed [9:0] m55_38;
   assign m55_38 =10'b0;

   // m55_39 = W*in
   wire signed [9:0] m55_39;
   assign m55_39 ={ {4{in55[5]}} , in55[5:0] };

   // m55_40 = W*in
   wire signed [9:0] m55_40;
   assign m55_40 =10'b0;

   // m55_41 = W*in
   wire signed [9:0] m55_41;
   assign m55_41 =10'b0;

   // m55_42 = W*in
   wire signed [9:0] m55_42;
   assign m55_42 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_43 = W*in
   wire signed [9:0] m55_43;
   assign m55_43 =10'b0;

   // m55_44 = W*in
   wire signed [9:0] m55_44;
   assign m55_44 =10'b0;

   // m55_45 = W*in
   wire signed [9:0] m55_45;
   assign m55_45 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_46 = W*in
   wire signed [9:0] m55_46;
   assign m55_46 ={ {4{in55[5]}} , in55[5:0] };

   // m55_47 = W*in
   wire signed [9:0] m55_47;
   assign m55_47 =10'b0;

   // m55_48 = W*in
   wire signed [9:0] m55_48;
   assign m55_48 =10'b0;

   // m55_49 = W*in
   wire signed [9:0] m55_49;
   assign m55_49 =10'b0;

   // m55_50 = W*in
   wire signed [9:0] m55_50;
   assign m55_50 =10'b0;

   // m55_51 = W*in
   wire signed [9:0] m55_51;
   assign m55_51 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_52 = W*in
   wire signed [9:0] m55_52;
   assign m55_52 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_53 = W*in
   wire signed [9:0] m55_53;
   assign m55_53 =10'b0;

   // m55_54 = W*in
   wire signed [9:0] m55_54;
   assign m55_54 =10'b0;

   // m55_55 = W*in
   wire signed [9:0] m55_55;
   assign m55_55 =10'b0;

   // m55_56 = W*in
   wire signed [9:0] m55_56;
   assign m55_56 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_57 = W*in
   wire signed [9:0] m55_57;
   assign m55_57 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_58 = W*in
   wire signed [9:0] m55_58;
   assign m55_58 ={ {4{in55[5]}} , in55[5:0] };

   // m55_59 = W*in
   wire signed [9:0] m55_59;
   assign m55_59 =10'b0;

   // m55_60 = W*in
   wire signed [9:0] m55_60;
   assign m55_60 =10'b0;

   // m55_61 = W*in
   wire signed [9:0] m55_61;
   assign m55_61 ={ {5{in55[5]}} , in55[5:1] };

   // m55_62 = W*in
   wire signed [9:0] m55_62;
   assign m55_62 =10'b0;

   // m55_63 = W*in
   wire signed [9:0] m55_63;
   assign m55_63 ={ {4{in55[5]}} , in55[5:0] };

   // m55_64 = W*in
   wire signed [9:0] m55_64;
   assign m55_64 =10'b0;

   // m55_65 = W*in
   wire signed [9:0] m55_65;
   assign m55_65 =10'b0;

   // m55_66 = W*in
   wire signed [9:0] m55_66;
   assign m55_66 =10'b0;

   // m55_67 = W*in
   wire signed [9:0] m55_67;
   assign m55_67 =10'b0;

   // m55_68 = W*in
   wire signed [9:0] m55_68;
   assign m55_68 =10'b0;

   // m55_69 = W*in
   wire signed [9:0] m55_69;
   assign m55_69 ={ {5{neg55[5]}} , neg55[5:1] };

   // m55_70 = W*in
   wire signed [9:0] m55_70;
   assign m55_70 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_71 = W*in
   wire signed [9:0] m55_71;
   assign m55_71 ={ {5{in55[5]}} , in55[5:1] };

   // m55_72 = W*in
   wire signed [9:0] m55_72;
   assign m55_72 =10'b0;

   // m55_73 = W*in
   wire signed [9:0] m55_73;
   assign m55_73 =10'b0;

   // m55_74 = W*in
   wire signed [9:0] m55_74;
   assign m55_74 =10'b0;

   // m55_75 = W*in
   wire signed [9:0] m55_75;
   assign m55_75 =10'b0;

   // m55_76 = W*in
   wire signed [9:0] m55_76;
   assign m55_76 =10'b0;

   // m55_77 = W*in
   wire signed [9:0] m55_77;
   assign m55_77 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_78 = W*in
   wire signed [9:0] m55_78;
   assign m55_78 =10'b0;

   // m55_79 = W*in
   wire signed [9:0] m55_79;
   assign m55_79 =10'b0;

   // m55_80 = W*in
   wire signed [9:0] m55_80;
   assign m55_80 =10'b0;

   // m55_81 = W*in
   wire signed [9:0] m55_81;
   assign m55_81 =10'b0;

   // m55_82 = W*in
   wire signed [9:0] m55_82;
   assign m55_82 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_83 = W*in
   wire signed [9:0] m55_83;
   assign m55_83 =10'b0;

   // m55_84 = W*in
   wire signed [9:0] m55_84;
   assign m55_84 =10'b0;

   // m55_85 = W*in
   wire signed [9:0] m55_85;
   assign m55_85 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_86 = W*in
   wire signed [9:0] m55_86;
   assign m55_86 =10'b0;

   // m55_87 = W*in
   wire signed [9:0] m55_87;
   assign m55_87 ={ {4{in55[5]}} , in55[5:0] };

   // m55_88 = W*in
   wire signed [9:0] m55_88;
   assign m55_88 =10'b0;

   // m55_89 = W*in
   wire signed [9:0] m55_89;
   assign m55_89 =10'b0;

   // m55_90 = W*in
   wire signed [9:0] m55_90;
   assign m55_90 =10'b0;

   // m55_91 = W*in
   wire signed [9:0] m55_91;
   assign m55_91 =10'b0;

   // m55_92 = W*in
   wire signed [9:0] m55_92;
   assign m55_92 =10'b0;

   // m55_93 = W*in
   wire signed [9:0] m55_93;
   assign m55_93 =10'b0;

   // m55_94 = W*in
   wire signed [9:0] m55_94;
   assign m55_94 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_95 = W*in
   wire signed [9:0] m55_95;
   assign m55_95 =10'b0;

   // m55_96 = W*in
   wire signed [9:0] m55_96;
   assign m55_96 =10'b0;

   // m55_97 = W*in
   wire signed [9:0] m55_97;
   assign m55_97 =10'b0;

   // m55_98 = W*in
   wire signed [9:0] m55_98;
   assign m55_98 =10'b0;

   // m55_99 = W*in
   wire signed [9:0] m55_99;
   assign m55_99 =10'b0;

   // m55_100 = W*in
   wire signed [9:0] m55_100;
   assign m55_100 =10'b0;

   // m55_101 = W*in
   wire signed [9:0] m55_101;
   assign m55_101 ={ {5{in55[5]}} , in55[5:1] };

   // m55_102 = W*in
   wire signed [9:0] m55_102;
   assign m55_102 ={ {5{neg55[5]}} , neg55[5:1] };

   // m55_103 = W*in
   wire signed [9:0] m55_103;
   assign m55_103 =10'b0;

   // m55_104 = W*in
   wire signed [9:0] m55_104;
   assign m55_104 =10'b0;

   // m55_105 = W*in
   wire signed [9:0] m55_105;
   assign m55_105 ={ {4{in55[5]}} , in55[5:0] };

   // m55_106 = W*in
   wire signed [9:0] m55_106;
   assign m55_106 ={ {5{neg55[5]}} , neg55[5:1] };

   // m55_107 = W*in
   wire signed [9:0] m55_107;
   assign m55_107 =10'b0;

   // m55_108 = W*in
   wire signed [9:0] m55_108;
   assign m55_108 =10'b0;

   // m55_109 = W*in
   wire signed [9:0] m55_109;
   assign m55_109 =10'b0;

   // m55_110 = W*in
   wire signed [9:0] m55_110;
   assign m55_110 =10'b0;

   // m55_111 = W*in
   wire signed [9:0] m55_111;
   assign m55_111 =10'b0;

   // m55_112 = W*in
   wire signed [9:0] m55_112;
   assign m55_112 ={ {4{neg55[5]}} , neg55[5:0] };

   // m55_113 = W*in
   wire signed [9:0] m55_113;
   assign m55_113 =10'b0;

   // m55_114 = W*in
   wire signed [9:0] m55_114;
   assign m55_114 =10'b0;

   // m55_115 = W*in
   wire signed [9:0] m55_115;
   assign m55_115 =10'b0;

   // m55_116 = W*in
   wire signed [9:0] m55_116;
   assign m55_116 =10'b0;

   // m55_117 = W*in
   wire signed [9:0] m55_117;
   assign m55_117 ={ {4{in55[5]}} , in55[5:0] };

   // m56_1 = W*in
   wire signed [9:0] m56_1;
   assign m56_1 =10'b0;

   // m56_2 = W*in
   wire signed [9:0] m56_2;
   assign m56_2 ={ {4{in56[5]}} , in56[5:0] };

   // m56_3 = W*in
   wire signed [9:0] m56_3;
   assign m56_3 =10'b0;

   // m56_4 = W*in
   wire signed [9:0] m56_4;
   assign m56_4 =10'b0;

   // m56_5 = W*in
   wire signed [9:0] m56_5;
   assign m56_5 =10'b0;

   // m56_6 = W*in
   wire signed [9:0] m56_6;
   assign m56_6 =10'b0;

   // m56_7 = W*in
   wire signed [9:0] m56_7;
   assign m56_7 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_8 = W*in
   wire signed [9:0] m56_8;
   assign m56_8 =10'b0;

   // m56_9 = W*in
   wire signed [9:0] m56_9;
   assign m56_9 =10'b0;

   // m56_10 = W*in
   wire signed [9:0] m56_10;
   assign m56_10 =10'b0;

   // m56_11 = W*in
   wire signed [9:0] m56_11;
   assign m56_11 =10'b0;

   // m56_12 = W*in
   wire signed [9:0] m56_12;
   assign m56_12 =10'b0;

   // m56_13 = W*in
   wire signed [9:0] m56_13;
   assign m56_13 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_14 = W*in
   wire signed [9:0] m56_14;
   assign m56_14 =10'b0;

   // m56_15 = W*in
   wire signed [9:0] m56_15;
   assign m56_15 ={ {4{in56[5]}} , in56[5:0] };

   // m56_16 = W*in
   wire signed [9:0] m56_16;
   assign m56_16 =10'b0;

   // m56_17 = W*in
   wire signed [9:0] m56_17;
   assign m56_17 =10'b0;

   // m56_18 = W*in
   wire signed [9:0] m56_18;
   assign m56_18 =10'b0;

   // m56_19 = W*in
   wire signed [9:0] m56_19;
   assign m56_19 =10'b0;

   // m56_20 = W*in
   wire signed [9:0] m56_20;
   assign m56_20 ={ {4{in56[5]}} , in56[5:0] };

   // m56_21 = W*in
   wire signed [9:0] m56_21;
   assign m56_21 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_22 = W*in
   wire signed [9:0] m56_22;
   assign m56_22 ={ {4{in56[5]}} , in56[5:0] };

   // m56_23 = W*in
   wire signed [9:0] m56_23;
   assign m56_23 =10'b0;

   // m56_24 = W*in
   wire signed [9:0] m56_24;
   assign m56_24 ={ {4{in56[5]}} , in56[5:0] };

   // m56_25 = W*in
   wire signed [9:0] m56_25;
   assign m56_25 =10'b0;

   // m56_26 = W*in
   wire signed [9:0] m56_26;
   assign m56_26 =10'b0;

   // m56_27 = W*in
   wire signed [9:0] m56_27;
   assign m56_27 =10'b0;

   // m56_28 = W*in
   wire signed [9:0] m56_28;
   assign m56_28 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_29 = W*in
   wire signed [9:0] m56_29;
   assign m56_29 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_30 = W*in
   wire signed [9:0] m56_30;
   assign m56_30 =10'b0;

   // m56_31 = W*in
   wire signed [9:0] m56_31;
   assign m56_31 =10'b0;

   // m56_32 = W*in
   wire signed [9:0] m56_32;
   assign m56_32 =10'b0;

   // m56_33 = W*in
   wire signed [9:0] m56_33;
   assign m56_33 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_34 = W*in
   wire signed [9:0] m56_34;
   assign m56_34 ={ {4{in56[5]}} , in56[5:0] };

   // m56_35 = W*in
   wire signed [9:0] m56_35;
   assign m56_35 ={ {4{in56[5]}} , in56[5:0] };

   // m56_36 = W*in
   wire signed [9:0] m56_36;
   assign m56_36 ={ {5{neg56[5]}} , neg56[5:1] };

   // m56_37 = W*in
   wire signed [9:0] m56_37;
   assign m56_37 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_38 = W*in
   wire signed [9:0] m56_38;
   assign m56_38 =10'b0;

   // m56_39 = W*in
   wire signed [9:0] m56_39;
   assign m56_39 =10'b0;

   // m56_40 = W*in
   wire signed [9:0] m56_40;
   assign m56_40 =10'b0;

   // m56_41 = W*in
   wire signed [9:0] m56_41;
   assign m56_41 =10'b0;

   // m56_42 = W*in
   wire signed [9:0] m56_42;
   assign m56_42 ={ {4{in56[5]}} , in56[5:0] };

   // m56_43 = W*in
   wire signed [9:0] m56_43;
   assign m56_43 =10'b0;

   // m56_44 = W*in
   wire signed [9:0] m56_44;
   assign m56_44 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_45 = W*in
   wire signed [9:0] m56_45;
   assign m56_45 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_46 = W*in
   wire signed [9:0] m56_46;
   assign m56_46 =10'b0;

   // m56_47 = W*in
   wire signed [9:0] m56_47;
   assign m56_47 =10'b0;

   // m56_48 = W*in
   wire signed [9:0] m56_48;
   assign m56_48 =10'b0;

   // m56_49 = W*in
   wire signed [9:0] m56_49;
   assign m56_49 =10'b0;

   // m56_50 = W*in
   wire signed [9:0] m56_50;
   assign m56_50 =10'b0;

   // m56_51 = W*in
   wire signed [9:0] m56_51;
   assign m56_51 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_52 = W*in
   wire signed [9:0] m56_52;
   assign m56_52 =10'b0;

   // m56_53 = W*in
   wire signed [9:0] m56_53;
   assign m56_53 =10'b0;

   // m56_54 = W*in
   wire signed [9:0] m56_54;
   assign m56_54 =10'b0;

   // m56_55 = W*in
   wire signed [9:0] m56_55;
   assign m56_55 =10'b0;

   // m56_56 = W*in
   wire signed [9:0] m56_56;
   assign m56_56 =10'b0;

   // m56_57 = W*in
   wire signed [9:0] m56_57;
   assign m56_57 =10'b0;

   // m56_58 = W*in
   wire signed [9:0] m56_58;
   assign m56_58 =10'b0;

   // m56_59 = W*in
   wire signed [9:0] m56_59;
   assign m56_59 =10'b0;

   // m56_60 = W*in
   wire signed [9:0] m56_60;
   assign m56_60 ={ {4{in56[5]}} , in56[5:0] };

   // m56_61 = W*in
   wire signed [9:0] m56_61;
   assign m56_61 =10'b0;

   // m56_62 = W*in
   wire signed [9:0] m56_62;
   assign m56_62 =10'b0;

   // m56_63 = W*in
   wire signed [9:0] m56_63;
   assign m56_63 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_64 = W*in
   wire signed [9:0] m56_64;
   assign m56_64 ={ {4{in56[5]}} , in56[5:0] };

   // m56_65 = W*in
   wire signed [9:0] m56_65;
   assign m56_65 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_66 = W*in
   wire signed [9:0] m56_66;
   assign m56_66 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_67 = W*in
   wire signed [9:0] m56_67;
   assign m56_67 =10'b0;

   // m56_68 = W*in
   wire signed [9:0] m56_68;
   assign m56_68 =10'b0;

   // m56_69 = W*in
   wire signed [9:0] m56_69;
   assign m56_69 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_70 = W*in
   wire signed [9:0] m56_70;
   assign m56_70 =10'b0;

   // m56_71 = W*in
   wire signed [9:0] m56_71;
   assign m56_71 =10'b0;

   // m56_72 = W*in
   wire signed [9:0] m56_72;
   assign m56_72 ={ {5{in56[5]}} , in56[5:1] };

   // m56_73 = W*in
   wire signed [9:0] m56_73;
   assign m56_73 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_74 = W*in
   wire signed [9:0] m56_74;
   assign m56_74 ={ {4{in56[5]}} , in56[5:0] };

   // m56_75 = W*in
   wire signed [9:0] m56_75;
   assign m56_75 =10'b0;

   // m56_76 = W*in
   wire signed [9:0] m56_76;
   assign m56_76 =10'b0;

   // m56_77 = W*in
   wire signed [9:0] m56_77;
   assign m56_77 =10'b0;

   // m56_78 = W*in
   wire signed [9:0] m56_78;
   assign m56_78 =10'b0;

   // m56_79 = W*in
   wire signed [9:0] m56_79;
   assign m56_79 =10'b0;

   // m56_80 = W*in
   wire signed [9:0] m56_80;
   assign m56_80 =10'b0;

   // m56_81 = W*in
   wire signed [9:0] m56_81;
   assign m56_81 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m56_82 = W*in
   wire signed [9:0] m56_82;
   assign m56_82 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_83 = W*in
   wire signed [9:0] m56_83;
   assign m56_83 =10'b0;

   // m56_84 = W*in
   wire signed [9:0] m56_84;
   assign m56_84 =10'b0;

   // m56_85 = W*in
   wire signed [9:0] m56_85;
   assign m56_85 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_86 = W*in
   wire signed [9:0] m56_86;
   assign m56_86 =10'b0;

   // m56_87 = W*in
   wire signed [9:0] m56_87;
   assign m56_87 ={ {4{in56[5]}} , in56[5:0] };

   // m56_88 = W*in
   wire signed [9:0] m56_88;
   assign m56_88 ={ {4{in56[5]}} , in56[5:0] };

   // m56_89 = W*in
   wire signed [9:0] m56_89;
   assign m56_89 =10'b0;

   // m56_90 = W*in
   wire signed [9:0] m56_90;
   assign m56_90 ={ {4{in56[5]}} , in56[5:0] };

   // m56_91 = W*in
   wire signed [9:0] m56_91;
   assign m56_91 =10'b0;

   // m56_92 = W*in
   wire signed [9:0] m56_92;
   assign m56_92 =10'b0;

   // m56_93 = W*in
   wire signed [9:0] m56_93;
   assign m56_93 ={ {3{neg56[5]}} , neg56 , {1{1'b0}} };

   // m56_94 = W*in
   wire signed [9:0] m56_94;
   assign m56_94 =10'b0;

   // m56_95 = W*in
   wire signed [9:0] m56_95;
   assign m56_95 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_96 = W*in
   wire signed [9:0] m56_96;
   assign m56_96 =10'b0;

   // m56_97 = W*in
   wire signed [9:0] m56_97;
   assign m56_97 =10'b0;

   // m56_98 = W*in
   wire signed [9:0] m56_98;
   assign m56_98 =10'b0;

   // m56_99 = W*in
   wire signed [9:0] m56_99;
   assign m56_99 =10'b0;

   // m56_100 = W*in
   wire signed [9:0] m56_100;
   assign m56_100 =10'b0;

   // m56_101 = W*in
   wire signed [9:0] m56_101;
   assign m56_101 =10'b0;

   // m56_102 = W*in
   wire signed [9:0] m56_102;
   assign m56_102 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_103 = W*in
   wire signed [9:0] m56_103;
   assign m56_103 =10'b0;

   // m56_104 = W*in
   wire signed [9:0] m56_104;
   assign m56_104 =10'b0;

   // m56_105 = W*in
   wire signed [9:0] m56_105;
   assign m56_105 =10'b0;

   // m56_106 = W*in
   wire signed [9:0] m56_106;
   assign m56_106 =10'b0;

   // m56_107 = W*in
   wire signed [9:0] m56_107;
   assign m56_107 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_108 = W*in
   wire signed [9:0] m56_108;
   assign m56_108 =10'b0;

   // m56_109 = W*in
   wire signed [9:0] m56_109;
   assign m56_109 =10'b0;

   // m56_110 = W*in
   wire signed [9:0] m56_110;
   assign m56_110 =10'b0;

   // m56_111 = W*in
   wire signed [9:0] m56_111;
   assign m56_111 =10'b0;

   // m56_112 = W*in
   wire signed [9:0] m56_112;
   assign m56_112 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_113 = W*in
   wire signed [9:0] m56_113;
   assign m56_113 =10'b0;

   // m56_114 = W*in
   wire signed [9:0] m56_114;
   assign m56_114 =10'b0;

   // m56_115 = W*in
   wire signed [9:0] m56_115;
   assign m56_115 ={ {4{in56[5]}} , in56[5:0] };

   // m56_116 = W*in
   wire signed [9:0] m56_116;
   assign m56_116 ={ {4{neg56[5]}} , neg56[5:0] };

   // m56_117 = W*in
   wire signed [9:0] m56_117;
   assign m56_117 ={ {3{in56[5]}} , in56 , {1{1'b0}} };

   // m57_1 = W*in
   wire signed [9:0] m57_1;
   assign m57_1 =10'b0;

   // m57_2 = W*in
   wire signed [9:0] m57_2;
   assign m57_2 =10'b0;

   // m57_3 = W*in
   wire signed [9:0] m57_3;
   assign m57_3 =10'b0;

   // m57_4 = W*in
   wire signed [9:0] m57_4;
   assign m57_4 =10'b0;

   // m57_5 = W*in
   wire signed [9:0] m57_5;
   assign m57_5 =10'b0;

   // m57_6 = W*in
   wire signed [9:0] m57_6;
   assign m57_6 =10'b0;

   // m57_7 = W*in
   wire signed [9:0] m57_7;
   assign m57_7 =10'b0;

   // m57_8 = W*in
   wire signed [9:0] m57_8;
   assign m57_8 =10'b0;

   // m57_9 = W*in
   wire signed [9:0] m57_9;
   assign m57_9 =10'b0;

   // m57_10 = W*in
   wire signed [9:0] m57_10;
   assign m57_10 =10'b0;

   // m57_11 = W*in
   wire signed [9:0] m57_11;
   assign m57_11 =10'b0;

   // m57_12 = W*in
   wire signed [9:0] m57_12;
   assign m57_12 =10'b0;

   // m57_13 = W*in
   wire signed [9:0] m57_13;
   assign m57_13 =10'b0;

   // m57_14 = W*in
   wire signed [9:0] m57_14;
   assign m57_14 =10'b0;

   // m57_15 = W*in
   wire signed [9:0] m57_15;
   assign m57_15 =10'b0;

   // m57_16 = W*in
   wire signed [9:0] m57_16;
   assign m57_16 =10'b0;

   // m57_17 = W*in
   wire signed [9:0] m57_17;
   assign m57_17 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_18 = W*in
   wire signed [9:0] m57_18;
   assign m57_18 =10'b0;

   // m57_19 = W*in
   wire signed [9:0] m57_19;
   assign m57_19 =10'b0;

   // m57_20 = W*in
   wire signed [9:0] m57_20;
   assign m57_20 =10'b0;

   // m57_21 = W*in
   wire signed [9:0] m57_21;
   assign m57_21 =10'b0;

   // m57_22 = W*in
   wire signed [9:0] m57_22;
   assign m57_22 =10'b0;

   // m57_23 = W*in
   wire signed [9:0] m57_23;
   assign m57_23 =10'b0;

   // m57_24 = W*in
   wire signed [9:0] m57_24;
   assign m57_24 =10'b0;

   // m57_25 = W*in
   wire signed [9:0] m57_25;
   assign m57_25 =10'b0;

   // m57_26 = W*in
   wire signed [9:0] m57_26;
   assign m57_26 =10'b0;

   // m57_27 = W*in
   wire signed [9:0] m57_27;
   assign m57_27 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_28 = W*in
   wire signed [9:0] m57_28;
   assign m57_28 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_29 = W*in
   wire signed [9:0] m57_29;
   assign m57_29 ={ {4{in57[5]}} , in57[5:0] };

   // m57_30 = W*in
   wire signed [9:0] m57_30;
   assign m57_30 =10'b0;

   // m57_31 = W*in
   wire signed [9:0] m57_31;
   assign m57_31 =10'b0;

   // m57_32 = W*in
   wire signed [9:0] m57_32;
   assign m57_32 =10'b0;

   // m57_33 = W*in
   wire signed [9:0] m57_33;
   assign m57_33 =10'b0;

   // m57_34 = W*in
   wire signed [9:0] m57_34;
   assign m57_34 =10'b0;

   // m57_35 = W*in
   wire signed [9:0] m57_35;
   assign m57_35 =10'b0;

   // m57_36 = W*in
   wire signed [9:0] m57_36;
   assign m57_36 =10'b0;

   // m57_37 = W*in
   wire signed [9:0] m57_37;
   assign m57_37 =10'b0;

   // m57_38 = W*in
   wire signed [9:0] m57_38;
   assign m57_38 =10'b0;

   // m57_39 = W*in
   wire signed [9:0] m57_39;
   assign m57_39 =10'b0;

   // m57_40 = W*in
   wire signed [9:0] m57_40;
   assign m57_40 =10'b0;

   // m57_41 = W*in
   wire signed [9:0] m57_41;
   assign m57_41 =10'b0;

   // m57_42 = W*in
   wire signed [9:0] m57_42;
   assign m57_42 =10'b0;

   // m57_43 = W*in
   wire signed [9:0] m57_43;
   assign m57_43 =10'b0;

   // m57_44 = W*in
   wire signed [9:0] m57_44;
   assign m57_44 =10'b0;

   // m57_45 = W*in
   wire signed [9:0] m57_45;
   assign m57_45 =10'b0;

   // m57_46 = W*in
   wire signed [9:0] m57_46;
   assign m57_46 =10'b0;

   // m57_47 = W*in
   wire signed [9:0] m57_47;
   assign m57_47 =10'b0;

   // m57_48 = W*in
   wire signed [9:0] m57_48;
   assign m57_48 =10'b0;

   // m57_49 = W*in
   wire signed [9:0] m57_49;
   assign m57_49 =10'b0;

   // m57_50 = W*in
   wire signed [9:0] m57_50;
   assign m57_50 =10'b0;

   // m57_51 = W*in
   wire signed [9:0] m57_51;
   assign m57_51 =10'b0;

   // m57_52 = W*in
   wire signed [9:0] m57_52;
   assign m57_52 =10'b0;

   // m57_53 = W*in
   wire signed [9:0] m57_53;
   assign m57_53 =10'b0;

   // m57_54 = W*in
   wire signed [9:0] m57_54;
   assign m57_54 =10'b0;

   // m57_55 = W*in
   wire signed [9:0] m57_55;
   assign m57_55 =10'b0;

   // m57_56 = W*in
   wire signed [9:0] m57_56;
   assign m57_56 =10'b0;

   // m57_57 = W*in
   wire signed [9:0] m57_57;
   assign m57_57 =10'b0;

   // m57_58 = W*in
   wire signed [9:0] m57_58;
   assign m57_58 =10'b0;

   // m57_59 = W*in
   wire signed [9:0] m57_59;
   assign m57_59 =10'b0;

   // m57_60 = W*in
   wire signed [9:0] m57_60;
   assign m57_60 ={ {4{neg57[5]}} , neg57[5:0] };

   // m57_61 = W*in
   wire signed [9:0] m57_61;
   assign m57_61 =10'b0;

   // m57_62 = W*in
   wire signed [9:0] m57_62;
   assign m57_62 =10'b0;

   // m57_63 = W*in
   wire signed [9:0] m57_63;
   assign m57_63 ={ {4{in57[5]}} , in57[5:0] };

   // m57_64 = W*in
   wire signed [9:0] m57_64;
   assign m57_64 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_65 = W*in
   wire signed [9:0] m57_65;
   assign m57_65 =10'b0;

   // m57_66 = W*in
   wire signed [9:0] m57_66;
   assign m57_66 =10'b0;

   // m57_67 = W*in
   wire signed [9:0] m57_67;
   assign m57_67 =10'b0;

   // m57_68 = W*in
   wire signed [9:0] m57_68;
   assign m57_68 =10'b0;

   // m57_69 = W*in
   wire signed [9:0] m57_69;
   assign m57_69 =10'b0;

   // m57_70 = W*in
   wire signed [9:0] m57_70;
   assign m57_70 =10'b0;

   // m57_71 = W*in
   wire signed [9:0] m57_71;
   assign m57_71 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_72 = W*in
   wire signed [9:0] m57_72;
   assign m57_72 =10'b0;

   // m57_73 = W*in
   wire signed [9:0] m57_73;
   assign m57_73 =10'b0;

   // m57_74 = W*in
   wire signed [9:0] m57_74;
   assign m57_74 =10'b0;

   // m57_75 = W*in
   wire signed [9:0] m57_75;
   assign m57_75 =10'b0;

   // m57_76 = W*in
   wire signed [9:0] m57_76;
   assign m57_76 =10'b0;

   // m57_77 = W*in
   wire signed [9:0] m57_77;
   assign m57_77 =10'b0;

   // m57_78 = W*in
   wire signed [9:0] m57_78;
   assign m57_78 =10'b0;

   // m57_79 = W*in
   wire signed [9:0] m57_79;
   assign m57_79 =10'b0;

   // m57_80 = W*in
   wire signed [9:0] m57_80;
   assign m57_80 =10'b0;

   // m57_81 = W*in
   wire signed [9:0] m57_81;
   assign m57_81 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_82 = W*in
   wire signed [9:0] m57_82;
   assign m57_82 =10'b0;

   // m57_83 = W*in
   wire signed [9:0] m57_83;
   assign m57_83 =10'b0;

   // m57_84 = W*in
   wire signed [9:0] m57_84;
   assign m57_84 =10'b0;

   // m57_85 = W*in
   wire signed [9:0] m57_85;
   assign m57_85 ={ {4{in57[5]}} , in57[5:0] };

   // m57_86 = W*in
   wire signed [9:0] m57_86;
   assign m57_86 =10'b0;

   // m57_87 = W*in
   wire signed [9:0] m57_87;
   assign m57_87 =10'b0;

   // m57_88 = W*in
   wire signed [9:0] m57_88;
   assign m57_88 =10'b0;

   // m57_89 = W*in
   wire signed [9:0] m57_89;
   assign m57_89 =10'b0;

   // m57_90 = W*in
   wire signed [9:0] m57_90;
   assign m57_90 =10'b0;

   // m57_91 = W*in
   wire signed [9:0] m57_91;
   assign m57_91 =10'b0;

   // m57_92 = W*in
   wire signed [9:0] m57_92;
   assign m57_92 =10'b0;

   // m57_93 = W*in
   wire signed [9:0] m57_93;
   assign m57_93 =10'b0;

   // m57_94 = W*in
   wire signed [9:0] m57_94;
   assign m57_94 =10'b0;

   // m57_95 = W*in
   wire signed [9:0] m57_95;
   assign m57_95 =10'b0;

   // m57_96 = W*in
   wire signed [9:0] m57_96;
   assign m57_96 =10'b0;

   // m57_97 = W*in
   wire signed [9:0] m57_97;
   assign m57_97 =10'b0;

   // m57_98 = W*in
   wire signed [9:0] m57_98;
   assign m57_98 =10'b0;

   // m57_99 = W*in
   wire signed [9:0] m57_99;
   assign m57_99 =10'b0;

   // m57_100 = W*in
   wire signed [9:0] m57_100;
   assign m57_100 =10'b0;

   // m57_101 = W*in
   wire signed [9:0] m57_101;
   assign m57_101 =10'b0;

   // m57_102 = W*in
   wire signed [9:0] m57_102;
   assign m57_102 =10'b0;

   // m57_103 = W*in
   wire signed [9:0] m57_103;
   assign m57_103 =10'b0;

   // m57_104 = W*in
   wire signed [9:0] m57_104;
   assign m57_104 ={ {4{neg57[5]}} , neg57[5:0] };

   // m57_105 = W*in
   wire signed [9:0] m57_105;
   assign m57_105 =10'b0;

   // m57_106 = W*in
   wire signed [9:0] m57_106;
   assign m57_106 =10'b0;

   // m57_107 = W*in
   wire signed [9:0] m57_107;
   assign m57_107 =10'b0;

   // m57_108 = W*in
   wire signed [9:0] m57_108;
   assign m57_108 =10'b0;

   // m57_109 = W*in
   wire signed [9:0] m57_109;
   assign m57_109 ={ {5{in57[5]}} , in57[5:1] };

   // m57_110 = W*in
   wire signed [9:0] m57_110;
   assign m57_110 =10'b0;

   // m57_111 = W*in
   wire signed [9:0] m57_111;
   assign m57_111 =10'b0;

   // m57_112 = W*in
   wire signed [9:0] m57_112;
   assign m57_112 =10'b0;

   // m57_113 = W*in
   wire signed [9:0] m57_113;
   assign m57_113 =10'b0;

   // m57_114 = W*in
   wire signed [9:0] m57_114;
   assign m57_114 =10'b0;

   // m57_115 = W*in
   wire signed [9:0] m57_115;
   assign m57_115 ={ {5{neg57[5]}} , neg57[5:1] };

   // m57_116 = W*in
   wire signed [9:0] m57_116;
   assign m57_116 ={ {4{in57[5]}} , in57[5:0] };

   // m57_117 = W*in
   wire signed [9:0] m57_117;
   assign m57_117 =10'b0;

   // m58_1 = W*in
   wire signed [9:0] m58_1;
   assign m58_1 =10'b0;

   // m58_2 = W*in
   wire signed [9:0] m58_2;
   assign m58_2 =10'b0;

   // m58_3 = W*in
   wire signed [9:0] m58_3;
   assign m58_3 =10'b0;

   // m58_4 = W*in
   wire signed [9:0] m58_4;
   assign m58_4 =10'b0;

   // m58_5 = W*in
   wire signed [9:0] m58_5;
   assign m58_5 =10'b0;

   // m58_6 = W*in
   wire signed [9:0] m58_6;
   assign m58_6 =10'b0;

   // m58_7 = W*in
   wire signed [9:0] m58_7;
   assign m58_7 =10'b0;

   // m58_8 = W*in
   wire signed [9:0] m58_8;
   assign m58_8 =10'b0;

   // m58_9 = W*in
   wire signed [9:0] m58_9;
   assign m58_9 =10'b0;

   // m58_10 = W*in
   wire signed [9:0] m58_10;
   assign m58_10 =10'b0;

   // m58_11 = W*in
   wire signed [9:0] m58_11;
   assign m58_11 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_12 = W*in
   wire signed [9:0] m58_12;
   assign m58_12 ={ {4{in58[5]}} , in58[5:0] };

   // m58_13 = W*in
   wire signed [9:0] m58_13;
   assign m58_13 =10'b0;

   // m58_14 = W*in
   wire signed [9:0] m58_14;
   assign m58_14 =10'b0;

   // m58_15 = W*in
   wire signed [9:0] m58_15;
   assign m58_15 =10'b0;

   // m58_16 = W*in
   wire signed [9:0] m58_16;
   assign m58_16 =10'b0;

   // m58_17 = W*in
   wire signed [9:0] m58_17;
   assign m58_17 ={ {5{neg58[5]}} , neg58[5:1] };

   // m58_18 = W*in
   wire signed [9:0] m58_18;
   assign m58_18 ={ {4{in58[5]}} , in58[5:0] };

   // m58_19 = W*in
   wire signed [9:0] m58_19;
   assign m58_19 ={ {5{neg58[5]}} , neg58[5:1] };

   // m58_20 = W*in
   wire signed [9:0] m58_20;
   assign m58_20 =10'b0;

   // m58_21 = W*in
   wire signed [9:0] m58_21;
   assign m58_21 =10'b0;

   // m58_22 = W*in
   wire signed [9:0] m58_22;
   assign m58_22 =10'b0;

   // m58_23 = W*in
   wire signed [9:0] m58_23;
   assign m58_23 ={ {4{in58[5]}} , in58[5:0] };

   // m58_24 = W*in
   wire signed [9:0] m58_24;
   assign m58_24 =10'b0;

   // m58_25 = W*in
   wire signed [9:0] m58_25;
   assign m58_25 =10'b0;

   // m58_26 = W*in
   wire signed [9:0] m58_26;
   assign m58_26 =10'b0;

   // m58_27 = W*in
   wire signed [9:0] m58_27;
   assign m58_27 =10'b0;

   // m58_28 = W*in
   wire signed [9:0] m58_28;
   assign m58_28 ={ {5{neg58[5]}} , neg58[5:1] };

   // m58_29 = W*in
   wire signed [9:0] m58_29;
   assign m58_29 ={ {4{in58[5]}} , in58[5:0] };

   // m58_30 = W*in
   wire signed [9:0] m58_30;
   assign m58_30 =10'b0;

   // m58_31 = W*in
   wire signed [9:0] m58_31;
   assign m58_31 =10'b0;

   // m58_32 = W*in
   wire signed [9:0] m58_32;
   assign m58_32 =10'b0;

   // m58_33 = W*in
   wire signed [9:0] m58_33;
   assign m58_33 =10'b0;

   // m58_34 = W*in
   wire signed [9:0] m58_34;
   assign m58_34 =10'b0;

   // m58_35 = W*in
   wire signed [9:0] m58_35;
   assign m58_35 =10'b0;

   // m58_36 = W*in
   wire signed [9:0] m58_36;
   assign m58_36 =10'b0;

   // m58_37 = W*in
   wire signed [9:0] m58_37;
   assign m58_37 =10'b0;

   // m58_38 = W*in
   wire signed [9:0] m58_38;
   assign m58_38 =10'b0;

   // m58_39 = W*in
   wire signed [9:0] m58_39;
   assign m58_39 =10'b0;

   // m58_40 = W*in
   wire signed [9:0] m58_40;
   assign m58_40 =10'b0;

   // m58_41 = W*in
   wire signed [9:0] m58_41;
   assign m58_41 =10'b0;

   // m58_42 = W*in
   wire signed [9:0] m58_42;
   assign m58_42 =10'b0;

   // m58_43 = W*in
   wire signed [9:0] m58_43;
   assign m58_43 =10'b0;

   // m58_44 = W*in
   wire signed [9:0] m58_44;
   assign m58_44 =10'b0;

   // m58_45 = W*in
   wire signed [9:0] m58_45;
   assign m58_45 =10'b0;

   // m58_46 = W*in
   wire signed [9:0] m58_46;
   assign m58_46 =10'b0;

   // m58_47 = W*in
   wire signed [9:0] m58_47;
   assign m58_47 =10'b0;

   // m58_48 = W*in
   wire signed [9:0] m58_48;
   assign m58_48 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_49 = W*in
   wire signed [9:0] m58_49;
   assign m58_49 =10'b0;

   // m58_50 = W*in
   wire signed [9:0] m58_50;
   assign m58_50 =10'b0;

   // m58_51 = W*in
   wire signed [9:0] m58_51;
   assign m58_51 =10'b0;

   // m58_52 = W*in
   wire signed [9:0] m58_52;
   assign m58_52 =10'b0;

   // m58_53 = W*in
   wire signed [9:0] m58_53;
   assign m58_53 =10'b0;

   // m58_54 = W*in
   wire signed [9:0] m58_54;
   assign m58_54 =10'b0;

   // m58_55 = W*in
   wire signed [9:0] m58_55;
   assign m58_55 =10'b0;

   // m58_56 = W*in
   wire signed [9:0] m58_56;
   assign m58_56 =10'b0;

   // m58_57 = W*in
   wire signed [9:0] m58_57;
   assign m58_57 =10'b0;

   // m58_58 = W*in
   wire signed [9:0] m58_58;
   assign m58_58 =10'b0;

   // m58_59 = W*in
   wire signed [9:0] m58_59;
   assign m58_59 =10'b0;

   // m58_60 = W*in
   wire signed [9:0] m58_60;
   assign m58_60 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_61 = W*in
   wire signed [9:0] m58_61;
   assign m58_61 =10'b0;

   // m58_62 = W*in
   wire signed [9:0] m58_62;
   assign m58_62 =10'b0;

   // m58_63 = W*in
   wire signed [9:0] m58_63;
   assign m58_63 =10'b0;

   // m58_64 = W*in
   wire signed [9:0] m58_64;
   assign m58_64 ={ {3{in58[5]}} , in58 , {1{1'b0}} };

   // m58_65 = W*in
   wire signed [9:0] m58_65;
   assign m58_65 ={ {5{in58[5]}} , in58[5:1] };

   // m58_66 = W*in
   wire signed [9:0] m58_66;
   assign m58_66 ={ {5{in58[5]}} , in58[5:1] };

   // m58_67 = W*in
   wire signed [9:0] m58_67;
   assign m58_67 =10'b0;

   // m58_68 = W*in
   wire signed [9:0] m58_68;
   assign m58_68 =10'b0;

   // m58_69 = W*in
   wire signed [9:0] m58_69;
   assign m58_69 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_70 = W*in
   wire signed [9:0] m58_70;
   assign m58_70 ={ {4{in58[5]}} , in58[5:0] };

   // m58_71 = W*in
   wire signed [9:0] m58_71;
   assign m58_71 =10'b0;

   // m58_72 = W*in
   wire signed [9:0] m58_72;
   assign m58_72 ={ {5{neg58[5]}} , neg58[5:1] };

   // m58_73 = W*in
   wire signed [9:0] m58_73;
   assign m58_73 =10'b0;

   // m58_74 = W*in
   wire signed [9:0] m58_74;
   assign m58_74 ={ {4{in58[5]}} , in58[5:0] };

   // m58_75 = W*in
   wire signed [9:0] m58_75;
   assign m58_75 =10'b0;

   // m58_76 = W*in
   wire signed [9:0] m58_76;
   assign m58_76 =10'b0;

   // m58_77 = W*in
   wire signed [9:0] m58_77;
   assign m58_77 =10'b0;

   // m58_78 = W*in
   wire signed [9:0] m58_78;
   assign m58_78 =10'b0;

   // m58_79 = W*in
   wire signed [9:0] m58_79;
   assign m58_79 =10'b0;

   // m58_80 = W*in
   wire signed [9:0] m58_80;
   assign m58_80 =10'b0;

   // m58_81 = W*in
   wire signed [9:0] m58_81;
   assign m58_81 ={ {4{in58[5]}} , in58[5:0] };

   // m58_82 = W*in
   wire signed [9:0] m58_82;
   assign m58_82 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_83 = W*in
   wire signed [9:0] m58_83;
   assign m58_83 =10'b0;

   // m58_84 = W*in
   wire signed [9:0] m58_84;
   assign m58_84 =10'b0;

   // m58_85 = W*in
   wire signed [9:0] m58_85;
   assign m58_85 =10'b0;

   // m58_86 = W*in
   wire signed [9:0] m58_86;
   assign m58_86 =10'b0;

   // m58_87 = W*in
   wire signed [9:0] m58_87;
   assign m58_87 =10'b0;

   // m58_88 = W*in
   wire signed [9:0] m58_88;
   assign m58_88 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_89 = W*in
   wire signed [9:0] m58_89;
   assign m58_89 =10'b0;

   // m58_90 = W*in
   wire signed [9:0] m58_90;
   assign m58_90 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_91 = W*in
   wire signed [9:0] m58_91;
   assign m58_91 =10'b0;

   // m58_92 = W*in
   wire signed [9:0] m58_92;
   assign m58_92 =10'b0;

   // m58_93 = W*in
   wire signed [9:0] m58_93;
   assign m58_93 =10'b0;

   // m58_94 = W*in
   wire signed [9:0] m58_94;
   assign m58_94 ={ {4{in58[5]}} , in58[5:0] };

   // m58_95 = W*in
   wire signed [9:0] m58_95;
   assign m58_95 =10'b0;

   // m58_96 = W*in
   wire signed [9:0] m58_96;
   assign m58_96 =10'b0;

   // m58_97 = W*in
   wire signed [9:0] m58_97;
   assign m58_97 =10'b0;

   // m58_98 = W*in
   wire signed [9:0] m58_98;
   assign m58_98 =10'b0;

   // m58_99 = W*in
   wire signed [9:0] m58_99;
   assign m58_99 =10'b0;

   // m58_100 = W*in
   wire signed [9:0] m58_100;
   assign m58_100 =10'b0;

   // m58_101 = W*in
   wire signed [9:0] m58_101;
   assign m58_101 =10'b0;

   // m58_102 = W*in
   wire signed [9:0] m58_102;
   assign m58_102 =10'b0;

   // m58_103 = W*in
   wire signed [9:0] m58_103;
   assign m58_103 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_104 = W*in
   wire signed [9:0] m58_104;
   assign m58_104 =10'b0;

   // m58_105 = W*in
   wire signed [9:0] m58_105;
   assign m58_105 =10'b0;

   // m58_106 = W*in
   wire signed [9:0] m58_106;
   assign m58_106 =10'b0;

   // m58_107 = W*in
   wire signed [9:0] m58_107;
   assign m58_107 =10'b0;

   // m58_108 = W*in
   wire signed [9:0] m58_108;
   assign m58_108 ={ {4{in58[5]}} , in58[5:0] };

   // m58_109 = W*in
   wire signed [9:0] m58_109;
   assign m58_109 ={ {4{in58[5]}} , in58[5:0] };

   // m58_110 = W*in
   wire signed [9:0] m58_110;
   assign m58_110 ={ {4{in58[5]}} , in58[5:0] };

   // m58_111 = W*in
   wire signed [9:0] m58_111;
   assign m58_111 =10'b0;

   // m58_112 = W*in
   wire signed [9:0] m58_112;
   assign m58_112 ={ {4{in58[5]}} , in58[5:0] };

   // m58_113 = W*in
   wire signed [9:0] m58_113;
   assign m58_113 ={ {4{neg58[5]}} , neg58[5:0] };

   // m58_114 = W*in
   wire signed [9:0] m58_114;
   assign m58_114 =10'b0;

   // m58_115 = W*in
   wire signed [9:0] m58_115;
   assign m58_115 ={ {5{neg58[5]}} , neg58[5:1] };

   // m58_116 = W*in
   wire signed [9:0] m58_116;
   assign m58_116 =10'b0;

   // m58_117 = W*in
   wire signed [9:0] m58_117;
   assign m58_117 =10'b0;

   // m59_1 = W*in
   wire signed [9:0] m59_1;
   assign m59_1 =10'b0;

   // m59_2 = W*in
   wire signed [9:0] m59_2;
   assign m59_2 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_3 = W*in
   wire signed [9:0] m59_3;
   assign m59_3 =10'b0;

   // m59_4 = W*in
   wire signed [9:0] m59_4;
   assign m59_4 =10'b0;

   // m59_5 = W*in
   wire signed [9:0] m59_5;
   assign m59_5 =10'b0;

   // m59_6 = W*in
   wire signed [9:0] m59_6;
   assign m59_6 =10'b0;

   // m59_7 = W*in
   wire signed [9:0] m59_7;
   assign m59_7 =10'b0;

   // m59_8 = W*in
   wire signed [9:0] m59_8;
   assign m59_8 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_9 = W*in
   wire signed [9:0] m59_9;
   assign m59_9 =10'b0;

   // m59_10 = W*in
   wire signed [9:0] m59_10;
   assign m59_10 ={ {4{in59[5]}} , in59[5:0] };

   // m59_11 = W*in
   wire signed [9:0] m59_11;
   assign m59_11 =10'b0;

   // m59_12 = W*in
   wire signed [9:0] m59_12;
   assign m59_12 =10'b0;

   // m59_13 = W*in
   wire signed [9:0] m59_13;
   assign m59_13 =10'b0;

   // m59_14 = W*in
   wire signed [9:0] m59_14;
   assign m59_14 =10'b0;

   // m59_15 = W*in
   wire signed [9:0] m59_15;
   assign m59_15 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_16 = W*in
   wire signed [9:0] m59_16;
   assign m59_16 =10'b0;

   // m59_17 = W*in
   wire signed [9:0] m59_17;
   assign m59_17 ={ {5{neg59[5]}} , neg59[5:1] };

   // m59_18 = W*in
   wire signed [9:0] m59_18;
   assign m59_18 ={ {5{neg59[5]}} , neg59[5:1] };

   // m59_19 = W*in
   wire signed [9:0] m59_19;
   assign m59_19 =10'b0;

   // m59_20 = W*in
   wire signed [9:0] m59_20;
   assign m59_20 =10'b0;

   // m59_21 = W*in
   wire signed [9:0] m59_21;
   assign m59_21 =10'b0;

   // m59_22 = W*in
   wire signed [9:0] m59_22;
   assign m59_22 =10'b0;

   // m59_23 = W*in
   wire signed [9:0] m59_23;
   assign m59_23 =10'b0;

   // m59_24 = W*in
   wire signed [9:0] m59_24;
   assign m59_24 =10'b0;

   // m59_25 = W*in
   wire signed [9:0] m59_25;
   assign m59_25 =10'b0;

   // m59_26 = W*in
   wire signed [9:0] m59_26;
   assign m59_26 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_27 = W*in
   wire signed [9:0] m59_27;
   assign m59_27 =10'b0;

   // m59_28 = W*in
   wire signed [9:0] m59_28;
   assign m59_28 =10'b0;

   // m59_29 = W*in
   wire signed [9:0] m59_29;
   assign m59_29 ={ {4{in59[5]}} , in59[5:0] };

   // m59_30 = W*in
   wire signed [9:0] m59_30;
   assign m59_30 =10'b0;

   // m59_31 = W*in
   wire signed [9:0] m59_31;
   assign m59_31 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_32 = W*in
   wire signed [9:0] m59_32;
   assign m59_32 =10'b0;

   // m59_33 = W*in
   wire signed [9:0] m59_33;
   assign m59_33 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_34 = W*in
   wire signed [9:0] m59_34;
   assign m59_34 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_35 = W*in
   wire signed [9:0] m59_35;
   assign m59_35 =10'b0;

   // m59_36 = W*in
   wire signed [9:0] m59_36;
   assign m59_36 =10'b0;

   // m59_37 = W*in
   wire signed [9:0] m59_37;
   assign m59_37 ={ {4{in59[5]}} , in59[5:0] };

   // m59_38 = W*in
   wire signed [9:0] m59_38;
   assign m59_38 =10'b0;

   // m59_39 = W*in
   wire signed [9:0] m59_39;
   assign m59_39 =10'b0;

   // m59_40 = W*in
   wire signed [9:0] m59_40;
   assign m59_40 ={ {5{in59[5]}} , in59[5:1] };

   // m59_41 = W*in
   wire signed [9:0] m59_41;
   assign m59_41 =10'b0;

   // m59_42 = W*in
   wire signed [9:0] m59_42;
   assign m59_42 =10'b0;

   // m59_43 = W*in
   wire signed [9:0] m59_43;
   assign m59_43 =10'b0;

   // m59_44 = W*in
   wire signed [9:0] m59_44;
   assign m59_44 =10'b0;

   // m59_45 = W*in
   wire signed [9:0] m59_45;
   assign m59_45 =10'b0;

   // m59_46 = W*in
   wire signed [9:0] m59_46;
   assign m59_46 =10'b0;

   // m59_47 = W*in
   wire signed [9:0] m59_47;
   assign m59_47 =10'b0;

   // m59_48 = W*in
   wire signed [9:0] m59_48;
   assign m59_48 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_49 = W*in
   wire signed [9:0] m59_49;
   assign m59_49 =10'b0;

   // m59_50 = W*in
   wire signed [9:0] m59_50;
   assign m59_50 =10'b0;

   // m59_51 = W*in
   wire signed [9:0] m59_51;
   assign m59_51 =10'b0;

   // m59_52 = W*in
   wire signed [9:0] m59_52;
   assign m59_52 =10'b0;

   // m59_53 = W*in
   wire signed [9:0] m59_53;
   assign m59_53 =10'b0;

   // m59_54 = W*in
   wire signed [9:0] m59_54;
   assign m59_54 ={ {4{in59[5]}} , in59[5:0] };

   // m59_55 = W*in
   wire signed [9:0] m59_55;
   assign m59_55 =10'b0;

   // m59_56 = W*in
   wire signed [9:0] m59_56;
   assign m59_56 =10'b0;

   // m59_57 = W*in
   wire signed [9:0] m59_57;
   assign m59_57 =10'b0;

   // m59_58 = W*in
   wire signed [9:0] m59_58;
   assign m59_58 =10'b0;

   // m59_59 = W*in
   wire signed [9:0] m59_59;
   assign m59_59 =10'b0;

   // m59_60 = W*in
   wire signed [9:0] m59_60;
   assign m59_60 ={ {4{in59[5]}} , in59[5:0] };

   // m59_61 = W*in
   wire signed [9:0] m59_61;
   assign m59_61 =10'b0;

   // m59_62 = W*in
   wire signed [9:0] m59_62;
   assign m59_62 =10'b0;

   // m59_63 = W*in
   wire signed [9:0] m59_63;
   assign m59_63 =10'b0;

   // m59_64 = W*in
   wire signed [9:0] m59_64;
   assign m59_64 ={ {4{in59[5]}} , in59[5:0] };

   // m59_65 = W*in
   wire signed [9:0] m59_65;
   assign m59_65 ={ {4{in59[5]}} , in59[5:0] };

   // m59_66 = W*in
   wire signed [9:0] m59_66;
   assign m59_66 ={ {4{in59[5]}} , in59[5:0] };

   // m59_67 = W*in
   wire signed [9:0] m59_67;
   assign m59_67 =10'b0;

   // m59_68 = W*in
   wire signed [9:0] m59_68;
   assign m59_68 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_69 = W*in
   wire signed [9:0] m59_69;
   assign m59_69 =10'b0;

   // m59_70 = W*in
   wire signed [9:0] m59_70;
   assign m59_70 ={ {4{in59[5]}} , in59[5:0] };

   // m59_71 = W*in
   wire signed [9:0] m59_71;
   assign m59_71 =10'b0;

   // m59_72 = W*in
   wire signed [9:0] m59_72;
   assign m59_72 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_73 = W*in
   wire signed [9:0] m59_73;
   assign m59_73 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_74 = W*in
   wire signed [9:0] m59_74;
   assign m59_74 =10'b0;

   // m59_75 = W*in
   wire signed [9:0] m59_75;
   assign m59_75 =10'b0;

   // m59_76 = W*in
   wire signed [9:0] m59_76;
   assign m59_76 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_77 = W*in
   wire signed [9:0] m59_77;
   assign m59_77 =10'b0;

   // m59_78 = W*in
   wire signed [9:0] m59_78;
   assign m59_78 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_79 = W*in
   wire signed [9:0] m59_79;
   assign m59_79 ={ {4{in59[5]}} , in59[5:0] };

   // m59_80 = W*in
   wire signed [9:0] m59_80;
   assign m59_80 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_81 = W*in
   wire signed [9:0] m59_81;
   assign m59_81 =10'b0;

   // m59_82 = W*in
   wire signed [9:0] m59_82;
   assign m59_82 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_83 = W*in
   wire signed [9:0] m59_83;
   assign m59_83 ={ {4{in59[5]}} , in59[5:0] };

   // m59_84 = W*in
   wire signed [9:0] m59_84;
   assign m59_84 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_85 = W*in
   wire signed [9:0] m59_85;
   assign m59_85 ={ {4{in59[5]}} , in59[5:0] };

   // m59_86 = W*in
   wire signed [9:0] m59_86;
   assign m59_86 =10'b0;

   // m59_87 = W*in
   wire signed [9:0] m59_87;
   assign m59_87 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_88 = W*in
   wire signed [9:0] m59_88;
   assign m59_88 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_89 = W*in
   wire signed [9:0] m59_89;
   assign m59_89 =10'b0;

   // m59_90 = W*in
   wire signed [9:0] m59_90;
   assign m59_90 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_91 = W*in
   wire signed [9:0] m59_91;
   assign m59_91 =10'b0;

   // m59_92 = W*in
   wire signed [9:0] m59_92;
   assign m59_92 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_93 = W*in
   wire signed [9:0] m59_93;
   assign m59_93 =10'b0;

   // m59_94 = W*in
   wire signed [9:0] m59_94;
   assign m59_94 ={ {4{in59[5]}} , in59[5:0] };

   // m59_95 = W*in
   wire signed [9:0] m59_95;
   assign m59_95 ={ {4{in59[5]}} , in59[5:0] };

   // m59_96 = W*in
   wire signed [9:0] m59_96;
   assign m59_96 =10'b0;

   // m59_97 = W*in
   wire signed [9:0] m59_97;
   assign m59_97 =10'b0;

   // m59_98 = W*in
   wire signed [9:0] m59_98;
   assign m59_98 =10'b0;

   // m59_99 = W*in
   wire signed [9:0] m59_99;
   assign m59_99 =10'b0;

   // m59_100 = W*in
   wire signed [9:0] m59_100;
   assign m59_100 ={ {4{in59[5]}} , in59[5:0] };

   // m59_101 = W*in
   wire signed [9:0] m59_101;
   assign m59_101 =10'b0;

   // m59_102 = W*in
   wire signed [9:0] m59_102;
   assign m59_102 =10'b0;

   // m59_103 = W*in
   wire signed [9:0] m59_103;
   assign m59_103 =10'b0;

   // m59_104 = W*in
   wire signed [9:0] m59_104;
   assign m59_104 =10'b0;

   // m59_105 = W*in
   wire signed [9:0] m59_105;
   assign m59_105 =10'b0;

   // m59_106 = W*in
   wire signed [9:0] m59_106;
   assign m59_106 =10'b0;

   // m59_107 = W*in
   wire signed [9:0] m59_107;
   assign m59_107 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_108 = W*in
   wire signed [9:0] m59_108;
   assign m59_108 ={ {4{in59[5]}} , in59[5:0] };

   // m59_109 = W*in
   wire signed [9:0] m59_109;
   assign m59_109 ={ {5{in59[5]}} , in59[5:1] };

   // m59_110 = W*in
   wire signed [9:0] m59_110;
   assign m59_110 =10'b0;

   // m59_111 = W*in
   wire signed [9:0] m59_111;
   assign m59_111 ={ {4{neg59[5]}} , neg59[5:0] };

   // m59_112 = W*in
   wire signed [9:0] m59_112;
   assign m59_112 ={ {4{in59[5]}} , in59[5:0] };

   // m59_113 = W*in
   wire signed [9:0] m59_113;
   assign m59_113 =10'b0;

   // m59_114 = W*in
   wire signed [9:0] m59_114;
   assign m59_114 =10'b0;

   // m59_115 = W*in
   wire signed [9:0] m59_115;
   assign m59_115 =10'b0;

   // m59_116 = W*in
   wire signed [9:0] m59_116;
   assign m59_116 ={ {5{in59[5]}} , in59[5:1] };

   // m59_117 = W*in
   wire signed [9:0] m59_117;
   assign m59_117 =10'b0;

   // m60_1 = W*in
   wire signed [9:0] m60_1;
   assign m60_1 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_2 = W*in
   wire signed [9:0] m60_2;
   assign m60_2 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_3 = W*in
   wire signed [9:0] m60_3;
   assign m60_3 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_4 = W*in
   wire signed [9:0] m60_4;
   assign m60_4 =10'b0;

   // m60_5 = W*in
   wire signed [9:0] m60_5;
   assign m60_5 =10'b0;

   // m60_6 = W*in
   wire signed [9:0] m60_6;
   assign m60_6 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_7 = W*in
   wire signed [9:0] m60_7;
   assign m60_7 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_8 = W*in
   wire signed [9:0] m60_8;
   assign m60_8 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_9 = W*in
   wire signed [9:0] m60_9;
   assign m60_9 =10'b0;

   // m60_10 = W*in
   wire signed [9:0] m60_10;
   assign m60_10 ={ {4{in60[5]}} , in60[5:0] };

   // m60_11 = W*in
   wire signed [9:0] m60_11;
   assign m60_11 =10'b0;

   // m60_12 = W*in
   wire signed [9:0] m60_12;
   assign m60_12 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_13 = W*in
   wire signed [9:0] m60_13;
   assign m60_13 =10'b0;

   // m60_14 = W*in
   wire signed [9:0] m60_14;
   assign m60_14 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_15 = W*in
   wire signed [9:0] m60_15;
   assign m60_15 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_16 = W*in
   wire signed [9:0] m60_16;
   assign m60_16 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_17 = W*in
   wire signed [9:0] m60_17;
   assign m60_17 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_18 = W*in
   wire signed [9:0] m60_18;
   assign m60_18 =10'b0;

   // m60_19 = W*in
   wire signed [9:0] m60_19;
   assign m60_19 ={ {4{in60[5]}} , in60[5:0] };

   // m60_20 = W*in
   wire signed [9:0] m60_20;
   assign m60_20 =10'b0;

   // m60_21 = W*in
   wire signed [9:0] m60_21;
   assign m60_21 ={ {4{in60[5]}} , in60[5:0] };

   // m60_22 = W*in
   wire signed [9:0] m60_22;
   assign m60_22 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_23 = W*in
   wire signed [9:0] m60_23;
   assign m60_23 =10'b0;

   // m60_24 = W*in
   wire signed [9:0] m60_24;
   assign m60_24 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_25 = W*in
   wire signed [9:0] m60_25;
   assign m60_25 =10'b0;

   // m60_26 = W*in
   wire signed [9:0] m60_26;
   assign m60_26 ={ {5{neg60[5]}} , neg60[5:1] };

   // m60_27 = W*in
   wire signed [9:0] m60_27;
   assign m60_27 =10'b0;

   // m60_28 = W*in
   wire signed [9:0] m60_28;
   assign m60_28 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_29 = W*in
   wire signed [9:0] m60_29;
   assign m60_29 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_30 = W*in
   wire signed [9:0] m60_30;
   assign m60_30 ={ {5{in60[5]}} , in60[5:1] };

   // m60_31 = W*in
   wire signed [9:0] m60_31;
   assign m60_31 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_32 = W*in
   wire signed [9:0] m60_32;
   assign m60_32 =10'b0;

   // m60_33 = W*in
   wire signed [9:0] m60_33;
   assign m60_33 =10'b0;

   // m60_34 = W*in
   wire signed [9:0] m60_34;
   assign m60_34 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_35 = W*in
   wire signed [9:0] m60_35;
   assign m60_35 =10'b0;

   // m60_36 = W*in
   wire signed [9:0] m60_36;
   assign m60_36 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_37 = W*in
   wire signed [9:0] m60_37;
   assign m60_37 =10'b0;

   // m60_38 = W*in
   wire signed [9:0] m60_38;
   assign m60_38 =10'b0;

   // m60_39 = W*in
   wire signed [9:0] m60_39;
   assign m60_39 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_40 = W*in
   wire signed [9:0] m60_40;
   assign m60_40 =10'b0;

   // m60_41 = W*in
   wire signed [9:0] m60_41;
   assign m60_41 ={ {4{in60[5]}} , in60[5:0] };

   // m60_42 = W*in
   wire signed [9:0] m60_42;
   assign m60_42 ={ {4{in60[5]}} , in60[5:0] };

   // m60_43 = W*in
   wire signed [9:0] m60_43;
   assign m60_43 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_44 = W*in
   wire signed [9:0] m60_44;
   assign m60_44 ={ {4{in60[5]}} , in60[5:0] };

   // m60_45 = W*in
   wire signed [9:0] m60_45;
   assign m60_45 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_46 = W*in
   wire signed [9:0] m60_46;
   assign m60_46 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_47 = W*in
   wire signed [9:0] m60_47;
   assign m60_47 =10'b0;

   // m60_48 = W*in
   wire signed [9:0] m60_48;
   assign m60_48 =10'b0;

   // m60_49 = W*in
   wire signed [9:0] m60_49;
   assign m60_49 =10'b0;

   // m60_50 = W*in
   wire signed [9:0] m60_50;
   assign m60_50 =10'b0;

   // m60_51 = W*in
   wire signed [9:0] m60_51;
   assign m60_51 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_52 = W*in
   wire signed [9:0] m60_52;
   assign m60_52 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_53 = W*in
   wire signed [9:0] m60_53;
   assign m60_53 =10'b0;

   // m60_54 = W*in
   wire signed [9:0] m60_54;
   assign m60_54 =10'b0;

   // m60_55 = W*in
   wire signed [9:0] m60_55;
   assign m60_55 =10'b0;

   // m60_56 = W*in
   wire signed [9:0] m60_56;
   assign m60_56 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_57 = W*in
   wire signed [9:0] m60_57;
   assign m60_57 =10'b0;

   // m60_58 = W*in
   wire signed [9:0] m60_58;
   assign m60_58 =10'b0;

   // m60_59 = W*in
   wire signed [9:0] m60_59;
   assign m60_59 =10'b0;

   // m60_60 = W*in
   wire signed [9:0] m60_60;
   assign m60_60 =10'b0;

   // m60_61 = W*in
   wire signed [9:0] m60_61;
   assign m60_61 =10'b0;

   // m60_62 = W*in
   wire signed [9:0] m60_62;
   assign m60_62 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_63 = W*in
   wire signed [9:0] m60_63;
   assign m60_63 =10'b0;

   // m60_64 = W*in
   wire signed [9:0] m60_64;
   assign m60_64 ={ {4{in60[5]}} , in60[5:0] };

   // m60_65 = W*in
   wire signed [9:0] m60_65;
   assign m60_65 =10'b0;

   // m60_66 = W*in
   wire signed [9:0] m60_66;
   assign m60_66 =10'b0;

   // m60_67 = W*in
   wire signed [9:0] m60_67;
   assign m60_67 ={ {4{in60[5]}} , in60[5:0] };

   // m60_68 = W*in
   wire signed [9:0] m60_68;
   assign m60_68 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_69 = W*in
   wire signed [9:0] m60_69;
   assign m60_69 ={ {4{in60[5]}} , in60[5:0] };

   // m60_70 = W*in
   wire signed [9:0] m60_70;
   assign m60_70 ={ {4{in60[5]}} , in60[5:0] };

   // m60_71 = W*in
   wire signed [9:0] m60_71;
   assign m60_71 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_72 = W*in
   wire signed [9:0] m60_72;
   assign m60_72 ={ {5{neg60[5]}} , neg60[5:1] };

   // m60_73 = W*in
   wire signed [9:0] m60_73;
   assign m60_73 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_74 = W*in
   wire signed [9:0] m60_74;
   assign m60_74 =10'b0;

   // m60_75 = W*in
   wire signed [9:0] m60_75;
   assign m60_75 ={ {4{in60[5]}} , in60[5:0] };

   // m60_76 = W*in
   wire signed [9:0] m60_76;
   assign m60_76 =10'b0;

   // m60_77 = W*in
   wire signed [9:0] m60_77;
   assign m60_77 =10'b0;

   // m60_78 = W*in
   wire signed [9:0] m60_78;
   assign m60_78 =10'b0;

   // m60_79 = W*in
   wire signed [9:0] m60_79;
   assign m60_79 ={ {3{in60[5]}} , in60 , {1{1'b0}} };

   // m60_80 = W*in
   wire signed [9:0] m60_80;
   assign m60_80 =10'b0;

   // m60_81 = W*in
   wire signed [9:0] m60_81;
   assign m60_81 ={ {4{in60[5]}} , in60[5:0] };

   // m60_82 = W*in
   wire signed [9:0] m60_82;
   assign m60_82 =10'b0;

   // m60_83 = W*in
   wire signed [9:0] m60_83;
   assign m60_83 =10'b0;

   // m60_84 = W*in
   wire signed [9:0] m60_84;
   assign m60_84 =10'b0;

   // m60_85 = W*in
   wire signed [9:0] m60_85;
   assign m60_85 ={ {4{in60[5]}} , in60[5:0] };

   // m60_86 = W*in
   wire signed [9:0] m60_86;
   assign m60_86 =10'b0;

   // m60_87 = W*in
   wire signed [9:0] m60_87;
   assign m60_87 =10'b0;

   // m60_88 = W*in
   wire signed [9:0] m60_88;
   assign m60_88 =10'b0;

   // m60_89 = W*in
   wire signed [9:0] m60_89;
   assign m60_89 =10'b0;

   // m60_90 = W*in
   wire signed [9:0] m60_90;
   assign m60_90 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_91 = W*in
   wire signed [9:0] m60_91;
   assign m60_91 ={ {4{in60[5]}} , in60[5:0] };

   // m60_92 = W*in
   wire signed [9:0] m60_92;
   assign m60_92 =10'b0;

   // m60_93 = W*in
   wire signed [9:0] m60_93;
   assign m60_93 =10'b0;

   // m60_94 = W*in
   wire signed [9:0] m60_94;
   assign m60_94 =10'b0;

   // m60_95 = W*in
   wire signed [9:0] m60_95;
   assign m60_95 =10'b0;

   // m60_96 = W*in
   wire signed [9:0] m60_96;
   assign m60_96 =10'b0;

   // m60_97 = W*in
   wire signed [9:0] m60_97;
   assign m60_97 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_98 = W*in
   wire signed [9:0] m60_98;
   assign m60_98 =10'b0;

   // m60_99 = W*in
   wire signed [9:0] m60_99;
   assign m60_99 =10'b0;

   // m60_100 = W*in
   wire signed [9:0] m60_100;
   assign m60_100 =10'b0;

   // m60_101 = W*in
   wire signed [9:0] m60_101;
   assign m60_101 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_102 = W*in
   wire signed [9:0] m60_102;
   assign m60_102 =10'b0;

   // m60_103 = W*in
   wire signed [9:0] m60_103;
   assign m60_103 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_104 = W*in
   wire signed [9:0] m60_104;
   assign m60_104 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_105 = W*in
   wire signed [9:0] m60_105;
   assign m60_105 =10'b0;

   // m60_106 = W*in
   wire signed [9:0] m60_106;
   assign m60_106 =10'b0;

   // m60_107 = W*in
   wire signed [9:0] m60_107;
   assign m60_107 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_108 = W*in
   wire signed [9:0] m60_108;
   assign m60_108 ={ {4{in60[5]}} , in60[5:0] };

   // m60_109 = W*in
   wire signed [9:0] m60_109;
   assign m60_109 =10'b0;

   // m60_110 = W*in
   wire signed [9:0] m60_110;
   assign m60_110 ={ {5{neg60[5]}} , neg60[5:1] };

   // m60_111 = W*in
   wire signed [9:0] m60_111;
   assign m60_111 =10'b0;

   // m60_112 = W*in
   wire signed [9:0] m60_112;
   assign m60_112 =10'b0;

   // m60_113 = W*in
   wire signed [9:0] m60_113;
   assign m60_113 =10'b0;

   // m60_114 = W*in
   wire signed [9:0] m60_114;
   assign m60_114 ={ {4{neg60[5]}} , neg60[5:0] };

   // m60_115 = W*in
   wire signed [9:0] m60_115;
   assign m60_115 =10'b0;

   // m60_116 = W*in
   wire signed [9:0] m60_116;
   assign m60_116 ={ {4{in60[5]}} , in60[5:0] };

   // m60_117 = W*in
   wire signed [9:0] m60_117;
   assign m60_117 ={ {5{neg60[5]}} , neg60[5:1] };

   // m61_1 = W*in
   wire signed [9:0] m61_1;
   assign m61_1 =10'b0;

   // m61_2 = W*in
   wire signed [9:0] m61_2;
   assign m61_2 =10'b0;

   // m61_3 = W*in
   wire signed [9:0] m61_3;
   assign m61_3 =10'b0;

   // m61_4 = W*in
   wire signed [9:0] m61_4;
   assign m61_4 =10'b0;

   // m61_5 = W*in
   wire signed [9:0] m61_5;
   assign m61_5 =10'b0;

   // m61_6 = W*in
   wire signed [9:0] m61_6;
   assign m61_6 ={ {5{in61[5]}} , in61[5:1] };

   // m61_7 = W*in
   wire signed [9:0] m61_7;
   assign m61_7 =10'b0;

   // m61_8 = W*in
   wire signed [9:0] m61_8;
   assign m61_8 =10'b0;

   // m61_9 = W*in
   wire signed [9:0] m61_9;
   assign m61_9 =10'b0;

   // m61_10 = W*in
   wire signed [9:0] m61_10;
   assign m61_10 =10'b0;

   // m61_11 = W*in
   wire signed [9:0] m61_11;
   assign m61_11 =10'b0;

   // m61_12 = W*in
   wire signed [9:0] m61_12;
   assign m61_12 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_13 = W*in
   wire signed [9:0] m61_13;
   assign m61_13 =10'b0;

   // m61_14 = W*in
   wire signed [9:0] m61_14;
   assign m61_14 ={ {4{in61[5]}} , in61[5:0] };

   // m61_15 = W*in
   wire signed [9:0] m61_15;
   assign m61_15 =10'b0;

   // m61_16 = W*in
   wire signed [9:0] m61_16;
   assign m61_16 ={ {4{in61[5]}} , in61[5:0] };

   // m61_17 = W*in
   wire signed [9:0] m61_17;
   assign m61_17 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_18 = W*in
   wire signed [9:0] m61_18;
   assign m61_18 =10'b0;

   // m61_19 = W*in
   wire signed [9:0] m61_19;
   assign m61_19 =10'b0;

   // m61_20 = W*in
   wire signed [9:0] m61_20;
   assign m61_20 =10'b0;

   // m61_21 = W*in
   wire signed [9:0] m61_21;
   assign m61_21 =10'b0;

   // m61_22 = W*in
   wire signed [9:0] m61_22;
   assign m61_22 ={ {4{in61[5]}} , in61[5:0] };

   // m61_23 = W*in
   wire signed [9:0] m61_23;
   assign m61_23 ={ {4{in61[5]}} , in61[5:0] };

   // m61_24 = W*in
   wire signed [9:0] m61_24;
   assign m61_24 =10'b0;

   // m61_25 = W*in
   wire signed [9:0] m61_25;
   assign m61_25 =10'b0;

   // m61_26 = W*in
   wire signed [9:0] m61_26;
   assign m61_26 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_27 = W*in
   wire signed [9:0] m61_27;
   assign m61_27 =10'b0;

   // m61_28 = W*in
   wire signed [9:0] m61_28;
   assign m61_28 =10'b0;

   // m61_29 = W*in
   wire signed [9:0] m61_29;
   assign m61_29 ={ {5{in61[5]}} , in61[5:1] };

   // m61_30 = W*in
   wire signed [9:0] m61_30;
   assign m61_30 =10'b0;

   // m61_31 = W*in
   wire signed [9:0] m61_31;
   assign m61_31 =10'b0;

   // m61_32 = W*in
   wire signed [9:0] m61_32;
   assign m61_32 =10'b0;

   // m61_33 = W*in
   wire signed [9:0] m61_33;
   assign m61_33 =10'b0;

   // m61_34 = W*in
   wire signed [9:0] m61_34;
   assign m61_34 =10'b0;

   // m61_35 = W*in
   wire signed [9:0] m61_35;
   assign m61_35 =10'b0;

   // m61_36 = W*in
   wire signed [9:0] m61_36;
   assign m61_36 ={ {5{neg61[5]}} , neg61[5:1] };

   // m61_37 = W*in
   wire signed [9:0] m61_37;
   assign m61_37 =10'b0;

   // m61_38 = W*in
   wire signed [9:0] m61_38;
   assign m61_38 =10'b0;

   // m61_39 = W*in
   wire signed [9:0] m61_39;
   assign m61_39 =10'b0;

   // m61_40 = W*in
   wire signed [9:0] m61_40;
   assign m61_40 =10'b0;

   // m61_41 = W*in
   wire signed [9:0] m61_41;
   assign m61_41 =10'b0;

   // m61_42 = W*in
   wire signed [9:0] m61_42;
   assign m61_42 =10'b0;

   // m61_43 = W*in
   wire signed [9:0] m61_43;
   assign m61_43 =10'b0;

   // m61_44 = W*in
   wire signed [9:0] m61_44;
   assign m61_44 =10'b0;

   // m61_45 = W*in
   wire signed [9:0] m61_45;
   assign m61_45 =10'b0;

   // m61_46 = W*in
   wire signed [9:0] m61_46;
   assign m61_46 =10'b0;

   // m61_47 = W*in
   wire signed [9:0] m61_47;
   assign m61_47 ={ {4{in61[5]}} , in61[5:0] };

   // m61_48 = W*in
   wire signed [9:0] m61_48;
   assign m61_48 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_49 = W*in
   wire signed [9:0] m61_49;
   assign m61_49 =10'b0;

   // m61_50 = W*in
   wire signed [9:0] m61_50;
   assign m61_50 =10'b0;

   // m61_51 = W*in
   wire signed [9:0] m61_51;
   assign m61_51 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_52 = W*in
   wire signed [9:0] m61_52;
   assign m61_52 =10'b0;

   // m61_53 = W*in
   wire signed [9:0] m61_53;
   assign m61_53 =10'b0;

   // m61_54 = W*in
   wire signed [9:0] m61_54;
   assign m61_54 =10'b0;

   // m61_55 = W*in
   wire signed [9:0] m61_55;
   assign m61_55 =10'b0;

   // m61_56 = W*in
   wire signed [9:0] m61_56;
   assign m61_56 =10'b0;

   // m61_57 = W*in
   wire signed [9:0] m61_57;
   assign m61_57 =10'b0;

   // m61_58 = W*in
   wire signed [9:0] m61_58;
   assign m61_58 =10'b0;

   // m61_59 = W*in
   wire signed [9:0] m61_59;
   assign m61_59 =10'b0;

   // m61_60 = W*in
   wire signed [9:0] m61_60;
   assign m61_60 =10'b0;

   // m61_61 = W*in
   wire signed [9:0] m61_61;
   assign m61_61 =10'b0;

   // m61_62 = W*in
   wire signed [9:0] m61_62;
   assign m61_62 =10'b0;

   // m61_63 = W*in
   wire signed [9:0] m61_63;
   assign m61_63 =10'b0;

   // m61_64 = W*in
   wire signed [9:0] m61_64;
   assign m61_64 ={ {4{in61[5]}} , in61[5:0] };

   // m61_65 = W*in
   wire signed [9:0] m61_65;
   assign m61_65 =10'b0;

   // m61_66 = W*in
   wire signed [9:0] m61_66;
   assign m61_66 =10'b0;

   // m61_67 = W*in
   wire signed [9:0] m61_67;
   assign m61_67 =10'b0;

   // m61_68 = W*in
   wire signed [9:0] m61_68;
   assign m61_68 =10'b0;

   // m61_69 = W*in
   wire signed [9:0] m61_69;
   assign m61_69 =10'b0;

   // m61_70 = W*in
   wire signed [9:0] m61_70;
   assign m61_70 ={ {5{in61[5]}} , in61[5:1] };

   // m61_71 = W*in
   wire signed [9:0] m61_71;
   assign m61_71 ={ {5{neg61[5]}} , neg61[5:1] };

   // m61_72 = W*in
   wire signed [9:0] m61_72;
   assign m61_72 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_73 = W*in
   wire signed [9:0] m61_73;
   assign m61_73 =10'b0;

   // m61_74 = W*in
   wire signed [9:0] m61_74;
   assign m61_74 =10'b0;

   // m61_75 = W*in
   wire signed [9:0] m61_75;
   assign m61_75 =10'b0;

   // m61_76 = W*in
   wire signed [9:0] m61_76;
   assign m61_76 =10'b0;

   // m61_77 = W*in
   wire signed [9:0] m61_77;
   assign m61_77 =10'b0;

   // m61_78 = W*in
   wire signed [9:0] m61_78;
   assign m61_78 =10'b0;

   // m61_79 = W*in
   wire signed [9:0] m61_79;
   assign m61_79 =10'b0;

   // m61_80 = W*in
   wire signed [9:0] m61_80;
   assign m61_80 =10'b0;

   // m61_81 = W*in
   wire signed [9:0] m61_81;
   assign m61_81 ={ {4{in61[5]}} , in61[5:0] };

   // m61_82 = W*in
   wire signed [9:0] m61_82;
   assign m61_82 =10'b0;

   // m61_83 = W*in
   wire signed [9:0] m61_83;
   assign m61_83 =10'b0;

   // m61_84 = W*in
   wire signed [9:0] m61_84;
   assign m61_84 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_85 = W*in
   wire signed [9:0] m61_85;
   assign m61_85 ={ {5{in61[5]}} , in61[5:1] };

   // m61_86 = W*in
   wire signed [9:0] m61_86;
   assign m61_86 =10'b0;

   // m61_87 = W*in
   wire signed [9:0] m61_87;
   assign m61_87 =10'b0;

   // m61_88 = W*in
   wire signed [9:0] m61_88;
   assign m61_88 =10'b0;

   // m61_89 = W*in
   wire signed [9:0] m61_89;
   assign m61_89 =10'b0;

   // m61_90 = W*in
   wire signed [9:0] m61_90;
   assign m61_90 =10'b0;

   // m61_91 = W*in
   wire signed [9:0] m61_91;
   assign m61_91 ={ {4{in61[5]}} , in61[5:0] };

   // m61_92 = W*in
   wire signed [9:0] m61_92;
   assign m61_92 =10'b0;

   // m61_93 = W*in
   wire signed [9:0] m61_93;
   assign m61_93 ={ {4{in61[5]}} , in61[5:0] };

   // m61_94 = W*in
   wire signed [9:0] m61_94;
   assign m61_94 =10'b0;

   // m61_95 = W*in
   wire signed [9:0] m61_95;
   assign m61_95 =10'b0;

   // m61_96 = W*in
   wire signed [9:0] m61_96;
   assign m61_96 =10'b0;

   // m61_97 = W*in
   wire signed [9:0] m61_97;
   assign m61_97 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_98 = W*in
   wire signed [9:0] m61_98;
   assign m61_98 =10'b0;

   // m61_99 = W*in
   wire signed [9:0] m61_99;
   assign m61_99 =10'b0;

   // m61_100 = W*in
   wire signed [9:0] m61_100;
   assign m61_100 =10'b0;

   // m61_101 = W*in
   wire signed [9:0] m61_101;
   assign m61_101 =10'b0;

   // m61_102 = W*in
   wire signed [9:0] m61_102;
   assign m61_102 =10'b0;

   // m61_103 = W*in
   wire signed [9:0] m61_103;
   assign m61_103 =10'b0;

   // m61_104 = W*in
   wire signed [9:0] m61_104;
   assign m61_104 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_105 = W*in
   wire signed [9:0] m61_105;
   assign m61_105 =10'b0;

   // m61_106 = W*in
   wire signed [9:0] m61_106;
   assign m61_106 =10'b0;

   // m61_107 = W*in
   wire signed [9:0] m61_107;
   assign m61_107 ={ {4{neg61[5]}} , neg61[5:0] };

   // m61_108 = W*in
   wire signed [9:0] m61_108;
   assign m61_108 =10'b0;

   // m61_109 = W*in
   wire signed [9:0] m61_109;
   assign m61_109 ={ {5{in61[5]}} , in61[5:1] };

   // m61_110 = W*in
   wire signed [9:0] m61_110;
   assign m61_110 =10'b0;

   // m61_111 = W*in
   wire signed [9:0] m61_111;
   assign m61_111 =10'b0;

   // m61_112 = W*in
   wire signed [9:0] m61_112;
   assign m61_112 =10'b0;

   // m61_113 = W*in
   wire signed [9:0] m61_113;
   assign m61_113 =10'b0;

   // m61_114 = W*in
   wire signed [9:0] m61_114;
   assign m61_114 =10'b0;

   // m61_115 = W*in
   wire signed [9:0] m61_115;
   assign m61_115 =10'b0;

   // m61_116 = W*in
   wire signed [9:0] m61_116;
   assign m61_116 =10'b0;

   // m61_117 = W*in
   wire signed [9:0] m61_117;
   assign m61_117 =10'b0;

   // m62_1 = W*in
   wire signed [9:0] m62_1;
   assign m62_1 =10'b0;

   // m62_2 = W*in
   wire signed [9:0] m62_2;
   assign m62_2 =10'b0;

   // m62_3 = W*in
   wire signed [9:0] m62_3;
   assign m62_3 =10'b0;

   // m62_4 = W*in
   wire signed [9:0] m62_4;
   assign m62_4 =10'b0;

   // m62_5 = W*in
   wire signed [9:0] m62_5;
   assign m62_5 =10'b0;

   // m62_6 = W*in
   wire signed [9:0] m62_6;
   assign m62_6 =10'b0;

   // m62_7 = W*in
   wire signed [9:0] m62_7;
   assign m62_7 =10'b0;

   // m62_8 = W*in
   wire signed [9:0] m62_8;
   assign m62_8 =10'b0;

   // m62_9 = W*in
   wire signed [9:0] m62_9;
   assign m62_9 =10'b0;

   // m62_10 = W*in
   wire signed [9:0] m62_10;
   assign m62_10 =10'b0;

   // m62_11 = W*in
   wire signed [9:0] m62_11;
   assign m62_11 =10'b0;

   // m62_12 = W*in
   wire signed [9:0] m62_12;
   assign m62_12 =10'b0;

   // m62_13 = W*in
   wire signed [9:0] m62_13;
   assign m62_13 =10'b0;

   // m62_14 = W*in
   wire signed [9:0] m62_14;
   assign m62_14 =10'b0;

   // m62_15 = W*in
   wire signed [9:0] m62_15;
   assign m62_15 =10'b0;

   // m62_16 = W*in
   wire signed [9:0] m62_16;
   assign m62_16 =10'b0;

   // m62_17 = W*in
   wire signed [9:0] m62_17;
   assign m62_17 =10'b0;

   // m62_18 = W*in
   wire signed [9:0] m62_18;
   assign m62_18 ={ {5{neg62[5]}} , neg62[5:1] };

   // m62_19 = W*in
   wire signed [9:0] m62_19;
   assign m62_19 =10'b0;

   // m62_20 = W*in
   wire signed [9:0] m62_20;
   assign m62_20 ={ {5{in62[5]}} , in62[5:1] };

   // m62_21 = W*in
   wire signed [9:0] m62_21;
   assign m62_21 =10'b0;

   // m62_22 = W*in
   wire signed [9:0] m62_22;
   assign m62_22 =10'b0;

   // m62_23 = W*in
   wire signed [9:0] m62_23;
   assign m62_23 =10'b0;

   // m62_24 = W*in
   wire signed [9:0] m62_24;
   assign m62_24 =10'b0;

   // m62_25 = W*in
   wire signed [9:0] m62_25;
   assign m62_25 =10'b0;

   // m62_26 = W*in
   wire signed [9:0] m62_26;
   assign m62_26 ={ {5{neg62[5]}} , neg62[5:1] };

   // m62_27 = W*in
   wire signed [9:0] m62_27;
   assign m62_27 =10'b0;

   // m62_28 = W*in
   wire signed [9:0] m62_28;
   assign m62_28 =10'b0;

   // m62_29 = W*in
   wire signed [9:0] m62_29;
   assign m62_29 ={ {5{in62[5]}} , in62[5:1] };

   // m62_30 = W*in
   wire signed [9:0] m62_30;
   assign m62_30 =10'b0;

   // m62_31 = W*in
   wire signed [9:0] m62_31;
   assign m62_31 =10'b0;

   // m62_32 = W*in
   wire signed [9:0] m62_32;
   assign m62_32 =10'b0;

   // m62_33 = W*in
   wire signed [9:0] m62_33;
   assign m62_33 =10'b0;

   // m62_34 = W*in
   wire signed [9:0] m62_34;
   assign m62_34 =10'b0;

   // m62_35 = W*in
   wire signed [9:0] m62_35;
   assign m62_35 =10'b0;

   // m62_36 = W*in
   wire signed [9:0] m62_36;
   assign m62_36 =10'b0;

   // m62_37 = W*in
   wire signed [9:0] m62_37;
   assign m62_37 =10'b0;

   // m62_38 = W*in
   wire signed [9:0] m62_38;
   assign m62_38 =10'b0;

   // m62_39 = W*in
   wire signed [9:0] m62_39;
   assign m62_39 =10'b0;

   // m62_40 = W*in
   wire signed [9:0] m62_40;
   assign m62_40 =10'b0;

   // m62_41 = W*in
   wire signed [9:0] m62_41;
   assign m62_41 =10'b0;

   // m62_42 = W*in
   wire signed [9:0] m62_42;
   assign m62_42 =10'b0;

   // m62_43 = W*in
   wire signed [9:0] m62_43;
   assign m62_43 =10'b0;

   // m62_44 = W*in
   wire signed [9:0] m62_44;
   assign m62_44 =10'b0;

   // m62_45 = W*in
   wire signed [9:0] m62_45;
   assign m62_45 =10'b0;

   // m62_46 = W*in
   wire signed [9:0] m62_46;
   assign m62_46 =10'b0;

   // m62_47 = W*in
   wire signed [9:0] m62_47;
   assign m62_47 =10'b0;

   // m62_48 = W*in
   wire signed [9:0] m62_48;
   assign m62_48 =10'b0;

   // m62_49 = W*in
   wire signed [9:0] m62_49;
   assign m62_49 =10'b0;

   // m62_50 = W*in
   wire signed [9:0] m62_50;
   assign m62_50 =10'b0;

   // m62_51 = W*in
   wire signed [9:0] m62_51;
   assign m62_51 =10'b0;

   // m62_52 = W*in
   wire signed [9:0] m62_52;
   assign m62_52 =10'b0;

   // m62_53 = W*in
   wire signed [9:0] m62_53;
   assign m62_53 =10'b0;

   // m62_54 = W*in
   wire signed [9:0] m62_54;
   assign m62_54 =10'b0;

   // m62_55 = W*in
   wire signed [9:0] m62_55;
   assign m62_55 =10'b0;

   // m62_56 = W*in
   wire signed [9:0] m62_56;
   assign m62_56 =10'b0;

   // m62_57 = W*in
   wire signed [9:0] m62_57;
   assign m62_57 =10'b0;

   // m62_58 = W*in
   wire signed [9:0] m62_58;
   assign m62_58 =10'b0;

   // m62_59 = W*in
   wire signed [9:0] m62_59;
   assign m62_59 =10'b0;

   // m62_60 = W*in
   wire signed [9:0] m62_60;
   assign m62_60 =10'b0;

   // m62_61 = W*in
   wire signed [9:0] m62_61;
   assign m62_61 =10'b0;

   // m62_62 = W*in
   wire signed [9:0] m62_62;
   assign m62_62 =10'b0;

   // m62_63 = W*in
   wire signed [9:0] m62_63;
   assign m62_63 =10'b0;

   // m62_64 = W*in
   wire signed [9:0] m62_64;
   assign m62_64 =10'b0;

   // m62_65 = W*in
   wire signed [9:0] m62_65;
   assign m62_65 =10'b0;

   // m62_66 = W*in
   wire signed [9:0] m62_66;
   assign m62_66 =10'b0;

   // m62_67 = W*in
   wire signed [9:0] m62_67;
   assign m62_67 =10'b0;

   // m62_68 = W*in
   wire signed [9:0] m62_68;
   assign m62_68 =10'b0;

   // m62_69 = W*in
   wire signed [9:0] m62_69;
   assign m62_69 ={ {5{in62[5]}} , in62[5:1] };

   // m62_70 = W*in
   wire signed [9:0] m62_70;
   assign m62_70 ={ {5{neg62[5]}} , neg62[5:1] };

   // m62_71 = W*in
   wire signed [9:0] m62_71;
   assign m62_71 =10'b0;

   // m62_72 = W*in
   wire signed [9:0] m62_72;
   assign m62_72 =10'b0;

   // m62_73 = W*in
   wire signed [9:0] m62_73;
   assign m62_73 =10'b0;

   // m62_74 = W*in
   wire signed [9:0] m62_74;
   assign m62_74 =10'b0;

   // m62_75 = W*in
   wire signed [9:0] m62_75;
   assign m62_75 =10'b0;

   // m62_76 = W*in
   wire signed [9:0] m62_76;
   assign m62_76 =10'b0;

   // m62_77 = W*in
   wire signed [9:0] m62_77;
   assign m62_77 =10'b0;

   // m62_78 = W*in
   wire signed [9:0] m62_78;
   assign m62_78 =10'b0;

   // m62_79 = W*in
   wire signed [9:0] m62_79;
   assign m62_79 ={ {4{in62[5]}} , in62[5:0] };

   // m62_80 = W*in
   wire signed [9:0] m62_80;
   assign m62_80 =10'b0;

   // m62_81 = W*in
   wire signed [9:0] m62_81;
   assign m62_81 =10'b0;

   // m62_82 = W*in
   wire signed [9:0] m62_82;
   assign m62_82 =10'b0;

   // m62_83 = W*in
   wire signed [9:0] m62_83;
   assign m62_83 =10'b0;

   // m62_84 = W*in
   wire signed [9:0] m62_84;
   assign m62_84 =10'b0;

   // m62_85 = W*in
   wire signed [9:0] m62_85;
   assign m62_85 =10'b0;

   // m62_86 = W*in
   wire signed [9:0] m62_86;
   assign m62_86 =10'b0;

   // m62_87 = W*in
   wire signed [9:0] m62_87;
   assign m62_87 =10'b0;

   // m62_88 = W*in
   wire signed [9:0] m62_88;
   assign m62_88 =10'b0;

   // m62_89 = W*in
   wire signed [9:0] m62_89;
   assign m62_89 =10'b0;

   // m62_90 = W*in
   wire signed [9:0] m62_90;
   assign m62_90 =10'b0;

   // m62_91 = W*in
   wire signed [9:0] m62_91;
   assign m62_91 =10'b0;

   // m62_92 = W*in
   wire signed [9:0] m62_92;
   assign m62_92 =10'b0;

   // m62_93 = W*in
   wire signed [9:0] m62_93;
   assign m62_93 =10'b0;

   // m62_94 = W*in
   wire signed [9:0] m62_94;
   assign m62_94 =10'b0;

   // m62_95 = W*in
   wire signed [9:0] m62_95;
   assign m62_95 =10'b0;

   // m62_96 = W*in
   wire signed [9:0] m62_96;
   assign m62_96 =10'b0;

   // m62_97 = W*in
   wire signed [9:0] m62_97;
   assign m62_97 =10'b0;

   // m62_98 = W*in
   wire signed [9:0] m62_98;
   assign m62_98 =10'b0;

   // m62_99 = W*in
   wire signed [9:0] m62_99;
   assign m62_99 =10'b0;

   // m62_100 = W*in
   wire signed [9:0] m62_100;
   assign m62_100 =10'b0;

   // m62_101 = W*in
   wire signed [9:0] m62_101;
   assign m62_101 =10'b0;

   // m62_102 = W*in
   wire signed [9:0] m62_102;
   assign m62_102 =10'b0;

   // m62_103 = W*in
   wire signed [9:0] m62_103;
   assign m62_103 =10'b0;

   // m62_104 = W*in
   wire signed [9:0] m62_104;
   assign m62_104 =10'b0;

   // m62_105 = W*in
   wire signed [9:0] m62_105;
   assign m62_105 =10'b0;

   // m62_106 = W*in
   wire signed [9:0] m62_106;
   assign m62_106 =10'b0;

   // m62_107 = W*in
   wire signed [9:0] m62_107;
   assign m62_107 ={ {4{neg62[5]}} , neg62[5:0] };

   // m62_108 = W*in
   wire signed [9:0] m62_108;
   assign m62_108 ={ {5{in62[5]}} , in62[5:1] };

   // m62_109 = W*in
   wire signed [9:0] m62_109;
   assign m62_109 =10'b0;

   // m62_110 = W*in
   wire signed [9:0] m62_110;
   assign m62_110 =10'b0;

   // m62_111 = W*in
   wire signed [9:0] m62_111;
   assign m62_111 =10'b0;

   // m62_112 = W*in
   wire signed [9:0] m62_112;
   assign m62_112 =10'b0;

   // m62_113 = W*in
   wire signed [9:0] m62_113;
   assign m62_113 =10'b0;

   // m62_114 = W*in
   wire signed [9:0] m62_114;
   assign m62_114 =10'b0;

   // m62_115 = W*in
   wire signed [9:0] m62_115;
   assign m62_115 =10'b0;

   // m62_116 = W*in
   wire signed [9:0] m62_116;
   assign m62_116 =10'b0;

   // m62_117 = W*in
   wire signed [9:0] m62_117;
   assign m62_117 =10'b0;

   // m63_1 = W*in
   wire signed [9:0] m63_1;
   assign m63_1 =10'b0;

   // m63_2 = W*in
   wire signed [9:0] m63_2;
   assign m63_2 =10'b0;

   // m63_3 = W*in
   wire signed [9:0] m63_3;
   assign m63_3 =10'b0;

   // m63_4 = W*in
   wire signed [9:0] m63_4;
   assign m63_4 =10'b0;

   // m63_5 = W*in
   wire signed [9:0] m63_5;
   assign m63_5 =10'b0;

   // m63_6 = W*in
   wire signed [9:0] m63_6;
   assign m63_6 ={ {4{in63[5]}} , in63[5:0] };

   // m63_7 = W*in
   wire signed [9:0] m63_7;
   assign m63_7 =10'b0;

   // m63_8 = W*in
   wire signed [9:0] m63_8;
   assign m63_8 =10'b0;

   // m63_9 = W*in
   wire signed [9:0] m63_9;
   assign m63_9 =10'b0;

   // m63_10 = W*in
   wire signed [9:0] m63_10;
   assign m63_10 =10'b0;

   // m63_11 = W*in
   wire signed [9:0] m63_11;
   assign m63_11 =10'b0;

   // m63_12 = W*in
   wire signed [9:0] m63_12;
   assign m63_12 =10'b0;

   // m63_13 = W*in
   wire signed [9:0] m63_13;
   assign m63_13 =10'b0;

   // m63_14 = W*in
   wire signed [9:0] m63_14;
   assign m63_14 =10'b0;

   // m63_15 = W*in
   wire signed [9:0] m63_15;
   assign m63_15 =10'b0;

   // m63_16 = W*in
   wire signed [9:0] m63_16;
   assign m63_16 =10'b0;

   // m63_17 = W*in
   wire signed [9:0] m63_17;
   assign m63_17 ={ {5{neg63[5]}} , neg63[5:1] };

   // m63_18 = W*in
   wire signed [9:0] m63_18;
   assign m63_18 =10'b0;

   // m63_19 = W*in
   wire signed [9:0] m63_19;
   assign m63_19 =10'b0;

   // m63_20 = W*in
   wire signed [9:0] m63_20;
   assign m63_20 =10'b0;

   // m63_21 = W*in
   wire signed [9:0] m63_21;
   assign m63_21 =10'b0;

   // m63_22 = W*in
   wire signed [9:0] m63_22;
   assign m63_22 ={ {4{in63[5]}} , in63[5:0] };

   // m63_23 = W*in
   wire signed [9:0] m63_23;
   assign m63_23 ={ {4{in63[5]}} , in63[5:0] };

   // m63_24 = W*in
   wire signed [9:0] m63_24;
   assign m63_24 ={ {4{in63[5]}} , in63[5:0] };

   // m63_25 = W*in
   wire signed [9:0] m63_25;
   assign m63_25 =10'b0;

   // m63_26 = W*in
   wire signed [9:0] m63_26;
   assign m63_26 ={ {4{neg63[5]}} , neg63[5:0] };

   // m63_27 = W*in
   wire signed [9:0] m63_27;
   assign m63_27 ={ {5{in63[5]}} , in63[5:1] };

   // m63_28 = W*in
   wire signed [9:0] m63_28;
   assign m63_28 =10'b0;

   // m63_29 = W*in
   wire signed [9:0] m63_29;
   assign m63_29 ={ {4{in63[5]}} , in63[5:0] };

   // m63_30 = W*in
   wire signed [9:0] m63_30;
   assign m63_30 =10'b0;

   // m63_31 = W*in
   wire signed [9:0] m63_31;
   assign m63_31 =10'b0;

   // m63_32 = W*in
   wire signed [9:0] m63_32;
   assign m63_32 =10'b0;

   // m63_33 = W*in
   wire signed [9:0] m63_33;
   assign m63_33 =10'b0;

   // m63_34 = W*in
   wire signed [9:0] m63_34;
   assign m63_34 =10'b0;

   // m63_35 = W*in
   wire signed [9:0] m63_35;
   assign m63_35 =10'b0;

   // m63_36 = W*in
   wire signed [9:0] m63_36;
   assign m63_36 =10'b0;

   // m63_37 = W*in
   wire signed [9:0] m63_37;
   assign m63_37 =10'b0;

   // m63_38 = W*in
   wire signed [9:0] m63_38;
   assign m63_38 =10'b0;

   // m63_39 = W*in
   wire signed [9:0] m63_39;
   assign m63_39 =10'b0;

   // m63_40 = W*in
   wire signed [9:0] m63_40;
   assign m63_40 =10'b0;

   // m63_41 = W*in
   wire signed [9:0] m63_41;
   assign m63_41 =10'b0;

   // m63_42 = W*in
   wire signed [9:0] m63_42;
   assign m63_42 =10'b0;

   // m63_43 = W*in
   wire signed [9:0] m63_43;
   assign m63_43 =10'b0;

   // m63_44 = W*in
   wire signed [9:0] m63_44;
   assign m63_44 =10'b0;

   // m63_45 = W*in
   wire signed [9:0] m63_45;
   assign m63_45 =10'b0;

   // m63_46 = W*in
   wire signed [9:0] m63_46;
   assign m63_46 =10'b0;

   // m63_47 = W*in
   wire signed [9:0] m63_47;
   assign m63_47 =10'b0;

   // m63_48 = W*in
   wire signed [9:0] m63_48;
   assign m63_48 ={ {4{neg63[5]}} , neg63[5:0] };

   // m63_49 = W*in
   wire signed [9:0] m63_49;
   assign m63_49 =10'b0;

   // m63_50 = W*in
   wire signed [9:0] m63_50;
   assign m63_50 =10'b0;

   // m63_51 = W*in
   wire signed [9:0] m63_51;
   assign m63_51 =10'b0;

   // m63_52 = W*in
   wire signed [9:0] m63_52;
   assign m63_52 =10'b0;

   // m63_53 = W*in
   wire signed [9:0] m63_53;
   assign m63_53 =10'b0;

   // m63_54 = W*in
   wire signed [9:0] m63_54;
   assign m63_54 =10'b0;

   // m63_55 = W*in
   wire signed [9:0] m63_55;
   assign m63_55 =10'b0;

   // m63_56 = W*in
   wire signed [9:0] m63_56;
   assign m63_56 =10'b0;

   // m63_57 = W*in
   wire signed [9:0] m63_57;
   assign m63_57 =10'b0;

   // m63_58 = W*in
   wire signed [9:0] m63_58;
   assign m63_58 ={ {5{in63[5]}} , in63[5:1] };

   // m63_59 = W*in
   wire signed [9:0] m63_59;
   assign m63_59 =10'b0;

   // m63_60 = W*in
   wire signed [9:0] m63_60;
   assign m63_60 =10'b0;

   // m63_61 = W*in
   wire signed [9:0] m63_61;
   assign m63_61 =10'b0;

   // m63_62 = W*in
   wire signed [9:0] m63_62;
   assign m63_62 =10'b0;

   // m63_63 = W*in
   wire signed [9:0] m63_63;
   assign m63_63 =10'b0;

   // m63_64 = W*in
   wire signed [9:0] m63_64;
   assign m63_64 =10'b0;

   // m63_65 = W*in
   wire signed [9:0] m63_65;
   assign m63_65 ={ {5{in63[5]}} , in63[5:1] };

   // m63_66 = W*in
   wire signed [9:0] m63_66;
   assign m63_66 =10'b0;

   // m63_67 = W*in
   wire signed [9:0] m63_67;
   assign m63_67 =10'b0;

   // m63_68 = W*in
   wire signed [9:0] m63_68;
   assign m63_68 =10'b0;

   // m63_69 = W*in
   wire signed [9:0] m63_69;
   assign m63_69 =10'b0;

   // m63_70 = W*in
   wire signed [9:0] m63_70;
   assign m63_70 =10'b0;

   // m63_71 = W*in
   wire signed [9:0] m63_71;
   assign m63_71 =10'b0;

   // m63_72 = W*in
   wire signed [9:0] m63_72;
   assign m63_72 =10'b0;

   // m63_73 = W*in
   wire signed [9:0] m63_73;
   assign m63_73 =10'b0;

   // m63_74 = W*in
   wire signed [9:0] m63_74;
   assign m63_74 ={ {5{neg63[5]}} , neg63[5:1] };

   // m63_75 = W*in
   wire signed [9:0] m63_75;
   assign m63_75 ={ {5{neg63[5]}} , neg63[5:1] };

   // m63_76 = W*in
   wire signed [9:0] m63_76;
   assign m63_76 =10'b0;

   // m63_77 = W*in
   wire signed [9:0] m63_77;
   assign m63_77 =10'b0;

   // m63_78 = W*in
   wire signed [9:0] m63_78;
   assign m63_78 ={ {4{neg63[5]}} , neg63[5:0] };

   // m63_79 = W*in
   wire signed [9:0] m63_79;
   assign m63_79 =10'b0;

   // m63_80 = W*in
   wire signed [9:0] m63_80;
   assign m63_80 =10'b0;

   // m63_81 = W*in
   wire signed [9:0] m63_81;
   assign m63_81 ={ {5{neg63[5]}} , neg63[5:1] };

   // m63_82 = W*in
   wire signed [9:0] m63_82;
   assign m63_82 =10'b0;

   // m63_83 = W*in
   wire signed [9:0] m63_83;
   assign m63_83 =10'b0;

   // m63_84 = W*in
   wire signed [9:0] m63_84;
   assign m63_84 =10'b0;

   // m63_85 = W*in
   wire signed [9:0] m63_85;
   assign m63_85 ={ {4{in63[5]}} , in63[5:0] };

   // m63_86 = W*in
   wire signed [9:0] m63_86;
   assign m63_86 =10'b0;

   // m63_87 = W*in
   wire signed [9:0] m63_87;
   assign m63_87 =10'b0;

   // m63_88 = W*in
   wire signed [9:0] m63_88;
   assign m63_88 ={ {4{neg63[5]}} , neg63[5:0] };

   // m63_89 = W*in
   wire signed [9:0] m63_89;
   assign m63_89 ={ {4{in63[5]}} , in63[5:0] };

   // m63_90 = W*in
   wire signed [9:0] m63_90;
   assign m63_90 =10'b0;

   // m63_91 = W*in
   wire signed [9:0] m63_91;
   assign m63_91 =10'b0;

   // m63_92 = W*in
   wire signed [9:0] m63_92;
   assign m63_92 ={ {4{neg63[5]}} , neg63[5:0] };

   // m63_93 = W*in
   wire signed [9:0] m63_93;
   assign m63_93 ={ {4{in63[5]}} , in63[5:0] };

   // m63_94 = W*in
   wire signed [9:0] m63_94;
   assign m63_94 =10'b0;

   // m63_95 = W*in
   wire signed [9:0] m63_95;
   assign m63_95 =10'b0;

   // m63_96 = W*in
   wire signed [9:0] m63_96;
   assign m63_96 =10'b0;

   // m63_97 = W*in
   wire signed [9:0] m63_97;
   assign m63_97 =10'b0;

   // m63_98 = W*in
   wire signed [9:0] m63_98;
   assign m63_98 =10'b0;

   // m63_99 = W*in
   wire signed [9:0] m63_99;
   assign m63_99 =10'b0;

   // m63_100 = W*in
   wire signed [9:0] m63_100;
   assign m63_100 =10'b0;

   // m63_101 = W*in
   wire signed [9:0] m63_101;
   assign m63_101 =10'b0;

   // m63_102 = W*in
   wire signed [9:0] m63_102;
   assign m63_102 =10'b0;

   // m63_103 = W*in
   wire signed [9:0] m63_103;
   assign m63_103 =10'b0;

   // m63_104 = W*in
   wire signed [9:0] m63_104;
   assign m63_104 =10'b0;

   // m63_105 = W*in
   wire signed [9:0] m63_105;
   assign m63_105 =10'b0;

   // m63_106 = W*in
   wire signed [9:0] m63_106;
   assign m63_106 =10'b0;

   // m63_107 = W*in
   wire signed [9:0] m63_107;
   assign m63_107 =10'b0;

   // m63_108 = W*in
   wire signed [9:0] m63_108;
   assign m63_108 ={ {4{in63[5]}} , in63[5:0] };

   // m63_109 = W*in
   wire signed [9:0] m63_109;
   assign m63_109 ={ {4{in63[5]}} , in63[5:0] };

   // m63_110 = W*in
   wire signed [9:0] m63_110;
   assign m63_110 =10'b0;

   // m63_111 = W*in
   wire signed [9:0] m63_111;
   assign m63_111 =10'b0;

   // m63_112 = W*in
   wire signed [9:0] m63_112;
   assign m63_112 =10'b0;

   // m63_113 = W*in
   wire signed [9:0] m63_113;
   assign m63_113 ={ {4{neg63[5]}} , neg63[5:0] };

   // m63_114 = W*in
   wire signed [9:0] m63_114;
   assign m63_114 =10'b0;

   // m63_115 = W*in
   wire signed [9:0] m63_115;
   assign m63_115 =10'b0;

   // m63_116 = W*in
   wire signed [9:0] m63_116;
   assign m63_116 =10'b0;

   // m63_117 = W*in
   wire signed [9:0] m63_117;
   assign m63_117 =10'b0;

   // m64_1 = W*in
   wire signed [9:0] m64_1;
   assign m64_1 =10'b0;

   // m64_2 = W*in
   wire signed [9:0] m64_2;
   assign m64_2 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_3 = W*in
   wire signed [9:0] m64_3;
   assign m64_3 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_4 = W*in
   wire signed [9:0] m64_4;
   assign m64_4 =10'b0;

   // m64_5 = W*in
   wire signed [9:0] m64_5;
   assign m64_5 =10'b0;

   // m64_6 = W*in
   wire signed [9:0] m64_6;
   assign m64_6 =10'b0;

   // m64_7 = W*in
   wire signed [9:0] m64_7;
   assign m64_7 =10'b0;

   // m64_8 = W*in
   wire signed [9:0] m64_8;
   assign m64_8 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_9 = W*in
   wire signed [9:0] m64_9;
   assign m64_9 =10'b0;

   // m64_10 = W*in
   wire signed [9:0] m64_10;
   assign m64_10 =10'b0;

   // m64_11 = W*in
   wire signed [9:0] m64_11;
   assign m64_11 =10'b0;

   // m64_12 = W*in
   wire signed [9:0] m64_12;
   assign m64_12 =10'b0;

   // m64_13 = W*in
   wire signed [9:0] m64_13;
   assign m64_13 ={ {4{in64[5]}} , in64[5:0] };

   // m64_14 = W*in
   wire signed [9:0] m64_14;
   assign m64_14 =10'b0;

   // m64_15 = W*in
   wire signed [9:0] m64_15;
   assign m64_15 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_16 = W*in
   wire signed [9:0] m64_16;
   assign m64_16 =10'b0;

   // m64_17 = W*in
   wire signed [9:0] m64_17;
   assign m64_17 ={ {5{neg64[5]}} , neg64[5:1] };

   // m64_18 = W*in
   wire signed [9:0] m64_18;
   assign m64_18 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_19 = W*in
   wire signed [9:0] m64_19;
   assign m64_19 =10'b0;

   // m64_20 = W*in
   wire signed [9:0] m64_20;
   assign m64_20 =10'b0;

   // m64_21 = W*in
   wire signed [9:0] m64_21;
   assign m64_21 =10'b0;

   // m64_22 = W*in
   wire signed [9:0] m64_22;
   assign m64_22 =10'b0;

   // m64_23 = W*in
   wire signed [9:0] m64_23;
   assign m64_23 =10'b0;

   // m64_24 = W*in
   wire signed [9:0] m64_24;
   assign m64_24 =10'b0;

   // m64_25 = W*in
   wire signed [9:0] m64_25;
   assign m64_25 =10'b0;

   // m64_26 = W*in
   wire signed [9:0] m64_26;
   assign m64_26 =10'b0;

   // m64_27 = W*in
   wire signed [9:0] m64_27;
   assign m64_27 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_28 = W*in
   wire signed [9:0] m64_28;
   assign m64_28 ={ {5{neg64[5]}} , neg64[5:1] };

   // m64_29 = W*in
   wire signed [9:0] m64_29;
   assign m64_29 ={ {4{in64[5]}} , in64[5:0] };

   // m64_30 = W*in
   wire signed [9:0] m64_30;
   assign m64_30 =10'b0;

   // m64_31 = W*in
   wire signed [9:0] m64_31;
   assign m64_31 ={ {5{neg64[5]}} , neg64[5:1] };

   // m64_32 = W*in
   wire signed [9:0] m64_32;
   assign m64_32 ={ {4{in64[5]}} , in64[5:0] };

   // m64_33 = W*in
   wire signed [9:0] m64_33;
   assign m64_33 =10'b0;

   // m64_34 = W*in
   wire signed [9:0] m64_34;
   assign m64_34 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_35 = W*in
   wire signed [9:0] m64_35;
   assign m64_35 =10'b0;

   // m64_36 = W*in
   wire signed [9:0] m64_36;
   assign m64_36 =10'b0;

   // m64_37 = W*in
   wire signed [9:0] m64_37;
   assign m64_37 ={ {4{in64[5]}} , in64[5:0] };

   // m64_38 = W*in
   wire signed [9:0] m64_38;
   assign m64_38 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_39 = W*in
   wire signed [9:0] m64_39;
   assign m64_39 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_40 = W*in
   wire signed [9:0] m64_40;
   assign m64_40 =10'b0;

   // m64_41 = W*in
   wire signed [9:0] m64_41;
   assign m64_41 =10'b0;

   // m64_42 = W*in
   wire signed [9:0] m64_42;
   assign m64_42 =10'b0;

   // m64_43 = W*in
   wire signed [9:0] m64_43;
   assign m64_43 =10'b0;

   // m64_44 = W*in
   wire signed [9:0] m64_44;
   assign m64_44 =10'b0;

   // m64_45 = W*in
   wire signed [9:0] m64_45;
   assign m64_45 =10'b0;

   // m64_46 = W*in
   wire signed [9:0] m64_46;
   assign m64_46 =10'b0;

   // m64_47 = W*in
   wire signed [9:0] m64_47;
   assign m64_47 =10'b0;

   // m64_48 = W*in
   wire signed [9:0] m64_48;
   assign m64_48 =10'b0;

   // m64_49 = W*in
   wire signed [9:0] m64_49;
   assign m64_49 =10'b0;

   // m64_50 = W*in
   wire signed [9:0] m64_50;
   assign m64_50 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_51 = W*in
   wire signed [9:0] m64_51;
   assign m64_51 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_52 = W*in
   wire signed [9:0] m64_52;
   assign m64_52 =10'b0;

   // m64_53 = W*in
   wire signed [9:0] m64_53;
   assign m64_53 =10'b0;

   // m64_54 = W*in
   wire signed [9:0] m64_54;
   assign m64_54 =10'b0;

   // m64_55 = W*in
   wire signed [9:0] m64_55;
   assign m64_55 =10'b0;

   // m64_56 = W*in
   wire signed [9:0] m64_56;
   assign m64_56 =10'b0;

   // m64_57 = W*in
   wire signed [9:0] m64_57;
   assign m64_57 =10'b0;

   // m64_58 = W*in
   wire signed [9:0] m64_58;
   assign m64_58 =10'b0;

   // m64_59 = W*in
   wire signed [9:0] m64_59;
   assign m64_59 =10'b0;

   // m64_60 = W*in
   wire signed [9:0] m64_60;
   assign m64_60 =10'b0;

   // m64_61 = W*in
   wire signed [9:0] m64_61;
   assign m64_61 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_62 = W*in
   wire signed [9:0] m64_62;
   assign m64_62 =10'b0;

   // m64_63 = W*in
   wire signed [9:0] m64_63;
   assign m64_63 =10'b0;

   // m64_64 = W*in
   wire signed [9:0] m64_64;
   assign m64_64 =10'b0;

   // m64_65 = W*in
   wire signed [9:0] m64_65;
   assign m64_65 ={ {4{in64[5]}} , in64[5:0] };

   // m64_66 = W*in
   wire signed [9:0] m64_66;
   assign m64_66 =10'b0;

   // m64_67 = W*in
   wire signed [9:0] m64_67;
   assign m64_67 =10'b0;

   // m64_68 = W*in
   wire signed [9:0] m64_68;
   assign m64_68 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_69 = W*in
   wire signed [9:0] m64_69;
   assign m64_69 =10'b0;

   // m64_70 = W*in
   wire signed [9:0] m64_70;
   assign m64_70 =10'b0;

   // m64_71 = W*in
   wire signed [9:0] m64_71;
   assign m64_71 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_72 = W*in
   wire signed [9:0] m64_72;
   assign m64_72 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_73 = W*in
   wire signed [9:0] m64_73;
   assign m64_73 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_74 = W*in
   wire signed [9:0] m64_74;
   assign m64_74 =10'b0;

   // m64_75 = W*in
   wire signed [9:0] m64_75;
   assign m64_75 =10'b0;

   // m64_76 = W*in
   wire signed [9:0] m64_76;
   assign m64_76 =10'b0;

   // m64_77 = W*in
   wire signed [9:0] m64_77;
   assign m64_77 =10'b0;

   // m64_78 = W*in
   wire signed [9:0] m64_78;
   assign m64_78 =10'b0;

   // m64_79 = W*in
   wire signed [9:0] m64_79;
   assign m64_79 =10'b0;

   // m64_80 = W*in
   wire signed [9:0] m64_80;
   assign m64_80 =10'b0;

   // m64_81 = W*in
   wire signed [9:0] m64_81;
   assign m64_81 =10'b0;

   // m64_82 = W*in
   wire signed [9:0] m64_82;
   assign m64_82 =10'b0;

   // m64_83 = W*in
   wire signed [9:0] m64_83;
   assign m64_83 =10'b0;

   // m64_84 = W*in
   wire signed [9:0] m64_84;
   assign m64_84 =10'b0;

   // m64_85 = W*in
   wire signed [9:0] m64_85;
   assign m64_85 ={ {4{in64[5]}} , in64[5:0] };

   // m64_86 = W*in
   wire signed [9:0] m64_86;
   assign m64_86 =10'b0;

   // m64_87 = W*in
   wire signed [9:0] m64_87;
   assign m64_87 =10'b0;

   // m64_88 = W*in
   wire signed [9:0] m64_88;
   assign m64_88 =10'b0;

   // m64_89 = W*in
   wire signed [9:0] m64_89;
   assign m64_89 =10'b0;

   // m64_90 = W*in
   wire signed [9:0] m64_90;
   assign m64_90 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_91 = W*in
   wire signed [9:0] m64_91;
   assign m64_91 =10'b0;

   // m64_92 = W*in
   wire signed [9:0] m64_92;
   assign m64_92 =10'b0;

   // m64_93 = W*in
   wire signed [9:0] m64_93;
   assign m64_93 ={ {4{in64[5]}} , in64[5:0] };

   // m64_94 = W*in
   wire signed [9:0] m64_94;
   assign m64_94 =10'b0;

   // m64_95 = W*in
   wire signed [9:0] m64_95;
   assign m64_95 =10'b0;

   // m64_96 = W*in
   wire signed [9:0] m64_96;
   assign m64_96 =10'b0;

   // m64_97 = W*in
   wire signed [9:0] m64_97;
   assign m64_97 =10'b0;

   // m64_98 = W*in
   wire signed [9:0] m64_98;
   assign m64_98 =10'b0;

   // m64_99 = W*in
   wire signed [9:0] m64_99;
   assign m64_99 =10'b0;

   // m64_100 = W*in
   wire signed [9:0] m64_100;
   assign m64_100 =10'b0;

   // m64_101 = W*in
   wire signed [9:0] m64_101;
   assign m64_101 =10'b0;

   // m64_102 = W*in
   wire signed [9:0] m64_102;
   assign m64_102 =10'b0;

   // m64_103 = W*in
   wire signed [9:0] m64_103;
   assign m64_103 =10'b0;

   // m64_104 = W*in
   wire signed [9:0] m64_104;
   assign m64_104 =10'b0;

   // m64_105 = W*in
   wire signed [9:0] m64_105;
   assign m64_105 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_106 = W*in
   wire signed [9:0] m64_106;
   assign m64_106 =10'b0;

   // m64_107 = W*in
   wire signed [9:0] m64_107;
   assign m64_107 ={ {4{neg64[5]}} , neg64[5:0] };

   // m64_108 = W*in
   wire signed [9:0] m64_108;
   assign m64_108 =10'b0;

   // m64_109 = W*in
   wire signed [9:0] m64_109;
   assign m64_109 ={ {4{in64[5]}} , in64[5:0] };

   // m64_110 = W*in
   wire signed [9:0] m64_110;
   assign m64_110 ={ {4{in64[5]}} , in64[5:0] };

   // m64_111 = W*in
   wire signed [9:0] m64_111;
   assign m64_111 =10'b0;

   // m64_112 = W*in
   wire signed [9:0] m64_112;
   assign m64_112 ={ {4{in64[5]}} , in64[5:0] };

   // m64_113 = W*in
   wire signed [9:0] m64_113;
   assign m64_113 =10'b0;

   // m64_114 = W*in
   wire signed [9:0] m64_114;
   assign m64_114 =10'b0;

   // m64_115 = W*in
   wire signed [9:0] m64_115;
   assign m64_115 =10'b0;

   // m64_116 = W*in
   wire signed [9:0] m64_116;
   assign m64_116 =10'b0;

   // m64_117 = W*in
   wire signed [9:0] m64_117;
   assign m64_117 =10'b0;

   // m65_1 = W*in
   wire signed [9:0] m65_1;
   assign m65_1 =10'b0;

   // m65_2 = W*in
   wire signed [9:0] m65_2;
   assign m65_2 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_3 = W*in
   wire signed [9:0] m65_3;
   assign m65_3 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_4 = W*in
   wire signed [9:0] m65_4;
   assign m65_4 =10'b0;

   // m65_5 = W*in
   wire signed [9:0] m65_5;
   assign m65_5 =10'b0;

   // m65_6 = W*in
   wire signed [9:0] m65_6;
   assign m65_6 ={ {4{in65[5]}} , in65[5:0] };

   // m65_7 = W*in
   wire signed [9:0] m65_7;
   assign m65_7 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_8 = W*in
   wire signed [9:0] m65_8;
   assign m65_8 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_9 = W*in
   wire signed [9:0] m65_9;
   assign m65_9 =10'b0;

   // m65_10 = W*in
   wire signed [9:0] m65_10;
   assign m65_10 ={ {4{in65[5]}} , in65[5:0] };

   // m65_11 = W*in
   wire signed [9:0] m65_11;
   assign m65_11 =10'b0;

   // m65_12 = W*in
   wire signed [9:0] m65_12;
   assign m65_12 =10'b0;

   // m65_13 = W*in
   wire signed [9:0] m65_13;
   assign m65_13 =10'b0;

   // m65_14 = W*in
   wire signed [9:0] m65_14;
   assign m65_14 =10'b0;

   // m65_15 = W*in
   wire signed [9:0] m65_15;
   assign m65_15 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_16 = W*in
   wire signed [9:0] m65_16;
   assign m65_16 =10'b0;

   // m65_17 = W*in
   wire signed [9:0] m65_17;
   assign m65_17 ={ {5{neg65[5]}} , neg65[5:1] };

   // m65_18 = W*in
   wire signed [9:0] m65_18;
   assign m65_18 ={ {5{neg65[5]}} , neg65[5:1] };

   // m65_19 = W*in
   wire signed [9:0] m65_19;
   assign m65_19 =10'b0;

   // m65_20 = W*in
   wire signed [9:0] m65_20;
   assign m65_20 =10'b0;

   // m65_21 = W*in
   wire signed [9:0] m65_21;
   assign m65_21 ={ {4{in65[5]}} , in65[5:0] };

   // m65_22 = W*in
   wire signed [9:0] m65_22;
   assign m65_22 ={ {5{neg65[5]}} , neg65[5:1] };

   // m65_23 = W*in
   wire signed [9:0] m65_23;
   assign m65_23 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_24 = W*in
   wire signed [9:0] m65_24;
   assign m65_24 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_25 = W*in
   wire signed [9:0] m65_25;
   assign m65_25 =10'b0;

   // m65_26 = W*in
   wire signed [9:0] m65_26;
   assign m65_26 =10'b0;

   // m65_27 = W*in
   wire signed [9:0] m65_27;
   assign m65_27 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_28 = W*in
   wire signed [9:0] m65_28;
   assign m65_28 =10'b0;

   // m65_29 = W*in
   wire signed [9:0] m65_29;
   assign m65_29 =10'b0;

   // m65_30 = W*in
   wire signed [9:0] m65_30;
   assign m65_30 =10'b0;

   // m65_31 = W*in
   wire signed [9:0] m65_31;
   assign m65_31 ={ {5{neg65[5]}} , neg65[5:1] };

   // m65_32 = W*in
   wire signed [9:0] m65_32;
   assign m65_32 ={ {4{in65[5]}} , in65[5:0] };

   // m65_33 = W*in
   wire signed [9:0] m65_33;
   assign m65_33 =10'b0;

   // m65_34 = W*in
   wire signed [9:0] m65_34;
   assign m65_34 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_35 = W*in
   wire signed [9:0] m65_35;
   assign m65_35 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_36 = W*in
   wire signed [9:0] m65_36;
   assign m65_36 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_37 = W*in
   wire signed [9:0] m65_37;
   assign m65_37 ={ {4{in65[5]}} , in65[5:0] };

   // m65_38 = W*in
   wire signed [9:0] m65_38;
   assign m65_38 ={ {5{in65[5]}} , in65[5:1] };

   // m65_39 = W*in
   wire signed [9:0] m65_39;
   assign m65_39 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_40 = W*in
   wire signed [9:0] m65_40;
   assign m65_40 =10'b0;

   // m65_41 = W*in
   wire signed [9:0] m65_41;
   assign m65_41 =10'b0;

   // m65_42 = W*in
   wire signed [9:0] m65_42;
   assign m65_42 ={ {4{in65[5]}} , in65[5:0] };

   // m65_43 = W*in
   wire signed [9:0] m65_43;
   assign m65_43 =10'b0;

   // m65_44 = W*in
   wire signed [9:0] m65_44;
   assign m65_44 =10'b0;

   // m65_45 = W*in
   wire signed [9:0] m65_45;
   assign m65_45 =10'b0;

   // m65_46 = W*in
   wire signed [9:0] m65_46;
   assign m65_46 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_47 = W*in
   wire signed [9:0] m65_47;
   assign m65_47 =10'b0;

   // m65_48 = W*in
   wire signed [9:0] m65_48;
   assign m65_48 =10'b0;

   // m65_49 = W*in
   wire signed [9:0] m65_49;
   assign m65_49 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_50 = W*in
   wire signed [9:0] m65_50;
   assign m65_50 =10'b0;

   // m65_51 = W*in
   wire signed [9:0] m65_51;
   assign m65_51 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_52 = W*in
   wire signed [9:0] m65_52;
   assign m65_52 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_53 = W*in
   wire signed [9:0] m65_53;
   assign m65_53 =10'b0;

   // m65_54 = W*in
   wire signed [9:0] m65_54;
   assign m65_54 ={ {4{in65[5]}} , in65[5:0] };

   // m65_55 = W*in
   wire signed [9:0] m65_55;
   assign m65_55 =10'b0;

   // m65_56 = W*in
   wire signed [9:0] m65_56;
   assign m65_56 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_57 = W*in
   wire signed [9:0] m65_57;
   assign m65_57 =10'b0;

   // m65_58 = W*in
   wire signed [9:0] m65_58;
   assign m65_58 =10'b0;

   // m65_59 = W*in
   wire signed [9:0] m65_59;
   assign m65_59 =10'b0;

   // m65_60 = W*in
   wire signed [9:0] m65_60;
   assign m65_60 =10'b0;

   // m65_61 = W*in
   wire signed [9:0] m65_61;
   assign m65_61 =10'b0;

   // m65_62 = W*in
   wire signed [9:0] m65_62;
   assign m65_62 =10'b0;

   // m65_63 = W*in
   wire signed [9:0] m65_63;
   assign m65_63 ={ {4{in65[5]}} , in65[5:0] };

   // m65_64 = W*in
   wire signed [9:0] m65_64;
   assign m65_64 ={ {4{in65[5]}} , in65[5:0] };

   // m65_65 = W*in
   wire signed [9:0] m65_65;
   assign m65_65 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_66 = W*in
   wire signed [9:0] m65_66;
   assign m65_66 ={ {4{in65[5]}} , in65[5:0] };

   // m65_67 = W*in
   wire signed [9:0] m65_67;
   assign m65_67 =10'b0;

   // m65_68 = W*in
   wire signed [9:0] m65_68;
   assign m65_68 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_69 = W*in
   wire signed [9:0] m65_69;
   assign m65_69 ={ {4{in65[5]}} , in65[5:0] };

   // m65_70 = W*in
   wire signed [9:0] m65_70;
   assign m65_70 =10'b0;

   // m65_71 = W*in
   wire signed [9:0] m65_71;
   assign m65_71 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_72 = W*in
   wire signed [9:0] m65_72;
   assign m65_72 =10'b0;

   // m65_73 = W*in
   wire signed [9:0] m65_73;
   assign m65_73 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_74 = W*in
   wire signed [9:0] m65_74;
   assign m65_74 =10'b0;

   // m65_75 = W*in
   wire signed [9:0] m65_75;
   assign m65_75 ={ {4{in65[5]}} , in65[5:0] };

   // m65_76 = W*in
   wire signed [9:0] m65_76;
   assign m65_76 =10'b0;

   // m65_77 = W*in
   wire signed [9:0] m65_77;
   assign m65_77 =10'b0;

   // m65_78 = W*in
   wire signed [9:0] m65_78;
   assign m65_78 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_79 = W*in
   wire signed [9:0] m65_79;
   assign m65_79 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_80 = W*in
   wire signed [9:0] m65_80;
   assign m65_80 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_81 = W*in
   wire signed [9:0] m65_81;
   assign m65_81 ={ {4{in65[5]}} , in65[5:0] };

   // m65_82 = W*in
   wire signed [9:0] m65_82;
   assign m65_82 ={ {4{in65[5]}} , in65[5:0] };

   // m65_83 = W*in
   wire signed [9:0] m65_83;
   assign m65_83 ={ {4{in65[5]}} , in65[5:0] };

   // m65_84 = W*in
   wire signed [9:0] m65_84;
   assign m65_84 =10'b0;

   // m65_85 = W*in
   wire signed [9:0] m65_85;
   assign m65_85 ={ {5{in65[5]}} , in65[5:1] };

   // m65_86 = W*in
   wire signed [9:0] m65_86;
   assign m65_86 =10'b0;

   // m65_87 = W*in
   wire signed [9:0] m65_87;
   assign m65_87 =10'b0;

   // m65_88 = W*in
   wire signed [9:0] m65_88;
   assign m65_88 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_89 = W*in
   wire signed [9:0] m65_89;
   assign m65_89 =10'b0;

   // m65_90 = W*in
   wire signed [9:0] m65_90;
   assign m65_90 ={ {3{neg65[5]}} , neg65 , {1{1'b0}} };

   // m65_91 = W*in
   wire signed [9:0] m65_91;
   assign m65_91 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_92 = W*in
   wire signed [9:0] m65_92;
   assign m65_92 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_93 = W*in
   wire signed [9:0] m65_93;
   assign m65_93 =10'b0;

   // m65_94 = W*in
   wire signed [9:0] m65_94;
   assign m65_94 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_95 = W*in
   wire signed [9:0] m65_95;
   assign m65_95 =10'b0;

   // m65_96 = W*in
   wire signed [9:0] m65_96;
   assign m65_96 =10'b0;

   // m65_97 = W*in
   wire signed [9:0] m65_97;
   assign m65_97 ={ {4{in65[5]}} , in65[5:0] };

   // m65_98 = W*in
   wire signed [9:0] m65_98;
   assign m65_98 =10'b0;

   // m65_99 = W*in
   wire signed [9:0] m65_99;
   assign m65_99 =10'b0;

   // m65_100 = W*in
   wire signed [9:0] m65_100;
   assign m65_100 ={ {4{in65[5]}} , in65[5:0] };

   // m65_101 = W*in
   wire signed [9:0] m65_101;
   assign m65_101 =10'b0;

   // m65_102 = W*in
   wire signed [9:0] m65_102;
   assign m65_102 =10'b0;

   // m65_103 = W*in
   wire signed [9:0] m65_103;
   assign m65_103 =10'b0;

   // m65_104 = W*in
   wire signed [9:0] m65_104;
   assign m65_104 =10'b0;

   // m65_105 = W*in
   wire signed [9:0] m65_105;
   assign m65_105 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_106 = W*in
   wire signed [9:0] m65_106;
   assign m65_106 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_107 = W*in
   wire signed [9:0] m65_107;
   assign m65_107 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_108 = W*in
   wire signed [9:0] m65_108;
   assign m65_108 =10'b0;

   // m65_109 = W*in
   wire signed [9:0] m65_109;
   assign m65_109 =10'b0;

   // m65_110 = W*in
   wire signed [9:0] m65_110;
   assign m65_110 =10'b0;

   // m65_111 = W*in
   wire signed [9:0] m65_111;
   assign m65_111 ={ {4{neg65[5]}} , neg65[5:0] };

   // m65_112 = W*in
   wire signed [9:0] m65_112;
   assign m65_112 ={ {3{in65[5]}} , in65 , {1{1'b0}} };

   // m65_113 = W*in
   wire signed [9:0] m65_113;
   assign m65_113 =10'b0;

   // m65_114 = W*in
   wire signed [9:0] m65_114;
   assign m65_114 =10'b0;

   // m65_115 = W*in
   wire signed [9:0] m65_115;
   assign m65_115 =10'b0;

   // m65_116 = W*in
   wire signed [9:0] m65_116;
   assign m65_116 =10'b0;

   // m65_117 = W*in
   wire signed [9:0] m65_117;
   assign m65_117 =10'b0;

   // m66_1 = W*in
   wire signed [9:0] m66_1;
   assign m66_1 =10'b0;

   // m66_2 = W*in
   wire signed [9:0] m66_2;
   assign m66_2 =10'b0;

   // m66_3 = W*in
   wire signed [9:0] m66_3;
   assign m66_3 ={ {3{neg66[5]}} , neg66 , {1{1'b0}} };

   // m66_4 = W*in
   wire signed [9:0] m66_4;
   assign m66_4 =10'b0;

   // m66_5 = W*in
   wire signed [9:0] m66_5;
   assign m66_5 =10'b0;

   // m66_6 = W*in
   wire signed [9:0] m66_6;
   assign m66_6 =10'b0;

   // m66_7 = W*in
   wire signed [9:0] m66_7;
   assign m66_7 =10'b0;

   // m66_8 = W*in
   wire signed [9:0] m66_8;
   assign m66_8 =10'b0;

   // m66_9 = W*in
   wire signed [9:0] m66_9;
   assign m66_9 =10'b0;

   // m66_10 = W*in
   wire signed [9:0] m66_10;
   assign m66_10 =10'b0;

   // m66_11 = W*in
   wire signed [9:0] m66_11;
   assign m66_11 =10'b0;

   // m66_12 = W*in
   wire signed [9:0] m66_12;
   assign m66_12 =10'b0;

   // m66_13 = W*in
   wire signed [9:0] m66_13;
   assign m66_13 =10'b0;

   // m66_14 = W*in
   wire signed [9:0] m66_14;
   assign m66_14 =10'b0;

   // m66_15 = W*in
   wire signed [9:0] m66_15;
   assign m66_15 =10'b0;

   // m66_16 = W*in
   wire signed [9:0] m66_16;
   assign m66_16 =10'b0;

   // m66_17 = W*in
   wire signed [9:0] m66_17;
   assign m66_17 ={ {5{neg66[5]}} , neg66[5:1] };

   // m66_18 = W*in
   wire signed [9:0] m66_18;
   assign m66_18 ={ {5{in66[5]}} , in66[5:1] };

   // m66_19 = W*in
   wire signed [9:0] m66_19;
   assign m66_19 =10'b0;

   // m66_20 = W*in
   wire signed [9:0] m66_20;
   assign m66_20 =10'b0;

   // m66_21 = W*in
   wire signed [9:0] m66_21;
   assign m66_21 =10'b0;

   // m66_22 = W*in
   wire signed [9:0] m66_22;
   assign m66_22 =10'b0;

   // m66_23 = W*in
   wire signed [9:0] m66_23;
   assign m66_23 ={ {5{neg66[5]}} , neg66[5:1] };

   // m66_24 = W*in
   wire signed [9:0] m66_24;
   assign m66_24 =10'b0;

   // m66_25 = W*in
   wire signed [9:0] m66_25;
   assign m66_25 ={ {4{in66[5]}} , in66[5:0] };

   // m66_26 = W*in
   wire signed [9:0] m66_26;
   assign m66_26 ={ {5{in66[5]}} , in66[5:1] };

   // m66_27 = W*in
   wire signed [9:0] m66_27;
   assign m66_27 =10'b0;

   // m66_28 = W*in
   wire signed [9:0] m66_28;
   assign m66_28 =10'b0;

   // m66_29 = W*in
   wire signed [9:0] m66_29;
   assign m66_29 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_30 = W*in
   wire signed [9:0] m66_30;
   assign m66_30 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_31 = W*in
   wire signed [9:0] m66_31;
   assign m66_31 ={ {5{neg66[5]}} , neg66[5:1] };

   // m66_32 = W*in
   wire signed [9:0] m66_32;
   assign m66_32 =10'b0;

   // m66_33 = W*in
   wire signed [9:0] m66_33;
   assign m66_33 =10'b0;

   // m66_34 = W*in
   wire signed [9:0] m66_34;
   assign m66_34 =10'b0;

   // m66_35 = W*in
   wire signed [9:0] m66_35;
   assign m66_35 =10'b0;

   // m66_36 = W*in
   wire signed [9:0] m66_36;
   assign m66_36 ={ {5{neg66[5]}} , neg66[5:1] };

   // m66_37 = W*in
   wire signed [9:0] m66_37;
   assign m66_37 ={ {4{in66[5]}} , in66[5:0] };

   // m66_38 = W*in
   wire signed [9:0] m66_38;
   assign m66_38 =10'b0;

   // m66_39 = W*in
   wire signed [9:0] m66_39;
   assign m66_39 =10'b0;

   // m66_40 = W*in
   wire signed [9:0] m66_40;
   assign m66_40 ={ {5{in66[5]}} , in66[5:1] };

   // m66_41 = W*in
   wire signed [9:0] m66_41;
   assign m66_41 =10'b0;

   // m66_42 = W*in
   wire signed [9:0] m66_42;
   assign m66_42 =10'b0;

   // m66_43 = W*in
   wire signed [9:0] m66_43;
   assign m66_43 =10'b0;

   // m66_44 = W*in
   wire signed [9:0] m66_44;
   assign m66_44 =10'b0;

   // m66_45 = W*in
   wire signed [9:0] m66_45;
   assign m66_45 =10'b0;

   // m66_46 = W*in
   wire signed [9:0] m66_46;
   assign m66_46 =10'b0;

   // m66_47 = W*in
   wire signed [9:0] m66_47;
   assign m66_47 =10'b0;

   // m66_48 = W*in
   wire signed [9:0] m66_48;
   assign m66_48 =10'b0;

   // m66_49 = W*in
   wire signed [9:0] m66_49;
   assign m66_49 =10'b0;

   // m66_50 = W*in
   wire signed [9:0] m66_50;
   assign m66_50 =10'b0;

   // m66_51 = W*in
   wire signed [9:0] m66_51;
   assign m66_51 =10'b0;

   // m66_52 = W*in
   wire signed [9:0] m66_52;
   assign m66_52 =10'b0;

   // m66_53 = W*in
   wire signed [9:0] m66_53;
   assign m66_53 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_54 = W*in
   wire signed [9:0] m66_54;
   assign m66_54 =10'b0;

   // m66_55 = W*in
   wire signed [9:0] m66_55;
   assign m66_55 =10'b0;

   // m66_56 = W*in
   wire signed [9:0] m66_56;
   assign m66_56 =10'b0;

   // m66_57 = W*in
   wire signed [9:0] m66_57;
   assign m66_57 =10'b0;

   // m66_58 = W*in
   wire signed [9:0] m66_58;
   assign m66_58 =10'b0;

   // m66_59 = W*in
   wire signed [9:0] m66_59;
   assign m66_59 =10'b0;

   // m66_60 = W*in
   wire signed [9:0] m66_60;
   assign m66_60 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_61 = W*in
   wire signed [9:0] m66_61;
   assign m66_61 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_62 = W*in
   wire signed [9:0] m66_62;
   assign m66_62 =10'b0;

   // m66_63 = W*in
   wire signed [9:0] m66_63;
   assign m66_63 =10'b0;

   // m66_64 = W*in
   wire signed [9:0] m66_64;
   assign m66_64 =10'b0;

   // m66_65 = W*in
   wire signed [9:0] m66_65;
   assign m66_65 ={ {4{in66[5]}} , in66[5:0] };

   // m66_66 = W*in
   wire signed [9:0] m66_66;
   assign m66_66 =10'b0;

   // m66_67 = W*in
   wire signed [9:0] m66_67;
   assign m66_67 =10'b0;

   // m66_68 = W*in
   wire signed [9:0] m66_68;
   assign m66_68 =10'b0;

   // m66_69 = W*in
   wire signed [9:0] m66_69;
   assign m66_69 ={ {5{in66[5]}} , in66[5:1] };

   // m66_70 = W*in
   wire signed [9:0] m66_70;
   assign m66_70 =10'b0;

   // m66_71 = W*in
   wire signed [9:0] m66_71;
   assign m66_71 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_72 = W*in
   wire signed [9:0] m66_72;
   assign m66_72 =10'b0;

   // m66_73 = W*in
   wire signed [9:0] m66_73;
   assign m66_73 =10'b0;

   // m66_74 = W*in
   wire signed [9:0] m66_74;
   assign m66_74 =10'b0;

   // m66_75 = W*in
   wire signed [9:0] m66_75;
   assign m66_75 =10'b0;

   // m66_76 = W*in
   wire signed [9:0] m66_76;
   assign m66_76 =10'b0;

   // m66_77 = W*in
   wire signed [9:0] m66_77;
   assign m66_77 ={ {4{in66[5]}} , in66[5:0] };

   // m66_78 = W*in
   wire signed [9:0] m66_78;
   assign m66_78 =10'b0;

   // m66_79 = W*in
   wire signed [9:0] m66_79;
   assign m66_79 =10'b0;

   // m66_80 = W*in
   wire signed [9:0] m66_80;
   assign m66_80 =10'b0;

   // m66_81 = W*in
   wire signed [9:0] m66_81;
   assign m66_81 ={ {4{in66[5]}} , in66[5:0] };

   // m66_82 = W*in
   wire signed [9:0] m66_82;
   assign m66_82 =10'b0;

   // m66_83 = W*in
   wire signed [9:0] m66_83;
   assign m66_83 =10'b0;

   // m66_84 = W*in
   wire signed [9:0] m66_84;
   assign m66_84 =10'b0;

   // m66_85 = W*in
   wire signed [9:0] m66_85;
   assign m66_85 =10'b0;

   // m66_86 = W*in
   wire signed [9:0] m66_86;
   assign m66_86 ={ {4{in66[5]}} , in66[5:0] };

   // m66_87 = W*in
   wire signed [9:0] m66_87;
   assign m66_87 =10'b0;

   // m66_88 = W*in
   wire signed [9:0] m66_88;
   assign m66_88 =10'b0;

   // m66_89 = W*in
   wire signed [9:0] m66_89;
   assign m66_89 =10'b0;

   // m66_90 = W*in
   wire signed [9:0] m66_90;
   assign m66_90 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_91 = W*in
   wire signed [9:0] m66_91;
   assign m66_91 ={ {3{in66[5]}} , in66 , {1{1'b0}} };

   // m66_92 = W*in
   wire signed [9:0] m66_92;
   assign m66_92 =10'b0;

   // m66_93 = W*in
   wire signed [9:0] m66_93;
   assign m66_93 =10'b0;

   // m66_94 = W*in
   wire signed [9:0] m66_94;
   assign m66_94 =10'b0;

   // m66_95 = W*in
   wire signed [9:0] m66_95;
   assign m66_95 =10'b0;

   // m66_96 = W*in
   wire signed [9:0] m66_96;
   assign m66_96 =10'b0;

   // m66_97 = W*in
   wire signed [9:0] m66_97;
   assign m66_97 =10'b0;

   // m66_98 = W*in
   wire signed [9:0] m66_98;
   assign m66_98 =10'b0;

   // m66_99 = W*in
   wire signed [9:0] m66_99;
   assign m66_99 =10'b0;

   // m66_100 = W*in
   wire signed [9:0] m66_100;
   assign m66_100 =10'b0;

   // m66_101 = W*in
   wire signed [9:0] m66_101;
   assign m66_101 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_102 = W*in
   wire signed [9:0] m66_102;
   assign m66_102 =10'b0;

   // m66_103 = W*in
   wire signed [9:0] m66_103;
   assign m66_103 =10'b0;

   // m66_104 = W*in
   wire signed [9:0] m66_104;
   assign m66_104 =10'b0;

   // m66_105 = W*in
   wire signed [9:0] m66_105;
   assign m66_105 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_106 = W*in
   wire signed [9:0] m66_106;
   assign m66_106 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_107 = W*in
   wire signed [9:0] m66_107;
   assign m66_107 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_108 = W*in
   wire signed [9:0] m66_108;
   assign m66_108 ={ {4{neg66[5]}} , neg66[5:0] };

   // m66_109 = W*in
   wire signed [9:0] m66_109;
   assign m66_109 ={ {5{neg66[5]}} , neg66[5:1] };

   // m66_110 = W*in
   wire signed [9:0] m66_110;
   assign m66_110 =10'b0;

   // m66_111 = W*in
   wire signed [9:0] m66_111;
   assign m66_111 =10'b0;

   // m66_112 = W*in
   wire signed [9:0] m66_112;
   assign m66_112 =10'b0;

   // m66_113 = W*in
   wire signed [9:0] m66_113;
   assign m66_113 =10'b0;

   // m66_114 = W*in
   wire signed [9:0] m66_114;
   assign m66_114 =10'b0;

   // m66_115 = W*in
   wire signed [9:0] m66_115;
   assign m66_115 =10'b0;

   // m66_116 = W*in
   wire signed [9:0] m66_116;
   assign m66_116 =10'b0;

   // m66_117 = W*in
   wire signed [9:0] m66_117;
   assign m66_117 ={ {4{neg66[5]}} , neg66[5:0] };

   // m67_1 = W*in
   wire signed [9:0] m67_1;
   assign m67_1 =10'b0;

   // m67_2 = W*in
   wire signed [9:0] m67_2;
   assign m67_2 =10'b0;

   // m67_3 = W*in
   wire signed [9:0] m67_3;
   assign m67_3 =10'b0;

   // m67_4 = W*in
   wire signed [9:0] m67_4;
   assign m67_4 =10'b0;

   // m67_5 = W*in
   wire signed [9:0] m67_5;
   assign m67_5 =10'b0;

   // m67_6 = W*in
   wire signed [9:0] m67_6;
   assign m67_6 =10'b0;

   // m67_7 = W*in
   wire signed [9:0] m67_7;
   assign m67_7 =10'b0;

   // m67_8 = W*in
   wire signed [9:0] m67_8;
   assign m67_8 =10'b0;

   // m67_9 = W*in
   wire signed [9:0] m67_9;
   assign m67_9 =10'b0;

   // m67_10 = W*in
   wire signed [9:0] m67_10;
   assign m67_10 =10'b0;

   // m67_11 = W*in
   wire signed [9:0] m67_11;
   assign m67_11 =10'b0;

   // m67_12 = W*in
   wire signed [9:0] m67_12;
   assign m67_12 =10'b0;

   // m67_13 = W*in
   wire signed [9:0] m67_13;
   assign m67_13 =10'b0;

   // m67_14 = W*in
   wire signed [9:0] m67_14;
   assign m67_14 =10'b0;

   // m67_15 = W*in
   wire signed [9:0] m67_15;
   assign m67_15 =10'b0;

   // m67_16 = W*in
   wire signed [9:0] m67_16;
   assign m67_16 =10'b0;

   // m67_17 = W*in
   wire signed [9:0] m67_17;
   assign m67_17 =10'b0;

   // m67_18 = W*in
   wire signed [9:0] m67_18;
   assign m67_18 ={ {5{in67[5]}} , in67[5:1] };

   // m67_19 = W*in
   wire signed [9:0] m67_19;
   assign m67_19 =10'b0;

   // m67_20 = W*in
   wire signed [9:0] m67_20;
   assign m67_20 ={ {5{in67[5]}} , in67[5:1] };

   // m67_21 = W*in
   wire signed [9:0] m67_21;
   assign m67_21 =10'b0;

   // m67_22 = W*in
   wire signed [9:0] m67_22;
   assign m67_22 =10'b0;

   // m67_23 = W*in
   wire signed [9:0] m67_23;
   assign m67_23 =10'b0;

   // m67_24 = W*in
   wire signed [9:0] m67_24;
   assign m67_24 =10'b0;

   // m67_25 = W*in
   wire signed [9:0] m67_25;
   assign m67_25 =10'b0;

   // m67_26 = W*in
   wire signed [9:0] m67_26;
   assign m67_26 =10'b0;

   // m67_27 = W*in
   wire signed [9:0] m67_27;
   assign m67_27 =10'b0;

   // m67_28 = W*in
   wire signed [9:0] m67_28;
   assign m67_28 =10'b0;

   // m67_29 = W*in
   wire signed [9:0] m67_29;
   assign m67_29 ={ {5{neg67[5]}} , neg67[5:1] };

   // m67_30 = W*in
   wire signed [9:0] m67_30;
   assign m67_30 =10'b0;

   // m67_31 = W*in
   wire signed [9:0] m67_31;
   assign m67_31 =10'b0;

   // m67_32 = W*in
   wire signed [9:0] m67_32;
   assign m67_32 =10'b0;

   // m67_33 = W*in
   wire signed [9:0] m67_33;
   assign m67_33 =10'b0;

   // m67_34 = W*in
   wire signed [9:0] m67_34;
   assign m67_34 =10'b0;

   // m67_35 = W*in
   wire signed [9:0] m67_35;
   assign m67_35 ={ {5{in67[5]}} , in67[5:1] };

   // m67_36 = W*in
   wire signed [9:0] m67_36;
   assign m67_36 =10'b0;

   // m67_37 = W*in
   wire signed [9:0] m67_37;
   assign m67_37 =10'b0;

   // m67_38 = W*in
   wire signed [9:0] m67_38;
   assign m67_38 =10'b0;

   // m67_39 = W*in
   wire signed [9:0] m67_39;
   assign m67_39 =10'b0;

   // m67_40 = W*in
   wire signed [9:0] m67_40;
   assign m67_40 =10'b0;

   // m67_41 = W*in
   wire signed [9:0] m67_41;
   assign m67_41 =10'b0;

   // m67_42 = W*in
   wire signed [9:0] m67_42;
   assign m67_42 =10'b0;

   // m67_43 = W*in
   wire signed [9:0] m67_43;
   assign m67_43 =10'b0;

   // m67_44 = W*in
   wire signed [9:0] m67_44;
   assign m67_44 =10'b0;

   // m67_45 = W*in
   wire signed [9:0] m67_45;
   assign m67_45 =10'b0;

   // m67_46 = W*in
   wire signed [9:0] m67_46;
   assign m67_46 =10'b0;

   // m67_47 = W*in
   wire signed [9:0] m67_47;
   assign m67_47 =10'b0;

   // m67_48 = W*in
   wire signed [9:0] m67_48;
   assign m67_48 =10'b0;

   // m67_49 = W*in
   wire signed [9:0] m67_49;
   assign m67_49 =10'b0;

   // m67_50 = W*in
   wire signed [9:0] m67_50;
   assign m67_50 =10'b0;

   // m67_51 = W*in
   wire signed [9:0] m67_51;
   assign m67_51 =10'b0;

   // m67_52 = W*in
   wire signed [9:0] m67_52;
   assign m67_52 =10'b0;

   // m67_53 = W*in
   wire signed [9:0] m67_53;
   assign m67_53 =10'b0;

   // m67_54 = W*in
   wire signed [9:0] m67_54;
   assign m67_54 =10'b0;

   // m67_55 = W*in
   wire signed [9:0] m67_55;
   assign m67_55 =10'b0;

   // m67_56 = W*in
   wire signed [9:0] m67_56;
   assign m67_56 =10'b0;

   // m67_57 = W*in
   wire signed [9:0] m67_57;
   assign m67_57 =10'b0;

   // m67_58 = W*in
   wire signed [9:0] m67_58;
   assign m67_58 =10'b0;

   // m67_59 = W*in
   wire signed [9:0] m67_59;
   assign m67_59 =10'b0;

   // m67_60 = W*in
   wire signed [9:0] m67_60;
   assign m67_60 =10'b0;

   // m67_61 = W*in
   wire signed [9:0] m67_61;
   assign m67_61 =10'b0;

   // m67_62 = W*in
   wire signed [9:0] m67_62;
   assign m67_62 =10'b0;

   // m67_63 = W*in
   wire signed [9:0] m67_63;
   assign m67_63 =10'b0;

   // m67_64 = W*in
   wire signed [9:0] m67_64;
   assign m67_64 ={ {5{in67[5]}} , in67[5:1] };

   // m67_65 = W*in
   wire signed [9:0] m67_65;
   assign m67_65 =10'b0;

   // m67_66 = W*in
   wire signed [9:0] m67_66;
   assign m67_66 =10'b0;

   // m67_67 = W*in
   wire signed [9:0] m67_67;
   assign m67_67 =10'b0;

   // m67_68 = W*in
   wire signed [9:0] m67_68;
   assign m67_68 =10'b0;

   // m67_69 = W*in
   wire signed [9:0] m67_69;
   assign m67_69 =10'b0;

   // m67_70 = W*in
   wire signed [9:0] m67_70;
   assign m67_70 =10'b0;

   // m67_71 = W*in
   wire signed [9:0] m67_71;
   assign m67_71 =10'b0;

   // m67_72 = W*in
   wire signed [9:0] m67_72;
   assign m67_72 ={ {5{in67[5]}} , in67[5:1] };

   // m67_73 = W*in
   wire signed [9:0] m67_73;
   assign m67_73 =10'b0;

   // m67_74 = W*in
   wire signed [9:0] m67_74;
   assign m67_74 =10'b0;

   // m67_75 = W*in
   wire signed [9:0] m67_75;
   assign m67_75 =10'b0;

   // m67_76 = W*in
   wire signed [9:0] m67_76;
   assign m67_76 =10'b0;

   // m67_77 = W*in
   wire signed [9:0] m67_77;
   assign m67_77 ={ {4{in67[5]}} , in67[5:0] };

   // m67_78 = W*in
   wire signed [9:0] m67_78;
   assign m67_78 =10'b0;

   // m67_79 = W*in
   wire signed [9:0] m67_79;
   assign m67_79 =10'b0;

   // m67_80 = W*in
   wire signed [9:0] m67_80;
   assign m67_80 =10'b0;

   // m67_81 = W*in
   wire signed [9:0] m67_81;
   assign m67_81 ={ {5{in67[5]}} , in67[5:1] };

   // m67_82 = W*in
   wire signed [9:0] m67_82;
   assign m67_82 =10'b0;

   // m67_83 = W*in
   wire signed [9:0] m67_83;
   assign m67_83 =10'b0;

   // m67_84 = W*in
   wire signed [9:0] m67_84;
   assign m67_84 =10'b0;

   // m67_85 = W*in
   wire signed [9:0] m67_85;
   assign m67_85 =10'b0;

   // m67_86 = W*in
   wire signed [9:0] m67_86;
   assign m67_86 =10'b0;

   // m67_87 = W*in
   wire signed [9:0] m67_87;
   assign m67_87 =10'b0;

   // m67_88 = W*in
   wire signed [9:0] m67_88;
   assign m67_88 =10'b0;

   // m67_89 = W*in
   wire signed [9:0] m67_89;
   assign m67_89 =10'b0;

   // m67_90 = W*in
   wire signed [9:0] m67_90;
   assign m67_90 =10'b0;

   // m67_91 = W*in
   wire signed [9:0] m67_91;
   assign m67_91 =10'b0;

   // m67_92 = W*in
   wire signed [9:0] m67_92;
   assign m67_92 =10'b0;

   // m67_93 = W*in
   wire signed [9:0] m67_93;
   assign m67_93 =10'b0;

   // m67_94 = W*in
   wire signed [9:0] m67_94;
   assign m67_94 =10'b0;

   // m67_95 = W*in
   wire signed [9:0] m67_95;
   assign m67_95 =10'b0;

   // m67_96 = W*in
   wire signed [9:0] m67_96;
   assign m67_96 =10'b0;

   // m67_97 = W*in
   wire signed [9:0] m67_97;
   assign m67_97 =10'b0;

   // m67_98 = W*in
   wire signed [9:0] m67_98;
   assign m67_98 =10'b0;

   // m67_99 = W*in
   wire signed [9:0] m67_99;
   assign m67_99 =10'b0;

   // m67_100 = W*in
   wire signed [9:0] m67_100;
   assign m67_100 =10'b0;

   // m67_101 = W*in
   wire signed [9:0] m67_101;
   assign m67_101 =10'b0;

   // m67_102 = W*in
   wire signed [9:0] m67_102;
   assign m67_102 =10'b0;

   // m67_103 = W*in
   wire signed [9:0] m67_103;
   assign m67_103 =10'b0;

   // m67_104 = W*in
   wire signed [9:0] m67_104;
   assign m67_104 =10'b0;

   // m67_105 = W*in
   wire signed [9:0] m67_105;
   assign m67_105 =10'b0;

   // m67_106 = W*in
   wire signed [9:0] m67_106;
   assign m67_106 =10'b0;

   // m67_107 = W*in
   wire signed [9:0] m67_107;
   assign m67_107 =10'b0;

   // m67_108 = W*in
   wire signed [9:0] m67_108;
   assign m67_108 =10'b0;

   // m67_109 = W*in
   wire signed [9:0] m67_109;
   assign m67_109 =10'b0;

   // m67_110 = W*in
   wire signed [9:0] m67_110;
   assign m67_110 =10'b0;

   // m67_111 = W*in
   wire signed [9:0] m67_111;
   assign m67_111 =10'b0;

   // m67_112 = W*in
   wire signed [9:0] m67_112;
   assign m67_112 =10'b0;

   // m67_113 = W*in
   wire signed [9:0] m67_113;
   assign m67_113 =10'b0;

   // m67_114 = W*in
   wire signed [9:0] m67_114;
   assign m67_114 =10'b0;

   // m67_115 = W*in
   wire signed [9:0] m67_115;
   assign m67_115 ={ {5{in67[5]}} , in67[5:1] };

   // m67_116 = W*in
   wire signed [9:0] m67_116;
   assign m67_116 =10'b0;

   // m67_117 = W*in
   wire signed [9:0] m67_117;
   assign m67_117 =10'b0;

   // m68_1 = W*in
   wire signed [9:0] m68_1;
   assign m68_1 =10'b0;

   // m68_2 = W*in
   wire signed [9:0] m68_2;
   assign m68_2 =10'b0;

   // m68_3 = W*in
   wire signed [9:0] m68_3;
   assign m68_3 =10'b0;

   // m68_4 = W*in
   wire signed [9:0] m68_4;
   assign m68_4 =10'b0;

   // m68_5 = W*in
   wire signed [9:0] m68_5;
   assign m68_5 =10'b0;

   // m68_6 = W*in
   wire signed [9:0] m68_6;
   assign m68_6 =10'b0;

   // m68_7 = W*in
   wire signed [9:0] m68_7;
   assign m68_7 =10'b0;

   // m68_8 = W*in
   wire signed [9:0] m68_8;
   assign m68_8 =10'b0;

   // m68_9 = W*in
   wire signed [9:0] m68_9;
   assign m68_9 =10'b0;

   // m68_10 = W*in
   wire signed [9:0] m68_10;
   assign m68_10 =10'b0;

   // m68_11 = W*in
   wire signed [9:0] m68_11;
   assign m68_11 =10'b0;

   // m68_12 = W*in
   wire signed [9:0] m68_12;
   assign m68_12 =10'b0;

   // m68_13 = W*in
   wire signed [9:0] m68_13;
   assign m68_13 =10'b0;

   // m68_14 = W*in
   wire signed [9:0] m68_14;
   assign m68_14 =10'b0;

   // m68_15 = W*in
   wire signed [9:0] m68_15;
   assign m68_15 =10'b0;

   // m68_16 = W*in
   wire signed [9:0] m68_16;
   assign m68_16 =10'b0;

   // m68_17 = W*in
   wire signed [9:0] m68_17;
   assign m68_17 =10'b0;

   // m68_18 = W*in
   wire signed [9:0] m68_18;
   assign m68_18 =10'b0;

   // m68_19 = W*in
   wire signed [9:0] m68_19;
   assign m68_19 ={ {4{in68[5]}} , in68[5:0] };

   // m68_20 = W*in
   wire signed [9:0] m68_20;
   assign m68_20 ={ {4{neg68[5]}} , neg68[5:0] };

   // m68_21 = W*in
   wire signed [9:0] m68_21;
   assign m68_21 =10'b0;

   // m68_22 = W*in
   wire signed [9:0] m68_22;
   assign m68_22 =10'b0;

   // m68_23 = W*in
   wire signed [9:0] m68_23;
   assign m68_23 =10'b0;

   // m68_24 = W*in
   wire signed [9:0] m68_24;
   assign m68_24 =10'b0;

   // m68_25 = W*in
   wire signed [9:0] m68_25;
   assign m68_25 =10'b0;

   // m68_26 = W*in
   wire signed [9:0] m68_26;
   assign m68_26 =10'b0;

   // m68_27 = W*in
   wire signed [9:0] m68_27;
   assign m68_27 ={ {4{neg68[5]}} , neg68[5:0] };

   // m68_28 = W*in
   wire signed [9:0] m68_28;
   assign m68_28 ={ {5{neg68[5]}} , neg68[5:1] };

   // m68_29 = W*in
   wire signed [9:0] m68_29;
   assign m68_29 =10'b0;

   // m68_30 = W*in
   wire signed [9:0] m68_30;
   assign m68_30 =10'b0;

   // m68_31 = W*in
   wire signed [9:0] m68_31;
   assign m68_31 ={ {5{neg68[5]}} , neg68[5:1] };

   // m68_32 = W*in
   wire signed [9:0] m68_32;
   assign m68_32 =10'b0;

   // m68_33 = W*in
   wire signed [9:0] m68_33;
   assign m68_33 =10'b0;

   // m68_34 = W*in
   wire signed [9:0] m68_34;
   assign m68_34 =10'b0;

   // m68_35 = W*in
   wire signed [9:0] m68_35;
   assign m68_35 ={ {5{neg68[5]}} , neg68[5:1] };

   // m68_36 = W*in
   wire signed [9:0] m68_36;
   assign m68_36 =10'b0;

   // m68_37 = W*in
   wire signed [9:0] m68_37;
   assign m68_37 =10'b0;

   // m68_38 = W*in
   wire signed [9:0] m68_38;
   assign m68_38 =10'b0;

   // m68_39 = W*in
   wire signed [9:0] m68_39;
   assign m68_39 =10'b0;

   // m68_40 = W*in
   wire signed [9:0] m68_40;
   assign m68_40 =10'b0;

   // m68_41 = W*in
   wire signed [9:0] m68_41;
   assign m68_41 =10'b0;

   // m68_42 = W*in
   wire signed [9:0] m68_42;
   assign m68_42 =10'b0;

   // m68_43 = W*in
   wire signed [9:0] m68_43;
   assign m68_43 =10'b0;

   // m68_44 = W*in
   wire signed [9:0] m68_44;
   assign m68_44 =10'b0;

   // m68_45 = W*in
   wire signed [9:0] m68_45;
   assign m68_45 =10'b0;

   // m68_46 = W*in
   wire signed [9:0] m68_46;
   assign m68_46 =10'b0;

   // m68_47 = W*in
   wire signed [9:0] m68_47;
   assign m68_47 =10'b0;

   // m68_48 = W*in
   wire signed [9:0] m68_48;
   assign m68_48 =10'b0;

   // m68_49 = W*in
   wire signed [9:0] m68_49;
   assign m68_49 =10'b0;

   // m68_50 = W*in
   wire signed [9:0] m68_50;
   assign m68_50 =10'b0;

   // m68_51 = W*in
   wire signed [9:0] m68_51;
   assign m68_51 =10'b0;

   // m68_52 = W*in
   wire signed [9:0] m68_52;
   assign m68_52 =10'b0;

   // m68_53 = W*in
   wire signed [9:0] m68_53;
   assign m68_53 =10'b0;

   // m68_54 = W*in
   wire signed [9:0] m68_54;
   assign m68_54 =10'b0;

   // m68_55 = W*in
   wire signed [9:0] m68_55;
   assign m68_55 =10'b0;

   // m68_56 = W*in
   wire signed [9:0] m68_56;
   assign m68_56 =10'b0;

   // m68_57 = W*in
   wire signed [9:0] m68_57;
   assign m68_57 =10'b0;

   // m68_58 = W*in
   wire signed [9:0] m68_58;
   assign m68_58 =10'b0;

   // m68_59 = W*in
   wire signed [9:0] m68_59;
   assign m68_59 =10'b0;

   // m68_60 = W*in
   wire signed [9:0] m68_60;
   assign m68_60 =10'b0;

   // m68_61 = W*in
   wire signed [9:0] m68_61;
   assign m68_61 =10'b0;

   // m68_62 = W*in
   wire signed [9:0] m68_62;
   assign m68_62 =10'b0;

   // m68_63 = W*in
   wire signed [9:0] m68_63;
   assign m68_63 ={ {4{in68[5]}} , in68[5:0] };

   // m68_64 = W*in
   wire signed [9:0] m68_64;
   assign m68_64 ={ {4{neg68[5]}} , neg68[5:0] };

   // m68_65 = W*in
   wire signed [9:0] m68_65;
   assign m68_65 =10'b0;

   // m68_66 = W*in
   wire signed [9:0] m68_66;
   assign m68_66 ={ {5{neg68[5]}} , neg68[5:1] };

   // m68_67 = W*in
   wire signed [9:0] m68_67;
   assign m68_67 ={ {4{in68[5]}} , in68[5:0] };

   // m68_68 = W*in
   wire signed [9:0] m68_68;
   assign m68_68 =10'b0;

   // m68_69 = W*in
   wire signed [9:0] m68_69;
   assign m68_69 ={ {4{neg68[5]}} , neg68[5:0] };

   // m68_70 = W*in
   wire signed [9:0] m68_70;
   assign m68_70 =10'b0;

   // m68_71 = W*in
   wire signed [9:0] m68_71;
   assign m68_71 =10'b0;

   // m68_72 = W*in
   wire signed [9:0] m68_72;
   assign m68_72 ={ {5{in68[5]}} , in68[5:1] };

   // m68_73 = W*in
   wire signed [9:0] m68_73;
   assign m68_73 =10'b0;

   // m68_74 = W*in
   wire signed [9:0] m68_74;
   assign m68_74 ={ {5{neg68[5]}} , neg68[5:1] };

   // m68_75 = W*in
   wire signed [9:0] m68_75;
   assign m68_75 =10'b0;

   // m68_76 = W*in
   wire signed [9:0] m68_76;
   assign m68_76 =10'b0;

   // m68_77 = W*in
   wire signed [9:0] m68_77;
   assign m68_77 =10'b0;

   // m68_78 = W*in
   wire signed [9:0] m68_78;
   assign m68_78 =10'b0;

   // m68_79 = W*in
   wire signed [9:0] m68_79;
   assign m68_79 =10'b0;

   // m68_80 = W*in
   wire signed [9:0] m68_80;
   assign m68_80 =10'b0;

   // m68_81 = W*in
   wire signed [9:0] m68_81;
   assign m68_81 ={ {5{neg68[5]}} , neg68[5:1] };

   // m68_82 = W*in
   wire signed [9:0] m68_82;
   assign m68_82 =10'b0;

   // m68_83 = W*in
   wire signed [9:0] m68_83;
   assign m68_83 =10'b0;

   // m68_84 = W*in
   wire signed [9:0] m68_84;
   assign m68_84 =10'b0;

   // m68_85 = W*in
   wire signed [9:0] m68_85;
   assign m68_85 =10'b0;

   // m68_86 = W*in
   wire signed [9:0] m68_86;
   assign m68_86 =10'b0;

   // m68_87 = W*in
   wire signed [9:0] m68_87;
   assign m68_87 =10'b0;

   // m68_88 = W*in
   wire signed [9:0] m68_88;
   assign m68_88 =10'b0;

   // m68_89 = W*in
   wire signed [9:0] m68_89;
   assign m68_89 =10'b0;

   // m68_90 = W*in
   wire signed [9:0] m68_90;
   assign m68_90 =10'b0;

   // m68_91 = W*in
   wire signed [9:0] m68_91;
   assign m68_91 =10'b0;

   // m68_92 = W*in
   wire signed [9:0] m68_92;
   assign m68_92 =10'b0;

   // m68_93 = W*in
   wire signed [9:0] m68_93;
   assign m68_93 =10'b0;

   // m68_94 = W*in
   wire signed [9:0] m68_94;
   assign m68_94 =10'b0;

   // m68_95 = W*in
   wire signed [9:0] m68_95;
   assign m68_95 =10'b0;

   // m68_96 = W*in
   wire signed [9:0] m68_96;
   assign m68_96 =10'b0;

   // m68_97 = W*in
   wire signed [9:0] m68_97;
   assign m68_97 =10'b0;

   // m68_98 = W*in
   wire signed [9:0] m68_98;
   assign m68_98 =10'b0;

   // m68_99 = W*in
   wire signed [9:0] m68_99;
   assign m68_99 =10'b0;

   // m68_100 = W*in
   wire signed [9:0] m68_100;
   assign m68_100 =10'b0;

   // m68_101 = W*in
   wire signed [9:0] m68_101;
   assign m68_101 =10'b0;

   // m68_102 = W*in
   wire signed [9:0] m68_102;
   assign m68_102 =10'b0;

   // m68_103 = W*in
   wire signed [9:0] m68_103;
   assign m68_103 =10'b0;

   // m68_104 = W*in
   wire signed [9:0] m68_104;
   assign m68_104 =10'b0;

   // m68_105 = W*in
   wire signed [9:0] m68_105;
   assign m68_105 =10'b0;

   // m68_106 = W*in
   wire signed [9:0] m68_106;
   assign m68_106 =10'b0;

   // m68_107 = W*in
   wire signed [9:0] m68_107;
   assign m68_107 =10'b0;

   // m68_108 = W*in
   wire signed [9:0] m68_108;
   assign m68_108 =10'b0;

   // m68_109 = W*in
   wire signed [9:0] m68_109;
   assign m68_109 =10'b0;

   // m68_110 = W*in
   wire signed [9:0] m68_110;
   assign m68_110 =10'b0;

   // m68_111 = W*in
   wire signed [9:0] m68_111;
   assign m68_111 =10'b0;

   // m68_112 = W*in
   wire signed [9:0] m68_112;
   assign m68_112 =10'b0;

   // m68_113 = W*in
   wire signed [9:0] m68_113;
   assign m68_113 =10'b0;

   // m68_114 = W*in
   wire signed [9:0] m68_114;
   assign m68_114 =10'b0;

   // m68_115 = W*in
   wire signed [9:0] m68_115;
   assign m68_115 =10'b0;

   // m68_116 = W*in
   wire signed [9:0] m68_116;
   assign m68_116 =10'b0;

   // m68_117 = W*in
   wire signed [9:0] m68_117;
   assign m68_117 =10'b0;

   // m69_1 = W*in
   wire signed [9:0] m69_1;
   assign m69_1 =10'b0;

   // m69_2 = W*in
   wire signed [9:0] m69_2;
   assign m69_2 =10'b0;

   // m69_3 = W*in
   wire signed [9:0] m69_3;
   assign m69_3 =10'b0;

   // m69_4 = W*in
   wire signed [9:0] m69_4;
   assign m69_4 =10'b0;

   // m69_5 = W*in
   wire signed [9:0] m69_5;
   assign m69_5 =10'b0;

   // m69_6 = W*in
   wire signed [9:0] m69_6;
   assign m69_6 =10'b0;

   // m69_7 = W*in
   wire signed [9:0] m69_7;
   assign m69_7 =10'b0;

   // m69_8 = W*in
   wire signed [9:0] m69_8;
   assign m69_8 =10'b0;

   // m69_9 = W*in
   wire signed [9:0] m69_9;
   assign m69_9 =10'b0;

   // m69_10 = W*in
   wire signed [9:0] m69_10;
   assign m69_10 =10'b0;

   // m69_11 = W*in
   wire signed [9:0] m69_11;
   assign m69_11 =10'b0;

   // m69_12 = W*in
   wire signed [9:0] m69_12;
   assign m69_12 =10'b0;

   // m69_13 = W*in
   wire signed [9:0] m69_13;
   assign m69_13 =10'b0;

   // m69_14 = W*in
   wire signed [9:0] m69_14;
   assign m69_14 =10'b0;

   // m69_15 = W*in
   wire signed [9:0] m69_15;
   assign m69_15 =10'b0;

   // m69_16 = W*in
   wire signed [9:0] m69_16;
   assign m69_16 =10'b0;

   // m69_17 = W*in
   wire signed [9:0] m69_17;
   assign m69_17 =10'b0;

   // m69_18 = W*in
   wire signed [9:0] m69_18;
   assign m69_18 =10'b0;

   // m69_19 = W*in
   wire signed [9:0] m69_19;
   assign m69_19 ={ {5{in69[5]}} , in69[5:1] };

   // m69_20 = W*in
   wire signed [9:0] m69_20;
   assign m69_20 ={ {4{neg69[5]}} , neg69[5:0] };

   // m69_21 = W*in
   wire signed [9:0] m69_21;
   assign m69_21 ={ {4{in69[5]}} , in69[5:0] };

   // m69_22 = W*in
   wire signed [9:0] m69_22;
   assign m69_22 =10'b0;

   // m69_23 = W*in
   wire signed [9:0] m69_23;
   assign m69_23 =10'b0;

   // m69_24 = W*in
   wire signed [9:0] m69_24;
   assign m69_24 =10'b0;

   // m69_25 = W*in
   wire signed [9:0] m69_25;
   assign m69_25 =10'b0;

   // m69_26 = W*in
   wire signed [9:0] m69_26;
   assign m69_26 ={ {5{neg69[5]}} , neg69[5:1] };

   // m69_27 = W*in
   wire signed [9:0] m69_27;
   assign m69_27 ={ {4{neg69[5]}} , neg69[5:0] };

   // m69_28 = W*in
   wire signed [9:0] m69_28;
   assign m69_28 ={ {5{neg69[5]}} , neg69[5:1] };

   // m69_29 = W*in
   wire signed [9:0] m69_29;
   assign m69_29 =10'b0;

   // m69_30 = W*in
   wire signed [9:0] m69_30;
   assign m69_30 =10'b0;

   // m69_31 = W*in
   wire signed [9:0] m69_31;
   assign m69_31 ={ {5{in69[5]}} , in69[5:1] };

   // m69_32 = W*in
   wire signed [9:0] m69_32;
   assign m69_32 =10'b0;

   // m69_33 = W*in
   wire signed [9:0] m69_33;
   assign m69_33 =10'b0;

   // m69_34 = W*in
   wire signed [9:0] m69_34;
   assign m69_34 =10'b0;

   // m69_35 = W*in
   wire signed [9:0] m69_35;
   assign m69_35 ={ {5{neg69[5]}} , neg69[5:1] };

   // m69_36 = W*in
   wire signed [9:0] m69_36;
   assign m69_36 =10'b0;

   // m69_37 = W*in
   wire signed [9:0] m69_37;
   assign m69_37 =10'b0;

   // m69_38 = W*in
   wire signed [9:0] m69_38;
   assign m69_38 =10'b0;

   // m69_39 = W*in
   wire signed [9:0] m69_39;
   assign m69_39 =10'b0;

   // m69_40 = W*in
   wire signed [9:0] m69_40;
   assign m69_40 =10'b0;

   // m69_41 = W*in
   wire signed [9:0] m69_41;
   assign m69_41 =10'b0;

   // m69_42 = W*in
   wire signed [9:0] m69_42;
   assign m69_42 =10'b0;

   // m69_43 = W*in
   wire signed [9:0] m69_43;
   assign m69_43 =10'b0;

   // m69_44 = W*in
   wire signed [9:0] m69_44;
   assign m69_44 =10'b0;

   // m69_45 = W*in
   wire signed [9:0] m69_45;
   assign m69_45 =10'b0;

   // m69_46 = W*in
   wire signed [9:0] m69_46;
   assign m69_46 =10'b0;

   // m69_47 = W*in
   wire signed [9:0] m69_47;
   assign m69_47 =10'b0;

   // m69_48 = W*in
   wire signed [9:0] m69_48;
   assign m69_48 =10'b0;

   // m69_49 = W*in
   wire signed [9:0] m69_49;
   assign m69_49 =10'b0;

   // m69_50 = W*in
   wire signed [9:0] m69_50;
   assign m69_50 =10'b0;

   // m69_51 = W*in
   wire signed [9:0] m69_51;
   assign m69_51 =10'b0;

   // m69_52 = W*in
   wire signed [9:0] m69_52;
   assign m69_52 =10'b0;

   // m69_53 = W*in
   wire signed [9:0] m69_53;
   assign m69_53 =10'b0;

   // m69_54 = W*in
   wire signed [9:0] m69_54;
   assign m69_54 =10'b0;

   // m69_55 = W*in
   wire signed [9:0] m69_55;
   assign m69_55 =10'b0;

   // m69_56 = W*in
   wire signed [9:0] m69_56;
   assign m69_56 =10'b0;

   // m69_57 = W*in
   wire signed [9:0] m69_57;
   assign m69_57 =10'b0;

   // m69_58 = W*in
   wire signed [9:0] m69_58;
   assign m69_58 =10'b0;

   // m69_59 = W*in
   wire signed [9:0] m69_59;
   assign m69_59 =10'b0;

   // m69_60 = W*in
   wire signed [9:0] m69_60;
   assign m69_60 =10'b0;

   // m69_61 = W*in
   wire signed [9:0] m69_61;
   assign m69_61 =10'b0;

   // m69_62 = W*in
   wire signed [9:0] m69_62;
   assign m69_62 =10'b0;

   // m69_63 = W*in
   wire signed [9:0] m69_63;
   assign m69_63 ={ {4{in69[5]}} , in69[5:0] };

   // m69_64 = W*in
   wire signed [9:0] m69_64;
   assign m69_64 ={ {5{neg69[5]}} , neg69[5:1] };

   // m69_65 = W*in
   wire signed [9:0] m69_65;
   assign m69_65 =10'b0;

   // m69_66 = W*in
   wire signed [9:0] m69_66;
   assign m69_66 =10'b0;

   // m69_67 = W*in
   wire signed [9:0] m69_67;
   assign m69_67 =10'b0;

   // m69_68 = W*in
   wire signed [9:0] m69_68;
   assign m69_68 =10'b0;

   // m69_69 = W*in
   wire signed [9:0] m69_69;
   assign m69_69 =10'b0;

   // m69_70 = W*in
   wire signed [9:0] m69_70;
   assign m69_70 =10'b0;

   // m69_71 = W*in
   wire signed [9:0] m69_71;
   assign m69_71 =10'b0;

   // m69_72 = W*in
   wire signed [9:0] m69_72;
   assign m69_72 =10'b0;

   // m69_73 = W*in
   wire signed [9:0] m69_73;
   assign m69_73 =10'b0;

   // m69_74 = W*in
   wire signed [9:0] m69_74;
   assign m69_74 =10'b0;

   // m69_75 = W*in
   wire signed [9:0] m69_75;
   assign m69_75 =10'b0;

   // m69_76 = W*in
   wire signed [9:0] m69_76;
   assign m69_76 ={ {4{neg69[5]}} , neg69[5:0] };

   // m69_77 = W*in
   wire signed [9:0] m69_77;
   assign m69_77 =10'b0;

   // m69_78 = W*in
   wire signed [9:0] m69_78;
   assign m69_78 =10'b0;

   // m69_79 = W*in
   wire signed [9:0] m69_79;
   assign m69_79 =10'b0;

   // m69_80 = W*in
   wire signed [9:0] m69_80;
   assign m69_80 =10'b0;

   // m69_81 = W*in
   wire signed [9:0] m69_81;
   assign m69_81 =10'b0;

   // m69_82 = W*in
   wire signed [9:0] m69_82;
   assign m69_82 ={ {4{in69[5]}} , in69[5:0] };

   // m69_83 = W*in
   wire signed [9:0] m69_83;
   assign m69_83 =10'b0;

   // m69_84 = W*in
   wire signed [9:0] m69_84;
   assign m69_84 =10'b0;

   // m69_85 = W*in
   wire signed [9:0] m69_85;
   assign m69_85 ={ {4{in69[5]}} , in69[5:0] };

   // m69_86 = W*in
   wire signed [9:0] m69_86;
   assign m69_86 =10'b0;

   // m69_87 = W*in
   wire signed [9:0] m69_87;
   assign m69_87 =10'b0;

   // m69_88 = W*in
   wire signed [9:0] m69_88;
   assign m69_88 =10'b0;

   // m69_89 = W*in
   wire signed [9:0] m69_89;
   assign m69_89 =10'b0;

   // m69_90 = W*in
   wire signed [9:0] m69_90;
   assign m69_90 =10'b0;

   // m69_91 = W*in
   wire signed [9:0] m69_91;
   assign m69_91 =10'b0;

   // m69_92 = W*in
   wire signed [9:0] m69_92;
   assign m69_92 =10'b0;

   // m69_93 = W*in
   wire signed [9:0] m69_93;
   assign m69_93 =10'b0;

   // m69_94 = W*in
   wire signed [9:0] m69_94;
   assign m69_94 =10'b0;

   // m69_95 = W*in
   wire signed [9:0] m69_95;
   assign m69_95 =10'b0;

   // m69_96 = W*in
   wire signed [9:0] m69_96;
   assign m69_96 =10'b0;

   // m69_97 = W*in
   wire signed [9:0] m69_97;
   assign m69_97 =10'b0;

   // m69_98 = W*in
   wire signed [9:0] m69_98;
   assign m69_98 ={ {4{in69[5]}} , in69[5:0] };

   // m69_99 = W*in
   wire signed [9:0] m69_99;
   assign m69_99 =10'b0;

   // m69_100 = W*in
   wire signed [9:0] m69_100;
   assign m69_100 =10'b0;

   // m69_101 = W*in
   wire signed [9:0] m69_101;
   assign m69_101 =10'b0;

   // m69_102 = W*in
   wire signed [9:0] m69_102;
   assign m69_102 ={ {5{neg69[5]}} , neg69[5:1] };

   // m69_103 = W*in
   wire signed [9:0] m69_103;
   assign m69_103 =10'b0;

   // m69_104 = W*in
   wire signed [9:0] m69_104;
   assign m69_104 =10'b0;

   // m69_105 = W*in
   wire signed [9:0] m69_105;
   assign m69_105 =10'b0;

   // m69_106 = W*in
   wire signed [9:0] m69_106;
   assign m69_106 =10'b0;

   // m69_107 = W*in
   wire signed [9:0] m69_107;
   assign m69_107 =10'b0;

   // m69_108 = W*in
   wire signed [9:0] m69_108;
   assign m69_108 =10'b0;

   // m69_109 = W*in
   wire signed [9:0] m69_109;
   assign m69_109 =10'b0;

   // m69_110 = W*in
   wire signed [9:0] m69_110;
   assign m69_110 =10'b0;

   // m69_111 = W*in
   wire signed [9:0] m69_111;
   assign m69_111 =10'b0;

   // m69_112 = W*in
   wire signed [9:0] m69_112;
   assign m69_112 =10'b0;

   // m69_113 = W*in
   wire signed [9:0] m69_113;
   assign m69_113 =10'b0;

   // m69_114 = W*in
   wire signed [9:0] m69_114;
   assign m69_114 =10'b0;

   // m69_115 = W*in
   wire signed [9:0] m69_115;
   assign m69_115 ={ {5{neg69[5]}} , neg69[5:1] };

   // m69_116 = W*in
   wire signed [9:0] m69_116;
   assign m69_116 =10'b0;

   // m69_117 = W*in
   wire signed [9:0] m69_117;
   assign m69_117 ={ {4{neg69[5]}} , neg69[5:0] };

   // m70_1 = W*in
   wire signed [9:0] m70_1;
   assign m70_1 =10'b0;

   // m70_2 = W*in
   wire signed [9:0] m70_2;
   assign m70_2 =10'b0;

   // m70_3 = W*in
   wire signed [9:0] m70_3;
   assign m70_3 =10'b0;

   // m70_4 = W*in
   wire signed [9:0] m70_4;
   assign m70_4 =10'b0;

   // m70_5 = W*in
   wire signed [9:0] m70_5;
   assign m70_5 =10'b0;

   // m70_6 = W*in
   wire signed [9:0] m70_6;
   assign m70_6 =10'b0;

   // m70_7 = W*in
   wire signed [9:0] m70_7;
   assign m70_7 =10'b0;

   // m70_8 = W*in
   wire signed [9:0] m70_8;
   assign m70_8 =10'b0;

   // m70_9 = W*in
   wire signed [9:0] m70_9;
   assign m70_9 =10'b0;

   // m70_10 = W*in
   wire signed [9:0] m70_10;
   assign m70_10 =10'b0;

   // m70_11 = W*in
   wire signed [9:0] m70_11;
   assign m70_11 =10'b0;

   // m70_12 = W*in
   wire signed [9:0] m70_12;
   assign m70_12 =10'b0;

   // m70_13 = W*in
   wire signed [9:0] m70_13;
   assign m70_13 =10'b0;

   // m70_14 = W*in
   wire signed [9:0] m70_14;
   assign m70_14 =10'b0;

   // m70_15 = W*in
   wire signed [9:0] m70_15;
   assign m70_15 =10'b0;

   // m70_16 = W*in
   wire signed [9:0] m70_16;
   assign m70_16 =10'b0;

   // m70_17 = W*in
   wire signed [9:0] m70_17;
   assign m70_17 =10'b0;

   // m70_18 = W*in
   wire signed [9:0] m70_18;
   assign m70_18 =10'b0;

   // m70_19 = W*in
   wire signed [9:0] m70_19;
   assign m70_19 =10'b0;

   // m70_20 = W*in
   wire signed [9:0] m70_20;
   assign m70_20 =10'b0;

   // m70_21 = W*in
   wire signed [9:0] m70_21;
   assign m70_21 =10'b0;

   // m70_22 = W*in
   wire signed [9:0] m70_22;
   assign m70_22 =10'b0;

   // m70_23 = W*in
   wire signed [9:0] m70_23;
   assign m70_23 =10'b0;

   // m70_24 = W*in
   wire signed [9:0] m70_24;
   assign m70_24 =10'b0;

   // m70_25 = W*in
   wire signed [9:0] m70_25;
   assign m70_25 =10'b0;

   // m70_26 = W*in
   wire signed [9:0] m70_26;
   assign m70_26 =10'b0;

   // m70_27 = W*in
   wire signed [9:0] m70_27;
   assign m70_27 =10'b0;

   // m70_28 = W*in
   wire signed [9:0] m70_28;
   assign m70_28 =10'b0;

   // m70_29 = W*in
   wire signed [9:0] m70_29;
   assign m70_29 ={ {5{neg70[5]}} , neg70[5:1] };

   // m70_30 = W*in
   wire signed [9:0] m70_30;
   assign m70_30 =10'b0;

   // m70_31 = W*in
   wire signed [9:0] m70_31;
   assign m70_31 =10'b0;

   // m70_32 = W*in
   wire signed [9:0] m70_32;
   assign m70_32 =10'b0;

   // m70_33 = W*in
   wire signed [9:0] m70_33;
   assign m70_33 =10'b0;

   // m70_34 = W*in
   wire signed [9:0] m70_34;
   assign m70_34 =10'b0;

   // m70_35 = W*in
   wire signed [9:0] m70_35;
   assign m70_35 =10'b0;

   // m70_36 = W*in
   wire signed [9:0] m70_36;
   assign m70_36 ={ {5{neg70[5]}} , neg70[5:1] };

   // m70_37 = W*in
   wire signed [9:0] m70_37;
   assign m70_37 =10'b0;

   // m70_38 = W*in
   wire signed [9:0] m70_38;
   assign m70_38 =10'b0;

   // m70_39 = W*in
   wire signed [9:0] m70_39;
   assign m70_39 =10'b0;

   // m70_40 = W*in
   wire signed [9:0] m70_40;
   assign m70_40 =10'b0;

   // m70_41 = W*in
   wire signed [9:0] m70_41;
   assign m70_41 =10'b0;

   // m70_42 = W*in
   wire signed [9:0] m70_42;
   assign m70_42 =10'b0;

   // m70_43 = W*in
   wire signed [9:0] m70_43;
   assign m70_43 =10'b0;

   // m70_44 = W*in
   wire signed [9:0] m70_44;
   assign m70_44 =10'b0;

   // m70_45 = W*in
   wire signed [9:0] m70_45;
   assign m70_45 =10'b0;

   // m70_46 = W*in
   wire signed [9:0] m70_46;
   assign m70_46 =10'b0;

   // m70_47 = W*in
   wire signed [9:0] m70_47;
   assign m70_47 =10'b0;

   // m70_48 = W*in
   wire signed [9:0] m70_48;
   assign m70_48 =10'b0;

   // m70_49 = W*in
   wire signed [9:0] m70_49;
   assign m70_49 =10'b0;

   // m70_50 = W*in
   wire signed [9:0] m70_50;
   assign m70_50 =10'b0;

   // m70_51 = W*in
   wire signed [9:0] m70_51;
   assign m70_51 =10'b0;

   // m70_52 = W*in
   wire signed [9:0] m70_52;
   assign m70_52 =10'b0;

   // m70_53 = W*in
   wire signed [9:0] m70_53;
   assign m70_53 =10'b0;

   // m70_54 = W*in
   wire signed [9:0] m70_54;
   assign m70_54 =10'b0;

   // m70_55 = W*in
   wire signed [9:0] m70_55;
   assign m70_55 =10'b0;

   // m70_56 = W*in
   wire signed [9:0] m70_56;
   assign m70_56 =10'b0;

   // m70_57 = W*in
   wire signed [9:0] m70_57;
   assign m70_57 =10'b0;

   // m70_58 = W*in
   wire signed [9:0] m70_58;
   assign m70_58 =10'b0;

   // m70_59 = W*in
   wire signed [9:0] m70_59;
   assign m70_59 =10'b0;

   // m70_60 = W*in
   wire signed [9:0] m70_60;
   assign m70_60 =10'b0;

   // m70_61 = W*in
   wire signed [9:0] m70_61;
   assign m70_61 =10'b0;

   // m70_62 = W*in
   wire signed [9:0] m70_62;
   assign m70_62 =10'b0;

   // m70_63 = W*in
   wire signed [9:0] m70_63;
   assign m70_63 ={ {4{in70[5]}} , in70[5:0] };

   // m70_64 = W*in
   wire signed [9:0] m70_64;
   assign m70_64 =10'b0;

   // m70_65 = W*in
   wire signed [9:0] m70_65;
   assign m70_65 =10'b0;

   // m70_66 = W*in
   wire signed [9:0] m70_66;
   assign m70_66 ={ {5{neg70[5]}} , neg70[5:1] };

   // m70_67 = W*in
   wire signed [9:0] m70_67;
   assign m70_67 =10'b0;

   // m70_68 = W*in
   wire signed [9:0] m70_68;
   assign m70_68 =10'b0;

   // m70_69 = W*in
   wire signed [9:0] m70_69;
   assign m70_69 ={ {5{in70[5]}} , in70[5:1] };

   // m70_70 = W*in
   wire signed [9:0] m70_70;
   assign m70_70 =10'b0;

   // m70_71 = W*in
   wire signed [9:0] m70_71;
   assign m70_71 =10'b0;

   // m70_72 = W*in
   wire signed [9:0] m70_72;
   assign m70_72 ={ {4{in70[5]}} , in70[5:0] };

   // m70_73 = W*in
   wire signed [9:0] m70_73;
   assign m70_73 ={ {5{neg70[5]}} , neg70[5:1] };

   // m70_74 = W*in
   wire signed [9:0] m70_74;
   assign m70_74 =10'b0;

   // m70_75 = W*in
   wire signed [9:0] m70_75;
   assign m70_75 =10'b0;

   // m70_76 = W*in
   wire signed [9:0] m70_76;
   assign m70_76 =10'b0;

   // m70_77 = W*in
   wire signed [9:0] m70_77;
   assign m70_77 =10'b0;

   // m70_78 = W*in
   wire signed [9:0] m70_78;
   assign m70_78 =10'b0;

   // m70_79 = W*in
   wire signed [9:0] m70_79;
   assign m70_79 ={ {4{neg70[5]}} , neg70[5:0] };

   // m70_80 = W*in
   wire signed [9:0] m70_80;
   assign m70_80 =10'b0;

   // m70_81 = W*in
   wire signed [9:0] m70_81;
   assign m70_81 =10'b0;

   // m70_82 = W*in
   wire signed [9:0] m70_82;
   assign m70_82 =10'b0;

   // m70_83 = W*in
   wire signed [9:0] m70_83;
   assign m70_83 =10'b0;

   // m70_84 = W*in
   wire signed [9:0] m70_84;
   assign m70_84 =10'b0;

   // m70_85 = W*in
   wire signed [9:0] m70_85;
   assign m70_85 =10'b0;

   // m70_86 = W*in
   wire signed [9:0] m70_86;
   assign m70_86 =10'b0;

   // m70_87 = W*in
   wire signed [9:0] m70_87;
   assign m70_87 =10'b0;

   // m70_88 = W*in
   wire signed [9:0] m70_88;
   assign m70_88 =10'b0;

   // m70_89 = W*in
   wire signed [9:0] m70_89;
   assign m70_89 =10'b0;

   // m70_90 = W*in
   wire signed [9:0] m70_90;
   assign m70_90 =10'b0;

   // m70_91 = W*in
   wire signed [9:0] m70_91;
   assign m70_91 =10'b0;

   // m70_92 = W*in
   wire signed [9:0] m70_92;
   assign m70_92 ={ {4{in70[5]}} , in70[5:0] };

   // m70_93 = W*in
   wire signed [9:0] m70_93;
   assign m70_93 =10'b0;

   // m70_94 = W*in
   wire signed [9:0] m70_94;
   assign m70_94 =10'b0;

   // m70_95 = W*in
   wire signed [9:0] m70_95;
   assign m70_95 =10'b0;

   // m70_96 = W*in
   wire signed [9:0] m70_96;
   assign m70_96 =10'b0;

   // m70_97 = W*in
   wire signed [9:0] m70_97;
   assign m70_97 =10'b0;

   // m70_98 = W*in
   wire signed [9:0] m70_98;
   assign m70_98 =10'b0;

   // m70_99 = W*in
   wire signed [9:0] m70_99;
   assign m70_99 =10'b0;

   // m70_100 = W*in
   wire signed [9:0] m70_100;
   assign m70_100 =10'b0;

   // m70_101 = W*in
   wire signed [9:0] m70_101;
   assign m70_101 =10'b0;

   // m70_102 = W*in
   wire signed [9:0] m70_102;
   assign m70_102 =10'b0;

   // m70_103 = W*in
   wire signed [9:0] m70_103;
   assign m70_103 =10'b0;

   // m70_104 = W*in
   wire signed [9:0] m70_104;
   assign m70_104 =10'b0;

   // m70_105 = W*in
   wire signed [9:0] m70_105;
   assign m70_105 =10'b0;

   // m70_106 = W*in
   wire signed [9:0] m70_106;
   assign m70_106 =10'b0;

   // m70_107 = W*in
   wire signed [9:0] m70_107;
   assign m70_107 =10'b0;

   // m70_108 = W*in
   wire signed [9:0] m70_108;
   assign m70_108 ={ {5{neg70[5]}} , neg70[5:1] };

   // m70_109 = W*in
   wire signed [9:0] m70_109;
   assign m70_109 ={ {4{neg70[5]}} , neg70[5:0] };

   // m70_110 = W*in
   wire signed [9:0] m70_110;
   assign m70_110 =10'b0;

   // m70_111 = W*in
   wire signed [9:0] m70_111;
   assign m70_111 =10'b0;

   // m70_112 = W*in
   wire signed [9:0] m70_112;
   assign m70_112 =10'b0;

   // m70_113 = W*in
   wire signed [9:0] m70_113;
   assign m70_113 =10'b0;

   // m70_114 = W*in
   wire signed [9:0] m70_114;
   assign m70_114 =10'b0;

   // m70_115 = W*in
   wire signed [9:0] m70_115;
   assign m70_115 =10'b0;

   // m70_116 = W*in
   wire signed [9:0] m70_116;
   assign m70_116 =10'b0;

   // m70_117 = W*in
   wire signed [9:0] m70_117;
   assign m70_117 =10'b0;

   // m71_1 = W*in
   wire signed [9:0] m71_1;
   assign m71_1 =10'b0;

   // m71_2 = W*in
   wire signed [9:0] m71_2;
   assign m71_2 =10'b0;

   // m71_3 = W*in
   wire signed [9:0] m71_3;
   assign m71_3 =10'b0;

   // m71_4 = W*in
   wire signed [9:0] m71_4;
   assign m71_4 =10'b0;

   // m71_5 = W*in
   wire signed [9:0] m71_5;
   assign m71_5 =10'b0;

   // m71_6 = W*in
   wire signed [9:0] m71_6;
   assign m71_6 =10'b0;

   // m71_7 = W*in
   wire signed [9:0] m71_7;
   assign m71_7 =10'b0;

   // m71_8 = W*in
   wire signed [9:0] m71_8;
   assign m71_8 =10'b0;

   // m71_9 = W*in
   wire signed [9:0] m71_9;
   assign m71_9 =10'b0;

   // m71_10 = W*in
   wire signed [9:0] m71_10;
   assign m71_10 =10'b0;

   // m71_11 = W*in
   wire signed [9:0] m71_11;
   assign m71_11 =10'b0;

   // m71_12 = W*in
   wire signed [9:0] m71_12;
   assign m71_12 =10'b0;

   // m71_13 = W*in
   wire signed [9:0] m71_13;
   assign m71_13 =10'b0;

   // m71_14 = W*in
   wire signed [9:0] m71_14;
   assign m71_14 =10'b0;

   // m71_15 = W*in
   wire signed [9:0] m71_15;
   assign m71_15 =10'b0;

   // m71_16 = W*in
   wire signed [9:0] m71_16;
   assign m71_16 =10'b0;

   // m71_17 = W*in
   wire signed [9:0] m71_17;
   assign m71_17 =10'b0;

   // m71_18 = W*in
   wire signed [9:0] m71_18;
   assign m71_18 =10'b0;

   // m71_19 = W*in
   wire signed [9:0] m71_19;
   assign m71_19 ={ {5{neg71[5]}} , neg71[5:1] };

   // m71_20 = W*in
   wire signed [9:0] m71_20;
   assign m71_20 =10'b0;

   // m71_21 = W*in
   wire signed [9:0] m71_21;
   assign m71_21 =10'b0;

   // m71_22 = W*in
   wire signed [9:0] m71_22;
   assign m71_22 =10'b0;

   // m71_23 = W*in
   wire signed [9:0] m71_23;
   assign m71_23 =10'b0;

   // m71_24 = W*in
   wire signed [9:0] m71_24;
   assign m71_24 =10'b0;

   // m71_25 = W*in
   wire signed [9:0] m71_25;
   assign m71_25 =10'b0;

   // m71_26 = W*in
   wire signed [9:0] m71_26;
   assign m71_26 =10'b0;

   // m71_27 = W*in
   wire signed [9:0] m71_27;
   assign m71_27 =10'b0;

   // m71_28 = W*in
   wire signed [9:0] m71_28;
   assign m71_28 =10'b0;

   // m71_29 = W*in
   wire signed [9:0] m71_29;
   assign m71_29 ={ {5{neg71[5]}} , neg71[5:1] };

   // m71_30 = W*in
   wire signed [9:0] m71_30;
   assign m71_30 =10'b0;

   // m71_31 = W*in
   wire signed [9:0] m71_31;
   assign m71_31 ={ {5{neg71[5]}} , neg71[5:1] };

   // m71_32 = W*in
   wire signed [9:0] m71_32;
   assign m71_32 =10'b0;

   // m71_33 = W*in
   wire signed [9:0] m71_33;
   assign m71_33 =10'b0;

   // m71_34 = W*in
   wire signed [9:0] m71_34;
   assign m71_34 =10'b0;

   // m71_35 = W*in
   wire signed [9:0] m71_35;
   assign m71_35 =10'b0;

   // m71_36 = W*in
   wire signed [9:0] m71_36;
   assign m71_36 ={ {5{neg71[5]}} , neg71[5:1] };

   // m71_37 = W*in
   wire signed [9:0] m71_37;
   assign m71_37 =10'b0;

   // m71_38 = W*in
   wire signed [9:0] m71_38;
   assign m71_38 =10'b0;

   // m71_39 = W*in
   wire signed [9:0] m71_39;
   assign m71_39 =10'b0;

   // m71_40 = W*in
   wire signed [9:0] m71_40;
   assign m71_40 =10'b0;

   // m71_41 = W*in
   wire signed [9:0] m71_41;
   assign m71_41 ={ {4{in71[5]}} , in71[5:0] };

   // m71_42 = W*in
   wire signed [9:0] m71_42;
   assign m71_42 =10'b0;

   // m71_43 = W*in
   wire signed [9:0] m71_43;
   assign m71_43 =10'b0;

   // m71_44 = W*in
   wire signed [9:0] m71_44;
   assign m71_44 ={ {4{neg71[5]}} , neg71[5:0] };

   // m71_45 = W*in
   wire signed [9:0] m71_45;
   assign m71_45 =10'b0;

   // m71_46 = W*in
   wire signed [9:0] m71_46;
   assign m71_46 =10'b0;

   // m71_47 = W*in
   wire signed [9:0] m71_47;
   assign m71_47 =10'b0;

   // m71_48 = W*in
   wire signed [9:0] m71_48;
   assign m71_48 =10'b0;

   // m71_49 = W*in
   wire signed [9:0] m71_49;
   assign m71_49 ={ {4{neg71[5]}} , neg71[5:0] };

   // m71_50 = W*in
   wire signed [9:0] m71_50;
   assign m71_50 =10'b0;

   // m71_51 = W*in
   wire signed [9:0] m71_51;
   assign m71_51 =10'b0;

   // m71_52 = W*in
   wire signed [9:0] m71_52;
   assign m71_52 =10'b0;

   // m71_53 = W*in
   wire signed [9:0] m71_53;
   assign m71_53 ={ {4{neg71[5]}} , neg71[5:0] };

   // m71_54 = W*in
   wire signed [9:0] m71_54;
   assign m71_54 ={ {4{neg71[5]}} , neg71[5:0] };

   // m71_55 = W*in
   wire signed [9:0] m71_55;
   assign m71_55 =10'b0;

   // m71_56 = W*in
   wire signed [9:0] m71_56;
   assign m71_56 =10'b0;

   // m71_57 = W*in
   wire signed [9:0] m71_57;
   assign m71_57 =10'b0;

   // m71_58 = W*in
   wire signed [9:0] m71_58;
   assign m71_58 =10'b0;

   // m71_59 = W*in
   wire signed [9:0] m71_59;
   assign m71_59 =10'b0;

   // m71_60 = W*in
   wire signed [9:0] m71_60;
   assign m71_60 =10'b0;

   // m71_61 = W*in
   wire signed [9:0] m71_61;
   assign m71_61 =10'b0;

   // m71_62 = W*in
   wire signed [9:0] m71_62;
   assign m71_62 =10'b0;

   // m71_63 = W*in
   wire signed [9:0] m71_63;
   assign m71_63 =10'b0;

   // m71_64 = W*in
   wire signed [9:0] m71_64;
   assign m71_64 =10'b0;

   // m71_65 = W*in
   wire signed [9:0] m71_65;
   assign m71_65 =10'b0;

   // m71_66 = W*in
   wire signed [9:0] m71_66;
   assign m71_66 =10'b0;

   // m71_67 = W*in
   wire signed [9:0] m71_67;
   assign m71_67 =10'b0;

   // m71_68 = W*in
   wire signed [9:0] m71_68;
   assign m71_68 =10'b0;

   // m71_69 = W*in
   wire signed [9:0] m71_69;
   assign m71_69 =10'b0;

   // m71_70 = W*in
   wire signed [9:0] m71_70;
   assign m71_70 ={ {5{in71[5]}} , in71[5:1] };

   // m71_71 = W*in
   wire signed [9:0] m71_71;
   assign m71_71 =10'b0;

   // m71_72 = W*in
   wire signed [9:0] m71_72;
   assign m71_72 ={ {4{in71[5]}} , in71[5:0] };

   // m71_73 = W*in
   wire signed [9:0] m71_73;
   assign m71_73 =10'b0;

   // m71_74 = W*in
   wire signed [9:0] m71_74;
   assign m71_74 =10'b0;

   // m71_75 = W*in
   wire signed [9:0] m71_75;
   assign m71_75 =10'b0;

   // m71_76 = W*in
   wire signed [9:0] m71_76;
   assign m71_76 =10'b0;

   // m71_77 = W*in
   wire signed [9:0] m71_77;
   assign m71_77 =10'b0;

   // m71_78 = W*in
   wire signed [9:0] m71_78;
   assign m71_78 =10'b0;

   // m71_79 = W*in
   wire signed [9:0] m71_79;
   assign m71_79 =10'b0;

   // m71_80 = W*in
   wire signed [9:0] m71_80;
   assign m71_80 =10'b0;

   // m71_81 = W*in
   wire signed [9:0] m71_81;
   assign m71_81 =10'b0;

   // m71_82 = W*in
   wire signed [9:0] m71_82;
   assign m71_82 =10'b0;

   // m71_83 = W*in
   wire signed [9:0] m71_83;
   assign m71_83 =10'b0;

   // m71_84 = W*in
   wire signed [9:0] m71_84;
   assign m71_84 =10'b0;

   // m71_85 = W*in
   wire signed [9:0] m71_85;
   assign m71_85 =10'b0;

   // m71_86 = W*in
   wire signed [9:0] m71_86;
   assign m71_86 ={ {4{in71[5]}} , in71[5:0] };

   // m71_87 = W*in
   wire signed [9:0] m71_87;
   assign m71_87 =10'b0;

   // m71_88 = W*in
   wire signed [9:0] m71_88;
   assign m71_88 =10'b0;

   // m71_89 = W*in
   wire signed [9:0] m71_89;
   assign m71_89 =10'b0;

   // m71_90 = W*in
   wire signed [9:0] m71_90;
   assign m71_90 =10'b0;

   // m71_91 = W*in
   wire signed [9:0] m71_91;
   assign m71_91 =10'b0;

   // m71_92 = W*in
   wire signed [9:0] m71_92;
   assign m71_92 =10'b0;

   // m71_93 = W*in
   wire signed [9:0] m71_93;
   assign m71_93 =10'b0;

   // m71_94 = W*in
   wire signed [9:0] m71_94;
   assign m71_94 =10'b0;

   // m71_95 = W*in
   wire signed [9:0] m71_95;
   assign m71_95 ={ {4{neg71[5]}} , neg71[5:0] };

   // m71_96 = W*in
   wire signed [9:0] m71_96;
   assign m71_96 =10'b0;

   // m71_97 = W*in
   wire signed [9:0] m71_97;
   assign m71_97 ={ {4{neg71[5]}} , neg71[5:0] };

   // m71_98 = W*in
   wire signed [9:0] m71_98;
   assign m71_98 =10'b0;

   // m71_99 = W*in
   wire signed [9:0] m71_99;
   assign m71_99 =10'b0;

   // m71_100 = W*in
   wire signed [9:0] m71_100;
   assign m71_100 =10'b0;

   // m71_101 = W*in
   wire signed [9:0] m71_101;
   assign m71_101 =10'b0;

   // m71_102 = W*in
   wire signed [9:0] m71_102;
   assign m71_102 =10'b0;

   // m71_103 = W*in
   wire signed [9:0] m71_103;
   assign m71_103 =10'b0;

   // m71_104 = W*in
   wire signed [9:0] m71_104;
   assign m71_104 =10'b0;

   // m71_105 = W*in
   wire signed [9:0] m71_105;
   assign m71_105 =10'b0;

   // m71_106 = W*in
   wire signed [9:0] m71_106;
   assign m71_106 =10'b0;

   // m71_107 = W*in
   wire signed [9:0] m71_107;
   assign m71_107 =10'b0;

   // m71_108 = W*in
   wire signed [9:0] m71_108;
   assign m71_108 ={ {4{in71[5]}} , in71[5:0] };

   // m71_109 = W*in
   wire signed [9:0] m71_109;
   assign m71_109 =10'b0;

   // m71_110 = W*in
   wire signed [9:0] m71_110;
   assign m71_110 =10'b0;

   // m71_111 = W*in
   wire signed [9:0] m71_111;
   assign m71_111 =10'b0;

   // m71_112 = W*in
   wire signed [9:0] m71_112;
   assign m71_112 =10'b0;

   // m71_113 = W*in
   wire signed [9:0] m71_113;
   assign m71_113 =10'b0;

   // m71_114 = W*in
   wire signed [9:0] m71_114;
   assign m71_114 =10'b0;

   // m71_115 = W*in
   wire signed [9:0] m71_115;
   assign m71_115 =10'b0;

   // m71_116 = W*in
   wire signed [9:0] m71_116;
   assign m71_116 ={ {4{in71[5]}} , in71[5:0] };

   // m71_117 = W*in
   wire signed [9:0] m71_117;
   assign m71_117 =10'b0;

   // m72_1 = W*in
   wire signed [9:0] m72_1;
   assign m72_1 =10'b0;

   // m72_2 = W*in
   wire signed [9:0] m72_2;
   assign m72_2 =10'b0;

   // m72_3 = W*in
   wire signed [9:0] m72_3;
   assign m72_3 =10'b0;

   // m72_4 = W*in
   wire signed [9:0] m72_4;
   assign m72_4 =10'b0;

   // m72_5 = W*in
   wire signed [9:0] m72_5;
   assign m72_5 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_6 = W*in
   wire signed [9:0] m72_6;
   assign m72_6 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_7 = W*in
   wire signed [9:0] m72_7;
   assign m72_7 =10'b0;

   // m72_8 = W*in
   wire signed [9:0] m72_8;
   assign m72_8 =10'b0;

   // m72_9 = W*in
   wire signed [9:0] m72_9;
   assign m72_9 =10'b0;

   // m72_10 = W*in
   wire signed [9:0] m72_10;
   assign m72_10 =10'b0;

   // m72_11 = W*in
   wire signed [9:0] m72_11;
   assign m72_11 =10'b0;

   // m72_12 = W*in
   wire signed [9:0] m72_12;
   assign m72_12 =10'b0;

   // m72_13 = W*in
   wire signed [9:0] m72_13;
   assign m72_13 ={ {4{in72[5]}} , in72[5:0] };

   // m72_14 = W*in
   wire signed [9:0] m72_14;
   assign m72_14 =10'b0;

   // m72_15 = W*in
   wire signed [9:0] m72_15;
   assign m72_15 =10'b0;

   // m72_16 = W*in
   wire signed [9:0] m72_16;
   assign m72_16 =10'b0;

   // m72_17 = W*in
   wire signed [9:0] m72_17;
   assign m72_17 ={ {5{in72[5]}} , in72[5:1] };

   // m72_18 = W*in
   wire signed [9:0] m72_18;
   assign m72_18 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_19 = W*in
   wire signed [9:0] m72_19;
   assign m72_19 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_20 = W*in
   wire signed [9:0] m72_20;
   assign m72_20 =10'b0;

   // m72_21 = W*in
   wire signed [9:0] m72_21;
   assign m72_21 =10'b0;

   // m72_22 = W*in
   wire signed [9:0] m72_22;
   assign m72_22 =10'b0;

   // m72_23 = W*in
   wire signed [9:0] m72_23;
   assign m72_23 =10'b0;

   // m72_24 = W*in
   wire signed [9:0] m72_24;
   assign m72_24 =10'b0;

   // m72_25 = W*in
   wire signed [9:0] m72_25;
   assign m72_25 =10'b0;

   // m72_26 = W*in
   wire signed [9:0] m72_26;
   assign m72_26 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_27 = W*in
   wire signed [9:0] m72_27;
   assign m72_27 =10'b0;

   // m72_28 = W*in
   wire signed [9:0] m72_28;
   assign m72_28 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_29 = W*in
   wire signed [9:0] m72_29;
   assign m72_29 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_30 = W*in
   wire signed [9:0] m72_30;
   assign m72_30 =10'b0;

   // m72_31 = W*in
   wire signed [9:0] m72_31;
   assign m72_31 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_32 = W*in
   wire signed [9:0] m72_32;
   assign m72_32 =10'b0;

   // m72_33 = W*in
   wire signed [9:0] m72_33;
   assign m72_33 =10'b0;

   // m72_34 = W*in
   wire signed [9:0] m72_34;
   assign m72_34 =10'b0;

   // m72_35 = W*in
   wire signed [9:0] m72_35;
   assign m72_35 =10'b0;

   // m72_36 = W*in
   wire signed [9:0] m72_36;
   assign m72_36 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_37 = W*in
   wire signed [9:0] m72_37;
   assign m72_37 ={ {4{in72[5]}} , in72[5:0] };

   // m72_38 = W*in
   wire signed [9:0] m72_38;
   assign m72_38 =10'b0;

   // m72_39 = W*in
   wire signed [9:0] m72_39;
   assign m72_39 =10'b0;

   // m72_40 = W*in
   wire signed [9:0] m72_40;
   assign m72_40 =10'b0;

   // m72_41 = W*in
   wire signed [9:0] m72_41;
   assign m72_41 ={ {4{in72[5]}} , in72[5:0] };

   // m72_42 = W*in
   wire signed [9:0] m72_42;
   assign m72_42 =10'b0;

   // m72_43 = W*in
   wire signed [9:0] m72_43;
   assign m72_43 =10'b0;

   // m72_44 = W*in
   wire signed [9:0] m72_44;
   assign m72_44 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_45 = W*in
   wire signed [9:0] m72_45;
   assign m72_45 =10'b0;

   // m72_46 = W*in
   wire signed [9:0] m72_46;
   assign m72_46 =10'b0;

   // m72_47 = W*in
   wire signed [9:0] m72_47;
   assign m72_47 =10'b0;

   // m72_48 = W*in
   wire signed [9:0] m72_48;
   assign m72_48 =10'b0;

   // m72_49 = W*in
   wire signed [9:0] m72_49;
   assign m72_49 ={ {3{neg72[5]}} , neg72 , {1{1'b0}} };

   // m72_50 = W*in
   wire signed [9:0] m72_50;
   assign m72_50 =10'b0;

   // m72_51 = W*in
   wire signed [9:0] m72_51;
   assign m72_51 =10'b0;

   // m72_52 = W*in
   wire signed [9:0] m72_52;
   assign m72_52 =10'b0;

   // m72_53 = W*in
   wire signed [9:0] m72_53;
   assign m72_53 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_54 = W*in
   wire signed [9:0] m72_54;
   assign m72_54 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_55 = W*in
   wire signed [9:0] m72_55;
   assign m72_55 =10'b0;

   // m72_56 = W*in
   wire signed [9:0] m72_56;
   assign m72_56 =10'b0;

   // m72_57 = W*in
   wire signed [9:0] m72_57;
   assign m72_57 =10'b0;

   // m72_58 = W*in
   wire signed [9:0] m72_58;
   assign m72_58 =10'b0;

   // m72_59 = W*in
   wire signed [9:0] m72_59;
   assign m72_59 =10'b0;

   // m72_60 = W*in
   wire signed [9:0] m72_60;
   assign m72_60 =10'b0;

   // m72_61 = W*in
   wire signed [9:0] m72_61;
   assign m72_61 =10'b0;

   // m72_62 = W*in
   wire signed [9:0] m72_62;
   assign m72_62 =10'b0;

   // m72_63 = W*in
   wire signed [9:0] m72_63;
   assign m72_63 =10'b0;

   // m72_64 = W*in
   wire signed [9:0] m72_64;
   assign m72_64 =10'b0;

   // m72_65 = W*in
   wire signed [9:0] m72_65;
   assign m72_65 ={ {5{in72[5]}} , in72[5:1] };

   // m72_66 = W*in
   wire signed [9:0] m72_66;
   assign m72_66 ={ {4{in72[5]}} , in72[5:0] };

   // m72_67 = W*in
   wire signed [9:0] m72_67;
   assign m72_67 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_68 = W*in
   wire signed [9:0] m72_68;
   assign m72_68 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_69 = W*in
   wire signed [9:0] m72_69;
   assign m72_69 ={ {4{in72[5]}} , in72[5:0] };

   // m72_70 = W*in
   wire signed [9:0] m72_70;
   assign m72_70 =10'b0;

   // m72_71 = W*in
   wire signed [9:0] m72_71;
   assign m72_71 =10'b0;

   // m72_72 = W*in
   wire signed [9:0] m72_72;
   assign m72_72 =10'b0;

   // m72_73 = W*in
   wire signed [9:0] m72_73;
   assign m72_73 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_74 = W*in
   wire signed [9:0] m72_74;
   assign m72_74 ={ {5{neg72[5]}} , neg72[5:1] };

   // m72_75 = W*in
   wire signed [9:0] m72_75;
   assign m72_75 =10'b0;

   // m72_76 = W*in
   wire signed [9:0] m72_76;
   assign m72_76 =10'b0;

   // m72_77 = W*in
   wire signed [9:0] m72_77;
   assign m72_77 =10'b0;

   // m72_78 = W*in
   wire signed [9:0] m72_78;
   assign m72_78 =10'b0;

   // m72_79 = W*in
   wire signed [9:0] m72_79;
   assign m72_79 =10'b0;

   // m72_80 = W*in
   wire signed [9:0] m72_80;
   assign m72_80 =10'b0;

   // m72_81 = W*in
   wire signed [9:0] m72_81;
   assign m72_81 ={ {4{in72[5]}} , in72[5:0] };

   // m72_82 = W*in
   wire signed [9:0] m72_82;
   assign m72_82 ={ {4{in72[5]}} , in72[5:0] };

   // m72_83 = W*in
   wire signed [9:0] m72_83;
   assign m72_83 =10'b0;

   // m72_84 = W*in
   wire signed [9:0] m72_84;
   assign m72_84 =10'b0;

   // m72_85 = W*in
   wire signed [9:0] m72_85;
   assign m72_85 ={ {4{in72[5]}} , in72[5:0] };

   // m72_86 = W*in
   wire signed [9:0] m72_86;
   assign m72_86 =10'b0;

   // m72_87 = W*in
   wire signed [9:0] m72_87;
   assign m72_87 =10'b0;

   // m72_88 = W*in
   wire signed [9:0] m72_88;
   assign m72_88 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_89 = W*in
   wire signed [9:0] m72_89;
   assign m72_89 ={ {4{in72[5]}} , in72[5:0] };

   // m72_90 = W*in
   wire signed [9:0] m72_90;
   assign m72_90 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_91 = W*in
   wire signed [9:0] m72_91;
   assign m72_91 =10'b0;

   // m72_92 = W*in
   wire signed [9:0] m72_92;
   assign m72_92 =10'b0;

   // m72_93 = W*in
   wire signed [9:0] m72_93;
   assign m72_93 =10'b0;

   // m72_94 = W*in
   wire signed [9:0] m72_94;
   assign m72_94 =10'b0;

   // m72_95 = W*in
   wire signed [9:0] m72_95;
   assign m72_95 =10'b0;

   // m72_96 = W*in
   wire signed [9:0] m72_96;
   assign m72_96 ={ {4{in72[5]}} , in72[5:0] };

   // m72_97 = W*in
   wire signed [9:0] m72_97;
   assign m72_97 ={ {4{neg72[5]}} , neg72[5:0] };

   // m72_98 = W*in
   wire signed [9:0] m72_98;
   assign m72_98 =10'b0;

   // m72_99 = W*in
   wire signed [9:0] m72_99;
   assign m72_99 =10'b0;

   // m72_100 = W*in
   wire signed [9:0] m72_100;
   assign m72_100 ={ {4{in72[5]}} , in72[5:0] };

   // m72_101 = W*in
   wire signed [9:0] m72_101;
   assign m72_101 =10'b0;

   // m72_102 = W*in
   wire signed [9:0] m72_102;
   assign m72_102 =10'b0;

   // m72_103 = W*in
   wire signed [9:0] m72_103;
   assign m72_103 =10'b0;

   // m72_104 = W*in
   wire signed [9:0] m72_104;
   assign m72_104 =10'b0;

   // m72_105 = W*in
   wire signed [9:0] m72_105;
   assign m72_105 =10'b0;

   // m72_106 = W*in
   wire signed [9:0] m72_106;
   assign m72_106 =10'b0;

   // m72_107 = W*in
   wire signed [9:0] m72_107;
   assign m72_107 =10'b0;

   // m72_108 = W*in
   wire signed [9:0] m72_108;
   assign m72_108 ={ {4{in72[5]}} , in72[5:0] };

   // m72_109 = W*in
   wire signed [9:0] m72_109;
   assign m72_109 ={ {4{in72[5]}} , in72[5:0] };

   // m72_110 = W*in
   wire signed [9:0] m72_110;
   assign m72_110 =10'b0;

   // m72_111 = W*in
   wire signed [9:0] m72_111;
   assign m72_111 =10'b0;

   // m72_112 = W*in
   wire signed [9:0] m72_112;
   assign m72_112 =10'b0;

   // m72_113 = W*in
   wire signed [9:0] m72_113;
   assign m72_113 =10'b0;

   // m72_114 = W*in
   wire signed [9:0] m72_114;
   assign m72_114 =10'b0;

   // m72_115 = W*in
   wire signed [9:0] m72_115;
   assign m72_115 =10'b0;

   // m72_116 = W*in
   wire signed [9:0] m72_116;
   assign m72_116 ={ {4{in72[5]}} , in72[5:0] };

   // m72_117 = W*in
   wire signed [9:0] m72_117;
   assign m72_117 =10'b0;

   // m73_1 = W*in
   wire signed [9:0] m73_1;
   assign m73_1 =10'b0;

   // m73_2 = W*in
   wire signed [9:0] m73_2;
   assign m73_2 =10'b0;

   // m73_3 = W*in
   wire signed [9:0] m73_3;
   assign m73_3 =10'b0;

   // m73_4 = W*in
   wire signed [9:0] m73_4;
   assign m73_4 =10'b0;

   // m73_5 = W*in
   wire signed [9:0] m73_5;
   assign m73_5 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_6 = W*in
   wire signed [9:0] m73_6;
   assign m73_6 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_7 = W*in
   wire signed [9:0] m73_7;
   assign m73_7 =10'b0;

   // m73_8 = W*in
   wire signed [9:0] m73_8;
   assign m73_8 =10'b0;

   // m73_9 = W*in
   wire signed [9:0] m73_9;
   assign m73_9 =10'b0;

   // m73_10 = W*in
   wire signed [9:0] m73_10;
   assign m73_10 =10'b0;

   // m73_11 = W*in
   wire signed [9:0] m73_11;
   assign m73_11 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_12 = W*in
   wire signed [9:0] m73_12;
   assign m73_12 =10'b0;

   // m73_13 = W*in
   wire signed [9:0] m73_13;
   assign m73_13 ={ {4{in73[5]}} , in73[5:0] };

   // m73_14 = W*in
   wire signed [9:0] m73_14;
   assign m73_14 =10'b0;

   // m73_15 = W*in
   wire signed [9:0] m73_15;
   assign m73_15 =10'b0;

   // m73_16 = W*in
   wire signed [9:0] m73_16;
   assign m73_16 =10'b0;

   // m73_17 = W*in
   wire signed [9:0] m73_17;
   assign m73_17 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_18 = W*in
   wire signed [9:0] m73_18;
   assign m73_18 =10'b0;

   // m73_19 = W*in
   wire signed [9:0] m73_19;
   assign m73_19 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_20 = W*in
   wire signed [9:0] m73_20;
   assign m73_20 =10'b0;

   // m73_21 = W*in
   wire signed [9:0] m73_21;
   assign m73_21 =10'b0;

   // m73_22 = W*in
   wire signed [9:0] m73_22;
   assign m73_22 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_23 = W*in
   wire signed [9:0] m73_23;
   assign m73_23 =10'b0;

   // m73_24 = W*in
   wire signed [9:0] m73_24;
   assign m73_24 =10'b0;

   // m73_25 = W*in
   wire signed [9:0] m73_25;
   assign m73_25 =10'b0;

   // m73_26 = W*in
   wire signed [9:0] m73_26;
   assign m73_26 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_27 = W*in
   wire signed [9:0] m73_27;
   assign m73_27 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_28 = W*in
   wire signed [9:0] m73_28;
   assign m73_28 =10'b0;

   // m73_29 = W*in
   wire signed [9:0] m73_29;
   assign m73_29 ={ {5{in73[5]}} , in73[5:1] };

   // m73_30 = W*in
   wire signed [9:0] m73_30;
   assign m73_30 ={ {4{in73[5]}} , in73[5:0] };

   // m73_31 = W*in
   wire signed [9:0] m73_31;
   assign m73_31 =10'b0;

   // m73_32 = W*in
   wire signed [9:0] m73_32;
   assign m73_32 =10'b0;

   // m73_33 = W*in
   wire signed [9:0] m73_33;
   assign m73_33 =10'b0;

   // m73_34 = W*in
   wire signed [9:0] m73_34;
   assign m73_34 =10'b0;

   // m73_35 = W*in
   wire signed [9:0] m73_35;
   assign m73_35 =10'b0;

   // m73_36 = W*in
   wire signed [9:0] m73_36;
   assign m73_36 =10'b0;

   // m73_37 = W*in
   wire signed [9:0] m73_37;
   assign m73_37 =10'b0;

   // m73_38 = W*in
   wire signed [9:0] m73_38;
   assign m73_38 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_39 = W*in
   wire signed [9:0] m73_39;
   assign m73_39 =10'b0;

   // m73_40 = W*in
   wire signed [9:0] m73_40;
   assign m73_40 =10'b0;

   // m73_41 = W*in
   wire signed [9:0] m73_41;
   assign m73_41 ={ {4{in73[5]}} , in73[5:0] };

   // m73_42 = W*in
   wire signed [9:0] m73_42;
   assign m73_42 =10'b0;

   // m73_43 = W*in
   wire signed [9:0] m73_43;
   assign m73_43 =10'b0;

   // m73_44 = W*in
   wire signed [9:0] m73_44;
   assign m73_44 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_45 = W*in
   wire signed [9:0] m73_45;
   assign m73_45 =10'b0;

   // m73_46 = W*in
   wire signed [9:0] m73_46;
   assign m73_46 =10'b0;

   // m73_47 = W*in
   wire signed [9:0] m73_47;
   assign m73_47 =10'b0;

   // m73_48 = W*in
   wire signed [9:0] m73_48;
   assign m73_48 =10'b0;

   // m73_49 = W*in
   wire signed [9:0] m73_49;
   assign m73_49 =10'b0;

   // m73_50 = W*in
   wire signed [9:0] m73_50;
   assign m73_50 =10'b0;

   // m73_51 = W*in
   wire signed [9:0] m73_51;
   assign m73_51 =10'b0;

   // m73_52 = W*in
   wire signed [9:0] m73_52;
   assign m73_52 =10'b0;

   // m73_53 = W*in
   wire signed [9:0] m73_53;
   assign m73_53 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_54 = W*in
   wire signed [9:0] m73_54;
   assign m73_54 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_55 = W*in
   wire signed [9:0] m73_55;
   assign m73_55 =10'b0;

   // m73_56 = W*in
   wire signed [9:0] m73_56;
   assign m73_56 =10'b0;

   // m73_57 = W*in
   wire signed [9:0] m73_57;
   assign m73_57 =10'b0;

   // m73_58 = W*in
   wire signed [9:0] m73_58;
   assign m73_58 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_59 = W*in
   wire signed [9:0] m73_59;
   assign m73_59 =10'b0;

   // m73_60 = W*in
   wire signed [9:0] m73_60;
   assign m73_60 =10'b0;

   // m73_61 = W*in
   wire signed [9:0] m73_61;
   assign m73_61 =10'b0;

   // m73_62 = W*in
   wire signed [9:0] m73_62;
   assign m73_62 =10'b0;

   // m73_63 = W*in
   wire signed [9:0] m73_63;
   assign m73_63 =10'b0;

   // m73_64 = W*in
   wire signed [9:0] m73_64;
   assign m73_64 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_65 = W*in
   wire signed [9:0] m73_65;
   assign m73_65 ={ {5{in73[5]}} , in73[5:1] };

   // m73_66 = W*in
   wire signed [9:0] m73_66;
   assign m73_66 ={ {5{in73[5]}} , in73[5:1] };

   // m73_67 = W*in
   wire signed [9:0] m73_67;
   assign m73_67 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_68 = W*in
   wire signed [9:0] m73_68;
   assign m73_68 =10'b0;

   // m73_69 = W*in
   wire signed [9:0] m73_69;
   assign m73_69 =10'b0;

   // m73_70 = W*in
   wire signed [9:0] m73_70;
   assign m73_70 =10'b0;

   // m73_71 = W*in
   wire signed [9:0] m73_71;
   assign m73_71 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_72 = W*in
   wire signed [9:0] m73_72;
   assign m73_72 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_73 = W*in
   wire signed [9:0] m73_73;
   assign m73_73 =10'b0;

   // m73_74 = W*in
   wire signed [9:0] m73_74;
   assign m73_74 ={ {5{neg73[5]}} , neg73[5:1] };

   // m73_75 = W*in
   wire signed [9:0] m73_75;
   assign m73_75 ={ {4{in73[5]}} , in73[5:0] };

   // m73_76 = W*in
   wire signed [9:0] m73_76;
   assign m73_76 =10'b0;

   // m73_77 = W*in
   wire signed [9:0] m73_77;
   assign m73_77 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_78 = W*in
   wire signed [9:0] m73_78;
   assign m73_78 =10'b0;

   // m73_79 = W*in
   wire signed [9:0] m73_79;
   assign m73_79 =10'b0;

   // m73_80 = W*in
   wire signed [9:0] m73_80;
   assign m73_80 =10'b0;

   // m73_81 = W*in
   wire signed [9:0] m73_81;
   assign m73_81 =10'b0;

   // m73_82 = W*in
   wire signed [9:0] m73_82;
   assign m73_82 =10'b0;

   // m73_83 = W*in
   wire signed [9:0] m73_83;
   assign m73_83 =10'b0;

   // m73_84 = W*in
   wire signed [9:0] m73_84;
   assign m73_84 =10'b0;

   // m73_85 = W*in
   wire signed [9:0] m73_85;
   assign m73_85 =10'b0;

   // m73_86 = W*in
   wire signed [9:0] m73_86;
   assign m73_86 =10'b0;

   // m73_87 = W*in
   wire signed [9:0] m73_87;
   assign m73_87 =10'b0;

   // m73_88 = W*in
   wire signed [9:0] m73_88;
   assign m73_88 =10'b0;

   // m73_89 = W*in
   wire signed [9:0] m73_89;
   assign m73_89 ={ {4{in73[5]}} , in73[5:0] };

   // m73_90 = W*in
   wire signed [9:0] m73_90;
   assign m73_90 =10'b0;

   // m73_91 = W*in
   wire signed [9:0] m73_91;
   assign m73_91 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_92 = W*in
   wire signed [9:0] m73_92;
   assign m73_92 =10'b0;

   // m73_93 = W*in
   wire signed [9:0] m73_93;
   assign m73_93 =10'b0;

   // m73_94 = W*in
   wire signed [9:0] m73_94;
   assign m73_94 ={ {4{in73[5]}} , in73[5:0] };

   // m73_95 = W*in
   wire signed [9:0] m73_95;
   assign m73_95 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_96 = W*in
   wire signed [9:0] m73_96;
   assign m73_96 ={ {4{in73[5]}} , in73[5:0] };

   // m73_97 = W*in
   wire signed [9:0] m73_97;
   assign m73_97 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_98 = W*in
   wire signed [9:0] m73_98;
   assign m73_98 =10'b0;

   // m73_99 = W*in
   wire signed [9:0] m73_99;
   assign m73_99 =10'b0;

   // m73_100 = W*in
   wire signed [9:0] m73_100;
   assign m73_100 =10'b0;

   // m73_101 = W*in
   wire signed [9:0] m73_101;
   assign m73_101 =10'b0;

   // m73_102 = W*in
   wire signed [9:0] m73_102;
   assign m73_102 =10'b0;

   // m73_103 = W*in
   wire signed [9:0] m73_103;
   assign m73_103 =10'b0;

   // m73_104 = W*in
   wire signed [9:0] m73_104;
   assign m73_104 =10'b0;

   // m73_105 = W*in
   wire signed [9:0] m73_105;
   assign m73_105 =10'b0;

   // m73_106 = W*in
   wire signed [9:0] m73_106;
   assign m73_106 =10'b0;

   // m73_107 = W*in
   wire signed [9:0] m73_107;
   assign m73_107 =10'b0;

   // m73_108 = W*in
   wire signed [9:0] m73_108;
   assign m73_108 ={ {4{in73[5]}} , in73[5:0] };

   // m73_109 = W*in
   wire signed [9:0] m73_109;
   assign m73_109 =10'b0;

   // m73_110 = W*in
   wire signed [9:0] m73_110;
   assign m73_110 ={ {4{neg73[5]}} , neg73[5:0] };

   // m73_111 = W*in
   wire signed [9:0] m73_111;
   assign m73_111 =10'b0;

   // m73_112 = W*in
   wire signed [9:0] m73_112;
   assign m73_112 =10'b0;

   // m73_113 = W*in
   wire signed [9:0] m73_113;
   assign m73_113 =10'b0;

   // m73_114 = W*in
   wire signed [9:0] m73_114;
   assign m73_114 =10'b0;

   // m73_115 = W*in
   wire signed [9:0] m73_115;
   assign m73_115 =10'b0;

   // m73_116 = W*in
   wire signed [9:0] m73_116;
   assign m73_116 ={ {4{in73[5]}} , in73[5:0] };

   // m73_117 = W*in
   wire signed [9:0] m73_117;
   assign m73_117 ={ {4{neg73[5]}} , neg73[5:0] };

   // m74_1 = W*in
   wire signed [9:0] m74_1;
   assign m74_1 =10'b0;

   // m74_2 = W*in
   wire signed [9:0] m74_2;
   assign m74_2 =10'b0;

   // m74_3 = W*in
   wire signed [9:0] m74_3;
   assign m74_3 =10'b0;

   // m74_4 = W*in
   wire signed [9:0] m74_4;
   assign m74_4 =10'b0;

   // m74_5 = W*in
   wire signed [9:0] m74_5;
   assign m74_5 =10'b0;

   // m74_6 = W*in
   wire signed [9:0] m74_6;
   assign m74_6 =10'b0;

   // m74_7 = W*in
   wire signed [9:0] m74_7;
   assign m74_7 =10'b0;

   // m74_8 = W*in
   wire signed [9:0] m74_8;
   assign m74_8 =10'b0;

   // m74_9 = W*in
   wire signed [9:0] m74_9;
   assign m74_9 =10'b0;

   // m74_10 = W*in
   wire signed [9:0] m74_10;
   assign m74_10 =10'b0;

   // m74_11 = W*in
   wire signed [9:0] m74_11;
   assign m74_11 =10'b0;

   // m74_12 = W*in
   wire signed [9:0] m74_12;
   assign m74_12 =10'b0;

   // m74_13 = W*in
   wire signed [9:0] m74_13;
   assign m74_13 =10'b0;

   // m74_14 = W*in
   wire signed [9:0] m74_14;
   assign m74_14 =10'b0;

   // m74_15 = W*in
   wire signed [9:0] m74_15;
   assign m74_15 =10'b0;

   // m74_16 = W*in
   wire signed [9:0] m74_16;
   assign m74_16 =10'b0;

   // m74_17 = W*in
   wire signed [9:0] m74_17;
   assign m74_17 ={ {5{neg74[5]}} , neg74[5:1] };

   // m74_18 = W*in
   wire signed [9:0] m74_18;
   assign m74_18 ={ {5{in74[5]}} , in74[5:1] };

   // m74_19 = W*in
   wire signed [9:0] m74_19;
   assign m74_19 ={ {5{neg74[5]}} , neg74[5:1] };

   // m74_20 = W*in
   wire signed [9:0] m74_20;
   assign m74_20 ={ {5{neg74[5]}} , neg74[5:1] };

   // m74_21 = W*in
   wire signed [9:0] m74_21;
   assign m74_21 =10'b0;

   // m74_22 = W*in
   wire signed [9:0] m74_22;
   assign m74_22 =10'b0;

   // m74_23 = W*in
   wire signed [9:0] m74_23;
   assign m74_23 =10'b0;

   // m74_24 = W*in
   wire signed [9:0] m74_24;
   assign m74_24 =10'b0;

   // m74_25 = W*in
   wire signed [9:0] m74_25;
   assign m74_25 =10'b0;

   // m74_26 = W*in
   wire signed [9:0] m74_26;
   assign m74_26 ={ {5{in74[5]}} , in74[5:1] };

   // m74_27 = W*in
   wire signed [9:0] m74_27;
   assign m74_27 =10'b0;

   // m74_28 = W*in
   wire signed [9:0] m74_28;
   assign m74_28 =10'b0;

   // m74_29 = W*in
   wire signed [9:0] m74_29;
   assign m74_29 ={ {5{in74[5]}} , in74[5:1] };

   // m74_30 = W*in
   wire signed [9:0] m74_30;
   assign m74_30 =10'b0;

   // m74_31 = W*in
   wire signed [9:0] m74_31;
   assign m74_31 =10'b0;

   // m74_32 = W*in
   wire signed [9:0] m74_32;
   assign m74_32 =10'b0;

   // m74_33 = W*in
   wire signed [9:0] m74_33;
   assign m74_33 =10'b0;

   // m74_34 = W*in
   wire signed [9:0] m74_34;
   assign m74_34 =10'b0;

   // m74_35 = W*in
   wire signed [9:0] m74_35;
   assign m74_35 =10'b0;

   // m74_36 = W*in
   wire signed [9:0] m74_36;
   assign m74_36 =10'b0;

   // m74_37 = W*in
   wire signed [9:0] m74_37;
   assign m74_37 =10'b0;

   // m74_38 = W*in
   wire signed [9:0] m74_38;
   assign m74_38 =10'b0;

   // m74_39 = W*in
   wire signed [9:0] m74_39;
   assign m74_39 =10'b0;

   // m74_40 = W*in
   wire signed [9:0] m74_40;
   assign m74_40 =10'b0;

   // m74_41 = W*in
   wire signed [9:0] m74_41;
   assign m74_41 =10'b0;

   // m74_42 = W*in
   wire signed [9:0] m74_42;
   assign m74_42 =10'b0;

   // m74_43 = W*in
   wire signed [9:0] m74_43;
   assign m74_43 =10'b0;

   // m74_44 = W*in
   wire signed [9:0] m74_44;
   assign m74_44 ={ {4{neg74[5]}} , neg74[5:0] };

   // m74_45 = W*in
   wire signed [9:0] m74_45;
   assign m74_45 =10'b0;

   // m74_46 = W*in
   wire signed [9:0] m74_46;
   assign m74_46 =10'b0;

   // m74_47 = W*in
   wire signed [9:0] m74_47;
   assign m74_47 =10'b0;

   // m74_48 = W*in
   wire signed [9:0] m74_48;
   assign m74_48 =10'b0;

   // m74_49 = W*in
   wire signed [9:0] m74_49;
   assign m74_49 =10'b0;

   // m74_50 = W*in
   wire signed [9:0] m74_50;
   assign m74_50 =10'b0;

   // m74_51 = W*in
   wire signed [9:0] m74_51;
   assign m74_51 =10'b0;

   // m74_52 = W*in
   wire signed [9:0] m74_52;
   assign m74_52 =10'b0;

   // m74_53 = W*in
   wire signed [9:0] m74_53;
   assign m74_53 =10'b0;

   // m74_54 = W*in
   wire signed [9:0] m74_54;
   assign m74_54 ={ {4{neg74[5]}} , neg74[5:0] };

   // m74_55 = W*in
   wire signed [9:0] m74_55;
   assign m74_55 =10'b0;

   // m74_56 = W*in
   wire signed [9:0] m74_56;
   assign m74_56 =10'b0;

   // m74_57 = W*in
   wire signed [9:0] m74_57;
   assign m74_57 =10'b0;

   // m74_58 = W*in
   wire signed [9:0] m74_58;
   assign m74_58 =10'b0;

   // m74_59 = W*in
   wire signed [9:0] m74_59;
   assign m74_59 =10'b0;

   // m74_60 = W*in
   wire signed [9:0] m74_60;
   assign m74_60 =10'b0;

   // m74_61 = W*in
   wire signed [9:0] m74_61;
   assign m74_61 =10'b0;

   // m74_62 = W*in
   wire signed [9:0] m74_62;
   assign m74_62 =10'b0;

   // m74_63 = W*in
   wire signed [9:0] m74_63;
   assign m74_63 =10'b0;

   // m74_64 = W*in
   wire signed [9:0] m74_64;
   assign m74_64 =10'b0;

   // m74_65 = W*in
   wire signed [9:0] m74_65;
   assign m74_65 =10'b0;

   // m74_66 = W*in
   wire signed [9:0] m74_66;
   assign m74_66 =10'b0;

   // m74_67 = W*in
   wire signed [9:0] m74_67;
   assign m74_67 =10'b0;

   // m74_68 = W*in
   wire signed [9:0] m74_68;
   assign m74_68 =10'b0;

   // m74_69 = W*in
   wire signed [9:0] m74_69;
   assign m74_69 =10'b0;

   // m74_70 = W*in
   wire signed [9:0] m74_70;
   assign m74_70 ={ {5{in74[5]}} , in74[5:1] };

   // m74_71 = W*in
   wire signed [9:0] m74_71;
   assign m74_71 =10'b0;

   // m74_72 = W*in
   wire signed [9:0] m74_72;
   assign m74_72 =10'b0;

   // m74_73 = W*in
   wire signed [9:0] m74_73;
   assign m74_73 =10'b0;

   // m74_74 = W*in
   wire signed [9:0] m74_74;
   assign m74_74 =10'b0;

   // m74_75 = W*in
   wire signed [9:0] m74_75;
   assign m74_75 ={ {5{neg74[5]}} , neg74[5:1] };

   // m74_76 = W*in
   wire signed [9:0] m74_76;
   assign m74_76 =10'b0;

   // m74_77 = W*in
   wire signed [9:0] m74_77;
   assign m74_77 =10'b0;

   // m74_78 = W*in
   wire signed [9:0] m74_78;
   assign m74_78 =10'b0;

   // m74_79 = W*in
   wire signed [9:0] m74_79;
   assign m74_79 =10'b0;

   // m74_80 = W*in
   wire signed [9:0] m74_80;
   assign m74_80 =10'b0;

   // m74_81 = W*in
   wire signed [9:0] m74_81;
   assign m74_81 =10'b0;

   // m74_82 = W*in
   wire signed [9:0] m74_82;
   assign m74_82 =10'b0;

   // m74_83 = W*in
   wire signed [9:0] m74_83;
   assign m74_83 =10'b0;

   // m74_84 = W*in
   wire signed [9:0] m74_84;
   assign m74_84 =10'b0;

   // m74_85 = W*in
   wire signed [9:0] m74_85;
   assign m74_85 =10'b0;

   // m74_86 = W*in
   wire signed [9:0] m74_86;
   assign m74_86 =10'b0;

   // m74_87 = W*in
   wire signed [9:0] m74_87;
   assign m74_87 =10'b0;

   // m74_88 = W*in
   wire signed [9:0] m74_88;
   assign m74_88 =10'b0;

   // m74_89 = W*in
   wire signed [9:0] m74_89;
   assign m74_89 =10'b0;

   // m74_90 = W*in
   wire signed [9:0] m74_90;
   assign m74_90 =10'b0;

   // m74_91 = W*in
   wire signed [9:0] m74_91;
   assign m74_91 =10'b0;

   // m74_92 = W*in
   wire signed [9:0] m74_92;
   assign m74_92 =10'b0;

   // m74_93 = W*in
   wire signed [9:0] m74_93;
   assign m74_93 =10'b0;

   // m74_94 = W*in
   wire signed [9:0] m74_94;
   assign m74_94 =10'b0;

   // m74_95 = W*in
   wire signed [9:0] m74_95;
   assign m74_95 =10'b0;

   // m74_96 = W*in
   wire signed [9:0] m74_96;
   assign m74_96 =10'b0;

   // m74_97 = W*in
   wire signed [9:0] m74_97;
   assign m74_97 =10'b0;

   // m74_98 = W*in
   wire signed [9:0] m74_98;
   assign m74_98 =10'b0;

   // m74_99 = W*in
   wire signed [9:0] m74_99;
   assign m74_99 =10'b0;

   // m74_100 = W*in
   wire signed [9:0] m74_100;
   assign m74_100 =10'b0;

   // m74_101 = W*in
   wire signed [9:0] m74_101;
   assign m74_101 =10'b0;

   // m74_102 = W*in
   wire signed [9:0] m74_102;
   assign m74_102 =10'b0;

   // m74_103 = W*in
   wire signed [9:0] m74_103;
   assign m74_103 =10'b0;

   // m74_104 = W*in
   wire signed [9:0] m74_104;
   assign m74_104 =10'b0;

   // m74_105 = W*in
   wire signed [9:0] m74_105;
   assign m74_105 =10'b0;

   // m74_106 = W*in
   wire signed [9:0] m74_106;
   assign m74_106 =10'b0;

   // m74_107 = W*in
   wire signed [9:0] m74_107;
   assign m74_107 =10'b0;

   // m74_108 = W*in
   wire signed [9:0] m74_108;
   assign m74_108 ={ {5{in74[5]}} , in74[5:1] };

   // m74_109 = W*in
   wire signed [9:0] m74_109;
   assign m74_109 =10'b0;

   // m74_110 = W*in
   wire signed [9:0] m74_110;
   assign m74_110 =10'b0;

   // m74_111 = W*in
   wire signed [9:0] m74_111;
   assign m74_111 =10'b0;

   // m74_112 = W*in
   wire signed [9:0] m74_112;
   assign m74_112 =10'b0;

   // m74_113 = W*in
   wire signed [9:0] m74_113;
   assign m74_113 =10'b0;

   // m74_114 = W*in
   wire signed [9:0] m74_114;
   assign m74_114 =10'b0;

   // m74_115 = W*in
   wire signed [9:0] m74_115;
   assign m74_115 =10'b0;

   // m74_116 = W*in
   wire signed [9:0] m74_116;
   assign m74_116 =10'b0;

   // m74_117 = W*in
   wire signed [9:0] m74_117;
   assign m74_117 =10'b0;

   // m75_1 = W*in
   wire signed [9:0] m75_1;
   assign m75_1 =10'b0;

   // m75_2 = W*in
   wire signed [9:0] m75_2;
   assign m75_2 =10'b0;

   // m75_3 = W*in
   wire signed [9:0] m75_3;
   assign m75_3 =10'b0;

   // m75_4 = W*in
   wire signed [9:0] m75_4;
   assign m75_4 =10'b0;

   // m75_5 = W*in
   wire signed [9:0] m75_5;
   assign m75_5 =10'b0;

   // m75_6 = W*in
   wire signed [9:0] m75_6;
   assign m75_6 =10'b0;

   // m75_7 = W*in
   wire signed [9:0] m75_7;
   assign m75_7 =10'b0;

   // m75_8 = W*in
   wire signed [9:0] m75_8;
   assign m75_8 =10'b0;

   // m75_9 = W*in
   wire signed [9:0] m75_9;
   assign m75_9 =10'b0;

   // m75_10 = W*in
   wire signed [9:0] m75_10;
   assign m75_10 =10'b0;

   // m75_11 = W*in
   wire signed [9:0] m75_11;
   assign m75_11 =10'b0;

   // m75_12 = W*in
   wire signed [9:0] m75_12;
   assign m75_12 =10'b0;

   // m75_13 = W*in
   wire signed [9:0] m75_13;
   assign m75_13 =10'b0;

   // m75_14 = W*in
   wire signed [9:0] m75_14;
   assign m75_14 =10'b0;

   // m75_15 = W*in
   wire signed [9:0] m75_15;
   assign m75_15 =10'b0;

   // m75_16 = W*in
   wire signed [9:0] m75_16;
   assign m75_16 =10'b0;

   // m75_17 = W*in
   wire signed [9:0] m75_17;
   assign m75_17 =10'b0;

   // m75_18 = W*in
   wire signed [9:0] m75_18;
   assign m75_18 =10'b0;

   // m75_19 = W*in
   wire signed [9:0] m75_19;
   assign m75_19 ={ {5{neg75[5]}} , neg75[5:1] };

   // m75_20 = W*in
   wire signed [9:0] m75_20;
   assign m75_20 =10'b0;

   // m75_21 = W*in
   wire signed [9:0] m75_21;
   assign m75_21 =10'b0;

   // m75_22 = W*in
   wire signed [9:0] m75_22;
   assign m75_22 =10'b0;

   // m75_23 = W*in
   wire signed [9:0] m75_23;
   assign m75_23 =10'b0;

   // m75_24 = W*in
   wire signed [9:0] m75_24;
   assign m75_24 =10'b0;

   // m75_25 = W*in
   wire signed [9:0] m75_25;
   assign m75_25 =10'b0;

   // m75_26 = W*in
   wire signed [9:0] m75_26;
   assign m75_26 =10'b0;

   // m75_27 = W*in
   wire signed [9:0] m75_27;
   assign m75_27 =10'b0;

   // m75_28 = W*in
   wire signed [9:0] m75_28;
   assign m75_28 ={ {5{neg75[5]}} , neg75[5:1] };

   // m75_29 = W*in
   wire signed [9:0] m75_29;
   assign m75_29 =10'b0;

   // m75_30 = W*in
   wire signed [9:0] m75_30;
   assign m75_30 =10'b0;

   // m75_31 = W*in
   wire signed [9:0] m75_31;
   assign m75_31 =10'b0;

   // m75_32 = W*in
   wire signed [9:0] m75_32;
   assign m75_32 =10'b0;

   // m75_33 = W*in
   wire signed [9:0] m75_33;
   assign m75_33 =10'b0;

   // m75_34 = W*in
   wire signed [9:0] m75_34;
   assign m75_34 =10'b0;

   // m75_35 = W*in
   wire signed [9:0] m75_35;
   assign m75_35 =10'b0;

   // m75_36 = W*in
   wire signed [9:0] m75_36;
   assign m75_36 =10'b0;

   // m75_37 = W*in
   wire signed [9:0] m75_37;
   assign m75_37 =10'b0;

   // m75_38 = W*in
   wire signed [9:0] m75_38;
   assign m75_38 =10'b0;

   // m75_39 = W*in
   wire signed [9:0] m75_39;
   assign m75_39 =10'b0;

   // m75_40 = W*in
   wire signed [9:0] m75_40;
   assign m75_40 =10'b0;

   // m75_41 = W*in
   wire signed [9:0] m75_41;
   assign m75_41 =10'b0;

   // m75_42 = W*in
   wire signed [9:0] m75_42;
   assign m75_42 =10'b0;

   // m75_43 = W*in
   wire signed [9:0] m75_43;
   assign m75_43 =10'b0;

   // m75_44 = W*in
   wire signed [9:0] m75_44;
   assign m75_44 =10'b0;

   // m75_45 = W*in
   wire signed [9:0] m75_45;
   assign m75_45 =10'b0;

   // m75_46 = W*in
   wire signed [9:0] m75_46;
   assign m75_46 =10'b0;

   // m75_47 = W*in
   wire signed [9:0] m75_47;
   assign m75_47 =10'b0;

   // m75_48 = W*in
   wire signed [9:0] m75_48;
   assign m75_48 =10'b0;

   // m75_49 = W*in
   wire signed [9:0] m75_49;
   assign m75_49 =10'b0;

   // m75_50 = W*in
   wire signed [9:0] m75_50;
   assign m75_50 =10'b0;

   // m75_51 = W*in
   wire signed [9:0] m75_51;
   assign m75_51 =10'b0;

   // m75_52 = W*in
   wire signed [9:0] m75_52;
   assign m75_52 =10'b0;

   // m75_53 = W*in
   wire signed [9:0] m75_53;
   assign m75_53 =10'b0;

   // m75_54 = W*in
   wire signed [9:0] m75_54;
   assign m75_54 =10'b0;

   // m75_55 = W*in
   wire signed [9:0] m75_55;
   assign m75_55 =10'b0;

   // m75_56 = W*in
   wire signed [9:0] m75_56;
   assign m75_56 =10'b0;

   // m75_57 = W*in
   wire signed [9:0] m75_57;
   assign m75_57 =10'b0;

   // m75_58 = W*in
   wire signed [9:0] m75_58;
   assign m75_58 =10'b0;

   // m75_59 = W*in
   wire signed [9:0] m75_59;
   assign m75_59 =10'b0;

   // m75_60 = W*in
   wire signed [9:0] m75_60;
   assign m75_60 =10'b0;

   // m75_61 = W*in
   wire signed [9:0] m75_61;
   assign m75_61 =10'b0;

   // m75_62 = W*in
   wire signed [9:0] m75_62;
   assign m75_62 =10'b0;

   // m75_63 = W*in
   wire signed [9:0] m75_63;
   assign m75_63 =10'b0;

   // m75_64 = W*in
   wire signed [9:0] m75_64;
   assign m75_64 =10'b0;

   // m75_65 = W*in
   wire signed [9:0] m75_65;
   assign m75_65 =10'b0;

   // m75_66 = W*in
   wire signed [9:0] m75_66;
   assign m75_66 =10'b0;

   // m75_67 = W*in
   wire signed [9:0] m75_67;
   assign m75_67 =10'b0;

   // m75_68 = W*in
   wire signed [9:0] m75_68;
   assign m75_68 =10'b0;

   // m75_69 = W*in
   wire signed [9:0] m75_69;
   assign m75_69 =10'b0;

   // m75_70 = W*in
   wire signed [9:0] m75_70;
   assign m75_70 =10'b0;

   // m75_71 = W*in
   wire signed [9:0] m75_71;
   assign m75_71 =10'b0;

   // m75_72 = W*in
   wire signed [9:0] m75_72;
   assign m75_72 ={ {5{in75[5]}} , in75[5:1] };

   // m75_73 = W*in
   wire signed [9:0] m75_73;
   assign m75_73 =10'b0;

   // m75_74 = W*in
   wire signed [9:0] m75_74;
   assign m75_74 =10'b0;

   // m75_75 = W*in
   wire signed [9:0] m75_75;
   assign m75_75 =10'b0;

   // m75_76 = W*in
   wire signed [9:0] m75_76;
   assign m75_76 =10'b0;

   // m75_77 = W*in
   wire signed [9:0] m75_77;
   assign m75_77 =10'b0;

   // m75_78 = W*in
   wire signed [9:0] m75_78;
   assign m75_78 =10'b0;

   // m75_79 = W*in
   wire signed [9:0] m75_79;
   assign m75_79 =10'b0;

   // m75_80 = W*in
   wire signed [9:0] m75_80;
   assign m75_80 =10'b0;

   // m75_81 = W*in
   wire signed [9:0] m75_81;
   assign m75_81 =10'b0;

   // m75_82 = W*in
   wire signed [9:0] m75_82;
   assign m75_82 =10'b0;

   // m75_83 = W*in
   wire signed [9:0] m75_83;
   assign m75_83 =10'b0;

   // m75_84 = W*in
   wire signed [9:0] m75_84;
   assign m75_84 =10'b0;

   // m75_85 = W*in
   wire signed [9:0] m75_85;
   assign m75_85 =10'b0;

   // m75_86 = W*in
   wire signed [9:0] m75_86;
   assign m75_86 =10'b0;

   // m75_87 = W*in
   wire signed [9:0] m75_87;
   assign m75_87 =10'b0;

   // m75_88 = W*in
   wire signed [9:0] m75_88;
   assign m75_88 =10'b0;

   // m75_89 = W*in
   wire signed [9:0] m75_89;
   assign m75_89 =10'b0;

   // m75_90 = W*in
   wire signed [9:0] m75_90;
   assign m75_90 =10'b0;

   // m75_91 = W*in
   wire signed [9:0] m75_91;
   assign m75_91 =10'b0;

   // m75_92 = W*in
   wire signed [9:0] m75_92;
   assign m75_92 =10'b0;

   // m75_93 = W*in
   wire signed [9:0] m75_93;
   assign m75_93 =10'b0;

   // m75_94 = W*in
   wire signed [9:0] m75_94;
   assign m75_94 =10'b0;

   // m75_95 = W*in
   wire signed [9:0] m75_95;
   assign m75_95 =10'b0;

   // m75_96 = W*in
   wire signed [9:0] m75_96;
   assign m75_96 =10'b0;

   // m75_97 = W*in
   wire signed [9:0] m75_97;
   assign m75_97 =10'b0;

   // m75_98 = W*in
   wire signed [9:0] m75_98;
   assign m75_98 =10'b0;

   // m75_99 = W*in
   wire signed [9:0] m75_99;
   assign m75_99 =10'b0;

   // m75_100 = W*in
   wire signed [9:0] m75_100;
   assign m75_100 =10'b0;

   // m75_101 = W*in
   wire signed [9:0] m75_101;
   assign m75_101 =10'b0;

   // m75_102 = W*in
   wire signed [9:0] m75_102;
   assign m75_102 =10'b0;

   // m75_103 = W*in
   wire signed [9:0] m75_103;
   assign m75_103 =10'b0;

   // m75_104 = W*in
   wire signed [9:0] m75_104;
   assign m75_104 =10'b0;

   // m75_105 = W*in
   wire signed [9:0] m75_105;
   assign m75_105 =10'b0;

   // m75_106 = W*in
   wire signed [9:0] m75_106;
   assign m75_106 =10'b0;

   // m75_107 = W*in
   wire signed [9:0] m75_107;
   assign m75_107 =10'b0;

   // m75_108 = W*in
   wire signed [9:0] m75_108;
   assign m75_108 =10'b0;

   // m75_109 = W*in
   wire signed [9:0] m75_109;
   assign m75_109 =10'b0;

   // m75_110 = W*in
   wire signed [9:0] m75_110;
   assign m75_110 =10'b0;

   // m75_111 = W*in
   wire signed [9:0] m75_111;
   assign m75_111 =10'b0;

   // m75_112 = W*in
   wire signed [9:0] m75_112;
   assign m75_112 =10'b0;

   // m75_113 = W*in
   wire signed [9:0] m75_113;
   assign m75_113 =10'b0;

   // m75_114 = W*in
   wire signed [9:0] m75_114;
   assign m75_114 =10'b0;

   // m75_115 = W*in
   wire signed [9:0] m75_115;
   assign m75_115 =10'b0;

   // m75_116 = W*in
   wire signed [9:0] m75_116;
   assign m75_116 =10'b0;

   // m75_117 = W*in
   wire signed [9:0] m75_117;
   assign m75_117 =10'b0;

   // m76_1 = W*in
   wire signed [9:0] m76_1;
   assign m76_1 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_2 = W*in
   wire signed [9:0] m76_2;
   assign m76_2 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_3 = W*in
   wire signed [9:0] m76_3;
   assign m76_3 =10'b0;

   // m76_4 = W*in
   wire signed [9:0] m76_4;
   assign m76_4 =10'b0;

   // m76_5 = W*in
   wire signed [9:0] m76_5;
   assign m76_5 =10'b0;

   // m76_6 = W*in
   wire signed [9:0] m76_6;
   assign m76_6 =10'b0;

   // m76_7 = W*in
   wire signed [9:0] m76_7;
   assign m76_7 =10'b0;

   // m76_8 = W*in
   wire signed [9:0] m76_8;
   assign m76_8 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_9 = W*in
   wire signed [9:0] m76_9;
   assign m76_9 =10'b0;

   // m76_10 = W*in
   wire signed [9:0] m76_10;
   assign m76_10 =10'b0;

   // m76_11 = W*in
   wire signed [9:0] m76_11;
   assign m76_11 =10'b0;

   // m76_12 = W*in
   wire signed [9:0] m76_12;
   assign m76_12 =10'b0;

   // m76_13 = W*in
   wire signed [9:0] m76_13;
   assign m76_13 =10'b0;

   // m76_14 = W*in
   wire signed [9:0] m76_14;
   assign m76_14 =10'b0;

   // m76_15 = W*in
   wire signed [9:0] m76_15;
   assign m76_15 =10'b0;

   // m76_16 = W*in
   wire signed [9:0] m76_16;
   assign m76_16 =10'b0;

   // m76_17 = W*in
   wire signed [9:0] m76_17;
   assign m76_17 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_18 = W*in
   wire signed [9:0] m76_18;
   assign m76_18 ={ {5{in76[5]}} , in76[5:1] };

   // m76_19 = W*in
   wire signed [9:0] m76_19;
   assign m76_19 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_20 = W*in
   wire signed [9:0] m76_20;
   assign m76_20 =10'b0;

   // m76_21 = W*in
   wire signed [9:0] m76_21;
   assign m76_21 =10'b0;

   // m76_22 = W*in
   wire signed [9:0] m76_22;
   assign m76_22 =10'b0;

   // m76_23 = W*in
   wire signed [9:0] m76_23;
   assign m76_23 =10'b0;

   // m76_24 = W*in
   wire signed [9:0] m76_24;
   assign m76_24 =10'b0;

   // m76_25 = W*in
   wire signed [9:0] m76_25;
   assign m76_25 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_26 = W*in
   wire signed [9:0] m76_26;
   assign m76_26 =10'b0;

   // m76_27 = W*in
   wire signed [9:0] m76_27;
   assign m76_27 =10'b0;

   // m76_28 = W*in
   wire signed [9:0] m76_28;
   assign m76_28 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_29 = W*in
   wire signed [9:0] m76_29;
   assign m76_29 =10'b0;

   // m76_30 = W*in
   wire signed [9:0] m76_30;
   assign m76_30 =10'b0;

   // m76_31 = W*in
   wire signed [9:0] m76_31;
   assign m76_31 =10'b0;

   // m76_32 = W*in
   wire signed [9:0] m76_32;
   assign m76_32 =10'b0;

   // m76_33 = W*in
   wire signed [9:0] m76_33;
   assign m76_33 =10'b0;

   // m76_34 = W*in
   wire signed [9:0] m76_34;
   assign m76_34 =10'b0;

   // m76_35 = W*in
   wire signed [9:0] m76_35;
   assign m76_35 =10'b0;

   // m76_36 = W*in
   wire signed [9:0] m76_36;
   assign m76_36 =10'b0;

   // m76_37 = W*in
   wire signed [9:0] m76_37;
   assign m76_37 =10'b0;

   // m76_38 = W*in
   wire signed [9:0] m76_38;
   assign m76_38 =10'b0;

   // m76_39 = W*in
   wire signed [9:0] m76_39;
   assign m76_39 =10'b0;

   // m76_40 = W*in
   wire signed [9:0] m76_40;
   assign m76_40 =10'b0;

   // m76_41 = W*in
   wire signed [9:0] m76_41;
   assign m76_41 =10'b0;

   // m76_42 = W*in
   wire signed [9:0] m76_42;
   assign m76_42 =10'b0;

   // m76_43 = W*in
   wire signed [9:0] m76_43;
   assign m76_43 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_44 = W*in
   wire signed [9:0] m76_44;
   assign m76_44 ={ {5{neg76[5]}} , neg76[5:1] };

   // m76_45 = W*in
   wire signed [9:0] m76_45;
   assign m76_45 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_46 = W*in
   wire signed [9:0] m76_46;
   assign m76_46 =10'b0;

   // m76_47 = W*in
   wire signed [9:0] m76_47;
   assign m76_47 =10'b0;

   // m76_48 = W*in
   wire signed [9:0] m76_48;
   assign m76_48 =10'b0;

   // m76_49 = W*in
   wire signed [9:0] m76_49;
   assign m76_49 =10'b0;

   // m76_50 = W*in
   wire signed [9:0] m76_50;
   assign m76_50 =10'b0;

   // m76_51 = W*in
   wire signed [9:0] m76_51;
   assign m76_51 =10'b0;

   // m76_52 = W*in
   wire signed [9:0] m76_52;
   assign m76_52 =10'b0;

   // m76_53 = W*in
   wire signed [9:0] m76_53;
   assign m76_53 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_54 = W*in
   wire signed [9:0] m76_54;
   assign m76_54 =10'b0;

   // m76_55 = W*in
   wire signed [9:0] m76_55;
   assign m76_55 =10'b0;

   // m76_56 = W*in
   wire signed [9:0] m76_56;
   assign m76_56 =10'b0;

   // m76_57 = W*in
   wire signed [9:0] m76_57;
   assign m76_57 =10'b0;

   // m76_58 = W*in
   wire signed [9:0] m76_58;
   assign m76_58 =10'b0;

   // m76_59 = W*in
   wire signed [9:0] m76_59;
   assign m76_59 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_60 = W*in
   wire signed [9:0] m76_60;
   assign m76_60 =10'b0;

   // m76_61 = W*in
   wire signed [9:0] m76_61;
   assign m76_61 =10'b0;

   // m76_62 = W*in
   wire signed [9:0] m76_62;
   assign m76_62 =10'b0;

   // m76_63 = W*in
   wire signed [9:0] m76_63;
   assign m76_63 =10'b0;

   // m76_64 = W*in
   wire signed [9:0] m76_64;
   assign m76_64 =10'b0;

   // m76_65 = W*in
   wire signed [9:0] m76_65;
   assign m76_65 ={ {5{in76[5]}} , in76[5:1] };

   // m76_66 = W*in
   wire signed [9:0] m76_66;
   assign m76_66 =10'b0;

   // m76_67 = W*in
   wire signed [9:0] m76_67;
   assign m76_67 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_68 = W*in
   wire signed [9:0] m76_68;
   assign m76_68 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_69 = W*in
   wire signed [9:0] m76_69;
   assign m76_69 =10'b0;

   // m76_70 = W*in
   wire signed [9:0] m76_70;
   assign m76_70 ={ {4{in76[5]}} , in76[5:0] };

   // m76_71 = W*in
   wire signed [9:0] m76_71;
   assign m76_71 =10'b0;

   // m76_72 = W*in
   wire signed [9:0] m76_72;
   assign m76_72 =10'b0;

   // m76_73 = W*in
   wire signed [9:0] m76_73;
   assign m76_73 =10'b0;

   // m76_74 = W*in
   wire signed [9:0] m76_74;
   assign m76_74 =10'b0;

   // m76_75 = W*in
   wire signed [9:0] m76_75;
   assign m76_75 =10'b0;

   // m76_76 = W*in
   wire signed [9:0] m76_76;
   assign m76_76 =10'b0;

   // m76_77 = W*in
   wire signed [9:0] m76_77;
   assign m76_77 =10'b0;

   // m76_78 = W*in
   wire signed [9:0] m76_78;
   assign m76_78 =10'b0;

   // m76_79 = W*in
   wire signed [9:0] m76_79;
   assign m76_79 =10'b0;

   // m76_80 = W*in
   wire signed [9:0] m76_80;
   assign m76_80 =10'b0;

   // m76_81 = W*in
   wire signed [9:0] m76_81;
   assign m76_81 =10'b0;

   // m76_82 = W*in
   wire signed [9:0] m76_82;
   assign m76_82 =10'b0;

   // m76_83 = W*in
   wire signed [9:0] m76_83;
   assign m76_83 =10'b0;

   // m76_84 = W*in
   wire signed [9:0] m76_84;
   assign m76_84 =10'b0;

   // m76_85 = W*in
   wire signed [9:0] m76_85;
   assign m76_85 =10'b0;

   // m76_86 = W*in
   wire signed [9:0] m76_86;
   assign m76_86 ={ {4{in76[5]}} , in76[5:0] };

   // m76_87 = W*in
   wire signed [9:0] m76_87;
   assign m76_87 =10'b0;

   // m76_88 = W*in
   wire signed [9:0] m76_88;
   assign m76_88 =10'b0;

   // m76_89 = W*in
   wire signed [9:0] m76_89;
   assign m76_89 =10'b0;

   // m76_90 = W*in
   wire signed [9:0] m76_90;
   assign m76_90 =10'b0;

   // m76_91 = W*in
   wire signed [9:0] m76_91;
   assign m76_91 =10'b0;

   // m76_92 = W*in
   wire signed [9:0] m76_92;
   assign m76_92 =10'b0;

   // m76_93 = W*in
   wire signed [9:0] m76_93;
   assign m76_93 =10'b0;

   // m76_94 = W*in
   wire signed [9:0] m76_94;
   assign m76_94 =10'b0;

   // m76_95 = W*in
   wire signed [9:0] m76_95;
   assign m76_95 =10'b0;

   // m76_96 = W*in
   wire signed [9:0] m76_96;
   assign m76_96 =10'b0;

   // m76_97 = W*in
   wire signed [9:0] m76_97;
   assign m76_97 =10'b0;

   // m76_98 = W*in
   wire signed [9:0] m76_98;
   assign m76_98 =10'b0;

   // m76_99 = W*in
   wire signed [9:0] m76_99;
   assign m76_99 =10'b0;

   // m76_100 = W*in
   wire signed [9:0] m76_100;
   assign m76_100 =10'b0;

   // m76_101 = W*in
   wire signed [9:0] m76_101;
   assign m76_101 =10'b0;

   // m76_102 = W*in
   wire signed [9:0] m76_102;
   assign m76_102 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_103 = W*in
   wire signed [9:0] m76_103;
   assign m76_103 ={ {4{neg76[5]}} , neg76[5:0] };

   // m76_104 = W*in
   wire signed [9:0] m76_104;
   assign m76_104 =10'b0;

   // m76_105 = W*in
   wire signed [9:0] m76_105;
   assign m76_105 =10'b0;

   // m76_106 = W*in
   wire signed [9:0] m76_106;
   assign m76_106 =10'b0;

   // m76_107 = W*in
   wire signed [9:0] m76_107;
   assign m76_107 =10'b0;

   // m76_108 = W*in
   wire signed [9:0] m76_108;
   assign m76_108 ={ {5{in76[5]}} , in76[5:1] };

   // m76_109 = W*in
   wire signed [9:0] m76_109;
   assign m76_109 ={ {4{in76[5]}} , in76[5:0] };

   // m76_110 = W*in
   wire signed [9:0] m76_110;
   assign m76_110 =10'b0;

   // m76_111 = W*in
   wire signed [9:0] m76_111;
   assign m76_111 =10'b0;

   // m76_112 = W*in
   wire signed [9:0] m76_112;
   assign m76_112 ={ {4{in76[5]}} , in76[5:0] };

   // m76_113 = W*in
   wire signed [9:0] m76_113;
   assign m76_113 =10'b0;

   // m76_114 = W*in
   wire signed [9:0] m76_114;
   assign m76_114 =10'b0;

   // m76_115 = W*in
   wire signed [9:0] m76_115;
   assign m76_115 =10'b0;

   // m76_116 = W*in
   wire signed [9:0] m76_116;
   assign m76_116 =10'b0;

   // m76_117 = W*in
   wire signed [9:0] m76_117;
   assign m76_117 =10'b0;

   // m77_1 = W*in
   wire signed [9:0] m77_1;
   assign m77_1 =10'b0;

   // m77_2 = W*in
   wire signed [9:0] m77_2;
   assign m77_2 =10'b0;

   // m77_3 = W*in
   wire signed [9:0] m77_3;
   assign m77_3 =10'b0;

   // m77_4 = W*in
   wire signed [9:0] m77_4;
   assign m77_4 =10'b0;

   // m77_5 = W*in
   wire signed [9:0] m77_5;
   assign m77_5 =10'b0;

   // m77_6 = W*in
   wire signed [9:0] m77_6;
   assign m77_6 =10'b0;

   // m77_7 = W*in
   wire signed [9:0] m77_7;
   assign m77_7 =10'b0;

   // m77_8 = W*in
   wire signed [9:0] m77_8;
   assign m77_8 =10'b0;

   // m77_9 = W*in
   wire signed [9:0] m77_9;
   assign m77_9 =10'b0;

   // m77_10 = W*in
   wire signed [9:0] m77_10;
   assign m77_10 =10'b0;

   // m77_11 = W*in
   wire signed [9:0] m77_11;
   assign m77_11 =10'b0;

   // m77_12 = W*in
   wire signed [9:0] m77_12;
   assign m77_12 =10'b0;

   // m77_13 = W*in
   wire signed [9:0] m77_13;
   assign m77_13 =10'b0;

   // m77_14 = W*in
   wire signed [9:0] m77_14;
   assign m77_14 =10'b0;

   // m77_15 = W*in
   wire signed [9:0] m77_15;
   assign m77_15 =10'b0;

   // m77_16 = W*in
   wire signed [9:0] m77_16;
   assign m77_16 =10'b0;

   // m77_17 = W*in
   wire signed [9:0] m77_17;
   assign m77_17 ={ {5{neg77[5]}} , neg77[5:1] };

   // m77_18 = W*in
   wire signed [9:0] m77_18;
   assign m77_18 ={ {5{neg77[5]}} , neg77[5:1] };

   // m77_19 = W*in
   wire signed [9:0] m77_19;
   assign m77_19 ={ {5{neg77[5]}} , neg77[5:1] };

   // m77_20 = W*in
   wire signed [9:0] m77_20;
   assign m77_20 =10'b0;

   // m77_21 = W*in
   wire signed [9:0] m77_21;
   assign m77_21 ={ {4{in77[5]}} , in77[5:0] };

   // m77_22 = W*in
   wire signed [9:0] m77_22;
   assign m77_22 =10'b0;

   // m77_23 = W*in
   wire signed [9:0] m77_23;
   assign m77_23 ={ {4{in77[5]}} , in77[5:0] };

   // m77_24 = W*in
   wire signed [9:0] m77_24;
   assign m77_24 =10'b0;

   // m77_25 = W*in
   wire signed [9:0] m77_25;
   assign m77_25 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_26 = W*in
   wire signed [9:0] m77_26;
   assign m77_26 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_27 = W*in
   wire signed [9:0] m77_27;
   assign m77_27 ={ {5{neg77[5]}} , neg77[5:1] };

   // m77_28 = W*in
   wire signed [9:0] m77_28;
   assign m77_28 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_29 = W*in
   wire signed [9:0] m77_29;
   assign m77_29 =10'b0;

   // m77_30 = W*in
   wire signed [9:0] m77_30;
   assign m77_30 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_31 = W*in
   wire signed [9:0] m77_31;
   assign m77_31 =10'b0;

   // m77_32 = W*in
   wire signed [9:0] m77_32;
   assign m77_32 =10'b0;

   // m77_33 = W*in
   wire signed [9:0] m77_33;
   assign m77_33 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_34 = W*in
   wire signed [9:0] m77_34;
   assign m77_34 =10'b0;

   // m77_35 = W*in
   wire signed [9:0] m77_35;
   assign m77_35 =10'b0;

   // m77_36 = W*in
   wire signed [9:0] m77_36;
   assign m77_36 =10'b0;

   // m77_37 = W*in
   wire signed [9:0] m77_37;
   assign m77_37 ={ {5{in77[5]}} , in77[5:1] };

   // m77_38 = W*in
   wire signed [9:0] m77_38;
   assign m77_38 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_39 = W*in
   wire signed [9:0] m77_39;
   assign m77_39 =10'b0;

   // m77_40 = W*in
   wire signed [9:0] m77_40;
   assign m77_40 =10'b0;

   // m77_41 = W*in
   wire signed [9:0] m77_41;
   assign m77_41 =10'b0;

   // m77_42 = W*in
   wire signed [9:0] m77_42;
   assign m77_42 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_43 = W*in
   wire signed [9:0] m77_43;
   assign m77_43 =10'b0;

   // m77_44 = W*in
   wire signed [9:0] m77_44;
   assign m77_44 =10'b0;

   // m77_45 = W*in
   wire signed [9:0] m77_45;
   assign m77_45 =10'b0;

   // m77_46 = W*in
   wire signed [9:0] m77_46;
   assign m77_46 =10'b0;

   // m77_47 = W*in
   wire signed [9:0] m77_47;
   assign m77_47 =10'b0;

   // m77_48 = W*in
   wire signed [9:0] m77_48;
   assign m77_48 =10'b0;

   // m77_49 = W*in
   wire signed [9:0] m77_49;
   assign m77_49 =10'b0;

   // m77_50 = W*in
   wire signed [9:0] m77_50;
   assign m77_50 =10'b0;

   // m77_51 = W*in
   wire signed [9:0] m77_51;
   assign m77_51 =10'b0;

   // m77_52 = W*in
   wire signed [9:0] m77_52;
   assign m77_52 =10'b0;

   // m77_53 = W*in
   wire signed [9:0] m77_53;
   assign m77_53 =10'b0;

   // m77_54 = W*in
   wire signed [9:0] m77_54;
   assign m77_54 =10'b0;

   // m77_55 = W*in
   wire signed [9:0] m77_55;
   assign m77_55 =10'b0;

   // m77_56 = W*in
   wire signed [9:0] m77_56;
   assign m77_56 =10'b0;

   // m77_57 = W*in
   wire signed [9:0] m77_57;
   assign m77_57 =10'b0;

   // m77_58 = W*in
   wire signed [9:0] m77_58;
   assign m77_58 =10'b0;

   // m77_59 = W*in
   wire signed [9:0] m77_59;
   assign m77_59 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_60 = W*in
   wire signed [9:0] m77_60;
   assign m77_60 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_61 = W*in
   wire signed [9:0] m77_61;
   assign m77_61 =10'b0;

   // m77_62 = W*in
   wire signed [9:0] m77_62;
   assign m77_62 =10'b0;

   // m77_63 = W*in
   wire signed [9:0] m77_63;
   assign m77_63 =10'b0;

   // m77_64 = W*in
   wire signed [9:0] m77_64;
   assign m77_64 =10'b0;

   // m77_65 = W*in
   wire signed [9:0] m77_65;
   assign m77_65 ={ {4{in77[5]}} , in77[5:0] };

   // m77_66 = W*in
   wire signed [9:0] m77_66;
   assign m77_66 =10'b0;

   // m77_67 = W*in
   wire signed [9:0] m77_67;
   assign m77_67 =10'b0;

   // m77_68 = W*in
   wire signed [9:0] m77_68;
   assign m77_68 =10'b0;

   // m77_69 = W*in
   wire signed [9:0] m77_69;
   assign m77_69 =10'b0;

   // m77_70 = W*in
   wire signed [9:0] m77_70;
   assign m77_70 ={ {5{in77[5]}} , in77[5:1] };

   // m77_71 = W*in
   wire signed [9:0] m77_71;
   assign m77_71 =10'b0;

   // m77_72 = W*in
   wire signed [9:0] m77_72;
   assign m77_72 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_73 = W*in
   wire signed [9:0] m77_73;
   assign m77_73 =10'b0;

   // m77_74 = W*in
   wire signed [9:0] m77_74;
   assign m77_74 =10'b0;

   // m77_75 = W*in
   wire signed [9:0] m77_75;
   assign m77_75 =10'b0;

   // m77_76 = W*in
   wire signed [9:0] m77_76;
   assign m77_76 ={ {4{in77[5]}} , in77[5:0] };

   // m77_77 = W*in
   wire signed [9:0] m77_77;
   assign m77_77 =10'b0;

   // m77_78 = W*in
   wire signed [9:0] m77_78;
   assign m77_78 =10'b0;

   // m77_79 = W*in
   wire signed [9:0] m77_79;
   assign m77_79 =10'b0;

   // m77_80 = W*in
   wire signed [9:0] m77_80;
   assign m77_80 =10'b0;

   // m77_81 = W*in
   wire signed [9:0] m77_81;
   assign m77_81 =10'b0;

   // m77_82 = W*in
   wire signed [9:0] m77_82;
   assign m77_82 ={ {4{in77[5]}} , in77[5:0] };

   // m77_83 = W*in
   wire signed [9:0] m77_83;
   assign m77_83 =10'b0;

   // m77_84 = W*in
   wire signed [9:0] m77_84;
   assign m77_84 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_85 = W*in
   wire signed [9:0] m77_85;
   assign m77_85 ={ {3{in77[5]}} , in77 , {1{1'b0}} };

   // m77_86 = W*in
   wire signed [9:0] m77_86;
   assign m77_86 =10'b0;

   // m77_87 = W*in
   wire signed [9:0] m77_87;
   assign m77_87 =10'b0;

   // m77_88 = W*in
   wire signed [9:0] m77_88;
   assign m77_88 =10'b0;

   // m77_89 = W*in
   wire signed [9:0] m77_89;
   assign m77_89 =10'b0;

   // m77_90 = W*in
   wire signed [9:0] m77_90;
   assign m77_90 =10'b0;

   // m77_91 = W*in
   wire signed [9:0] m77_91;
   assign m77_91 =10'b0;

   // m77_92 = W*in
   wire signed [9:0] m77_92;
   assign m77_92 =10'b0;

   // m77_93 = W*in
   wire signed [9:0] m77_93;
   assign m77_93 ={ {4{in77[5]}} , in77[5:0] };

   // m77_94 = W*in
   wire signed [9:0] m77_94;
   assign m77_94 =10'b0;

   // m77_95 = W*in
   wire signed [9:0] m77_95;
   assign m77_95 =10'b0;

   // m77_96 = W*in
   wire signed [9:0] m77_96;
   assign m77_96 =10'b0;

   // m77_97 = W*in
   wire signed [9:0] m77_97;
   assign m77_97 ={ {4{in77[5]}} , in77[5:0] };

   // m77_98 = W*in
   wire signed [9:0] m77_98;
   assign m77_98 =10'b0;

   // m77_99 = W*in
   wire signed [9:0] m77_99;
   assign m77_99 =10'b0;

   // m77_100 = W*in
   wire signed [9:0] m77_100;
   assign m77_100 ={ {4{in77[5]}} , in77[5:0] };

   // m77_101 = W*in
   wire signed [9:0] m77_101;
   assign m77_101 =10'b0;

   // m77_102 = W*in
   wire signed [9:0] m77_102;
   assign m77_102 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_103 = W*in
   wire signed [9:0] m77_103;
   assign m77_103 =10'b0;

   // m77_104 = W*in
   wire signed [9:0] m77_104;
   assign m77_104 =10'b0;

   // m77_105 = W*in
   wire signed [9:0] m77_105;
   assign m77_105 =10'b0;

   // m77_106 = W*in
   wire signed [9:0] m77_106;
   assign m77_106 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_107 = W*in
   wire signed [9:0] m77_107;
   assign m77_107 =10'b0;

   // m77_108 = W*in
   wire signed [9:0] m77_108;
   assign m77_108 =10'b0;

   // m77_109 = W*in
   wire signed [9:0] m77_109;
   assign m77_109 =10'b0;

   // m77_110 = W*in
   wire signed [9:0] m77_110;
   assign m77_110 =10'b0;

   // m77_111 = W*in
   wire signed [9:0] m77_111;
   assign m77_111 =10'b0;

   // m77_112 = W*in
   wire signed [9:0] m77_112;
   assign m77_112 ={ {4{in77[5]}} , in77[5:0] };

   // m77_113 = W*in
   wire signed [9:0] m77_113;
   assign m77_113 =10'b0;

   // m77_114 = W*in
   wire signed [9:0] m77_114;
   assign m77_114 =10'b0;

   // m77_115 = W*in
   wire signed [9:0] m77_115;
   assign m77_115 =10'b0;

   // m77_116 = W*in
   wire signed [9:0] m77_116;
   assign m77_116 ={ {4{neg77[5]}} , neg77[5:0] };

   // m77_117 = W*in
   wire signed [9:0] m77_117;
   assign m77_117 =10'b0;

   // m78_1 = W*in
   wire signed [9:0] m78_1;
   assign m78_1 =10'b0;

   // m78_2 = W*in
   wire signed [9:0] m78_2;
   assign m78_2 =10'b0;

   // m78_3 = W*in
   wire signed [9:0] m78_3;
   assign m78_3 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_4 = W*in
   wire signed [9:0] m78_4;
   assign m78_4 =10'b0;

   // m78_5 = W*in
   wire signed [9:0] m78_5;
   assign m78_5 =10'b0;

   // m78_6 = W*in
   wire signed [9:0] m78_6;
   assign m78_6 =10'b0;

   // m78_7 = W*in
   wire signed [9:0] m78_7;
   assign m78_7 =10'b0;

   // m78_8 = W*in
   wire signed [9:0] m78_8;
   assign m78_8 =10'b0;

   // m78_9 = W*in
   wire signed [9:0] m78_9;
   assign m78_9 =10'b0;

   // m78_10 = W*in
   wire signed [9:0] m78_10;
   assign m78_10 =10'b0;

   // m78_11 = W*in
   wire signed [9:0] m78_11;
   assign m78_11 =10'b0;

   // m78_12 = W*in
   wire signed [9:0] m78_12;
   assign m78_12 =10'b0;

   // m78_13 = W*in
   wire signed [9:0] m78_13;
   assign m78_13 =10'b0;

   // m78_14 = W*in
   wire signed [9:0] m78_14;
   assign m78_14 =10'b0;

   // m78_15 = W*in
   wire signed [9:0] m78_15;
   assign m78_15 =10'b0;

   // m78_16 = W*in
   wire signed [9:0] m78_16;
   assign m78_16 =10'b0;

   // m78_17 = W*in
   wire signed [9:0] m78_17;
   assign m78_17 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_18 = W*in
   wire signed [9:0] m78_18;
   assign m78_18 =10'b0;

   // m78_19 = W*in
   wire signed [9:0] m78_19;
   assign m78_19 ={ {5{neg78[5]}} , neg78[5:1] };

   // m78_20 = W*in
   wire signed [9:0] m78_20;
   assign m78_20 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_21 = W*in
   wire signed [9:0] m78_21;
   assign m78_21 ={ {4{in78[5]}} , in78[5:0] };

   // m78_22 = W*in
   wire signed [9:0] m78_22;
   assign m78_22 ={ {5{neg78[5]}} , neg78[5:1] };

   // m78_23 = W*in
   wire signed [9:0] m78_23;
   assign m78_23 =10'b0;

   // m78_24 = W*in
   wire signed [9:0] m78_24;
   assign m78_24 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_25 = W*in
   wire signed [9:0] m78_25;
   assign m78_25 =10'b0;

   // m78_26 = W*in
   wire signed [9:0] m78_26;
   assign m78_26 =10'b0;

   // m78_27 = W*in
   wire signed [9:0] m78_27;
   assign m78_27 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_28 = W*in
   wire signed [9:0] m78_28;
   assign m78_28 =10'b0;

   // m78_29 = W*in
   wire signed [9:0] m78_29;
   assign m78_29 ={ {3{in78[5]}} , in78 , {1{1'b0}} };

   // m78_30 = W*in
   wire signed [9:0] m78_30;
   assign m78_30 =10'b0;

   // m78_31 = W*in
   wire signed [9:0] m78_31;
   assign m78_31 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_32 = W*in
   wire signed [9:0] m78_32;
   assign m78_32 =10'b0;

   // m78_33 = W*in
   wire signed [9:0] m78_33;
   assign m78_33 =10'b0;

   // m78_34 = W*in
   wire signed [9:0] m78_34;
   assign m78_34 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_35 = W*in
   wire signed [9:0] m78_35;
   assign m78_35 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_36 = W*in
   wire signed [9:0] m78_36;
   assign m78_36 ={ {5{neg78[5]}} , neg78[5:1] };

   // m78_37 = W*in
   wire signed [9:0] m78_37;
   assign m78_37 =10'b0;

   // m78_38 = W*in
   wire signed [9:0] m78_38;
   assign m78_38 =10'b0;

   // m78_39 = W*in
   wire signed [9:0] m78_39;
   assign m78_39 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_40 = W*in
   wire signed [9:0] m78_40;
   assign m78_40 =10'b0;

   // m78_41 = W*in
   wire signed [9:0] m78_41;
   assign m78_41 =10'b0;

   // m78_42 = W*in
   wire signed [9:0] m78_42;
   assign m78_42 =10'b0;

   // m78_43 = W*in
   wire signed [9:0] m78_43;
   assign m78_43 =10'b0;

   // m78_44 = W*in
   wire signed [9:0] m78_44;
   assign m78_44 =10'b0;

   // m78_45 = W*in
   wire signed [9:0] m78_45;
   assign m78_45 =10'b0;

   // m78_46 = W*in
   wire signed [9:0] m78_46;
   assign m78_46 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_47 = W*in
   wire signed [9:0] m78_47;
   assign m78_47 =10'b0;

   // m78_48 = W*in
   wire signed [9:0] m78_48;
   assign m78_48 =10'b0;

   // m78_49 = W*in
   wire signed [9:0] m78_49;
   assign m78_49 =10'b0;

   // m78_50 = W*in
   wire signed [9:0] m78_50;
   assign m78_50 =10'b0;

   // m78_51 = W*in
   wire signed [9:0] m78_51;
   assign m78_51 =10'b0;

   // m78_52 = W*in
   wire signed [9:0] m78_52;
   assign m78_52 =10'b0;

   // m78_53 = W*in
   wire signed [9:0] m78_53;
   assign m78_53 =10'b0;

   // m78_54 = W*in
   wire signed [9:0] m78_54;
   assign m78_54 =10'b0;

   // m78_55 = W*in
   wire signed [9:0] m78_55;
   assign m78_55 =10'b0;

   // m78_56 = W*in
   wire signed [9:0] m78_56;
   assign m78_56 =10'b0;

   // m78_57 = W*in
   wire signed [9:0] m78_57;
   assign m78_57 =10'b0;

   // m78_58 = W*in
   wire signed [9:0] m78_58;
   assign m78_58 ={ {5{neg78[5]}} , neg78[5:1] };

   // m78_59 = W*in
   wire signed [9:0] m78_59;
   assign m78_59 =10'b0;

   // m78_60 = W*in
   wire signed [9:0] m78_60;
   assign m78_60 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_61 = W*in
   wire signed [9:0] m78_61;
   assign m78_61 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_62 = W*in
   wire signed [9:0] m78_62;
   assign m78_62 =10'b0;

   // m78_63 = W*in
   wire signed [9:0] m78_63;
   assign m78_63 ={ {4{in78[5]}} , in78[5:0] };

   // m78_64 = W*in
   wire signed [9:0] m78_64;
   assign m78_64 =10'b0;

   // m78_65 = W*in
   wire signed [9:0] m78_65;
   assign m78_65 ={ {4{in78[5]}} , in78[5:0] };

   // m78_66 = W*in
   wire signed [9:0] m78_66;
   assign m78_66 =10'b0;

   // m78_67 = W*in
   wire signed [9:0] m78_67;
   assign m78_67 =10'b0;

   // m78_68 = W*in
   wire signed [9:0] m78_68;
   assign m78_68 =10'b0;

   // m78_69 = W*in
   wire signed [9:0] m78_69;
   assign m78_69 ={ {4{in78[5]}} , in78[5:0] };

   // m78_70 = W*in
   wire signed [9:0] m78_70;
   assign m78_70 ={ {4{in78[5]}} , in78[5:0] };

   // m78_71 = W*in
   wire signed [9:0] m78_71;
   assign m78_71 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_72 = W*in
   wire signed [9:0] m78_72;
   assign m78_72 =10'b0;

   // m78_73 = W*in
   wire signed [9:0] m78_73;
   assign m78_73 ={ {5{neg78[5]}} , neg78[5:1] };

   // m78_74 = W*in
   wire signed [9:0] m78_74;
   assign m78_74 =10'b0;

   // m78_75 = W*in
   wire signed [9:0] m78_75;
   assign m78_75 =10'b0;

   // m78_76 = W*in
   wire signed [9:0] m78_76;
   assign m78_76 =10'b0;

   // m78_77 = W*in
   wire signed [9:0] m78_77;
   assign m78_77 ={ {4{in78[5]}} , in78[5:0] };

   // m78_78 = W*in
   wire signed [9:0] m78_78;
   assign m78_78 =10'b0;

   // m78_79 = W*in
   wire signed [9:0] m78_79;
   assign m78_79 ={ {4{in78[5]}} , in78[5:0] };

   // m78_80 = W*in
   wire signed [9:0] m78_80;
   assign m78_80 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_81 = W*in
   wire signed [9:0] m78_81;
   assign m78_81 =10'b0;

   // m78_82 = W*in
   wire signed [9:0] m78_82;
   assign m78_82 =10'b0;

   // m78_83 = W*in
   wire signed [9:0] m78_83;
   assign m78_83 =10'b0;

   // m78_84 = W*in
   wire signed [9:0] m78_84;
   assign m78_84 =10'b0;

   // m78_85 = W*in
   wire signed [9:0] m78_85;
   assign m78_85 ={ {4{in78[5]}} , in78[5:0] };

   // m78_86 = W*in
   wire signed [9:0] m78_86;
   assign m78_86 ={ {4{in78[5]}} , in78[5:0] };

   // m78_87 = W*in
   wire signed [9:0] m78_87;
   assign m78_87 =10'b0;

   // m78_88 = W*in
   wire signed [9:0] m78_88;
   assign m78_88 =10'b0;

   // m78_89 = W*in
   wire signed [9:0] m78_89;
   assign m78_89 =10'b0;

   // m78_90 = W*in
   wire signed [9:0] m78_90;
   assign m78_90 =10'b0;

   // m78_91 = W*in
   wire signed [9:0] m78_91;
   assign m78_91 ={ {4{in78[5]}} , in78[5:0] };

   // m78_92 = W*in
   wire signed [9:0] m78_92;
   assign m78_92 =10'b0;

   // m78_93 = W*in
   wire signed [9:0] m78_93;
   assign m78_93 ={ {4{in78[5]}} , in78[5:0] };

   // m78_94 = W*in
   wire signed [9:0] m78_94;
   assign m78_94 ={ {4{in78[5]}} , in78[5:0] };

   // m78_95 = W*in
   wire signed [9:0] m78_95;
   assign m78_95 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_96 = W*in
   wire signed [9:0] m78_96;
   assign m78_96 =10'b0;

   // m78_97 = W*in
   wire signed [9:0] m78_97;
   assign m78_97 =10'b0;

   // m78_98 = W*in
   wire signed [9:0] m78_98;
   assign m78_98 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_99 = W*in
   wire signed [9:0] m78_99;
   assign m78_99 =10'b0;

   // m78_100 = W*in
   wire signed [9:0] m78_100;
   assign m78_100 =10'b0;

   // m78_101 = W*in
   wire signed [9:0] m78_101;
   assign m78_101 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_102 = W*in
   wire signed [9:0] m78_102;
   assign m78_102 =10'b0;

   // m78_103 = W*in
   wire signed [9:0] m78_103;
   assign m78_103 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_104 = W*in
   wire signed [9:0] m78_104;
   assign m78_104 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_105 = W*in
   wire signed [9:0] m78_105;
   assign m78_105 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_106 = W*in
   wire signed [9:0] m78_106;
   assign m78_106 =10'b0;

   // m78_107 = W*in
   wire signed [9:0] m78_107;
   assign m78_107 ={ {4{neg78[5]}} , neg78[5:0] };

   // m78_108 = W*in
   wire signed [9:0] m78_108;
   assign m78_108 =10'b0;

   // m78_109 = W*in
   wire signed [9:0] m78_109;
   assign m78_109 =10'b0;

   // m78_110 = W*in
   wire signed [9:0] m78_110;
   assign m78_110 =10'b0;

   // m78_111 = W*in
   wire signed [9:0] m78_111;
   assign m78_111 =10'b0;

   // m78_112 = W*in
   wire signed [9:0] m78_112;
   assign m78_112 =10'b0;

   // m78_113 = W*in
   wire signed [9:0] m78_113;
   assign m78_113 =10'b0;

   // m78_114 = W*in
   wire signed [9:0] m78_114;
   assign m78_114 =10'b0;

   // m78_115 = W*in
   wire signed [9:0] m78_115;
   assign m78_115 =10'b0;

   // m78_116 = W*in
   wire signed [9:0] m78_116;
   assign m78_116 ={ {4{in78[5]}} , in78[5:0] };

   // m78_117 = W*in
   wire signed [9:0] m78_117;
   assign m78_117 ={ {4{neg78[5]}} , neg78[5:0] };

   // m79_1 = W*in
   wire signed [9:0] m79_1;
   assign m79_1 =10'b0;

   // m79_2 = W*in
   wire signed [9:0] m79_2;
   assign m79_2 =10'b0;

   // m79_3 = W*in
   wire signed [9:0] m79_3;
   assign m79_3 =10'b0;

   // m79_4 = W*in
   wire signed [9:0] m79_4;
   assign m79_4 =10'b0;

   // m79_5 = W*in
   wire signed [9:0] m79_5;
   assign m79_5 =10'b0;

   // m79_6 = W*in
   wire signed [9:0] m79_6;
   assign m79_6 =10'b0;

   // m79_7 = W*in
   wire signed [9:0] m79_7;
   assign m79_7 ={ {4{in79[5]}} , in79[5:0] };

   // m79_8 = W*in
   wire signed [9:0] m79_8;
   assign m79_8 =10'b0;

   // m79_9 = W*in
   wire signed [9:0] m79_9;
   assign m79_9 =10'b0;

   // m79_10 = W*in
   wire signed [9:0] m79_10;
   assign m79_10 =10'b0;

   // m79_11 = W*in
   wire signed [9:0] m79_11;
   assign m79_11 =10'b0;

   // m79_12 = W*in
   wire signed [9:0] m79_12;
   assign m79_12 =10'b0;

   // m79_13 = W*in
   wire signed [9:0] m79_13;
   assign m79_13 ={ {4{in79[5]}} , in79[5:0] };

   // m79_14 = W*in
   wire signed [9:0] m79_14;
   assign m79_14 =10'b0;

   // m79_15 = W*in
   wire signed [9:0] m79_15;
   assign m79_15 =10'b0;

   // m79_16 = W*in
   wire signed [9:0] m79_16;
   assign m79_16 =10'b0;

   // m79_17 = W*in
   wire signed [9:0] m79_17;
   assign m79_17 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_18 = W*in
   wire signed [9:0] m79_18;
   assign m79_18 =10'b0;

   // m79_19 = W*in
   wire signed [9:0] m79_19;
   assign m79_19 ={ {5{in79[5]}} , in79[5:1] };

   // m79_20 = W*in
   wire signed [9:0] m79_20;
   assign m79_20 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_21 = W*in
   wire signed [9:0] m79_21;
   assign m79_21 ={ {5{in79[5]}} , in79[5:1] };

   // m79_22 = W*in
   wire signed [9:0] m79_22;
   assign m79_22 =10'b0;

   // m79_23 = W*in
   wire signed [9:0] m79_23;
   assign m79_23 =10'b0;

   // m79_24 = W*in
   wire signed [9:0] m79_24;
   assign m79_24 =10'b0;

   // m79_25 = W*in
   wire signed [9:0] m79_25;
   assign m79_25 =10'b0;

   // m79_26 = W*in
   wire signed [9:0] m79_26;
   assign m79_26 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_27 = W*in
   wire signed [9:0] m79_27;
   assign m79_27 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_28 = W*in
   wire signed [9:0] m79_28;
   assign m79_28 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_29 = W*in
   wire signed [9:0] m79_29;
   assign m79_29 ={ {4{in79[5]}} , in79[5:0] };

   // m79_30 = W*in
   wire signed [9:0] m79_30;
   assign m79_30 =10'b0;

   // m79_31 = W*in
   wire signed [9:0] m79_31;
   assign m79_31 =10'b0;

   // m79_32 = W*in
   wire signed [9:0] m79_32;
   assign m79_32 =10'b0;

   // m79_33 = W*in
   wire signed [9:0] m79_33;
   assign m79_33 =10'b0;

   // m79_34 = W*in
   wire signed [9:0] m79_34;
   assign m79_34 =10'b0;

   // m79_35 = W*in
   wire signed [9:0] m79_35;
   assign m79_35 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_36 = W*in
   wire signed [9:0] m79_36;
   assign m79_36 =10'b0;

   // m79_37 = W*in
   wire signed [9:0] m79_37;
   assign m79_37 =10'b0;

   // m79_38 = W*in
   wire signed [9:0] m79_38;
   assign m79_38 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_39 = W*in
   wire signed [9:0] m79_39;
   assign m79_39 =10'b0;

   // m79_40 = W*in
   wire signed [9:0] m79_40;
   assign m79_40 =10'b0;

   // m79_41 = W*in
   wire signed [9:0] m79_41;
   assign m79_41 ={ {4{in79[5]}} , in79[5:0] };

   // m79_42 = W*in
   wire signed [9:0] m79_42;
   assign m79_42 =10'b0;

   // m79_43 = W*in
   wire signed [9:0] m79_43;
   assign m79_43 =10'b0;

   // m79_44 = W*in
   wire signed [9:0] m79_44;
   assign m79_44 =10'b0;

   // m79_45 = W*in
   wire signed [9:0] m79_45;
   assign m79_45 ={ {4{in79[5]}} , in79[5:0] };

   // m79_46 = W*in
   wire signed [9:0] m79_46;
   assign m79_46 =10'b0;

   // m79_47 = W*in
   wire signed [9:0] m79_47;
   assign m79_47 =10'b0;

   // m79_48 = W*in
   wire signed [9:0] m79_48;
   assign m79_48 =10'b0;

   // m79_49 = W*in
   wire signed [9:0] m79_49;
   assign m79_49 =10'b0;

   // m79_50 = W*in
   wire signed [9:0] m79_50;
   assign m79_50 =10'b0;

   // m79_51 = W*in
   wire signed [9:0] m79_51;
   assign m79_51 =10'b0;

   // m79_52 = W*in
   wire signed [9:0] m79_52;
   assign m79_52 =10'b0;

   // m79_53 = W*in
   wire signed [9:0] m79_53;
   assign m79_53 =10'b0;

   // m79_54 = W*in
   wire signed [9:0] m79_54;
   assign m79_54 =10'b0;

   // m79_55 = W*in
   wire signed [9:0] m79_55;
   assign m79_55 =10'b0;

   // m79_56 = W*in
   wire signed [9:0] m79_56;
   assign m79_56 =10'b0;

   // m79_57 = W*in
   wire signed [9:0] m79_57;
   assign m79_57 =10'b0;

   // m79_58 = W*in
   wire signed [9:0] m79_58;
   assign m79_58 =10'b0;

   // m79_59 = W*in
   wire signed [9:0] m79_59;
   assign m79_59 =10'b0;

   // m79_60 = W*in
   wire signed [9:0] m79_60;
   assign m79_60 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_61 = W*in
   wire signed [9:0] m79_61;
   assign m79_61 =10'b0;

   // m79_62 = W*in
   wire signed [9:0] m79_62;
   assign m79_62 =10'b0;

   // m79_63 = W*in
   wire signed [9:0] m79_63;
   assign m79_63 ={ {4{in79[5]}} , in79[5:0] };

   // m79_64 = W*in
   wire signed [9:0] m79_64;
   assign m79_64 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_65 = W*in
   wire signed [9:0] m79_65;
   assign m79_65 ={ {4{in79[5]}} , in79[5:0] };

   // m79_66 = W*in
   wire signed [9:0] m79_66;
   assign m79_66 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_67 = W*in
   wire signed [9:0] m79_67;
   assign m79_67 =10'b0;

   // m79_68 = W*in
   wire signed [9:0] m79_68;
   assign m79_68 =10'b0;

   // m79_69 = W*in
   wire signed [9:0] m79_69;
   assign m79_69 =10'b0;

   // m79_70 = W*in
   wire signed [9:0] m79_70;
   assign m79_70 =10'b0;

   // m79_71 = W*in
   wire signed [9:0] m79_71;
   assign m79_71 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_72 = W*in
   wire signed [9:0] m79_72;
   assign m79_72 =10'b0;

   // m79_73 = W*in
   wire signed [9:0] m79_73;
   assign m79_73 ={ {5{in79[5]}} , in79[5:1] };

   // m79_74 = W*in
   wire signed [9:0] m79_74;
   assign m79_74 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_75 = W*in
   wire signed [9:0] m79_75;
   assign m79_75 =10'b0;

   // m79_76 = W*in
   wire signed [9:0] m79_76;
   assign m79_76 =10'b0;

   // m79_77 = W*in
   wire signed [9:0] m79_77;
   assign m79_77 =10'b0;

   // m79_78 = W*in
   wire signed [9:0] m79_78;
   assign m79_78 =10'b0;

   // m79_79 = W*in
   wire signed [9:0] m79_79;
   assign m79_79 ={ {4{in79[5]}} , in79[5:0] };

   // m79_80 = W*in
   wire signed [9:0] m79_80;
   assign m79_80 =10'b0;

   // m79_81 = W*in
   wire signed [9:0] m79_81;
   assign m79_81 ={ {5{neg79[5]}} , neg79[5:1] };

   // m79_82 = W*in
   wire signed [9:0] m79_82;
   assign m79_82 =10'b0;

   // m79_83 = W*in
   wire signed [9:0] m79_83;
   assign m79_83 =10'b0;

   // m79_84 = W*in
   wire signed [9:0] m79_84;
   assign m79_84 =10'b0;

   // m79_85 = W*in
   wire signed [9:0] m79_85;
   assign m79_85 ={ {4{in79[5]}} , in79[5:0] };

   // m79_86 = W*in
   wire signed [9:0] m79_86;
   assign m79_86 ={ {4{in79[5]}} , in79[5:0] };

   // m79_87 = W*in
   wire signed [9:0] m79_87;
   assign m79_87 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_88 = W*in
   wire signed [9:0] m79_88;
   assign m79_88 =10'b0;

   // m79_89 = W*in
   wire signed [9:0] m79_89;
   assign m79_89 =10'b0;

   // m79_90 = W*in
   wire signed [9:0] m79_90;
   assign m79_90 =10'b0;

   // m79_91 = W*in
   wire signed [9:0] m79_91;
   assign m79_91 =10'b0;

   // m79_92 = W*in
   wire signed [9:0] m79_92;
   assign m79_92 =10'b0;

   // m79_93 = W*in
   wire signed [9:0] m79_93;
   assign m79_93 ={ {4{in79[5]}} , in79[5:0] };

   // m79_94 = W*in
   wire signed [9:0] m79_94;
   assign m79_94 =10'b0;

   // m79_95 = W*in
   wire signed [9:0] m79_95;
   assign m79_95 =10'b0;

   // m79_96 = W*in
   wire signed [9:0] m79_96;
   assign m79_96 =10'b0;

   // m79_97 = W*in
   wire signed [9:0] m79_97;
   assign m79_97 =10'b0;

   // m79_98 = W*in
   wire signed [9:0] m79_98;
   assign m79_98 =10'b0;

   // m79_99 = W*in
   wire signed [9:0] m79_99;
   assign m79_99 =10'b0;

   // m79_100 = W*in
   wire signed [9:0] m79_100;
   assign m79_100 =10'b0;

   // m79_101 = W*in
   wire signed [9:0] m79_101;
   assign m79_101 =10'b0;

   // m79_102 = W*in
   wire signed [9:0] m79_102;
   assign m79_102 =10'b0;

   // m79_103 = W*in
   wire signed [9:0] m79_103;
   assign m79_103 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_104 = W*in
   wire signed [9:0] m79_104;
   assign m79_104 ={ {4{neg79[5]}} , neg79[5:0] };

   // m79_105 = W*in
   wire signed [9:0] m79_105;
   assign m79_105 =10'b0;

   // m79_106 = W*in
   wire signed [9:0] m79_106;
   assign m79_106 =10'b0;

   // m79_107 = W*in
   wire signed [9:0] m79_107;
   assign m79_107 =10'b0;

   // m79_108 = W*in
   wire signed [9:0] m79_108;
   assign m79_108 ={ {4{in79[5]}} , in79[5:0] };

   // m79_109 = W*in
   wire signed [9:0] m79_109;
   assign m79_109 ={ {4{in79[5]}} , in79[5:0] };

   // m79_110 = W*in
   wire signed [9:0] m79_110;
   assign m79_110 =10'b0;

   // m79_111 = W*in
   wire signed [9:0] m79_111;
   assign m79_111 =10'b0;

   // m79_112 = W*in
   wire signed [9:0] m79_112;
   assign m79_112 =10'b0;

   // m79_113 = W*in
   wire signed [9:0] m79_113;
   assign m79_113 =10'b0;

   // m79_114 = W*in
   wire signed [9:0] m79_114;
   assign m79_114 =10'b0;

   // m79_115 = W*in
   wire signed [9:0] m79_115;
   assign m79_115 =10'b0;

   // m79_116 = W*in
   wire signed [9:0] m79_116;
   assign m79_116 ={ {4{in79[5]}} , in79[5:0] };

   // m79_117 = W*in
   wire signed [9:0] m79_117;
   assign m79_117 ={ {4{neg79[5]}} , neg79[5:0] };

   // m80_1 = W*in
   wire signed [9:0] m80_1;
   assign m80_1 =10'b0;

   // m80_2 = W*in
   wire signed [9:0] m80_2;
   assign m80_2 =10'b0;

   // m80_3 = W*in
   wire signed [9:0] m80_3;
   assign m80_3 =10'b0;

   // m80_4 = W*in
   wire signed [9:0] m80_4;
   assign m80_4 =10'b0;

   // m80_5 = W*in
   wire signed [9:0] m80_5;
   assign m80_5 =10'b0;

   // m80_6 = W*in
   wire signed [9:0] m80_6;
   assign m80_6 =10'b0;

   // m80_7 = W*in
   wire signed [9:0] m80_7;
   assign m80_7 =10'b0;

   // m80_8 = W*in
   wire signed [9:0] m80_8;
   assign m80_8 =10'b0;

   // m80_9 = W*in
   wire signed [9:0] m80_9;
   assign m80_9 =10'b0;

   // m80_10 = W*in
   wire signed [9:0] m80_10;
   assign m80_10 =10'b0;

   // m80_11 = W*in
   wire signed [9:0] m80_11;
   assign m80_11 =10'b0;

   // m80_12 = W*in
   wire signed [9:0] m80_12;
   assign m80_12 =10'b0;

   // m80_13 = W*in
   wire signed [9:0] m80_13;
   assign m80_13 =10'b0;

   // m80_14 = W*in
   wire signed [9:0] m80_14;
   assign m80_14 =10'b0;

   // m80_15 = W*in
   wire signed [9:0] m80_15;
   assign m80_15 =10'b0;

   // m80_16 = W*in
   wire signed [9:0] m80_16;
   assign m80_16 =10'b0;

   // m80_17 = W*in
   wire signed [9:0] m80_17;
   assign m80_17 =10'b0;

   // m80_18 = W*in
   wire signed [9:0] m80_18;
   assign m80_18 =10'b0;

   // m80_19 = W*in
   wire signed [9:0] m80_19;
   assign m80_19 ={ {4{neg80[5]}} , neg80[5:0] };

   // m80_20 = W*in
   wire signed [9:0] m80_20;
   assign m80_20 =10'b0;

   // m80_21 = W*in
   wire signed [9:0] m80_21;
   assign m80_21 =10'b0;

   // m80_22 = W*in
   wire signed [9:0] m80_22;
   assign m80_22 =10'b0;

   // m80_23 = W*in
   wire signed [9:0] m80_23;
   assign m80_23 =10'b0;

   // m80_24 = W*in
   wire signed [9:0] m80_24;
   assign m80_24 =10'b0;

   // m80_25 = W*in
   wire signed [9:0] m80_25;
   assign m80_25 =10'b0;

   // m80_26 = W*in
   wire signed [9:0] m80_26;
   assign m80_26 =10'b0;

   // m80_27 = W*in
   wire signed [9:0] m80_27;
   assign m80_27 =10'b0;

   // m80_28 = W*in
   wire signed [9:0] m80_28;
   assign m80_28 ={ {5{in80[5]}} , in80[5:1] };

   // m80_29 = W*in
   wire signed [9:0] m80_29;
   assign m80_29 ={ {4{neg80[5]}} , neg80[5:0] };

   // m80_30 = W*in
   wire signed [9:0] m80_30;
   assign m80_30 =10'b0;

   // m80_31 = W*in
   wire signed [9:0] m80_31;
   assign m80_31 =10'b0;

   // m80_32 = W*in
   wire signed [9:0] m80_32;
   assign m80_32 =10'b0;

   // m80_33 = W*in
   wire signed [9:0] m80_33;
   assign m80_33 =10'b0;

   // m80_34 = W*in
   wire signed [9:0] m80_34;
   assign m80_34 =10'b0;

   // m80_35 = W*in
   wire signed [9:0] m80_35;
   assign m80_35 =10'b0;

   // m80_36 = W*in
   wire signed [9:0] m80_36;
   assign m80_36 =10'b0;

   // m80_37 = W*in
   wire signed [9:0] m80_37;
   assign m80_37 =10'b0;

   // m80_38 = W*in
   wire signed [9:0] m80_38;
   assign m80_38 =10'b0;

   // m80_39 = W*in
   wire signed [9:0] m80_39;
   assign m80_39 =10'b0;

   // m80_40 = W*in
   wire signed [9:0] m80_40;
   assign m80_40 =10'b0;

   // m80_41 = W*in
   wire signed [9:0] m80_41;
   assign m80_41 =10'b0;

   // m80_42 = W*in
   wire signed [9:0] m80_42;
   assign m80_42 =10'b0;

   // m80_43 = W*in
   wire signed [9:0] m80_43;
   assign m80_43 =10'b0;

   // m80_44 = W*in
   wire signed [9:0] m80_44;
   assign m80_44 =10'b0;

   // m80_45 = W*in
   wire signed [9:0] m80_45;
   assign m80_45 =10'b0;

   // m80_46 = W*in
   wire signed [9:0] m80_46;
   assign m80_46 =10'b0;

   // m80_47 = W*in
   wire signed [9:0] m80_47;
   assign m80_47 =10'b0;

   // m80_48 = W*in
   wire signed [9:0] m80_48;
   assign m80_48 =10'b0;

   // m80_49 = W*in
   wire signed [9:0] m80_49;
   assign m80_49 =10'b0;

   // m80_50 = W*in
   wire signed [9:0] m80_50;
   assign m80_50 =10'b0;

   // m80_51 = W*in
   wire signed [9:0] m80_51;
   assign m80_51 =10'b0;

   // m80_52 = W*in
   wire signed [9:0] m80_52;
   assign m80_52 =10'b0;

   // m80_53 = W*in
   wire signed [9:0] m80_53;
   assign m80_53 =10'b0;

   // m80_54 = W*in
   wire signed [9:0] m80_54;
   assign m80_54 =10'b0;

   // m80_55 = W*in
   wire signed [9:0] m80_55;
   assign m80_55 =10'b0;

   // m80_56 = W*in
   wire signed [9:0] m80_56;
   assign m80_56 =10'b0;

   // m80_57 = W*in
   wire signed [9:0] m80_57;
   assign m80_57 =10'b0;

   // m80_58 = W*in
   wire signed [9:0] m80_58;
   assign m80_58 =10'b0;

   // m80_59 = W*in
   wire signed [9:0] m80_59;
   assign m80_59 =10'b0;

   // m80_60 = W*in
   wire signed [9:0] m80_60;
   assign m80_60 =10'b0;

   // m80_61 = W*in
   wire signed [9:0] m80_61;
   assign m80_61 =10'b0;

   // m80_62 = W*in
   wire signed [9:0] m80_62;
   assign m80_62 =10'b0;

   // m80_63 = W*in
   wire signed [9:0] m80_63;
   assign m80_63 =10'b0;

   // m80_64 = W*in
   wire signed [9:0] m80_64;
   assign m80_64 =10'b0;

   // m80_65 = W*in
   wire signed [9:0] m80_65;
   assign m80_65 =10'b0;

   // m80_66 = W*in
   wire signed [9:0] m80_66;
   assign m80_66 =10'b0;

   // m80_67 = W*in
   wire signed [9:0] m80_67;
   assign m80_67 ={ {4{neg80[5]}} , neg80[5:0] };

   // m80_68 = W*in
   wire signed [9:0] m80_68;
   assign m80_68 =10'b0;

   // m80_69 = W*in
   wire signed [9:0] m80_69;
   assign m80_69 ={ {5{neg80[5]}} , neg80[5:1] };

   // m80_70 = W*in
   wire signed [9:0] m80_70;
   assign m80_70 =10'b0;

   // m80_71 = W*in
   wire signed [9:0] m80_71;
   assign m80_71 =10'b0;

   // m80_72 = W*in
   wire signed [9:0] m80_72;
   assign m80_72 ={ {5{in80[5]}} , in80[5:1] };

   // m80_73 = W*in
   wire signed [9:0] m80_73;
   assign m80_73 =10'b0;

   // m80_74 = W*in
   wire signed [9:0] m80_74;
   assign m80_74 =10'b0;

   // m80_75 = W*in
   wire signed [9:0] m80_75;
   assign m80_75 =10'b0;

   // m80_76 = W*in
   wire signed [9:0] m80_76;
   assign m80_76 =10'b0;

   // m80_77 = W*in
   wire signed [9:0] m80_77;
   assign m80_77 =10'b0;

   // m80_78 = W*in
   wire signed [9:0] m80_78;
   assign m80_78 =10'b0;

   // m80_79 = W*in
   wire signed [9:0] m80_79;
   assign m80_79 =10'b0;

   // m80_80 = W*in
   wire signed [9:0] m80_80;
   assign m80_80 =10'b0;

   // m80_81 = W*in
   wire signed [9:0] m80_81;
   assign m80_81 =10'b0;

   // m80_82 = W*in
   wire signed [9:0] m80_82;
   assign m80_82 =10'b0;

   // m80_83 = W*in
   wire signed [9:0] m80_83;
   assign m80_83 =10'b0;

   // m80_84 = W*in
   wire signed [9:0] m80_84;
   assign m80_84 =10'b0;

   // m80_85 = W*in
   wire signed [9:0] m80_85;
   assign m80_85 =10'b0;

   // m80_86 = W*in
   wire signed [9:0] m80_86;
   assign m80_86 =10'b0;

   // m80_87 = W*in
   wire signed [9:0] m80_87;
   assign m80_87 =10'b0;

   // m80_88 = W*in
   wire signed [9:0] m80_88;
   assign m80_88 =10'b0;

   // m80_89 = W*in
   wire signed [9:0] m80_89;
   assign m80_89 =10'b0;

   // m80_90 = W*in
   wire signed [9:0] m80_90;
   assign m80_90 =10'b0;

   // m80_91 = W*in
   wire signed [9:0] m80_91;
   assign m80_91 =10'b0;

   // m80_92 = W*in
   wire signed [9:0] m80_92;
   assign m80_92 =10'b0;

   // m80_93 = W*in
   wire signed [9:0] m80_93;
   assign m80_93 =10'b0;

   // m80_94 = W*in
   wire signed [9:0] m80_94;
   assign m80_94 =10'b0;

   // m80_95 = W*in
   wire signed [9:0] m80_95;
   assign m80_95 =10'b0;

   // m80_96 = W*in
   wire signed [9:0] m80_96;
   assign m80_96 =10'b0;

   // m80_97 = W*in
   wire signed [9:0] m80_97;
   assign m80_97 =10'b0;

   // m80_98 = W*in
   wire signed [9:0] m80_98;
   assign m80_98 =10'b0;

   // m80_99 = W*in
   wire signed [9:0] m80_99;
   assign m80_99 =10'b0;

   // m80_100 = W*in
   wire signed [9:0] m80_100;
   assign m80_100 =10'b0;

   // m80_101 = W*in
   wire signed [9:0] m80_101;
   assign m80_101 =10'b0;

   // m80_102 = W*in
   wire signed [9:0] m80_102;
   assign m80_102 =10'b0;

   // m80_103 = W*in
   wire signed [9:0] m80_103;
   assign m80_103 =10'b0;

   // m80_104 = W*in
   wire signed [9:0] m80_104;
   assign m80_104 =10'b0;

   // m80_105 = W*in
   wire signed [9:0] m80_105;
   assign m80_105 =10'b0;

   // m80_106 = W*in
   wire signed [9:0] m80_106;
   assign m80_106 =10'b0;

   // m80_107 = W*in
   wire signed [9:0] m80_107;
   assign m80_107 =10'b0;

   // m80_108 = W*in
   wire signed [9:0] m80_108;
   assign m80_108 =10'b0;

   // m80_109 = W*in
   wire signed [9:0] m80_109;
   assign m80_109 =10'b0;

   // m80_110 = W*in
   wire signed [9:0] m80_110;
   assign m80_110 =10'b0;

   // m80_111 = W*in
   wire signed [9:0] m80_111;
   assign m80_111 =10'b0;

   // m80_112 = W*in
   wire signed [9:0] m80_112;
   assign m80_112 =10'b0;

   // m80_113 = W*in
   wire signed [9:0] m80_113;
   assign m80_113 =10'b0;

   // m80_114 = W*in
   wire signed [9:0] m80_114;
   assign m80_114 =10'b0;

   // m80_115 = W*in
   wire signed [9:0] m80_115;
   assign m80_115 =10'b0;

   // m80_116 = W*in
   wire signed [9:0] m80_116;
   assign m80_116 =10'b0;

   // m80_117 = W*in
   wire signed [9:0] m80_117;
   assign m80_117 =10'b0;

   // m81_1 = W*in
   wire signed [9:0] m81_1;
   assign m81_1 =10'b0;

   // m81_2 = W*in
   wire signed [9:0] m81_2;
   assign m81_2 =10'b0;

   // m81_3 = W*in
   wire signed [9:0] m81_3;
   assign m81_3 =10'b0;

   // m81_4 = W*in
   wire signed [9:0] m81_4;
   assign m81_4 =10'b0;

   // m81_5 = W*in
   wire signed [9:0] m81_5;
   assign m81_5 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_6 = W*in
   wire signed [9:0] m81_6;
   assign m81_6 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_7 = W*in
   wire signed [9:0] m81_7;
   assign m81_7 ={ {4{in81[5]}} , in81[5:0] };

   // m81_8 = W*in
   wire signed [9:0] m81_8;
   assign m81_8 =10'b0;

   // m81_9 = W*in
   wire signed [9:0] m81_9;
   assign m81_9 =10'b0;

   // m81_10 = W*in
   wire signed [9:0] m81_10;
   assign m81_10 =10'b0;

   // m81_11 = W*in
   wire signed [9:0] m81_11;
   assign m81_11 =10'b0;

   // m81_12 = W*in
   wire signed [9:0] m81_12;
   assign m81_12 =10'b0;

   // m81_13 = W*in
   wire signed [9:0] m81_13;
   assign m81_13 =10'b0;

   // m81_14 = W*in
   wire signed [9:0] m81_14;
   assign m81_14 =10'b0;

   // m81_15 = W*in
   wire signed [9:0] m81_15;
   assign m81_15 =10'b0;

   // m81_16 = W*in
   wire signed [9:0] m81_16;
   assign m81_16 =10'b0;

   // m81_17 = W*in
   wire signed [9:0] m81_17;
   assign m81_17 =10'b0;

   // m81_18 = W*in
   wire signed [9:0] m81_18;
   assign m81_18 =10'b0;

   // m81_19 = W*in
   wire signed [9:0] m81_19;
   assign m81_19 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_20 = W*in
   wire signed [9:0] m81_20;
   assign m81_20 =10'b0;

   // m81_21 = W*in
   wire signed [9:0] m81_21;
   assign m81_21 =10'b0;

   // m81_22 = W*in
   wire signed [9:0] m81_22;
   assign m81_22 =10'b0;

   // m81_23 = W*in
   wire signed [9:0] m81_23;
   assign m81_23 =10'b0;

   // m81_24 = W*in
   wire signed [9:0] m81_24;
   assign m81_24 =10'b0;

   // m81_25 = W*in
   wire signed [9:0] m81_25;
   assign m81_25 ={ {4{in81[5]}} , in81[5:0] };

   // m81_26 = W*in
   wire signed [9:0] m81_26;
   assign m81_26 ={ {4{in81[5]}} , in81[5:0] };

   // m81_27 = W*in
   wire signed [9:0] m81_27;
   assign m81_27 ={ {5{in81[5]}} , in81[5:1] };

   // m81_28 = W*in
   wire signed [9:0] m81_28;
   assign m81_28 ={ {5{in81[5]}} , in81[5:1] };

   // m81_29 = W*in
   wire signed [9:0] m81_29;
   assign m81_29 ={ {5{neg81[5]}} , neg81[5:1] };

   // m81_30 = W*in
   wire signed [9:0] m81_30;
   assign m81_30 =10'b0;

   // m81_31 = W*in
   wire signed [9:0] m81_31;
   assign m81_31 ={ {5{neg81[5]}} , neg81[5:1] };

   // m81_32 = W*in
   wire signed [9:0] m81_32;
   assign m81_32 =10'b0;

   // m81_33 = W*in
   wire signed [9:0] m81_33;
   assign m81_33 ={ {4{in81[5]}} , in81[5:0] };

   // m81_34 = W*in
   wire signed [9:0] m81_34;
   assign m81_34 =10'b0;

   // m81_35 = W*in
   wire signed [9:0] m81_35;
   assign m81_35 =10'b0;

   // m81_36 = W*in
   wire signed [9:0] m81_36;
   assign m81_36 ={ {5{in81[5]}} , in81[5:1] };

   // m81_37 = W*in
   wire signed [9:0] m81_37;
   assign m81_37 =10'b0;

   // m81_38 = W*in
   wire signed [9:0] m81_38;
   assign m81_38 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_39 = W*in
   wire signed [9:0] m81_39;
   assign m81_39 =10'b0;

   // m81_40 = W*in
   wire signed [9:0] m81_40;
   assign m81_40 =10'b0;

   // m81_41 = W*in
   wire signed [9:0] m81_41;
   assign m81_41 =10'b0;

   // m81_42 = W*in
   wire signed [9:0] m81_42;
   assign m81_42 =10'b0;

   // m81_43 = W*in
   wire signed [9:0] m81_43;
   assign m81_43 =10'b0;

   // m81_44 = W*in
   wire signed [9:0] m81_44;
   assign m81_44 =10'b0;

   // m81_45 = W*in
   wire signed [9:0] m81_45;
   assign m81_45 =10'b0;

   // m81_46 = W*in
   wire signed [9:0] m81_46;
   assign m81_46 =10'b0;

   // m81_47 = W*in
   wire signed [9:0] m81_47;
   assign m81_47 =10'b0;

   // m81_48 = W*in
   wire signed [9:0] m81_48;
   assign m81_48 =10'b0;

   // m81_49 = W*in
   wire signed [9:0] m81_49;
   assign m81_49 =10'b0;

   // m81_50 = W*in
   wire signed [9:0] m81_50;
   assign m81_50 =10'b0;

   // m81_51 = W*in
   wire signed [9:0] m81_51;
   assign m81_51 =10'b0;

   // m81_52 = W*in
   wire signed [9:0] m81_52;
   assign m81_52 =10'b0;

   // m81_53 = W*in
   wire signed [9:0] m81_53;
   assign m81_53 =10'b0;

   // m81_54 = W*in
   wire signed [9:0] m81_54;
   assign m81_54 =10'b0;

   // m81_55 = W*in
   wire signed [9:0] m81_55;
   assign m81_55 =10'b0;

   // m81_56 = W*in
   wire signed [9:0] m81_56;
   assign m81_56 =10'b0;

   // m81_57 = W*in
   wire signed [9:0] m81_57;
   assign m81_57 =10'b0;

   // m81_58 = W*in
   wire signed [9:0] m81_58;
   assign m81_58 =10'b0;

   // m81_59 = W*in
   wire signed [9:0] m81_59;
   assign m81_59 ={ {4{in81[5]}} , in81[5:0] };

   // m81_60 = W*in
   wire signed [9:0] m81_60;
   assign m81_60 =10'b0;

   // m81_61 = W*in
   wire signed [9:0] m81_61;
   assign m81_61 =10'b0;

   // m81_62 = W*in
   wire signed [9:0] m81_62;
   assign m81_62 =10'b0;

   // m81_63 = W*in
   wire signed [9:0] m81_63;
   assign m81_63 ={ {3{neg81[5]}} , neg81 , {1{1'b0}} };

   // m81_64 = W*in
   wire signed [9:0] m81_64;
   assign m81_64 =10'b0;

   // m81_65 = W*in
   wire signed [9:0] m81_65;
   assign m81_65 ={ {4{in81[5]}} , in81[5:0] };

   // m81_66 = W*in
   wire signed [9:0] m81_66;
   assign m81_66 ={ {4{in81[5]}} , in81[5:0] };

   // m81_67 = W*in
   wire signed [9:0] m81_67;
   assign m81_67 =10'b0;

   // m81_68 = W*in
   wire signed [9:0] m81_68;
   assign m81_68 =10'b0;

   // m81_69 = W*in
   wire signed [9:0] m81_69;
   assign m81_69 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_70 = W*in
   wire signed [9:0] m81_70;
   assign m81_70 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_71 = W*in
   wire signed [9:0] m81_71;
   assign m81_71 =10'b0;

   // m81_72 = W*in
   wire signed [9:0] m81_72;
   assign m81_72 =10'b0;

   // m81_73 = W*in
   wire signed [9:0] m81_73;
   assign m81_73 =10'b0;

   // m81_74 = W*in
   wire signed [9:0] m81_74;
   assign m81_74 ={ {5{neg81[5]}} , neg81[5:1] };

   // m81_75 = W*in
   wire signed [9:0] m81_75;
   assign m81_75 ={ {5{in81[5]}} , in81[5:1] };

   // m81_76 = W*in
   wire signed [9:0] m81_76;
   assign m81_76 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_77 = W*in
   wire signed [9:0] m81_77;
   assign m81_77 =10'b0;

   // m81_78 = W*in
   wire signed [9:0] m81_78;
   assign m81_78 =10'b0;

   // m81_79 = W*in
   wire signed [9:0] m81_79;
   assign m81_79 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_80 = W*in
   wire signed [9:0] m81_80;
   assign m81_80 =10'b0;

   // m81_81 = W*in
   wire signed [9:0] m81_81;
   assign m81_81 ={ {5{in81[5]}} , in81[5:1] };

   // m81_82 = W*in
   wire signed [9:0] m81_82;
   assign m81_82 =10'b0;

   // m81_83 = W*in
   wire signed [9:0] m81_83;
   assign m81_83 =10'b0;

   // m81_84 = W*in
   wire signed [9:0] m81_84;
   assign m81_84 =10'b0;

   // m81_85 = W*in
   wire signed [9:0] m81_85;
   assign m81_85 =10'b0;

   // m81_86 = W*in
   wire signed [9:0] m81_86;
   assign m81_86 =10'b0;

   // m81_87 = W*in
   wire signed [9:0] m81_87;
   assign m81_87 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_88 = W*in
   wire signed [9:0] m81_88;
   assign m81_88 =10'b0;

   // m81_89 = W*in
   wire signed [9:0] m81_89;
   assign m81_89 =10'b0;

   // m81_90 = W*in
   wire signed [9:0] m81_90;
   assign m81_90 =10'b0;

   // m81_91 = W*in
   wire signed [9:0] m81_91;
   assign m81_91 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_92 = W*in
   wire signed [9:0] m81_92;
   assign m81_92 =10'b0;

   // m81_93 = W*in
   wire signed [9:0] m81_93;
   assign m81_93 =10'b0;

   // m81_94 = W*in
   wire signed [9:0] m81_94;
   assign m81_94 =10'b0;

   // m81_95 = W*in
   wire signed [9:0] m81_95;
   assign m81_95 =10'b0;

   // m81_96 = W*in
   wire signed [9:0] m81_96;
   assign m81_96 =10'b0;

   // m81_97 = W*in
   wire signed [9:0] m81_97;
   assign m81_97 =10'b0;

   // m81_98 = W*in
   wire signed [9:0] m81_98;
   assign m81_98 =10'b0;

   // m81_99 = W*in
   wire signed [9:0] m81_99;
   assign m81_99 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_100 = W*in
   wire signed [9:0] m81_100;
   assign m81_100 =10'b0;

   // m81_101 = W*in
   wire signed [9:0] m81_101;
   assign m81_101 =10'b0;

   // m81_102 = W*in
   wire signed [9:0] m81_102;
   assign m81_102 =10'b0;

   // m81_103 = W*in
   wire signed [9:0] m81_103;
   assign m81_103 =10'b0;

   // m81_104 = W*in
   wire signed [9:0] m81_104;
   assign m81_104 =10'b0;

   // m81_105 = W*in
   wire signed [9:0] m81_105;
   assign m81_105 =10'b0;

   // m81_106 = W*in
   wire signed [9:0] m81_106;
   assign m81_106 =10'b0;

   // m81_107 = W*in
   wire signed [9:0] m81_107;
   assign m81_107 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_108 = W*in
   wire signed [9:0] m81_108;
   assign m81_108 =10'b0;

   // m81_109 = W*in
   wire signed [9:0] m81_109;
   assign m81_109 =10'b0;

   // m81_110 = W*in
   wire signed [9:0] m81_110;
   assign m81_110 =10'b0;

   // m81_111 = W*in
   wire signed [9:0] m81_111;
   assign m81_111 ={ {4{in81[5]}} , in81[5:0] };

   // m81_112 = W*in
   wire signed [9:0] m81_112;
   assign m81_112 =10'b0;

   // m81_113 = W*in
   wire signed [9:0] m81_113;
   assign m81_113 =10'b0;

   // m81_114 = W*in
   wire signed [9:0] m81_114;
   assign m81_114 =10'b0;

   // m81_115 = W*in
   wire signed [9:0] m81_115;
   assign m81_115 =10'b0;

   // m81_116 = W*in
   wire signed [9:0] m81_116;
   assign m81_116 ={ {4{neg81[5]}} , neg81[5:0] };

   // m81_117 = W*in
   wire signed [9:0] m81_117;
   assign m81_117 =10'b0;

   // m82_1 = W*in
   wire signed [9:0] m82_1;
   assign m82_1 =10'b0;

   // m82_2 = W*in
   wire signed [9:0] m82_2;
   assign m82_2 =10'b0;

   // m82_3 = W*in
   wire signed [9:0] m82_3;
   assign m82_3 =10'b0;

   // m82_4 = W*in
   wire signed [9:0] m82_4;
   assign m82_4 =10'b0;

   // m82_5 = W*in
   wire signed [9:0] m82_5;
   assign m82_5 =10'b0;

   // m82_6 = W*in
   wire signed [9:0] m82_6;
   assign m82_6 =10'b0;

   // m82_7 = W*in
   wire signed [9:0] m82_7;
   assign m82_7 =10'b0;

   // m82_8 = W*in
   wire signed [9:0] m82_8;
   assign m82_8 =10'b0;

   // m82_9 = W*in
   wire signed [9:0] m82_9;
   assign m82_9 =10'b0;

   // m82_10 = W*in
   wire signed [9:0] m82_10;
   assign m82_10 =10'b0;

   // m82_11 = W*in
   wire signed [9:0] m82_11;
   assign m82_11 =10'b0;

   // m82_12 = W*in
   wire signed [9:0] m82_12;
   assign m82_12 =10'b0;

   // m82_13 = W*in
   wire signed [9:0] m82_13;
   assign m82_13 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_14 = W*in
   wire signed [9:0] m82_14;
   assign m82_14 =10'b0;

   // m82_15 = W*in
   wire signed [9:0] m82_15;
   assign m82_15 =10'b0;

   // m82_16 = W*in
   wire signed [9:0] m82_16;
   assign m82_16 =10'b0;

   // m82_17 = W*in
   wire signed [9:0] m82_17;
   assign m82_17 =10'b0;

   // m82_18 = W*in
   wire signed [9:0] m82_18;
   assign m82_18 ={ {4{in82[5]}} , in82[5:0] };

   // m82_19 = W*in
   wire signed [9:0] m82_19;
   assign m82_19 ={ {5{in82[5]}} , in82[5:1] };

   // m82_20 = W*in
   wire signed [9:0] m82_20;
   assign m82_20 ={ {5{neg82[5]}} , neg82[5:1] };

   // m82_21 = W*in
   wire signed [9:0] m82_21;
   assign m82_21 =10'b0;

   // m82_22 = W*in
   wire signed [9:0] m82_22;
   assign m82_22 =10'b0;

   // m82_23 = W*in
   wire signed [9:0] m82_23;
   assign m82_23 =10'b0;

   // m82_24 = W*in
   wire signed [9:0] m82_24;
   assign m82_24 =10'b0;

   // m82_25 = W*in
   wire signed [9:0] m82_25;
   assign m82_25 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_26 = W*in
   wire signed [9:0] m82_26;
   assign m82_26 ={ {5{in82[5]}} , in82[5:1] };

   // m82_27 = W*in
   wire signed [9:0] m82_27;
   assign m82_27 ={ {5{neg82[5]}} , neg82[5:1] };

   // m82_28 = W*in
   wire signed [9:0] m82_28;
   assign m82_28 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_29 = W*in
   wire signed [9:0] m82_29;
   assign m82_29 =10'b0;

   // m82_30 = W*in
   wire signed [9:0] m82_30;
   assign m82_30 =10'b0;

   // m82_31 = W*in
   wire signed [9:0] m82_31;
   assign m82_31 =10'b0;

   // m82_32 = W*in
   wire signed [9:0] m82_32;
   assign m82_32 =10'b0;

   // m82_33 = W*in
   wire signed [9:0] m82_33;
   assign m82_33 =10'b0;

   // m82_34 = W*in
   wire signed [9:0] m82_34;
   assign m82_34 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_35 = W*in
   wire signed [9:0] m82_35;
   assign m82_35 ={ {5{neg82[5]}} , neg82[5:1] };

   // m82_36 = W*in
   wire signed [9:0] m82_36;
   assign m82_36 =10'b0;

   // m82_37 = W*in
   wire signed [9:0] m82_37;
   assign m82_37 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_38 = W*in
   wire signed [9:0] m82_38;
   assign m82_38 =10'b0;

   // m82_39 = W*in
   wire signed [9:0] m82_39;
   assign m82_39 =10'b0;

   // m82_40 = W*in
   wire signed [9:0] m82_40;
   assign m82_40 =10'b0;

   // m82_41 = W*in
   wire signed [9:0] m82_41;
   assign m82_41 =10'b0;

   // m82_42 = W*in
   wire signed [9:0] m82_42;
   assign m82_42 ={ {4{in82[5]}} , in82[5:0] };

   // m82_43 = W*in
   wire signed [9:0] m82_43;
   assign m82_43 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_44 = W*in
   wire signed [9:0] m82_44;
   assign m82_44 =10'b0;

   // m82_45 = W*in
   wire signed [9:0] m82_45;
   assign m82_45 =10'b0;

   // m82_46 = W*in
   wire signed [9:0] m82_46;
   assign m82_46 =10'b0;

   // m82_47 = W*in
   wire signed [9:0] m82_47;
   assign m82_47 =10'b0;

   // m82_48 = W*in
   wire signed [9:0] m82_48;
   assign m82_48 =10'b0;

   // m82_49 = W*in
   wire signed [9:0] m82_49;
   assign m82_49 =10'b0;

   // m82_50 = W*in
   wire signed [9:0] m82_50;
   assign m82_50 =10'b0;

   // m82_51 = W*in
   wire signed [9:0] m82_51;
   assign m82_51 =10'b0;

   // m82_52 = W*in
   wire signed [9:0] m82_52;
   assign m82_52 =10'b0;

   // m82_53 = W*in
   wire signed [9:0] m82_53;
   assign m82_53 =10'b0;

   // m82_54 = W*in
   wire signed [9:0] m82_54;
   assign m82_54 =10'b0;

   // m82_55 = W*in
   wire signed [9:0] m82_55;
   assign m82_55 =10'b0;

   // m82_56 = W*in
   wire signed [9:0] m82_56;
   assign m82_56 =10'b0;

   // m82_57 = W*in
   wire signed [9:0] m82_57;
   assign m82_57 =10'b0;

   // m82_58 = W*in
   wire signed [9:0] m82_58;
   assign m82_58 =10'b0;

   // m82_59 = W*in
   wire signed [9:0] m82_59;
   assign m82_59 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_60 = W*in
   wire signed [9:0] m82_60;
   assign m82_60 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_61 = W*in
   wire signed [9:0] m82_61;
   assign m82_61 =10'b0;

   // m82_62 = W*in
   wire signed [9:0] m82_62;
   assign m82_62 =10'b0;

   // m82_63 = W*in
   wire signed [9:0] m82_63;
   assign m82_63 =10'b0;

   // m82_64 = W*in
   wire signed [9:0] m82_64;
   assign m82_64 ={ {4{in82[5]}} , in82[5:0] };

   // m82_65 = W*in
   wire signed [9:0] m82_65;
   assign m82_65 ={ {4{in82[5]}} , in82[5:0] };

   // m82_66 = W*in
   wire signed [9:0] m82_66;
   assign m82_66 ={ {4{in82[5]}} , in82[5:0] };

   // m82_67 = W*in
   wire signed [9:0] m82_67;
   assign m82_67 ={ {4{in82[5]}} , in82[5:0] };

   // m82_68 = W*in
   wire signed [9:0] m82_68;
   assign m82_68 =10'b0;

   // m82_69 = W*in
   wire signed [9:0] m82_69;
   assign m82_69 =10'b0;

   // m82_70 = W*in
   wire signed [9:0] m82_70;
   assign m82_70 =10'b0;

   // m82_71 = W*in
   wire signed [9:0] m82_71;
   assign m82_71 =10'b0;

   // m82_72 = W*in
   wire signed [9:0] m82_72;
   assign m82_72 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_73 = W*in
   wire signed [9:0] m82_73;
   assign m82_73 =10'b0;

   // m82_74 = W*in
   wire signed [9:0] m82_74;
   assign m82_74 =10'b0;

   // m82_75 = W*in
   wire signed [9:0] m82_75;
   assign m82_75 =10'b0;

   // m82_76 = W*in
   wire signed [9:0] m82_76;
   assign m82_76 =10'b0;

   // m82_77 = W*in
   wire signed [9:0] m82_77;
   assign m82_77 ={ {4{in82[5]}} , in82[5:0] };

   // m82_78 = W*in
   wire signed [9:0] m82_78;
   assign m82_78 =10'b0;

   // m82_79 = W*in
   wire signed [9:0] m82_79;
   assign m82_79 =10'b0;

   // m82_80 = W*in
   wire signed [9:0] m82_80;
   assign m82_80 =10'b0;

   // m82_81 = W*in
   wire signed [9:0] m82_81;
   assign m82_81 ={ {4{in82[5]}} , in82[5:0] };

   // m82_82 = W*in
   wire signed [9:0] m82_82;
   assign m82_82 =10'b0;

   // m82_83 = W*in
   wire signed [9:0] m82_83;
   assign m82_83 =10'b0;

   // m82_84 = W*in
   wire signed [9:0] m82_84;
   assign m82_84 =10'b0;

   // m82_85 = W*in
   wire signed [9:0] m82_85;
   assign m82_85 =10'b0;

   // m82_86 = W*in
   wire signed [9:0] m82_86;
   assign m82_86 ={ {4{in82[5]}} , in82[5:0] };

   // m82_87 = W*in
   wire signed [9:0] m82_87;
   assign m82_87 =10'b0;

   // m82_88 = W*in
   wire signed [9:0] m82_88;
   assign m82_88 =10'b0;

   // m82_89 = W*in
   wire signed [9:0] m82_89;
   assign m82_89 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_90 = W*in
   wire signed [9:0] m82_90;
   assign m82_90 =10'b0;

   // m82_91 = W*in
   wire signed [9:0] m82_91;
   assign m82_91 ={ {4{in82[5]}} , in82[5:0] };

   // m82_92 = W*in
   wire signed [9:0] m82_92;
   assign m82_92 =10'b0;

   // m82_93 = W*in
   wire signed [9:0] m82_93;
   assign m82_93 =10'b0;

   // m82_94 = W*in
   wire signed [9:0] m82_94;
   assign m82_94 ={ {4{in82[5]}} , in82[5:0] };

   // m82_95 = W*in
   wire signed [9:0] m82_95;
   assign m82_95 =10'b0;

   // m82_96 = W*in
   wire signed [9:0] m82_96;
   assign m82_96 =10'b0;

   // m82_97 = W*in
   wire signed [9:0] m82_97;
   assign m82_97 ={ {4{in82[5]}} , in82[5:0] };

   // m82_98 = W*in
   wire signed [9:0] m82_98;
   assign m82_98 =10'b0;

   // m82_99 = W*in
   wire signed [9:0] m82_99;
   assign m82_99 =10'b0;

   // m82_100 = W*in
   wire signed [9:0] m82_100;
   assign m82_100 =10'b0;

   // m82_101 = W*in
   wire signed [9:0] m82_101;
   assign m82_101 =10'b0;

   // m82_102 = W*in
   wire signed [9:0] m82_102;
   assign m82_102 =10'b0;

   // m82_103 = W*in
   wire signed [9:0] m82_103;
   assign m82_103 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_104 = W*in
   wire signed [9:0] m82_104;
   assign m82_104 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_105 = W*in
   wire signed [9:0] m82_105;
   assign m82_105 =10'b0;

   // m82_106 = W*in
   wire signed [9:0] m82_106;
   assign m82_106 =10'b0;

   // m82_107 = W*in
   wire signed [9:0] m82_107;
   assign m82_107 =10'b0;

   // m82_108 = W*in
   wire signed [9:0] m82_108;
   assign m82_108 =10'b0;

   // m82_109 = W*in
   wire signed [9:0] m82_109;
   assign m82_109 ={ {4{neg82[5]}} , neg82[5:0] };

   // m82_110 = W*in
   wire signed [9:0] m82_110;
   assign m82_110 ={ {4{in82[5]}} , in82[5:0] };

   // m82_111 = W*in
   wire signed [9:0] m82_111;
   assign m82_111 =10'b0;

   // m82_112 = W*in
   wire signed [9:0] m82_112;
   assign m82_112 =10'b0;

   // m82_113 = W*in
   wire signed [9:0] m82_113;
   assign m82_113 =10'b0;

   // m82_114 = W*in
   wire signed [9:0] m82_114;
   assign m82_114 ={ {5{neg82[5]}} , neg82[5:1] };

   // m82_115 = W*in
   wire signed [9:0] m82_115;
   assign m82_115 =10'b0;

   // m82_116 = W*in
   wire signed [9:0] m82_116;
   assign m82_116 =10'b0;

   // m82_117 = W*in
   wire signed [9:0] m82_117;
   assign m82_117 ={ {4{neg82[5]}} , neg82[5:0] };

   // m83_1 = W*in
   wire signed [9:0] m83_1;
   assign m83_1 =10'b0;

   // m83_2 = W*in
   wire signed [9:0] m83_2;
   assign m83_2 =10'b0;

   // m83_3 = W*in
   wire signed [9:0] m83_3;
   assign m83_3 =10'b0;

   // m83_4 = W*in
   wire signed [9:0] m83_4;
   assign m83_4 =10'b0;

   // m83_5 = W*in
   wire signed [9:0] m83_5;
   assign m83_5 ={ {4{in83[5]}} , in83[5:0] };

   // m83_6 = W*in
   wire signed [9:0] m83_6;
   assign m83_6 ={ {4{in83[5]}} , in83[5:0] };

   // m83_7 = W*in
   wire signed [9:0] m83_7;
   assign m83_7 =10'b0;

   // m83_8 = W*in
   wire signed [9:0] m83_8;
   assign m83_8 =10'b0;

   // m83_9 = W*in
   wire signed [9:0] m83_9;
   assign m83_9 =10'b0;

   // m83_10 = W*in
   wire signed [9:0] m83_10;
   assign m83_10 =10'b0;

   // m83_11 = W*in
   wire signed [9:0] m83_11;
   assign m83_11 =10'b0;

   // m83_12 = W*in
   wire signed [9:0] m83_12;
   assign m83_12 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_13 = W*in
   wire signed [9:0] m83_13;
   assign m83_13 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_14 = W*in
   wire signed [9:0] m83_14;
   assign m83_14 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_15 = W*in
   wire signed [9:0] m83_15;
   assign m83_15 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_16 = W*in
   wire signed [9:0] m83_16;
   assign m83_16 =10'b0;

   // m83_17 = W*in
   wire signed [9:0] m83_17;
   assign m83_17 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_18 = W*in
   wire signed [9:0] m83_18;
   assign m83_18 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_19 = W*in
   wire signed [9:0] m83_19;
   assign m83_19 ={ {4{in83[5]}} , in83[5:0] };

   // m83_20 = W*in
   wire signed [9:0] m83_20;
   assign m83_20 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_21 = W*in
   wire signed [9:0] m83_21;
   assign m83_21 =10'b0;

   // m83_22 = W*in
   wire signed [9:0] m83_22;
   assign m83_22 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_23 = W*in
   wire signed [9:0] m83_23;
   assign m83_23 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_24 = W*in
   wire signed [9:0] m83_24;
   assign m83_24 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_25 = W*in
   wire signed [9:0] m83_25;
   assign m83_25 =10'b0;

   // m83_26 = W*in
   wire signed [9:0] m83_26;
   assign m83_26 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_27 = W*in
   wire signed [9:0] m83_27;
   assign m83_27 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_28 = W*in
   wire signed [9:0] m83_28;
   assign m83_28 ={ {5{in83[5]}} , in83[5:1] };

   // m83_29 = W*in
   wire signed [9:0] m83_29;
   assign m83_29 ={ {5{in83[5]}} , in83[5:1] };

   // m83_30 = W*in
   wire signed [9:0] m83_30;
   assign m83_30 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_31 = W*in
   wire signed [9:0] m83_31;
   assign m83_31 ={ {5{neg83[5]}} , neg83[5:1] };

   // m83_32 = W*in
   wire signed [9:0] m83_32;
   assign m83_32 =10'b0;

   // m83_33 = W*in
   wire signed [9:0] m83_33;
   assign m83_33 ={ {4{in83[5]}} , in83[5:0] };

   // m83_34 = W*in
   wire signed [9:0] m83_34;
   assign m83_34 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_35 = W*in
   wire signed [9:0] m83_35;
   assign m83_35 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_36 = W*in
   wire signed [9:0] m83_36;
   assign m83_36 ={ {4{in83[5]}} , in83[5:0] };

   // m83_37 = W*in
   wire signed [9:0] m83_37;
   assign m83_37 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_38 = W*in
   wire signed [9:0] m83_38;
   assign m83_38 ={ {4{in83[5]}} , in83[5:0] };

   // m83_39 = W*in
   wire signed [9:0] m83_39;
   assign m83_39 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_40 = W*in
   wire signed [9:0] m83_40;
   assign m83_40 =10'b0;

   // m83_41 = W*in
   wire signed [9:0] m83_41;
   assign m83_41 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_42 = W*in
   wire signed [9:0] m83_42;
   assign m83_42 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_43 = W*in
   wire signed [9:0] m83_43;
   assign m83_43 =10'b0;

   // m83_44 = W*in
   wire signed [9:0] m83_44;
   assign m83_44 ={ {4{in83[5]}} , in83[5:0] };

   // m83_45 = W*in
   wire signed [9:0] m83_45;
   assign m83_45 =10'b0;

   // m83_46 = W*in
   wire signed [9:0] m83_46;
   assign m83_46 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_47 = W*in
   wire signed [9:0] m83_47;
   assign m83_47 =10'b0;

   // m83_48 = W*in
   wire signed [9:0] m83_48;
   assign m83_48 =10'b0;

   // m83_49 = W*in
   wire signed [9:0] m83_49;
   assign m83_49 =10'b0;

   // m83_50 = W*in
   wire signed [9:0] m83_50;
   assign m83_50 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_51 = W*in
   wire signed [9:0] m83_51;
   assign m83_51 =10'b0;

   // m83_52 = W*in
   wire signed [9:0] m83_52;
   assign m83_52 =10'b0;

   // m83_53 = W*in
   wire signed [9:0] m83_53;
   assign m83_53 ={ {4{in83[5]}} , in83[5:0] };

   // m83_54 = W*in
   wire signed [9:0] m83_54;
   assign m83_54 ={ {4{in83[5]}} , in83[5:0] };

   // m83_55 = W*in
   wire signed [9:0] m83_55;
   assign m83_55 =10'b0;

   // m83_56 = W*in
   wire signed [9:0] m83_56;
   assign m83_56 =10'b0;

   // m83_57 = W*in
   wire signed [9:0] m83_57;
   assign m83_57 =10'b0;

   // m83_58 = W*in
   wire signed [9:0] m83_58;
   assign m83_58 ={ {5{neg83[5]}} , neg83[5:1] };

   // m83_59 = W*in
   wire signed [9:0] m83_59;
   assign m83_59 ={ {4{in83[5]}} , in83[5:0] };

   // m83_60 = W*in
   wire signed [9:0] m83_60;
   assign m83_60 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_61 = W*in
   wire signed [9:0] m83_61;
   assign m83_61 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_62 = W*in
   wire signed [9:0] m83_62;
   assign m83_62 =10'b0;

   // m83_63 = W*in
   wire signed [9:0] m83_63;
   assign m83_63 =10'b0;

   // m83_64 = W*in
   wire signed [9:0] m83_64;
   assign m83_64 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_65 = W*in
   wire signed [9:0] m83_65;
   assign m83_65 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_66 = W*in
   wire signed [9:0] m83_66;
   assign m83_66 ={ {4{in83[5]}} , in83[5:0] };

   // m83_67 = W*in
   wire signed [9:0] m83_67;
   assign m83_67 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_68 = W*in
   wire signed [9:0] m83_68;
   assign m83_68 =10'b0;

   // m83_69 = W*in
   wire signed [9:0] m83_69;
   assign m83_69 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_70 = W*in
   wire signed [9:0] m83_70;
   assign m83_70 =10'b0;

   // m83_71 = W*in
   wire signed [9:0] m83_71;
   assign m83_71 =10'b0;

   // m83_72 = W*in
   wire signed [9:0] m83_72;
   assign m83_72 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_73 = W*in
   wire signed [9:0] m83_73;
   assign m83_73 ={ {4{in83[5]}} , in83[5:0] };

   // m83_74 = W*in
   wire signed [9:0] m83_74;
   assign m83_74 =10'b0;

   // m83_75 = W*in
   wire signed [9:0] m83_75;
   assign m83_75 ={ {4{in83[5]}} , in83[5:0] };

   // m83_76 = W*in
   wire signed [9:0] m83_76;
   assign m83_76 =10'b0;

   // m83_77 = W*in
   wire signed [9:0] m83_77;
   assign m83_77 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_78 = W*in
   wire signed [9:0] m83_78;
   assign m83_78 ={ {4{in83[5]}} , in83[5:0] };

   // m83_79 = W*in
   wire signed [9:0] m83_79;
   assign m83_79 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_80 = W*in
   wire signed [9:0] m83_80;
   assign m83_80 =10'b0;

   // m83_81 = W*in
   wire signed [9:0] m83_81;
   assign m83_81 ={ {5{in83[5]}} , in83[5:1] };

   // m83_82 = W*in
   wire signed [9:0] m83_82;
   assign m83_82 =10'b0;

   // m83_83 = W*in
   wire signed [9:0] m83_83;
   assign m83_83 ={ {5{neg83[5]}} , neg83[5:1] };

   // m83_84 = W*in
   wire signed [9:0] m83_84;
   assign m83_84 =10'b0;

   // m83_85 = W*in
   wire signed [9:0] m83_85;
   assign m83_85 =10'b0;

   // m83_86 = W*in
   wire signed [9:0] m83_86;
   assign m83_86 =10'b0;

   // m83_87 = W*in
   wire signed [9:0] m83_87;
   assign m83_87 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_88 = W*in
   wire signed [9:0] m83_88;
   assign m83_88 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_89 = W*in
   wire signed [9:0] m83_89;
   assign m83_89 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_90 = W*in
   wire signed [9:0] m83_90;
   assign m83_90 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_91 = W*in
   wire signed [9:0] m83_91;
   assign m83_91 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_92 = W*in
   wire signed [9:0] m83_92;
   assign m83_92 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_93 = W*in
   wire signed [9:0] m83_93;
   assign m83_93 ={ {4{in83[5]}} , in83[5:0] };

   // m83_94 = W*in
   wire signed [9:0] m83_94;
   assign m83_94 ={ {4{in83[5]}} , in83[5:0] };

   // m83_95 = W*in
   wire signed [9:0] m83_95;
   assign m83_95 =10'b0;

   // m83_96 = W*in
   wire signed [9:0] m83_96;
   assign m83_96 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_97 = W*in
   wire signed [9:0] m83_97;
   assign m83_97 ={ {3{in83[5]}} , in83 , {1{1'b0}} };

   // m83_98 = W*in
   wire signed [9:0] m83_98;
   assign m83_98 =10'b0;

   // m83_99 = W*in
   wire signed [9:0] m83_99;
   assign m83_99 =10'b0;

   // m83_100 = W*in
   wire signed [9:0] m83_100;
   assign m83_100 ={ {4{in83[5]}} , in83[5:0] };

   // m83_101 = W*in
   wire signed [9:0] m83_101;
   assign m83_101 =10'b0;

   // m83_102 = W*in
   wire signed [9:0] m83_102;
   assign m83_102 =10'b0;

   // m83_103 = W*in
   wire signed [9:0] m83_103;
   assign m83_103 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_104 = W*in
   wire signed [9:0] m83_104;
   assign m83_104 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_105 = W*in
   wire signed [9:0] m83_105;
   assign m83_105 =10'b0;

   // m83_106 = W*in
   wire signed [9:0] m83_106;
   assign m83_106 =10'b0;

   // m83_107 = W*in
   wire signed [9:0] m83_107;
   assign m83_107 =10'b0;

   // m83_108 = W*in
   wire signed [9:0] m83_108;
   assign m83_108 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_109 = W*in
   wire signed [9:0] m83_109;
   assign m83_109 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_110 = W*in
   wire signed [9:0] m83_110;
   assign m83_110 ={ {4{in83[5]}} , in83[5:0] };

   // m83_111 = W*in
   wire signed [9:0] m83_111;
   assign m83_111 =10'b0;

   // m83_112 = W*in
   wire signed [9:0] m83_112;
   assign m83_112 ={ {4{in83[5]}} , in83[5:0] };

   // m83_113 = W*in
   wire signed [9:0] m83_113;
   assign m83_113 =10'b0;

   // m83_114 = W*in
   wire signed [9:0] m83_114;
   assign m83_114 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_115 = W*in
   wire signed [9:0] m83_115;
   assign m83_115 ={ {4{neg83[5]}} , neg83[5:0] };

   // m83_116 = W*in
   wire signed [9:0] m83_116;
   assign m83_116 ={ {3{neg83[5]}} , neg83 , {1{1'b0}} };

   // m83_117 = W*in
   wire signed [9:0] m83_117;
   assign m83_117 ={ {4{neg83[5]}} , neg83[5:0] };

   // m84_1 = W*in
   wire signed [9:0] m84_1;
   assign m84_1 =10'b0;

   // m84_2 = W*in
   wire signed [9:0] m84_2;
   assign m84_2 =10'b0;

   // m84_3 = W*in
   wire signed [9:0] m84_3;
   assign m84_3 =10'b0;

   // m84_4 = W*in
   wire signed [9:0] m84_4;
   assign m84_4 =10'b0;

   // m84_5 = W*in
   wire signed [9:0] m84_5;
   assign m84_5 =10'b0;

   // m84_6 = W*in
   wire signed [9:0] m84_6;
   assign m84_6 =10'b0;

   // m84_7 = W*in
   wire signed [9:0] m84_7;
   assign m84_7 =10'b0;

   // m84_8 = W*in
   wire signed [9:0] m84_8;
   assign m84_8 =10'b0;

   // m84_9 = W*in
   wire signed [9:0] m84_9;
   assign m84_9 =10'b0;

   // m84_10 = W*in
   wire signed [9:0] m84_10;
   assign m84_10 =10'b0;

   // m84_11 = W*in
   wire signed [9:0] m84_11;
   assign m84_11 =10'b0;

   // m84_12 = W*in
   wire signed [9:0] m84_12;
   assign m84_12 =10'b0;

   // m84_13 = W*in
   wire signed [9:0] m84_13;
   assign m84_13 =10'b0;

   // m84_14 = W*in
   wire signed [9:0] m84_14;
   assign m84_14 =10'b0;

   // m84_15 = W*in
   wire signed [9:0] m84_15;
   assign m84_15 =10'b0;

   // m84_16 = W*in
   wire signed [9:0] m84_16;
   assign m84_16 =10'b0;

   // m84_17 = W*in
   wire signed [9:0] m84_17;
   assign m84_17 =10'b0;

   // m84_18 = W*in
   wire signed [9:0] m84_18;
   assign m84_18 ={ {5{in84[5]}} , in84[5:1] };

   // m84_19 = W*in
   wire signed [9:0] m84_19;
   assign m84_19 ={ {5{in84[5]}} , in84[5:1] };

   // m84_20 = W*in
   wire signed [9:0] m84_20;
   assign m84_20 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_21 = W*in
   wire signed [9:0] m84_21;
   assign m84_21 =10'b0;

   // m84_22 = W*in
   wire signed [9:0] m84_22;
   assign m84_22 ={ {5{neg84[5]}} , neg84[5:1] };

   // m84_23 = W*in
   wire signed [9:0] m84_23;
   assign m84_23 =10'b0;

   // m84_24 = W*in
   wire signed [9:0] m84_24;
   assign m84_24 =10'b0;

   // m84_25 = W*in
   wire signed [9:0] m84_25;
   assign m84_25 =10'b0;

   // m84_26 = W*in
   wire signed [9:0] m84_26;
   assign m84_26 =10'b0;

   // m84_27 = W*in
   wire signed [9:0] m84_27;
   assign m84_27 =10'b0;

   // m84_28 = W*in
   wire signed [9:0] m84_28;
   assign m84_28 ={ {5{in84[5]}} , in84[5:1] };

   // m84_29 = W*in
   wire signed [9:0] m84_29;
   assign m84_29 =10'b0;

   // m84_30 = W*in
   wire signed [9:0] m84_30;
   assign m84_30 =10'b0;

   // m84_31 = W*in
   wire signed [9:0] m84_31;
   assign m84_31 =10'b0;

   // m84_32 = W*in
   wire signed [9:0] m84_32;
   assign m84_32 =10'b0;

   // m84_33 = W*in
   wire signed [9:0] m84_33;
   assign m84_33 =10'b0;

   // m84_34 = W*in
   wire signed [9:0] m84_34;
   assign m84_34 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_35 = W*in
   wire signed [9:0] m84_35;
   assign m84_35 =10'b0;

   // m84_36 = W*in
   wire signed [9:0] m84_36;
   assign m84_36 ={ {5{in84[5]}} , in84[5:1] };

   // m84_37 = W*in
   wire signed [9:0] m84_37;
   assign m84_37 =10'b0;

   // m84_38 = W*in
   wire signed [9:0] m84_38;
   assign m84_38 =10'b0;

   // m84_39 = W*in
   wire signed [9:0] m84_39;
   assign m84_39 =10'b0;

   // m84_40 = W*in
   wire signed [9:0] m84_40;
   assign m84_40 =10'b0;

   // m84_41 = W*in
   wire signed [9:0] m84_41;
   assign m84_41 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_42 = W*in
   wire signed [9:0] m84_42;
   assign m84_42 ={ {4{in84[5]}} , in84[5:0] };

   // m84_43 = W*in
   wire signed [9:0] m84_43;
   assign m84_43 =10'b0;

   // m84_44 = W*in
   wire signed [9:0] m84_44;
   assign m84_44 =10'b0;

   // m84_45 = W*in
   wire signed [9:0] m84_45;
   assign m84_45 ={ {4{in84[5]}} , in84[5:0] };

   // m84_46 = W*in
   wire signed [9:0] m84_46;
   assign m84_46 =10'b0;

   // m84_47 = W*in
   wire signed [9:0] m84_47;
   assign m84_47 =10'b0;

   // m84_48 = W*in
   wire signed [9:0] m84_48;
   assign m84_48 =10'b0;

   // m84_49 = W*in
   wire signed [9:0] m84_49;
   assign m84_49 =10'b0;

   // m84_50 = W*in
   wire signed [9:0] m84_50;
   assign m84_50 =10'b0;

   // m84_51 = W*in
   wire signed [9:0] m84_51;
   assign m84_51 =10'b0;

   // m84_52 = W*in
   wire signed [9:0] m84_52;
   assign m84_52 =10'b0;

   // m84_53 = W*in
   wire signed [9:0] m84_53;
   assign m84_53 =10'b0;

   // m84_54 = W*in
   wire signed [9:0] m84_54;
   assign m84_54 =10'b0;

   // m84_55 = W*in
   wire signed [9:0] m84_55;
   assign m84_55 =10'b0;

   // m84_56 = W*in
   wire signed [9:0] m84_56;
   assign m84_56 =10'b0;

   // m84_57 = W*in
   wire signed [9:0] m84_57;
   assign m84_57 =10'b0;

   // m84_58 = W*in
   wire signed [9:0] m84_58;
   assign m84_58 =10'b0;

   // m84_59 = W*in
   wire signed [9:0] m84_59;
   assign m84_59 =10'b0;

   // m84_60 = W*in
   wire signed [9:0] m84_60;
   assign m84_60 =10'b0;

   // m84_61 = W*in
   wire signed [9:0] m84_61;
   assign m84_61 =10'b0;

   // m84_62 = W*in
   wire signed [9:0] m84_62;
   assign m84_62 =10'b0;

   // m84_63 = W*in
   wire signed [9:0] m84_63;
   assign m84_63 =10'b0;

   // m84_64 = W*in
   wire signed [9:0] m84_64;
   assign m84_64 =10'b0;

   // m84_65 = W*in
   wire signed [9:0] m84_65;
   assign m84_65 =10'b0;

   // m84_66 = W*in
   wire signed [9:0] m84_66;
   assign m84_66 ={ {5{in84[5]}} , in84[5:1] };

   // m84_67 = W*in
   wire signed [9:0] m84_67;
   assign m84_67 =10'b0;

   // m84_68 = W*in
   wire signed [9:0] m84_68;
   assign m84_68 =10'b0;

   // m84_69 = W*in
   wire signed [9:0] m84_69;
   assign m84_69 =10'b0;

   // m84_70 = W*in
   wire signed [9:0] m84_70;
   assign m84_70 =10'b0;

   // m84_71 = W*in
   wire signed [9:0] m84_71;
   assign m84_71 ={ {5{in84[5]}} , in84[5:1] };

   // m84_72 = W*in
   wire signed [9:0] m84_72;
   assign m84_72 =10'b0;

   // m84_73 = W*in
   wire signed [9:0] m84_73;
   assign m84_73 ={ {5{in84[5]}} , in84[5:1] };

   // m84_74 = W*in
   wire signed [9:0] m84_74;
   assign m84_74 =10'b0;

   // m84_75 = W*in
   wire signed [9:0] m84_75;
   assign m84_75 =10'b0;

   // m84_76 = W*in
   wire signed [9:0] m84_76;
   assign m84_76 =10'b0;

   // m84_77 = W*in
   wire signed [9:0] m84_77;
   assign m84_77 ={ {4{in84[5]}} , in84[5:0] };

   // m84_78 = W*in
   wire signed [9:0] m84_78;
   assign m84_78 =10'b0;

   // m84_79 = W*in
   wire signed [9:0] m84_79;
   assign m84_79 =10'b0;

   // m84_80 = W*in
   wire signed [9:0] m84_80;
   assign m84_80 =10'b0;

   // m84_81 = W*in
   wire signed [9:0] m84_81;
   assign m84_81 =10'b0;

   // m84_82 = W*in
   wire signed [9:0] m84_82;
   assign m84_82 =10'b0;

   // m84_83 = W*in
   wire signed [9:0] m84_83;
   assign m84_83 =10'b0;

   // m84_84 = W*in
   wire signed [9:0] m84_84;
   assign m84_84 =10'b0;

   // m84_85 = W*in
   wire signed [9:0] m84_85;
   assign m84_85 =10'b0;

   // m84_86 = W*in
   wire signed [9:0] m84_86;
   assign m84_86 =10'b0;

   // m84_87 = W*in
   wire signed [9:0] m84_87;
   assign m84_87 =10'b0;

   // m84_88 = W*in
   wire signed [9:0] m84_88;
   assign m84_88 =10'b0;

   // m84_89 = W*in
   wire signed [9:0] m84_89;
   assign m84_89 =10'b0;

   // m84_90 = W*in
   wire signed [9:0] m84_90;
   assign m84_90 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_91 = W*in
   wire signed [9:0] m84_91;
   assign m84_91 =10'b0;

   // m84_92 = W*in
   wire signed [9:0] m84_92;
   assign m84_92 =10'b0;

   // m84_93 = W*in
   wire signed [9:0] m84_93;
   assign m84_93 =10'b0;

   // m84_94 = W*in
   wire signed [9:0] m84_94;
   assign m84_94 =10'b0;

   // m84_95 = W*in
   wire signed [9:0] m84_95;
   assign m84_95 =10'b0;

   // m84_96 = W*in
   wire signed [9:0] m84_96;
   assign m84_96 =10'b0;

   // m84_97 = W*in
   wire signed [9:0] m84_97;
   assign m84_97 ={ {4{in84[5]}} , in84[5:0] };

   // m84_98 = W*in
   wire signed [9:0] m84_98;
   assign m84_98 =10'b0;

   // m84_99 = W*in
   wire signed [9:0] m84_99;
   assign m84_99 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_100 = W*in
   wire signed [9:0] m84_100;
   assign m84_100 =10'b0;

   // m84_101 = W*in
   wire signed [9:0] m84_101;
   assign m84_101 =10'b0;

   // m84_102 = W*in
   wire signed [9:0] m84_102;
   assign m84_102 =10'b0;

   // m84_103 = W*in
   wire signed [9:0] m84_103;
   assign m84_103 =10'b0;

   // m84_104 = W*in
   wire signed [9:0] m84_104;
   assign m84_104 =10'b0;

   // m84_105 = W*in
   wire signed [9:0] m84_105;
   assign m84_105 =10'b0;

   // m84_106 = W*in
   wire signed [9:0] m84_106;
   assign m84_106 =10'b0;

   // m84_107 = W*in
   wire signed [9:0] m84_107;
   assign m84_107 =10'b0;

   // m84_108 = W*in
   wire signed [9:0] m84_108;
   assign m84_108 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_109 = W*in
   wire signed [9:0] m84_109;
   assign m84_109 ={ {4{neg84[5]}} , neg84[5:0] };

   // m84_110 = W*in
   wire signed [9:0] m84_110;
   assign m84_110 ={ {4{in84[5]}} , in84[5:0] };

   // m84_111 = W*in
   wire signed [9:0] m84_111;
   assign m84_111 =10'b0;

   // m84_112 = W*in
   wire signed [9:0] m84_112;
   assign m84_112 =10'b0;

   // m84_113 = W*in
   wire signed [9:0] m84_113;
   assign m84_113 =10'b0;

   // m84_114 = W*in
   wire signed [9:0] m84_114;
   assign m84_114 ={ {5{neg84[5]}} , neg84[5:1] };

   // m84_115 = W*in
   wire signed [9:0] m84_115;
   assign m84_115 =10'b0;

   // m84_116 = W*in
   wire signed [9:0] m84_116;
   assign m84_116 =10'b0;

   // m84_117 = W*in
   wire signed [9:0] m84_117;
   assign m84_117 =10'b0;

   // m85_1 = W*in
   wire signed [9:0] m85_1;
   assign m85_1 =10'b0;

   // m85_2 = W*in
   wire signed [9:0] m85_2;
   assign m85_2 =10'b0;

   // m85_3 = W*in
   wire signed [9:0] m85_3;
   assign m85_3 =10'b0;

   // m85_4 = W*in
   wire signed [9:0] m85_4;
   assign m85_4 =10'b0;

   // m85_5 = W*in
   wire signed [9:0] m85_5;
   assign m85_5 =10'b0;

   // m85_6 = W*in
   wire signed [9:0] m85_6;
   assign m85_6 =10'b0;

   // m85_7 = W*in
   wire signed [9:0] m85_7;
   assign m85_7 =10'b0;

   // m85_8 = W*in
   wire signed [9:0] m85_8;
   assign m85_8 =10'b0;

   // m85_9 = W*in
   wire signed [9:0] m85_9;
   assign m85_9 =10'b0;

   // m85_10 = W*in
   wire signed [9:0] m85_10;
   assign m85_10 =10'b0;

   // m85_11 = W*in
   wire signed [9:0] m85_11;
   assign m85_11 =10'b0;

   // m85_12 = W*in
   wire signed [9:0] m85_12;
   assign m85_12 =10'b0;

   // m85_13 = W*in
   wire signed [9:0] m85_13;
   assign m85_13 =10'b0;

   // m85_14 = W*in
   wire signed [9:0] m85_14;
   assign m85_14 =10'b0;

   // m85_15 = W*in
   wire signed [9:0] m85_15;
   assign m85_15 =10'b0;

   // m85_16 = W*in
   wire signed [9:0] m85_16;
   assign m85_16 =10'b0;

   // m85_17 = W*in
   wire signed [9:0] m85_17;
   assign m85_17 =10'b0;

   // m85_18 = W*in
   wire signed [9:0] m85_18;
   assign m85_18 =10'b0;

   // m85_19 = W*in
   wire signed [9:0] m85_19;
   assign m85_19 ={ {5{neg85[5]}} , neg85[5:1] };

   // m85_20 = W*in
   wire signed [9:0] m85_20;
   assign m85_20 =10'b0;

   // m85_21 = W*in
   wire signed [9:0] m85_21;
   assign m85_21 =10'b0;

   // m85_22 = W*in
   wire signed [9:0] m85_22;
   assign m85_22 =10'b0;

   // m85_23 = W*in
   wire signed [9:0] m85_23;
   assign m85_23 =10'b0;

   // m85_24 = W*in
   wire signed [9:0] m85_24;
   assign m85_24 =10'b0;

   // m85_25 = W*in
   wire signed [9:0] m85_25;
   assign m85_25 =10'b0;

   // m85_26 = W*in
   wire signed [9:0] m85_26;
   assign m85_26 =10'b0;

   // m85_27 = W*in
   wire signed [9:0] m85_27;
   assign m85_27 =10'b0;

   // m85_28 = W*in
   wire signed [9:0] m85_28;
   assign m85_28 ={ {5{in85[5]}} , in85[5:1] };

   // m85_29 = W*in
   wire signed [9:0] m85_29;
   assign m85_29 ={ {5{neg85[5]}} , neg85[5:1] };

   // m85_30 = W*in
   wire signed [9:0] m85_30;
   assign m85_30 =10'b0;

   // m85_31 = W*in
   wire signed [9:0] m85_31;
   assign m85_31 =10'b0;

   // m85_32 = W*in
   wire signed [9:0] m85_32;
   assign m85_32 =10'b0;

   // m85_33 = W*in
   wire signed [9:0] m85_33;
   assign m85_33 =10'b0;

   // m85_34 = W*in
   wire signed [9:0] m85_34;
   assign m85_34 =10'b0;

   // m85_35 = W*in
   wire signed [9:0] m85_35;
   assign m85_35 =10'b0;

   // m85_36 = W*in
   wire signed [9:0] m85_36;
   assign m85_36 ={ {5{in85[5]}} , in85[5:1] };

   // m85_37 = W*in
   wire signed [9:0] m85_37;
   assign m85_37 =10'b0;

   // m85_38 = W*in
   wire signed [9:0] m85_38;
   assign m85_38 =10'b0;

   // m85_39 = W*in
   wire signed [9:0] m85_39;
   assign m85_39 =10'b0;

   // m85_40 = W*in
   wire signed [9:0] m85_40;
   assign m85_40 =10'b0;

   // m85_41 = W*in
   wire signed [9:0] m85_41;
   assign m85_41 =10'b0;

   // m85_42 = W*in
   wire signed [9:0] m85_42;
   assign m85_42 =10'b0;

   // m85_43 = W*in
   wire signed [9:0] m85_43;
   assign m85_43 =10'b0;

   // m85_44 = W*in
   wire signed [9:0] m85_44;
   assign m85_44 =10'b0;

   // m85_45 = W*in
   wire signed [9:0] m85_45;
   assign m85_45 =10'b0;

   // m85_46 = W*in
   wire signed [9:0] m85_46;
   assign m85_46 =10'b0;

   // m85_47 = W*in
   wire signed [9:0] m85_47;
   assign m85_47 =10'b0;

   // m85_48 = W*in
   wire signed [9:0] m85_48;
   assign m85_48 =10'b0;

   // m85_49 = W*in
   wire signed [9:0] m85_49;
   assign m85_49 =10'b0;

   // m85_50 = W*in
   wire signed [9:0] m85_50;
   assign m85_50 =10'b0;

   // m85_51 = W*in
   wire signed [9:0] m85_51;
   assign m85_51 =10'b0;

   // m85_52 = W*in
   wire signed [9:0] m85_52;
   assign m85_52 =10'b0;

   // m85_53 = W*in
   wire signed [9:0] m85_53;
   assign m85_53 =10'b0;

   // m85_54 = W*in
   wire signed [9:0] m85_54;
   assign m85_54 =10'b0;

   // m85_55 = W*in
   wire signed [9:0] m85_55;
   assign m85_55 =10'b0;

   // m85_56 = W*in
   wire signed [9:0] m85_56;
   assign m85_56 =10'b0;

   // m85_57 = W*in
   wire signed [9:0] m85_57;
   assign m85_57 =10'b0;

   // m85_58 = W*in
   wire signed [9:0] m85_58;
   assign m85_58 =10'b0;

   // m85_59 = W*in
   wire signed [9:0] m85_59;
   assign m85_59 =10'b0;

   // m85_60 = W*in
   wire signed [9:0] m85_60;
   assign m85_60 =10'b0;

   // m85_61 = W*in
   wire signed [9:0] m85_61;
   assign m85_61 =10'b0;

   // m85_62 = W*in
   wire signed [9:0] m85_62;
   assign m85_62 =10'b0;

   // m85_63 = W*in
   wire signed [9:0] m85_63;
   assign m85_63 =10'b0;

   // m85_64 = W*in
   wire signed [9:0] m85_64;
   assign m85_64 ={ {5{in85[5]}} , in85[5:1] };

   // m85_65 = W*in
   wire signed [9:0] m85_65;
   assign m85_65 =10'b0;

   // m85_66 = W*in
   wire signed [9:0] m85_66;
   assign m85_66 ={ {5{in85[5]}} , in85[5:1] };

   // m85_67 = W*in
   wire signed [9:0] m85_67;
   assign m85_67 ={ {4{neg85[5]}} , neg85[5:0] };

   // m85_68 = W*in
   wire signed [9:0] m85_68;
   assign m85_68 =10'b0;

   // m85_69 = W*in
   wire signed [9:0] m85_69;
   assign m85_69 ={ {5{neg85[5]}} , neg85[5:1] };

   // m85_70 = W*in
   wire signed [9:0] m85_70;
   assign m85_70 =10'b0;

   // m85_71 = W*in
   wire signed [9:0] m85_71;
   assign m85_71 ={ {5{in85[5]}} , in85[5:1] };

   // m85_72 = W*in
   wire signed [9:0] m85_72;
   assign m85_72 ={ {5{in85[5]}} , in85[5:1] };

   // m85_73 = W*in
   wire signed [9:0] m85_73;
   assign m85_73 =10'b0;

   // m85_74 = W*in
   wire signed [9:0] m85_74;
   assign m85_74 =10'b0;

   // m85_75 = W*in
   wire signed [9:0] m85_75;
   assign m85_75 =10'b0;

   // m85_76 = W*in
   wire signed [9:0] m85_76;
   assign m85_76 =10'b0;

   // m85_77 = W*in
   wire signed [9:0] m85_77;
   assign m85_77 =10'b0;

   // m85_78 = W*in
   wire signed [9:0] m85_78;
   assign m85_78 =10'b0;

   // m85_79 = W*in
   wire signed [9:0] m85_79;
   assign m85_79 =10'b0;

   // m85_80 = W*in
   wire signed [9:0] m85_80;
   assign m85_80 =10'b0;

   // m85_81 = W*in
   wire signed [9:0] m85_81;
   assign m85_81 ={ {5{in85[5]}} , in85[5:1] };

   // m85_82 = W*in
   wire signed [9:0] m85_82;
   assign m85_82 ={ {5{neg85[5]}} , neg85[5:1] };

   // m85_83 = W*in
   wire signed [9:0] m85_83;
   assign m85_83 =10'b0;

   // m85_84 = W*in
   wire signed [9:0] m85_84;
   assign m85_84 =10'b0;

   // m85_85 = W*in
   wire signed [9:0] m85_85;
   assign m85_85 =10'b0;

   // m85_86 = W*in
   wire signed [9:0] m85_86;
   assign m85_86 =10'b0;

   // m85_87 = W*in
   wire signed [9:0] m85_87;
   assign m85_87 =10'b0;

   // m85_88 = W*in
   wire signed [9:0] m85_88;
   assign m85_88 =10'b0;

   // m85_89 = W*in
   wire signed [9:0] m85_89;
   assign m85_89 =10'b0;

   // m85_90 = W*in
   wire signed [9:0] m85_90;
   assign m85_90 =10'b0;

   // m85_91 = W*in
   wire signed [9:0] m85_91;
   assign m85_91 =10'b0;

   // m85_92 = W*in
   wire signed [9:0] m85_92;
   assign m85_92 =10'b0;

   // m85_93 = W*in
   wire signed [9:0] m85_93;
   assign m85_93 ={ {4{neg85[5]}} , neg85[5:0] };

   // m85_94 = W*in
   wire signed [9:0] m85_94;
   assign m85_94 =10'b0;

   // m85_95 = W*in
   wire signed [9:0] m85_95;
   assign m85_95 =10'b0;

   // m85_96 = W*in
   wire signed [9:0] m85_96;
   assign m85_96 =10'b0;

   // m85_97 = W*in
   wire signed [9:0] m85_97;
   assign m85_97 =10'b0;

   // m85_98 = W*in
   wire signed [9:0] m85_98;
   assign m85_98 =10'b0;

   // m85_99 = W*in
   wire signed [9:0] m85_99;
   assign m85_99 =10'b0;

   // m85_100 = W*in
   wire signed [9:0] m85_100;
   assign m85_100 =10'b0;

   // m85_101 = W*in
   wire signed [9:0] m85_101;
   assign m85_101 =10'b0;

   // m85_102 = W*in
   wire signed [9:0] m85_102;
   assign m85_102 =10'b0;

   // m85_103 = W*in
   wire signed [9:0] m85_103;
   assign m85_103 =10'b0;

   // m85_104 = W*in
   wire signed [9:0] m85_104;
   assign m85_104 =10'b0;

   // m85_105 = W*in
   wire signed [9:0] m85_105;
   assign m85_105 =10'b0;

   // m85_106 = W*in
   wire signed [9:0] m85_106;
   assign m85_106 =10'b0;

   // m85_107 = W*in
   wire signed [9:0] m85_107;
   assign m85_107 =10'b0;

   // m85_108 = W*in
   wire signed [9:0] m85_108;
   assign m85_108 =10'b0;

   // m85_109 = W*in
   wire signed [9:0] m85_109;
   assign m85_109 =10'b0;

   // m85_110 = W*in
   wire signed [9:0] m85_110;
   assign m85_110 =10'b0;

   // m85_111 = W*in
   wire signed [9:0] m85_111;
   assign m85_111 =10'b0;

   // m85_112 = W*in
   wire signed [9:0] m85_112;
   assign m85_112 =10'b0;

   // m85_113 = W*in
   wire signed [9:0] m85_113;
   assign m85_113 =10'b0;

   // m85_114 = W*in
   wire signed [9:0] m85_114;
   assign m85_114 =10'b0;

   // m85_115 = W*in
   wire signed [9:0] m85_115;
   assign m85_115 =10'b0;

   // m85_116 = W*in
   wire signed [9:0] m85_116;
   assign m85_116 =10'b0;

   // m85_117 = W*in
   wire signed [9:0] m85_117;
   assign m85_117 =10'b0;

   // m86_1 = W*in
   wire signed [9:0] m86_1;
   assign m86_1 =10'b0;

   // m86_2 = W*in
   wire signed [9:0] m86_2;
   assign m86_2 =10'b0;

   // m86_3 = W*in
   wire signed [9:0] m86_3;
   assign m86_3 =10'b0;

   // m86_4 = W*in
   wire signed [9:0] m86_4;
   assign m86_4 =10'b0;

   // m86_5 = W*in
   wire signed [9:0] m86_5;
   assign m86_5 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_6 = W*in
   wire signed [9:0] m86_6;
   assign m86_6 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_7 = W*in
   wire signed [9:0] m86_7;
   assign m86_7 =10'b0;

   // m86_8 = W*in
   wire signed [9:0] m86_8;
   assign m86_8 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_9 = W*in
   wire signed [9:0] m86_9;
   assign m86_9 =10'b0;

   // m86_10 = W*in
   wire signed [9:0] m86_10;
   assign m86_10 =10'b0;

   // m86_11 = W*in
   wire signed [9:0] m86_11;
   assign m86_11 =10'b0;

   // m86_12 = W*in
   wire signed [9:0] m86_12;
   assign m86_12 ={ {4{in86[5]}} , in86[5:0] };

   // m86_13 = W*in
   wire signed [9:0] m86_13;
   assign m86_13 =10'b0;

   // m86_14 = W*in
   wire signed [9:0] m86_14;
   assign m86_14 =10'b0;

   // m86_15 = W*in
   wire signed [9:0] m86_15;
   assign m86_15 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_16 = W*in
   wire signed [9:0] m86_16;
   assign m86_16 =10'b0;

   // m86_17 = W*in
   wire signed [9:0] m86_17;
   assign m86_17 ={ {4{in86[5]}} , in86[5:0] };

   // m86_18 = W*in
   wire signed [9:0] m86_18;
   assign m86_18 =10'b0;

   // m86_19 = W*in
   wire signed [9:0] m86_19;
   assign m86_19 =10'b0;

   // m86_20 = W*in
   wire signed [9:0] m86_20;
   assign m86_20 ={ {5{neg86[5]}} , neg86[5:1] };

   // m86_21 = W*in
   wire signed [9:0] m86_21;
   assign m86_21 =10'b0;

   // m86_22 = W*in
   wire signed [9:0] m86_22;
   assign m86_22 =10'b0;

   // m86_23 = W*in
   wire signed [9:0] m86_23;
   assign m86_23 =10'b0;

   // m86_24 = W*in
   wire signed [9:0] m86_24;
   assign m86_24 =10'b0;

   // m86_25 = W*in
   wire signed [9:0] m86_25;
   assign m86_25 =10'b0;

   // m86_26 = W*in
   wire signed [9:0] m86_26;
   assign m86_26 =10'b0;

   // m86_27 = W*in
   wire signed [9:0] m86_27;
   assign m86_27 =10'b0;

   // m86_28 = W*in
   wire signed [9:0] m86_28;
   assign m86_28 ={ {5{in86[5]}} , in86[5:1] };

   // m86_29 = W*in
   wire signed [9:0] m86_29;
   assign m86_29 =10'b0;

   // m86_30 = W*in
   wire signed [9:0] m86_30;
   assign m86_30 =10'b0;

   // m86_31 = W*in
   wire signed [9:0] m86_31;
   assign m86_31 ={ {5{neg86[5]}} , neg86[5:1] };

   // m86_32 = W*in
   wire signed [9:0] m86_32;
   assign m86_32 =10'b0;

   // m86_33 = W*in
   wire signed [9:0] m86_33;
   assign m86_33 =10'b0;

   // m86_34 = W*in
   wire signed [9:0] m86_34;
   assign m86_34 =10'b0;

   // m86_35 = W*in
   wire signed [9:0] m86_35;
   assign m86_35 =10'b0;

   // m86_36 = W*in
   wire signed [9:0] m86_36;
   assign m86_36 ={ {4{in86[5]}} , in86[5:0] };

   // m86_37 = W*in
   wire signed [9:0] m86_37;
   assign m86_37 =10'b0;

   // m86_38 = W*in
   wire signed [9:0] m86_38;
   assign m86_38 =10'b0;

   // m86_39 = W*in
   wire signed [9:0] m86_39;
   assign m86_39 =10'b0;

   // m86_40 = W*in
   wire signed [9:0] m86_40;
   assign m86_40 =10'b0;

   // m86_41 = W*in
   wire signed [9:0] m86_41;
   assign m86_41 =10'b0;

   // m86_42 = W*in
   wire signed [9:0] m86_42;
   assign m86_42 ={ {4{in86[5]}} , in86[5:0] };

   // m86_43 = W*in
   wire signed [9:0] m86_43;
   assign m86_43 ={ {4{in86[5]}} , in86[5:0] };

   // m86_44 = W*in
   wire signed [9:0] m86_44;
   assign m86_44 =10'b0;

   // m86_45 = W*in
   wire signed [9:0] m86_45;
   assign m86_45 =10'b0;

   // m86_46 = W*in
   wire signed [9:0] m86_46;
   assign m86_46 =10'b0;

   // m86_47 = W*in
   wire signed [9:0] m86_47;
   assign m86_47 =10'b0;

   // m86_48 = W*in
   wire signed [9:0] m86_48;
   assign m86_48 =10'b0;

   // m86_49 = W*in
   wire signed [9:0] m86_49;
   assign m86_49 =10'b0;

   // m86_50 = W*in
   wire signed [9:0] m86_50;
   assign m86_50 =10'b0;

   // m86_51 = W*in
   wire signed [9:0] m86_51;
   assign m86_51 =10'b0;

   // m86_52 = W*in
   wire signed [9:0] m86_52;
   assign m86_52 =10'b0;

   // m86_53 = W*in
   wire signed [9:0] m86_53;
   assign m86_53 =10'b0;

   // m86_54 = W*in
   wire signed [9:0] m86_54;
   assign m86_54 =10'b0;

   // m86_55 = W*in
   wire signed [9:0] m86_55;
   assign m86_55 =10'b0;

   // m86_56 = W*in
   wire signed [9:0] m86_56;
   assign m86_56 =10'b0;

   // m86_57 = W*in
   wire signed [9:0] m86_57;
   assign m86_57 =10'b0;

   // m86_58 = W*in
   wire signed [9:0] m86_58;
   assign m86_58 =10'b0;

   // m86_59 = W*in
   wire signed [9:0] m86_59;
   assign m86_59 =10'b0;

   // m86_60 = W*in
   wire signed [9:0] m86_60;
   assign m86_60 =10'b0;

   // m86_61 = W*in
   wire signed [9:0] m86_61;
   assign m86_61 ={ {4{in86[5]}} , in86[5:0] };

   // m86_62 = W*in
   wire signed [9:0] m86_62;
   assign m86_62 =10'b0;

   // m86_63 = W*in
   wire signed [9:0] m86_63;
   assign m86_63 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_64 = W*in
   wire signed [9:0] m86_64;
   assign m86_64 =10'b0;

   // m86_65 = W*in
   wire signed [9:0] m86_65;
   assign m86_65 ={ {5{in86[5]}} , in86[5:1] };

   // m86_66 = W*in
   wire signed [9:0] m86_66;
   assign m86_66 ={ {4{in86[5]}} , in86[5:0] };

   // m86_67 = W*in
   wire signed [9:0] m86_67;
   assign m86_67 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_68 = W*in
   wire signed [9:0] m86_68;
   assign m86_68 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_69 = W*in
   wire signed [9:0] m86_69;
   assign m86_69 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_70 = W*in
   wire signed [9:0] m86_70;
   assign m86_70 =10'b0;

   // m86_71 = W*in
   wire signed [9:0] m86_71;
   assign m86_71 ={ {5{in86[5]}} , in86[5:1] };

   // m86_72 = W*in
   wire signed [9:0] m86_72;
   assign m86_72 =10'b0;

   // m86_73 = W*in
   wire signed [9:0] m86_73;
   assign m86_73 ={ {5{neg86[5]}} , neg86[5:1] };

   // m86_74 = W*in
   wire signed [9:0] m86_74;
   assign m86_74 =10'b0;

   // m86_75 = W*in
   wire signed [9:0] m86_75;
   assign m86_75 ={ {5{in86[5]}} , in86[5:1] };

   // m86_76 = W*in
   wire signed [9:0] m86_76;
   assign m86_76 =10'b0;

   // m86_77 = W*in
   wire signed [9:0] m86_77;
   assign m86_77 ={ {4{in86[5]}} , in86[5:0] };

   // m86_78 = W*in
   wire signed [9:0] m86_78;
   assign m86_78 =10'b0;

   // m86_79 = W*in
   wire signed [9:0] m86_79;
   assign m86_79 =10'b0;

   // m86_80 = W*in
   wire signed [9:0] m86_80;
   assign m86_80 =10'b0;

   // m86_81 = W*in
   wire signed [9:0] m86_81;
   assign m86_81 ={ {5{in86[5]}} , in86[5:1] };

   // m86_82 = W*in
   wire signed [9:0] m86_82;
   assign m86_82 =10'b0;

   // m86_83 = W*in
   wire signed [9:0] m86_83;
   assign m86_83 ={ {5{in86[5]}} , in86[5:1] };

   // m86_84 = W*in
   wire signed [9:0] m86_84;
   assign m86_84 =10'b0;

   // m86_85 = W*in
   wire signed [9:0] m86_85;
   assign m86_85 =10'b0;

   // m86_86 = W*in
   wire signed [9:0] m86_86;
   assign m86_86 =10'b0;

   // m86_87 = W*in
   wire signed [9:0] m86_87;
   assign m86_87 =10'b0;

   // m86_88 = W*in
   wire signed [9:0] m86_88;
   assign m86_88 =10'b0;

   // m86_89 = W*in
   wire signed [9:0] m86_89;
   assign m86_89 =10'b0;

   // m86_90 = W*in
   wire signed [9:0] m86_90;
   assign m86_90 =10'b0;

   // m86_91 = W*in
   wire signed [9:0] m86_91;
   assign m86_91 =10'b0;

   // m86_92 = W*in
   wire signed [9:0] m86_92;
   assign m86_92 =10'b0;

   // m86_93 = W*in
   wire signed [9:0] m86_93;
   assign m86_93 ={ {4{neg86[5]}} , neg86[5:0] };

   // m86_94 = W*in
   wire signed [9:0] m86_94;
   assign m86_94 =10'b0;

   // m86_95 = W*in
   wire signed [9:0] m86_95;
   assign m86_95 ={ {4{in86[5]}} , in86[5:0] };

   // m86_96 = W*in
   wire signed [9:0] m86_96;
   assign m86_96 =10'b0;

   // m86_97 = W*in
   wire signed [9:0] m86_97;
   assign m86_97 ={ {4{in86[5]}} , in86[5:0] };

   // m86_98 = W*in
   wire signed [9:0] m86_98;
   assign m86_98 =10'b0;

   // m86_99 = W*in
   wire signed [9:0] m86_99;
   assign m86_99 =10'b0;

   // m86_100 = W*in
   wire signed [9:0] m86_100;
   assign m86_100 ={ {4{in86[5]}} , in86[5:0] };

   // m86_101 = W*in
   wire signed [9:0] m86_101;
   assign m86_101 =10'b0;

   // m86_102 = W*in
   wire signed [9:0] m86_102;
   assign m86_102 =10'b0;

   // m86_103 = W*in
   wire signed [9:0] m86_103;
   assign m86_103 =10'b0;

   // m86_104 = W*in
   wire signed [9:0] m86_104;
   assign m86_104 ={ {4{in86[5]}} , in86[5:0] };

   // m86_105 = W*in
   wire signed [9:0] m86_105;
   assign m86_105 =10'b0;

   // m86_106 = W*in
   wire signed [9:0] m86_106;
   assign m86_106 =10'b0;

   // m86_107 = W*in
   wire signed [9:0] m86_107;
   assign m86_107 ={ {4{in86[5]}} , in86[5:0] };

   // m86_108 = W*in
   wire signed [9:0] m86_108;
   assign m86_108 =10'b0;

   // m86_109 = W*in
   wire signed [9:0] m86_109;
   assign m86_109 =10'b0;

   // m86_110 = W*in
   wire signed [9:0] m86_110;
   assign m86_110 ={ {5{in86[5]}} , in86[5:1] };

   // m86_111 = W*in
   wire signed [9:0] m86_111;
   assign m86_111 =10'b0;

   // m86_112 = W*in
   wire signed [9:0] m86_112;
   assign m86_112 =10'b0;

   // m86_113 = W*in
   wire signed [9:0] m86_113;
   assign m86_113 =10'b0;

   // m86_114 = W*in
   wire signed [9:0] m86_114;
   assign m86_114 =10'b0;

   // m86_115 = W*in
   wire signed [9:0] m86_115;
   assign m86_115 =10'b0;

   // m86_116 = W*in
   wire signed [9:0] m86_116;
   assign m86_116 =10'b0;

   // m86_117 = W*in
   wire signed [9:0] m86_117;
   assign m86_117 =10'b0;

   // m87_1 = W*in
   wire signed [9:0] m87_1;
   assign m87_1 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_2 = W*in
   wire signed [9:0] m87_2;
   assign m87_2 ={ {4{in87[5]}} , in87[5:0] };

   // m87_3 = W*in
   wire signed [9:0] m87_3;
   assign m87_3 ={ {4{in87[5]}} , in87[5:0] };

   // m87_4 = W*in
   wire signed [9:0] m87_4;
   assign m87_4 =10'b0;

   // m87_5 = W*in
   wire signed [9:0] m87_5;
   assign m87_5 =10'b0;

   // m87_6 = W*in
   wire signed [9:0] m87_6;
   assign m87_6 =10'b0;

   // m87_7 = W*in
   wire signed [9:0] m87_7;
   assign m87_7 =10'b0;

   // m87_8 = W*in
   wire signed [9:0] m87_8;
   assign m87_8 ={ {4{in87[5]}} , in87[5:0] };

   // m87_9 = W*in
   wire signed [9:0] m87_9;
   assign m87_9 =10'b0;

   // m87_10 = W*in
   wire signed [9:0] m87_10;
   assign m87_10 =10'b0;

   // m87_11 = W*in
   wire signed [9:0] m87_11;
   assign m87_11 =10'b0;

   // m87_12 = W*in
   wire signed [9:0] m87_12;
   assign m87_12 ={ {4{in87[5]}} , in87[5:0] };

   // m87_13 = W*in
   wire signed [9:0] m87_13;
   assign m87_13 =10'b0;

   // m87_14 = W*in
   wire signed [9:0] m87_14;
   assign m87_14 ={ {4{in87[5]}} , in87[5:0] };

   // m87_15 = W*in
   wire signed [9:0] m87_15;
   assign m87_15 =10'b0;

   // m87_16 = W*in
   wire signed [9:0] m87_16;
   assign m87_16 =10'b0;

   // m87_17 = W*in
   wire signed [9:0] m87_17;
   assign m87_17 ={ {4{in87[5]}} , in87[5:0] };

   // m87_18 = W*in
   wire signed [9:0] m87_18;
   assign m87_18 ={ {4{in87[5]}} , in87[5:0] };

   // m87_19 = W*in
   wire signed [9:0] m87_19;
   assign m87_19 ={ {4{in87[5]}} , in87[5:0] };

   // m87_20 = W*in
   wire signed [9:0] m87_20;
   assign m87_20 =10'b0;

   // m87_21 = W*in
   wire signed [9:0] m87_21;
   assign m87_21 =10'b0;

   // m87_22 = W*in
   wire signed [9:0] m87_22;
   assign m87_22 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_23 = W*in
   wire signed [9:0] m87_23;
   assign m87_23 =10'b0;

   // m87_24 = W*in
   wire signed [9:0] m87_24;
   assign m87_24 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_25 = W*in
   wire signed [9:0] m87_25;
   assign m87_25 =10'b0;

   // m87_26 = W*in
   wire signed [9:0] m87_26;
   assign m87_26 ={ {4{in87[5]}} , in87[5:0] };

   // m87_27 = W*in
   wire signed [9:0] m87_27;
   assign m87_27 =10'b0;

   // m87_28 = W*in
   wire signed [9:0] m87_28;
   assign m87_28 =10'b0;

   // m87_29 = W*in
   wire signed [9:0] m87_29;
   assign m87_29 ={ {5{neg87[5]}} , neg87[5:1] };

   // m87_30 = W*in
   wire signed [9:0] m87_30;
   assign m87_30 =10'b0;

   // m87_31 = W*in
   wire signed [9:0] m87_31;
   assign m87_31 =10'b0;

   // m87_32 = W*in
   wire signed [9:0] m87_32;
   assign m87_32 =10'b0;

   // m87_33 = W*in
   wire signed [9:0] m87_33;
   assign m87_33 =10'b0;

   // m87_34 = W*in
   wire signed [9:0] m87_34;
   assign m87_34 =10'b0;

   // m87_35 = W*in
   wire signed [9:0] m87_35;
   assign m87_35 =10'b0;

   // m87_36 = W*in
   wire signed [9:0] m87_36;
   assign m87_36 ={ {4{in87[5]}} , in87[5:0] };

   // m87_37 = W*in
   wire signed [9:0] m87_37;
   assign m87_37 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_38 = W*in
   wire signed [9:0] m87_38;
   assign m87_38 =10'b0;

   // m87_39 = W*in
   wire signed [9:0] m87_39;
   assign m87_39 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_40 = W*in
   wire signed [9:0] m87_40;
   assign m87_40 =10'b0;

   // m87_41 = W*in
   wire signed [9:0] m87_41;
   assign m87_41 =10'b0;

   // m87_42 = W*in
   wire signed [9:0] m87_42;
   assign m87_42 =10'b0;

   // m87_43 = W*in
   wire signed [9:0] m87_43;
   assign m87_43 =10'b0;

   // m87_44 = W*in
   wire signed [9:0] m87_44;
   assign m87_44 =10'b0;

   // m87_45 = W*in
   wire signed [9:0] m87_45;
   assign m87_45 =10'b0;

   // m87_46 = W*in
   wire signed [9:0] m87_46;
   assign m87_46 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_47 = W*in
   wire signed [9:0] m87_47;
   assign m87_47 =10'b0;

   // m87_48 = W*in
   wire signed [9:0] m87_48;
   assign m87_48 =10'b0;

   // m87_49 = W*in
   wire signed [9:0] m87_49;
   assign m87_49 =10'b0;

   // m87_50 = W*in
   wire signed [9:0] m87_50;
   assign m87_50 =10'b0;

   // m87_51 = W*in
   wire signed [9:0] m87_51;
   assign m87_51 =10'b0;

   // m87_52 = W*in
   wire signed [9:0] m87_52;
   assign m87_52 =10'b0;

   // m87_53 = W*in
   wire signed [9:0] m87_53;
   assign m87_53 =10'b0;

   // m87_54 = W*in
   wire signed [9:0] m87_54;
   assign m87_54 =10'b0;

   // m87_55 = W*in
   wire signed [9:0] m87_55;
   assign m87_55 =10'b0;

   // m87_56 = W*in
   wire signed [9:0] m87_56;
   assign m87_56 =10'b0;

   // m87_57 = W*in
   wire signed [9:0] m87_57;
   assign m87_57 =10'b0;

   // m87_58 = W*in
   wire signed [9:0] m87_58;
   assign m87_58 =10'b0;

   // m87_59 = W*in
   wire signed [9:0] m87_59;
   assign m87_59 =10'b0;

   // m87_60 = W*in
   wire signed [9:0] m87_60;
   assign m87_60 =10'b0;

   // m87_61 = W*in
   wire signed [9:0] m87_61;
   assign m87_61 ={ {4{in87[5]}} , in87[5:0] };

   // m87_62 = W*in
   wire signed [9:0] m87_62;
   assign m87_62 =10'b0;

   // m87_63 = W*in
   wire signed [9:0] m87_63;
   assign m87_63 =10'b0;

   // m87_64 = W*in
   wire signed [9:0] m87_64;
   assign m87_64 =10'b0;

   // m87_65 = W*in
   wire signed [9:0] m87_65;
   assign m87_65 =10'b0;

   // m87_66 = W*in
   wire signed [9:0] m87_66;
   assign m87_66 =10'b0;

   // m87_67 = W*in
   wire signed [9:0] m87_67;
   assign m87_67 =10'b0;

   // m87_68 = W*in
   wire signed [9:0] m87_68;
   assign m87_68 ={ {4{in87[5]}} , in87[5:0] };

   // m87_69 = W*in
   wire signed [9:0] m87_69;
   assign m87_69 ={ {5{neg87[5]}} , neg87[5:1] };

   // m87_70 = W*in
   wire signed [9:0] m87_70;
   assign m87_70 =10'b0;

   // m87_71 = W*in
   wire signed [9:0] m87_71;
   assign m87_71 =10'b0;

   // m87_72 = W*in
   wire signed [9:0] m87_72;
   assign m87_72 =10'b0;

   // m87_73 = W*in
   wire signed [9:0] m87_73;
   assign m87_73 =10'b0;

   // m87_74 = W*in
   wire signed [9:0] m87_74;
   assign m87_74 =10'b0;

   // m87_75 = W*in
   wire signed [9:0] m87_75;
   assign m87_75 =10'b0;

   // m87_76 = W*in
   wire signed [9:0] m87_76;
   assign m87_76 =10'b0;

   // m87_77 = W*in
   wire signed [9:0] m87_77;
   assign m87_77 =10'b0;

   // m87_78 = W*in
   wire signed [9:0] m87_78;
   assign m87_78 =10'b0;

   // m87_79 = W*in
   wire signed [9:0] m87_79;
   assign m87_79 =10'b0;

   // m87_80 = W*in
   wire signed [9:0] m87_80;
   assign m87_80 =10'b0;

   // m87_81 = W*in
   wire signed [9:0] m87_81;
   assign m87_81 ={ {5{in87[5]}} , in87[5:1] };

   // m87_82 = W*in
   wire signed [9:0] m87_82;
   assign m87_82 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_83 = W*in
   wire signed [9:0] m87_83;
   assign m87_83 =10'b0;

   // m87_84 = W*in
   wire signed [9:0] m87_84;
   assign m87_84 =10'b0;

   // m87_85 = W*in
   wire signed [9:0] m87_85;
   assign m87_85 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_86 = W*in
   wire signed [9:0] m87_86;
   assign m87_86 =10'b0;

   // m87_87 = W*in
   wire signed [9:0] m87_87;
   assign m87_87 =10'b0;

   // m87_88 = W*in
   wire signed [9:0] m87_88;
   assign m87_88 =10'b0;

   // m87_89 = W*in
   wire signed [9:0] m87_89;
   assign m87_89 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_90 = W*in
   wire signed [9:0] m87_90;
   assign m87_90 =10'b0;

   // m87_91 = W*in
   wire signed [9:0] m87_91;
   assign m87_91 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_92 = W*in
   wire signed [9:0] m87_92;
   assign m87_92 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_93 = W*in
   wire signed [9:0] m87_93;
   assign m87_93 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_94 = W*in
   wire signed [9:0] m87_94;
   assign m87_94 ={ {4{in87[5]}} , in87[5:0] };

   // m87_95 = W*in
   wire signed [9:0] m87_95;
   assign m87_95 =10'b0;

   // m87_96 = W*in
   wire signed [9:0] m87_96;
   assign m87_96 =10'b0;

   // m87_97 = W*in
   wire signed [9:0] m87_97;
   assign m87_97 =10'b0;

   // m87_98 = W*in
   wire signed [9:0] m87_98;
   assign m87_98 =10'b0;

   // m87_99 = W*in
   wire signed [9:0] m87_99;
   assign m87_99 =10'b0;

   // m87_100 = W*in
   wire signed [9:0] m87_100;
   assign m87_100 =10'b0;

   // m87_101 = W*in
   wire signed [9:0] m87_101;
   assign m87_101 =10'b0;

   // m87_102 = W*in
   wire signed [9:0] m87_102;
   assign m87_102 =10'b0;

   // m87_103 = W*in
   wire signed [9:0] m87_103;
   assign m87_103 =10'b0;

   // m87_104 = W*in
   wire signed [9:0] m87_104;
   assign m87_104 =10'b0;

   // m87_105 = W*in
   wire signed [9:0] m87_105;
   assign m87_105 =10'b0;

   // m87_106 = W*in
   wire signed [9:0] m87_106;
   assign m87_106 =10'b0;

   // m87_107 = W*in
   wire signed [9:0] m87_107;
   assign m87_107 ={ {4{in87[5]}} , in87[5:0] };

   // m87_108 = W*in
   wire signed [9:0] m87_108;
   assign m87_108 =10'b0;

   // m87_109 = W*in
   wire signed [9:0] m87_109;
   assign m87_109 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_110 = W*in
   wire signed [9:0] m87_110;
   assign m87_110 =10'b0;

   // m87_111 = W*in
   wire signed [9:0] m87_111;
   assign m87_111 =10'b0;

   // m87_112 = W*in
   wire signed [9:0] m87_112;
   assign m87_112 =10'b0;

   // m87_113 = W*in
   wire signed [9:0] m87_113;
   assign m87_113 ={ {4{neg87[5]}} , neg87[5:0] };

   // m87_114 = W*in
   wire signed [9:0] m87_114;
   assign m87_114 ={ {5{neg87[5]}} , neg87[5:1] };

   // m87_115 = W*in
   wire signed [9:0] m87_115;
   assign m87_115 =10'b0;

   // m87_116 = W*in
   wire signed [9:0] m87_116;
   assign m87_116 =10'b0;

   // m87_117 = W*in
   wire signed [9:0] m87_117;
   assign m87_117 =10'b0;

   // m88_1 = W*in
   wire signed [9:0] m88_1;
   assign m88_1 =10'b0;

   // m88_2 = W*in
   wire signed [9:0] m88_2;
   assign m88_2 ={ {4{in88[5]}} , in88[5:0] };

   // m88_3 = W*in
   wire signed [9:0] m88_3;
   assign m88_3 =10'b0;

   // m88_4 = W*in
   wire signed [9:0] m88_4;
   assign m88_4 =10'b0;

   // m88_5 = W*in
   wire signed [9:0] m88_5;
   assign m88_5 =10'b0;

   // m88_6 = W*in
   wire signed [9:0] m88_6;
   assign m88_6 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_7 = W*in
   wire signed [9:0] m88_7;
   assign m88_7 ={ {4{in88[5]}} , in88[5:0] };

   // m88_8 = W*in
   wire signed [9:0] m88_8;
   assign m88_8 ={ {4{in88[5]}} , in88[5:0] };

   // m88_9 = W*in
   wire signed [9:0] m88_9;
   assign m88_9 =10'b0;

   // m88_10 = W*in
   wire signed [9:0] m88_10;
   assign m88_10 =10'b0;

   // m88_11 = W*in
   wire signed [9:0] m88_11;
   assign m88_11 =10'b0;

   // m88_12 = W*in
   wire signed [9:0] m88_12;
   assign m88_12 ={ {4{in88[5]}} , in88[5:0] };

   // m88_13 = W*in
   wire signed [9:0] m88_13;
   assign m88_13 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_14 = W*in
   wire signed [9:0] m88_14;
   assign m88_14 =10'b0;

   // m88_15 = W*in
   wire signed [9:0] m88_15;
   assign m88_15 =10'b0;

   // m88_16 = W*in
   wire signed [9:0] m88_16;
   assign m88_16 =10'b0;

   // m88_17 = W*in
   wire signed [9:0] m88_17;
   assign m88_17 ={ {5{in88[5]}} , in88[5:1] };

   // m88_18 = W*in
   wire signed [9:0] m88_18;
   assign m88_18 =10'b0;

   // m88_19 = W*in
   wire signed [9:0] m88_19;
   assign m88_19 ={ {4{in88[5]}} , in88[5:0] };

   // m88_20 = W*in
   wire signed [9:0] m88_20;
   assign m88_20 =10'b0;

   // m88_21 = W*in
   wire signed [9:0] m88_21;
   assign m88_21 =10'b0;

   // m88_22 = W*in
   wire signed [9:0] m88_22;
   assign m88_22 ={ {5{neg88[5]}} , neg88[5:1] };

   // m88_23 = W*in
   wire signed [9:0] m88_23;
   assign m88_23 =10'b0;

   // m88_24 = W*in
   wire signed [9:0] m88_24;
   assign m88_24 =10'b0;

   // m88_25 = W*in
   wire signed [9:0] m88_25;
   assign m88_25 =10'b0;

   // m88_26 = W*in
   wire signed [9:0] m88_26;
   assign m88_26 ={ {5{neg88[5]}} , neg88[5:1] };

   // m88_27 = W*in
   wire signed [9:0] m88_27;
   assign m88_27 =10'b0;

   // m88_28 = W*in
   wire signed [9:0] m88_28;
   assign m88_28 ={ {5{in88[5]}} , in88[5:1] };

   // m88_29 = W*in
   wire signed [9:0] m88_29;
   assign m88_29 =10'b0;

   // m88_30 = W*in
   wire signed [9:0] m88_30;
   assign m88_30 =10'b0;

   // m88_31 = W*in
   wire signed [9:0] m88_31;
   assign m88_31 =10'b0;

   // m88_32 = W*in
   wire signed [9:0] m88_32;
   assign m88_32 =10'b0;

   // m88_33 = W*in
   wire signed [9:0] m88_33;
   assign m88_33 =10'b0;

   // m88_34 = W*in
   wire signed [9:0] m88_34;
   assign m88_34 =10'b0;

   // m88_35 = W*in
   wire signed [9:0] m88_35;
   assign m88_35 =10'b0;

   // m88_36 = W*in
   wire signed [9:0] m88_36;
   assign m88_36 ={ {4{in88[5]}} , in88[5:0] };

   // m88_37 = W*in
   wire signed [9:0] m88_37;
   assign m88_37 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_38 = W*in
   wire signed [9:0] m88_38;
   assign m88_38 =10'b0;

   // m88_39 = W*in
   wire signed [9:0] m88_39;
   assign m88_39 =10'b0;

   // m88_40 = W*in
   wire signed [9:0] m88_40;
   assign m88_40 =10'b0;

   // m88_41 = W*in
   wire signed [9:0] m88_41;
   assign m88_41 =10'b0;

   // m88_42 = W*in
   wire signed [9:0] m88_42;
   assign m88_42 =10'b0;

   // m88_43 = W*in
   wire signed [9:0] m88_43;
   assign m88_43 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_44 = W*in
   wire signed [9:0] m88_44;
   assign m88_44 =10'b0;

   // m88_45 = W*in
   wire signed [9:0] m88_45;
   assign m88_45 =10'b0;

   // m88_46 = W*in
   wire signed [9:0] m88_46;
   assign m88_46 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_47 = W*in
   wire signed [9:0] m88_47;
   assign m88_47 =10'b0;

   // m88_48 = W*in
   wire signed [9:0] m88_48;
   assign m88_48 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_49 = W*in
   wire signed [9:0] m88_49;
   assign m88_49 =10'b0;

   // m88_50 = W*in
   wire signed [9:0] m88_50;
   assign m88_50 =10'b0;

   // m88_51 = W*in
   wire signed [9:0] m88_51;
   assign m88_51 =10'b0;

   // m88_52 = W*in
   wire signed [9:0] m88_52;
   assign m88_52 =10'b0;

   // m88_53 = W*in
   wire signed [9:0] m88_53;
   assign m88_53 ={ {4{in88[5]}} , in88[5:0] };

   // m88_54 = W*in
   wire signed [9:0] m88_54;
   assign m88_54 =10'b0;

   // m88_55 = W*in
   wire signed [9:0] m88_55;
   assign m88_55 =10'b0;

   // m88_56 = W*in
   wire signed [9:0] m88_56;
   assign m88_56 =10'b0;

   // m88_57 = W*in
   wire signed [9:0] m88_57;
   assign m88_57 =10'b0;

   // m88_58 = W*in
   wire signed [9:0] m88_58;
   assign m88_58 =10'b0;

   // m88_59 = W*in
   wire signed [9:0] m88_59;
   assign m88_59 =10'b0;

   // m88_60 = W*in
   wire signed [9:0] m88_60;
   assign m88_60 =10'b0;

   // m88_61 = W*in
   wire signed [9:0] m88_61;
   assign m88_61 =10'b0;

   // m88_62 = W*in
   wire signed [9:0] m88_62;
   assign m88_62 =10'b0;

   // m88_63 = W*in
   wire signed [9:0] m88_63;
   assign m88_63 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_64 = W*in
   wire signed [9:0] m88_64;
   assign m88_64 =10'b0;

   // m88_65 = W*in
   wire signed [9:0] m88_65;
   assign m88_65 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_66 = W*in
   wire signed [9:0] m88_66;
   assign m88_66 =10'b0;

   // m88_67 = W*in
   wire signed [9:0] m88_67;
   assign m88_67 =10'b0;

   // m88_68 = W*in
   wire signed [9:0] m88_68;
   assign m88_68 =10'b0;

   // m88_69 = W*in
   wire signed [9:0] m88_69;
   assign m88_69 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_70 = W*in
   wire signed [9:0] m88_70;
   assign m88_70 =10'b0;

   // m88_71 = W*in
   wire signed [9:0] m88_71;
   assign m88_71 ={ {4{in88[5]}} , in88[5:0] };

   // m88_72 = W*in
   wire signed [9:0] m88_72;
   assign m88_72 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_73 = W*in
   wire signed [9:0] m88_73;
   assign m88_73 ={ {4{in88[5]}} , in88[5:0] };

   // m88_74 = W*in
   wire signed [9:0] m88_74;
   assign m88_74 =10'b0;

   // m88_75 = W*in
   wire signed [9:0] m88_75;
   assign m88_75 =10'b0;

   // m88_76 = W*in
   wire signed [9:0] m88_76;
   assign m88_76 =10'b0;

   // m88_77 = W*in
   wire signed [9:0] m88_77;
   assign m88_77 =10'b0;

   // m88_78 = W*in
   wire signed [9:0] m88_78;
   assign m88_78 =10'b0;

   // m88_79 = W*in
   wire signed [9:0] m88_79;
   assign m88_79 =10'b0;

   // m88_80 = W*in
   wire signed [9:0] m88_80;
   assign m88_80 ={ {5{in88[5]}} , in88[5:1] };

   // m88_81 = W*in
   wire signed [9:0] m88_81;
   assign m88_81 =10'b0;

   // m88_82 = W*in
   wire signed [9:0] m88_82;
   assign m88_82 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_83 = W*in
   wire signed [9:0] m88_83;
   assign m88_83 ={ {5{neg88[5]}} , neg88[5:1] };

   // m88_84 = W*in
   wire signed [9:0] m88_84;
   assign m88_84 =10'b0;

   // m88_85 = W*in
   wire signed [9:0] m88_85;
   assign m88_85 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_86 = W*in
   wire signed [9:0] m88_86;
   assign m88_86 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_87 = W*in
   wire signed [9:0] m88_87;
   assign m88_87 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_88 = W*in
   wire signed [9:0] m88_88;
   assign m88_88 ={ {4{in88[5]}} , in88[5:0] };

   // m88_89 = W*in
   wire signed [9:0] m88_89;
   assign m88_89 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_90 = W*in
   wire signed [9:0] m88_90;
   assign m88_90 =10'b0;

   // m88_91 = W*in
   wire signed [9:0] m88_91;
   assign m88_91 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_92 = W*in
   wire signed [9:0] m88_92;
   assign m88_92 =10'b0;

   // m88_93 = W*in
   wire signed [9:0] m88_93;
   assign m88_93 =10'b0;

   // m88_94 = W*in
   wire signed [9:0] m88_94;
   assign m88_94 =10'b0;

   // m88_95 = W*in
   wire signed [9:0] m88_95;
   assign m88_95 =10'b0;

   // m88_96 = W*in
   wire signed [9:0] m88_96;
   assign m88_96 =10'b0;

   // m88_97 = W*in
   wire signed [9:0] m88_97;
   assign m88_97 =10'b0;

   // m88_98 = W*in
   wire signed [9:0] m88_98;
   assign m88_98 =10'b0;

   // m88_99 = W*in
   wire signed [9:0] m88_99;
   assign m88_99 =10'b0;

   // m88_100 = W*in
   wire signed [9:0] m88_100;
   assign m88_100 =10'b0;

   // m88_101 = W*in
   wire signed [9:0] m88_101;
   assign m88_101 =10'b0;

   // m88_102 = W*in
   wire signed [9:0] m88_102;
   assign m88_102 =10'b0;

   // m88_103 = W*in
   wire signed [9:0] m88_103;
   assign m88_103 =10'b0;

   // m88_104 = W*in
   wire signed [9:0] m88_104;
   assign m88_104 =10'b0;

   // m88_105 = W*in
   wire signed [9:0] m88_105;
   assign m88_105 =10'b0;

   // m88_106 = W*in
   wire signed [9:0] m88_106;
   assign m88_106 ={ {4{in88[5]}} , in88[5:0] };

   // m88_107 = W*in
   wire signed [9:0] m88_107;
   assign m88_107 =10'b0;

   // m88_108 = W*in
   wire signed [9:0] m88_108;
   assign m88_108 =10'b0;

   // m88_109 = W*in
   wire signed [9:0] m88_109;
   assign m88_109 ={ {4{neg88[5]}} , neg88[5:0] };

   // m88_110 = W*in
   wire signed [9:0] m88_110;
   assign m88_110 =10'b0;

   // m88_111 = W*in
   wire signed [9:0] m88_111;
   assign m88_111 =10'b0;

   // m88_112 = W*in
   wire signed [9:0] m88_112;
   assign m88_112 =10'b0;

   // m88_113 = W*in
   wire signed [9:0] m88_113;
   assign m88_113 =10'b0;

   // m88_114 = W*in
   wire signed [9:0] m88_114;
   assign m88_114 =10'b0;

   // m88_115 = W*in
   wire signed [9:0] m88_115;
   assign m88_115 =10'b0;

   // m88_116 = W*in
   wire signed [9:0] m88_116;
   assign m88_116 =10'b0;

   // m88_117 = W*in
   wire signed [9:0] m88_117;
   assign m88_117 =10'b0;

   // m89_1 = W*in
   wire signed [9:0] m89_1;
   assign m89_1 =10'b0;

   // m89_2 = W*in
   wire signed [9:0] m89_2;
   assign m89_2 =10'b0;

   // m89_3 = W*in
   wire signed [9:0] m89_3;
   assign m89_3 =10'b0;

   // m89_4 = W*in
   wire signed [9:0] m89_4;
   assign m89_4 =10'b0;

   // m89_5 = W*in
   wire signed [9:0] m89_5;
   assign m89_5 =10'b0;

   // m89_6 = W*in
   wire signed [9:0] m89_6;
   assign m89_6 =10'b0;

   // m89_7 = W*in
   wire signed [9:0] m89_7;
   assign m89_7 =10'b0;

   // m89_8 = W*in
   wire signed [9:0] m89_8;
   assign m89_8 =10'b0;

   // m89_9 = W*in
   wire signed [9:0] m89_9;
   assign m89_9 =10'b0;

   // m89_10 = W*in
   wire signed [9:0] m89_10;
   assign m89_10 =10'b0;

   // m89_11 = W*in
   wire signed [9:0] m89_11;
   assign m89_11 =10'b0;

   // m89_12 = W*in
   wire signed [9:0] m89_12;
   assign m89_12 =10'b0;

   // m89_13 = W*in
   wire signed [9:0] m89_13;
   assign m89_13 =10'b0;

   // m89_14 = W*in
   wire signed [9:0] m89_14;
   assign m89_14 =10'b0;

   // m89_15 = W*in
   wire signed [9:0] m89_15;
   assign m89_15 =10'b0;

   // m89_16 = W*in
   wire signed [9:0] m89_16;
   assign m89_16 =10'b0;

   // m89_17 = W*in
   wire signed [9:0] m89_17;
   assign m89_17 ={ {5{in89[5]}} , in89[5:1] };

   // m89_18 = W*in
   wire signed [9:0] m89_18;
   assign m89_18 =10'b0;

   // m89_19 = W*in
   wire signed [9:0] m89_19;
   assign m89_19 =10'b0;

   // m89_20 = W*in
   wire signed [9:0] m89_20;
   assign m89_20 =10'b0;

   // m89_21 = W*in
   wire signed [9:0] m89_21;
   assign m89_21 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_22 = W*in
   wire signed [9:0] m89_22;
   assign m89_22 =10'b0;

   // m89_23 = W*in
   wire signed [9:0] m89_23;
   assign m89_23 =10'b0;

   // m89_24 = W*in
   wire signed [9:0] m89_24;
   assign m89_24 =10'b0;

   // m89_25 = W*in
   wire signed [9:0] m89_25;
   assign m89_25 =10'b0;

   // m89_26 = W*in
   wire signed [9:0] m89_26;
   assign m89_26 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_27 = W*in
   wire signed [9:0] m89_27;
   assign m89_27 ={ {4{in89[5]}} , in89[5:0] };

   // m89_28 = W*in
   wire signed [9:0] m89_28;
   assign m89_28 ={ {5{in89[5]}} , in89[5:1] };

   // m89_29 = W*in
   wire signed [9:0] m89_29;
   assign m89_29 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_30 = W*in
   wire signed [9:0] m89_30;
   assign m89_30 =10'b0;

   // m89_31 = W*in
   wire signed [9:0] m89_31;
   assign m89_31 ={ {5{in89[5]}} , in89[5:1] };

   // m89_32 = W*in
   wire signed [9:0] m89_32;
   assign m89_32 =10'b0;

   // m89_33 = W*in
   wire signed [9:0] m89_33;
   assign m89_33 =10'b0;

   // m89_34 = W*in
   wire signed [9:0] m89_34;
   assign m89_34 =10'b0;

   // m89_35 = W*in
   wire signed [9:0] m89_35;
   assign m89_35 ={ {5{in89[5]}} , in89[5:1] };

   // m89_36 = W*in
   wire signed [9:0] m89_36;
   assign m89_36 =10'b0;

   // m89_37 = W*in
   wire signed [9:0] m89_37;
   assign m89_37 =10'b0;

   // m89_38 = W*in
   wire signed [9:0] m89_38;
   assign m89_38 =10'b0;

   // m89_39 = W*in
   wire signed [9:0] m89_39;
   assign m89_39 =10'b0;

   // m89_40 = W*in
   wire signed [9:0] m89_40;
   assign m89_40 =10'b0;

   // m89_41 = W*in
   wire signed [9:0] m89_41;
   assign m89_41 =10'b0;

   // m89_42 = W*in
   wire signed [9:0] m89_42;
   assign m89_42 =10'b0;

   // m89_43 = W*in
   wire signed [9:0] m89_43;
   assign m89_43 =10'b0;

   // m89_44 = W*in
   wire signed [9:0] m89_44;
   assign m89_44 =10'b0;

   // m89_45 = W*in
   wire signed [9:0] m89_45;
   assign m89_45 =10'b0;

   // m89_46 = W*in
   wire signed [9:0] m89_46;
   assign m89_46 =10'b0;

   // m89_47 = W*in
   wire signed [9:0] m89_47;
   assign m89_47 =10'b0;

   // m89_48 = W*in
   wire signed [9:0] m89_48;
   assign m89_48 =10'b0;

   // m89_49 = W*in
   wire signed [9:0] m89_49;
   assign m89_49 =10'b0;

   // m89_50 = W*in
   wire signed [9:0] m89_50;
   assign m89_50 =10'b0;

   // m89_51 = W*in
   wire signed [9:0] m89_51;
   assign m89_51 =10'b0;

   // m89_52 = W*in
   wire signed [9:0] m89_52;
   assign m89_52 =10'b0;

   // m89_53 = W*in
   wire signed [9:0] m89_53;
   assign m89_53 =10'b0;

   // m89_54 = W*in
   wire signed [9:0] m89_54;
   assign m89_54 =10'b0;

   // m89_55 = W*in
   wire signed [9:0] m89_55;
   assign m89_55 =10'b0;

   // m89_56 = W*in
   wire signed [9:0] m89_56;
   assign m89_56 =10'b0;

   // m89_57 = W*in
   wire signed [9:0] m89_57;
   assign m89_57 =10'b0;

   // m89_58 = W*in
   wire signed [9:0] m89_58;
   assign m89_58 =10'b0;

   // m89_59 = W*in
   wire signed [9:0] m89_59;
   assign m89_59 =10'b0;

   // m89_60 = W*in
   wire signed [9:0] m89_60;
   assign m89_60 ={ {4{in89[5]}} , in89[5:0] };

   // m89_61 = W*in
   wire signed [9:0] m89_61;
   assign m89_61 =10'b0;

   // m89_62 = W*in
   wire signed [9:0] m89_62;
   assign m89_62 =10'b0;

   // m89_63 = W*in
   wire signed [9:0] m89_63;
   assign m89_63 ={ {4{neg89[5]}} , neg89[5:0] };

   // m89_64 = W*in
   wire signed [9:0] m89_64;
   assign m89_64 =10'b0;

   // m89_65 = W*in
   wire signed [9:0] m89_65;
   assign m89_65 ={ {4{neg89[5]}} , neg89[5:0] };

   // m89_66 = W*in
   wire signed [9:0] m89_66;
   assign m89_66 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_67 = W*in
   wire signed [9:0] m89_67;
   assign m89_67 =10'b0;

   // m89_68 = W*in
   wire signed [9:0] m89_68;
   assign m89_68 =10'b0;

   // m89_69 = W*in
   wire signed [9:0] m89_69;
   assign m89_69 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_70 = W*in
   wire signed [9:0] m89_70;
   assign m89_70 ={ {4{neg89[5]}} , neg89[5:0] };

   // m89_71 = W*in
   wire signed [9:0] m89_71;
   assign m89_71 ={ {4{in89[5]}} , in89[5:0] };

   // m89_72 = W*in
   wire signed [9:0] m89_72;
   assign m89_72 =10'b0;

   // m89_73 = W*in
   wire signed [9:0] m89_73;
   assign m89_73 =10'b0;

   // m89_74 = W*in
   wire signed [9:0] m89_74;
   assign m89_74 =10'b0;

   // m89_75 = W*in
   wire signed [9:0] m89_75;
   assign m89_75 =10'b0;

   // m89_76 = W*in
   wire signed [9:0] m89_76;
   assign m89_76 =10'b0;

   // m89_77 = W*in
   wire signed [9:0] m89_77;
   assign m89_77 =10'b0;

   // m89_78 = W*in
   wire signed [9:0] m89_78;
   assign m89_78 =10'b0;

   // m89_79 = W*in
   wire signed [9:0] m89_79;
   assign m89_79 =10'b0;

   // m89_80 = W*in
   wire signed [9:0] m89_80;
   assign m89_80 =10'b0;

   // m89_81 = W*in
   wire signed [9:0] m89_81;
   assign m89_81 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_82 = W*in
   wire signed [9:0] m89_82;
   assign m89_82 ={ {5{neg89[5]}} , neg89[5:1] };

   // m89_83 = W*in
   wire signed [9:0] m89_83;
   assign m89_83 =10'b0;

   // m89_84 = W*in
   wire signed [9:0] m89_84;
   assign m89_84 =10'b0;

   // m89_85 = W*in
   wire signed [9:0] m89_85;
   assign m89_85 =10'b0;

   // m89_86 = W*in
   wire signed [9:0] m89_86;
   assign m89_86 ={ {4{neg89[5]}} , neg89[5:0] };

   // m89_87 = W*in
   wire signed [9:0] m89_87;
   assign m89_87 =10'b0;

   // m89_88 = W*in
   wire signed [9:0] m89_88;
   assign m89_88 =10'b0;

   // m89_89 = W*in
   wire signed [9:0] m89_89;
   assign m89_89 =10'b0;

   // m89_90 = W*in
   wire signed [9:0] m89_90;
   assign m89_90 =10'b0;

   // m89_91 = W*in
   wire signed [9:0] m89_91;
   assign m89_91 =10'b0;

   // m89_92 = W*in
   wire signed [9:0] m89_92;
   assign m89_92 =10'b0;

   // m89_93 = W*in
   wire signed [9:0] m89_93;
   assign m89_93 =10'b0;

   // m89_94 = W*in
   wire signed [9:0] m89_94;
   assign m89_94 =10'b0;

   // m89_95 = W*in
   wire signed [9:0] m89_95;
   assign m89_95 =10'b0;

   // m89_96 = W*in
   wire signed [9:0] m89_96;
   assign m89_96 =10'b0;

   // m89_97 = W*in
   wire signed [9:0] m89_97;
   assign m89_97 =10'b0;

   // m89_98 = W*in
   wire signed [9:0] m89_98;
   assign m89_98 =10'b0;

   // m89_99 = W*in
   wire signed [9:0] m89_99;
   assign m89_99 =10'b0;

   // m89_100 = W*in
   wire signed [9:0] m89_100;
   assign m89_100 =10'b0;

   // m89_101 = W*in
   wire signed [9:0] m89_101;
   assign m89_101 =10'b0;

   // m89_102 = W*in
   wire signed [9:0] m89_102;
   assign m89_102 =10'b0;

   // m89_103 = W*in
   wire signed [9:0] m89_103;
   assign m89_103 =10'b0;

   // m89_104 = W*in
   wire signed [9:0] m89_104;
   assign m89_104 =10'b0;

   // m89_105 = W*in
   wire signed [9:0] m89_105;
   assign m89_105 =10'b0;

   // m89_106 = W*in
   wire signed [9:0] m89_106;
   assign m89_106 =10'b0;

   // m89_107 = W*in
   wire signed [9:0] m89_107;
   assign m89_107 =10'b0;

   // m89_108 = W*in
   wire signed [9:0] m89_108;
   assign m89_108 =10'b0;

   // m89_109 = W*in
   wire signed [9:0] m89_109;
   assign m89_109 =10'b0;

   // m89_110 = W*in
   wire signed [9:0] m89_110;
   assign m89_110 =10'b0;

   // m89_111 = W*in
   wire signed [9:0] m89_111;
   assign m89_111 =10'b0;

   // m89_112 = W*in
   wire signed [9:0] m89_112;
   assign m89_112 =10'b0;

   // m89_113 = W*in
   wire signed [9:0] m89_113;
   assign m89_113 =10'b0;

   // m89_114 = W*in
   wire signed [9:0] m89_114;
   assign m89_114 =10'b0;

   // m89_115 = W*in
   wire signed [9:0] m89_115;
   assign m89_115 =10'b0;

   // m89_116 = W*in
   wire signed [9:0] m89_116;
   assign m89_116 =10'b0;

   // m89_117 = W*in
   wire signed [9:0] m89_117;
   assign m89_117 ={ {4{in89[5]}} , in89[5:0] };

   // m90_1 = W*in
   wire signed [9:0] m90_1;
   assign m90_1 =10'b0;

   // m90_2 = W*in
   wire signed [9:0] m90_2;
   assign m90_2 =10'b0;

   // m90_3 = W*in
   wire signed [9:0] m90_3;
   assign m90_3 =10'b0;

   // m90_4 = W*in
   wire signed [9:0] m90_4;
   assign m90_4 =10'b0;

   // m90_5 = W*in
   wire signed [9:0] m90_5;
   assign m90_5 =10'b0;

   // m90_6 = W*in
   wire signed [9:0] m90_6;
   assign m90_6 =10'b0;

   // m90_7 = W*in
   wire signed [9:0] m90_7;
   assign m90_7 =10'b0;

   // m90_8 = W*in
   wire signed [9:0] m90_8;
   assign m90_8 =10'b0;

   // m90_9 = W*in
   wire signed [9:0] m90_9;
   assign m90_9 =10'b0;

   // m90_10 = W*in
   wire signed [9:0] m90_10;
   assign m90_10 =10'b0;

   // m90_11 = W*in
   wire signed [9:0] m90_11;
   assign m90_11 =10'b0;

   // m90_12 = W*in
   wire signed [9:0] m90_12;
   assign m90_12 =10'b0;

   // m90_13 = W*in
   wire signed [9:0] m90_13;
   assign m90_13 =10'b0;

   // m90_14 = W*in
   wire signed [9:0] m90_14;
   assign m90_14 =10'b0;

   // m90_15 = W*in
   wire signed [9:0] m90_15;
   assign m90_15 =10'b0;

   // m90_16 = W*in
   wire signed [9:0] m90_16;
   assign m90_16 =10'b0;

   // m90_17 = W*in
   wire signed [9:0] m90_17;
   assign m90_17 =10'b0;

   // m90_18 = W*in
   wire signed [9:0] m90_18;
   assign m90_18 ={ {5{in90[5]}} , in90[5:1] };

   // m90_19 = W*in
   wire signed [9:0] m90_19;
   assign m90_19 =10'b0;

   // m90_20 = W*in
   wire signed [9:0] m90_20;
   assign m90_20 =10'b0;

   // m90_21 = W*in
   wire signed [9:0] m90_21;
   assign m90_21 ={ {5{neg90[5]}} , neg90[5:1] };

   // m90_22 = W*in
   wire signed [9:0] m90_22;
   assign m90_22 =10'b0;

   // m90_23 = W*in
   wire signed [9:0] m90_23;
   assign m90_23 =10'b0;

   // m90_24 = W*in
   wire signed [9:0] m90_24;
   assign m90_24 =10'b0;

   // m90_25 = W*in
   wire signed [9:0] m90_25;
   assign m90_25 =10'b0;

   // m90_26 = W*in
   wire signed [9:0] m90_26;
   assign m90_26 =10'b0;

   // m90_27 = W*in
   wire signed [9:0] m90_27;
   assign m90_27 =10'b0;

   // m90_28 = W*in
   wire signed [9:0] m90_28;
   assign m90_28 =10'b0;

   // m90_29 = W*in
   wire signed [9:0] m90_29;
   assign m90_29 =10'b0;

   // m90_30 = W*in
   wire signed [9:0] m90_30;
   assign m90_30 =10'b0;

   // m90_31 = W*in
   wire signed [9:0] m90_31;
   assign m90_31 =10'b0;

   // m90_32 = W*in
   wire signed [9:0] m90_32;
   assign m90_32 =10'b0;

   // m90_33 = W*in
   wire signed [9:0] m90_33;
   assign m90_33 =10'b0;

   // m90_34 = W*in
   wire signed [9:0] m90_34;
   assign m90_34 =10'b0;

   // m90_35 = W*in
   wire signed [9:0] m90_35;
   assign m90_35 =10'b0;

   // m90_36 = W*in
   wire signed [9:0] m90_36;
   assign m90_36 =10'b0;

   // m90_37 = W*in
   wire signed [9:0] m90_37;
   assign m90_37 =10'b0;

   // m90_38 = W*in
   wire signed [9:0] m90_38;
   assign m90_38 =10'b0;

   // m90_39 = W*in
   wire signed [9:0] m90_39;
   assign m90_39 =10'b0;

   // m90_40 = W*in
   wire signed [9:0] m90_40;
   assign m90_40 =10'b0;

   // m90_41 = W*in
   wire signed [9:0] m90_41;
   assign m90_41 =10'b0;

   // m90_42 = W*in
   wire signed [9:0] m90_42;
   assign m90_42 =10'b0;

   // m90_43 = W*in
   wire signed [9:0] m90_43;
   assign m90_43 =10'b0;

   // m90_44 = W*in
   wire signed [9:0] m90_44;
   assign m90_44 =10'b0;

   // m90_45 = W*in
   wire signed [9:0] m90_45;
   assign m90_45 =10'b0;

   // m90_46 = W*in
   wire signed [9:0] m90_46;
   assign m90_46 =10'b0;

   // m90_47 = W*in
   wire signed [9:0] m90_47;
   assign m90_47 =10'b0;

   // m90_48 = W*in
   wire signed [9:0] m90_48;
   assign m90_48 =10'b0;

   // m90_49 = W*in
   wire signed [9:0] m90_49;
   assign m90_49 =10'b0;

   // m90_50 = W*in
   wire signed [9:0] m90_50;
   assign m90_50 =10'b0;

   // m90_51 = W*in
   wire signed [9:0] m90_51;
   assign m90_51 =10'b0;

   // m90_52 = W*in
   wire signed [9:0] m90_52;
   assign m90_52 =10'b0;

   // m90_53 = W*in
   wire signed [9:0] m90_53;
   assign m90_53 =10'b0;

   // m90_54 = W*in
   wire signed [9:0] m90_54;
   assign m90_54 =10'b0;

   // m90_55 = W*in
   wire signed [9:0] m90_55;
   assign m90_55 =10'b0;

   // m90_56 = W*in
   wire signed [9:0] m90_56;
   assign m90_56 =10'b0;

   // m90_57 = W*in
   wire signed [9:0] m90_57;
   assign m90_57 =10'b0;

   // m90_58 = W*in
   wire signed [9:0] m90_58;
   assign m90_58 =10'b0;

   // m90_59 = W*in
   wire signed [9:0] m90_59;
   assign m90_59 =10'b0;

   // m90_60 = W*in
   wire signed [9:0] m90_60;
   assign m90_60 =10'b0;

   // m90_61 = W*in
   wire signed [9:0] m90_61;
   assign m90_61 =10'b0;

   // m90_62 = W*in
   wire signed [9:0] m90_62;
   assign m90_62 =10'b0;

   // m90_63 = W*in
   wire signed [9:0] m90_63;
   assign m90_63 =10'b0;

   // m90_64 = W*in
   wire signed [9:0] m90_64;
   assign m90_64 =10'b0;

   // m90_65 = W*in
   wire signed [9:0] m90_65;
   assign m90_65 ={ {5{neg90[5]}} , neg90[5:1] };

   // m90_66 = W*in
   wire signed [9:0] m90_66;
   assign m90_66 =10'b0;

   // m90_67 = W*in
   wire signed [9:0] m90_67;
   assign m90_67 =10'b0;

   // m90_68 = W*in
   wire signed [9:0] m90_68;
   assign m90_68 =10'b0;

   // m90_69 = W*in
   wire signed [9:0] m90_69;
   assign m90_69 =10'b0;

   // m90_70 = W*in
   wire signed [9:0] m90_70;
   assign m90_70 =10'b0;

   // m90_71 = W*in
   wire signed [9:0] m90_71;
   assign m90_71 ={ {5{in90[5]}} , in90[5:1] };

   // m90_72 = W*in
   wire signed [9:0] m90_72;
   assign m90_72 =10'b0;

   // m90_73 = W*in
   wire signed [9:0] m90_73;
   assign m90_73 =10'b0;

   // m90_74 = W*in
   wire signed [9:0] m90_74;
   assign m90_74 =10'b0;

   // m90_75 = W*in
   wire signed [9:0] m90_75;
   assign m90_75 =10'b0;

   // m90_76 = W*in
   wire signed [9:0] m90_76;
   assign m90_76 =10'b0;

   // m90_77 = W*in
   wire signed [9:0] m90_77;
   assign m90_77 =10'b0;

   // m90_78 = W*in
   wire signed [9:0] m90_78;
   assign m90_78 =10'b0;

   // m90_79 = W*in
   wire signed [9:0] m90_79;
   assign m90_79 =10'b0;

   // m90_80 = W*in
   wire signed [9:0] m90_80;
   assign m90_80 =10'b0;

   // m90_81 = W*in
   wire signed [9:0] m90_81;
   assign m90_81 ={ {5{in90[5]}} , in90[5:1] };

   // m90_82 = W*in
   wire signed [9:0] m90_82;
   assign m90_82 =10'b0;

   // m90_83 = W*in
   wire signed [9:0] m90_83;
   assign m90_83 =10'b0;

   // m90_84 = W*in
   wire signed [9:0] m90_84;
   assign m90_84 =10'b0;

   // m90_85 = W*in
   wire signed [9:0] m90_85;
   assign m90_85 =10'b0;

   // m90_86 = W*in
   wire signed [9:0] m90_86;
   assign m90_86 =10'b0;

   // m90_87 = W*in
   wire signed [9:0] m90_87;
   assign m90_87 =10'b0;

   // m90_88 = W*in
   wire signed [9:0] m90_88;
   assign m90_88 =10'b0;

   // m90_89 = W*in
   wire signed [9:0] m90_89;
   assign m90_89 =10'b0;

   // m90_90 = W*in
   wire signed [9:0] m90_90;
   assign m90_90 =10'b0;

   // m90_91 = W*in
   wire signed [9:0] m90_91;
   assign m90_91 =10'b0;

   // m90_92 = W*in
   wire signed [9:0] m90_92;
   assign m90_92 =10'b0;

   // m90_93 = W*in
   wire signed [9:0] m90_93;
   assign m90_93 =10'b0;

   // m90_94 = W*in
   wire signed [9:0] m90_94;
   assign m90_94 =10'b0;

   // m90_95 = W*in
   wire signed [9:0] m90_95;
   assign m90_95 =10'b0;

   // m90_96 = W*in
   wire signed [9:0] m90_96;
   assign m90_96 =10'b0;

   // m90_97 = W*in
   wire signed [9:0] m90_97;
   assign m90_97 =10'b0;

   // m90_98 = W*in
   wire signed [9:0] m90_98;
   assign m90_98 =10'b0;

   // m90_99 = W*in
   wire signed [9:0] m90_99;
   assign m90_99 =10'b0;

   // m90_100 = W*in
   wire signed [9:0] m90_100;
   assign m90_100 =10'b0;

   // m90_101 = W*in
   wire signed [9:0] m90_101;
   assign m90_101 =10'b0;

   // m90_102 = W*in
   wire signed [9:0] m90_102;
   assign m90_102 =10'b0;

   // m90_103 = W*in
   wire signed [9:0] m90_103;
   assign m90_103 =10'b0;

   // m90_104 = W*in
   wire signed [9:0] m90_104;
   assign m90_104 =10'b0;

   // m90_105 = W*in
   wire signed [9:0] m90_105;
   assign m90_105 =10'b0;

   // m90_106 = W*in
   wire signed [9:0] m90_106;
   assign m90_106 =10'b0;

   // m90_107 = W*in
   wire signed [9:0] m90_107;
   assign m90_107 =10'b0;

   // m90_108 = W*in
   wire signed [9:0] m90_108;
   assign m90_108 ={ {4{neg90[5]}} , neg90[5:0] };

   // m90_109 = W*in
   wire signed [9:0] m90_109;
   assign m90_109 ={ {4{neg90[5]}} , neg90[5:0] };

   // m90_110 = W*in
   wire signed [9:0] m90_110;
   assign m90_110 =10'b0;

   // m90_111 = W*in
   wire signed [9:0] m90_111;
   assign m90_111 =10'b0;

   // m90_112 = W*in
   wire signed [9:0] m90_112;
   assign m90_112 =10'b0;

   // m90_113 = W*in
   wire signed [9:0] m90_113;
   assign m90_113 =10'b0;

   // m90_114 = W*in
   wire signed [9:0] m90_114;
   assign m90_114 =10'b0;

   // m90_115 = W*in
   wire signed [9:0] m90_115;
   assign m90_115 =10'b0;

   // m90_116 = W*in
   wire signed [9:0] m90_116;
   assign m90_116 =10'b0;

   // m90_117 = W*in
   wire signed [9:0] m90_117;
   assign m90_117 =10'b0;

   // m91_1 = W*in
   wire signed [9:0] m91_1;
   assign m91_1 =10'b0;

   // m91_2 = W*in
   wire signed [9:0] m91_2;
   assign m91_2 =10'b0;

   // m91_3 = W*in
   wire signed [9:0] m91_3;
   assign m91_3 =10'b0;

   // m91_4 = W*in
   wire signed [9:0] m91_4;
   assign m91_4 =10'b0;

   // m91_5 = W*in
   wire signed [9:0] m91_5;
   assign m91_5 =10'b0;

   // m91_6 = W*in
   wire signed [9:0] m91_6;
   assign m91_6 ={ {5{in91[5]}} , in91[5:1] };

   // m91_7 = W*in
   wire signed [9:0] m91_7;
   assign m91_7 =10'b0;

   // m91_8 = W*in
   wire signed [9:0] m91_8;
   assign m91_8 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_9 = W*in
   wire signed [9:0] m91_9;
   assign m91_9 =10'b0;

   // m91_10 = W*in
   wire signed [9:0] m91_10;
   assign m91_10 =10'b0;

   // m91_11 = W*in
   wire signed [9:0] m91_11;
   assign m91_11 ={ {4{in91[5]}} , in91[5:0] };

   // m91_12 = W*in
   wire signed [9:0] m91_12;
   assign m91_12 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_13 = W*in
   wire signed [9:0] m91_13;
   assign m91_13 =10'b0;

   // m91_14 = W*in
   wire signed [9:0] m91_14;
   assign m91_14 =10'b0;

   // m91_15 = W*in
   wire signed [9:0] m91_15;
   assign m91_15 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_16 = W*in
   wire signed [9:0] m91_16;
   assign m91_16 =10'b0;

   // m91_17 = W*in
   wire signed [9:0] m91_17;
   assign m91_17 ={ {5{in91[5]}} , in91[5:1] };

   // m91_18 = W*in
   wire signed [9:0] m91_18;
   assign m91_18 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_19 = W*in
   wire signed [9:0] m91_19;
   assign m91_19 ={ {5{in91[5]}} , in91[5:1] };

   // m91_20 = W*in
   wire signed [9:0] m91_20;
   assign m91_20 =10'b0;

   // m91_21 = W*in
   wire signed [9:0] m91_21;
   assign m91_21 =10'b0;

   // m91_22 = W*in
   wire signed [9:0] m91_22;
   assign m91_22 ={ {4{in91[5]}} , in91[5:0] };

   // m91_23 = W*in
   wire signed [9:0] m91_23;
   assign m91_23 =10'b0;

   // m91_24 = W*in
   wire signed [9:0] m91_24;
   assign m91_24 ={ {4{in91[5]}} , in91[5:0] };

   // m91_25 = W*in
   wire signed [9:0] m91_25;
   assign m91_25 =10'b0;

   // m91_26 = W*in
   wire signed [9:0] m91_26;
   assign m91_26 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_27 = W*in
   wire signed [9:0] m91_27;
   assign m91_27 ={ {5{in91[5]}} , in91[5:1] };

   // m91_28 = W*in
   wire signed [9:0] m91_28;
   assign m91_28 =10'b0;

   // m91_29 = W*in
   wire signed [9:0] m91_29;
   assign m91_29 ={ {5{in91[5]}} , in91[5:1] };

   // m91_30 = W*in
   wire signed [9:0] m91_30;
   assign m91_30 =10'b0;

   // m91_31 = W*in
   wire signed [9:0] m91_31;
   assign m91_31 ={ {5{neg91[5]}} , neg91[5:1] };

   // m91_32 = W*in
   wire signed [9:0] m91_32;
   assign m91_32 =10'b0;

   // m91_33 = W*in
   wire signed [9:0] m91_33;
   assign m91_33 =10'b0;

   // m91_34 = W*in
   wire signed [9:0] m91_34;
   assign m91_34 =10'b0;

   // m91_35 = W*in
   wire signed [9:0] m91_35;
   assign m91_35 =10'b0;

   // m91_36 = W*in
   wire signed [9:0] m91_36;
   assign m91_36 =10'b0;

   // m91_37 = W*in
   wire signed [9:0] m91_37;
   assign m91_37 =10'b0;

   // m91_38 = W*in
   wire signed [9:0] m91_38;
   assign m91_38 =10'b0;

   // m91_39 = W*in
   wire signed [9:0] m91_39;
   assign m91_39 =10'b0;

   // m91_40 = W*in
   wire signed [9:0] m91_40;
   assign m91_40 =10'b0;

   // m91_41 = W*in
   wire signed [9:0] m91_41;
   assign m91_41 =10'b0;

   // m91_42 = W*in
   wire signed [9:0] m91_42;
   assign m91_42 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_43 = W*in
   wire signed [9:0] m91_43;
   assign m91_43 =10'b0;

   // m91_44 = W*in
   wire signed [9:0] m91_44;
   assign m91_44 ={ {4{in91[5]}} , in91[5:0] };

   // m91_45 = W*in
   wire signed [9:0] m91_45;
   assign m91_45 =10'b0;

   // m91_46 = W*in
   wire signed [9:0] m91_46;
   assign m91_46 =10'b0;

   // m91_47 = W*in
   wire signed [9:0] m91_47;
   assign m91_47 =10'b0;

   // m91_48 = W*in
   wire signed [9:0] m91_48;
   assign m91_48 =10'b0;

   // m91_49 = W*in
   wire signed [9:0] m91_49;
   assign m91_49 =10'b0;

   // m91_50 = W*in
   wire signed [9:0] m91_50;
   assign m91_50 =10'b0;

   // m91_51 = W*in
   wire signed [9:0] m91_51;
   assign m91_51 =10'b0;

   // m91_52 = W*in
   wire signed [9:0] m91_52;
   assign m91_52 =10'b0;

   // m91_53 = W*in
   wire signed [9:0] m91_53;
   assign m91_53 =10'b0;

   // m91_54 = W*in
   wire signed [9:0] m91_54;
   assign m91_54 ={ {4{in91[5]}} , in91[5:0] };

   // m91_55 = W*in
   wire signed [9:0] m91_55;
   assign m91_55 =10'b0;

   // m91_56 = W*in
   wire signed [9:0] m91_56;
   assign m91_56 =10'b0;

   // m91_57 = W*in
   wire signed [9:0] m91_57;
   assign m91_57 =10'b0;

   // m91_58 = W*in
   wire signed [9:0] m91_58;
   assign m91_58 =10'b0;

   // m91_59 = W*in
   wire signed [9:0] m91_59;
   assign m91_59 =10'b0;

   // m91_60 = W*in
   wire signed [9:0] m91_60;
   assign m91_60 =10'b0;

   // m91_61 = W*in
   wire signed [9:0] m91_61;
   assign m91_61 ={ {4{in91[5]}} , in91[5:0] };

   // m91_62 = W*in
   wire signed [9:0] m91_62;
   assign m91_62 =10'b0;

   // m91_63 = W*in
   wire signed [9:0] m91_63;
   assign m91_63 =10'b0;

   // m91_64 = W*in
   wire signed [9:0] m91_64;
   assign m91_64 ={ {5{neg91[5]}} , neg91[5:1] };

   // m91_65 = W*in
   wire signed [9:0] m91_65;
   assign m91_65 =10'b0;

   // m91_66 = W*in
   wire signed [9:0] m91_66;
   assign m91_66 =10'b0;

   // m91_67 = W*in
   wire signed [9:0] m91_67;
   assign m91_67 =10'b0;

   // m91_68 = W*in
   wire signed [9:0] m91_68;
   assign m91_68 =10'b0;

   // m91_69 = W*in
   wire signed [9:0] m91_69;
   assign m91_69 =10'b0;

   // m91_70 = W*in
   wire signed [9:0] m91_70;
   assign m91_70 =10'b0;

   // m91_71 = W*in
   wire signed [9:0] m91_71;
   assign m91_71 =10'b0;

   // m91_72 = W*in
   wire signed [9:0] m91_72;
   assign m91_72 ={ {5{neg91[5]}} , neg91[5:1] };

   // m91_73 = W*in
   wire signed [9:0] m91_73;
   assign m91_73 =10'b0;

   // m91_74 = W*in
   wire signed [9:0] m91_74;
   assign m91_74 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_75 = W*in
   wire signed [9:0] m91_75;
   assign m91_75 ={ {5{neg91[5]}} , neg91[5:1] };

   // m91_76 = W*in
   wire signed [9:0] m91_76;
   assign m91_76 =10'b0;

   // m91_77 = W*in
   wire signed [9:0] m91_77;
   assign m91_77 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_78 = W*in
   wire signed [9:0] m91_78;
   assign m91_78 ={ {5{neg91[5]}} , neg91[5:1] };

   // m91_79 = W*in
   wire signed [9:0] m91_79;
   assign m91_79 ={ {4{in91[5]}} , in91[5:0] };

   // m91_80 = W*in
   wire signed [9:0] m91_80;
   assign m91_80 =10'b0;

   // m91_81 = W*in
   wire signed [9:0] m91_81;
   assign m91_81 ={ {5{neg91[5]}} , neg91[5:1] };

   // m91_82 = W*in
   wire signed [9:0] m91_82;
   assign m91_82 =10'b0;

   // m91_83 = W*in
   wire signed [9:0] m91_83;
   assign m91_83 ={ {5{in91[5]}} , in91[5:1] };

   // m91_84 = W*in
   wire signed [9:0] m91_84;
   assign m91_84 =10'b0;

   // m91_85 = W*in
   wire signed [9:0] m91_85;
   assign m91_85 ={ {4{in91[5]}} , in91[5:0] };

   // m91_86 = W*in
   wire signed [9:0] m91_86;
   assign m91_86 =10'b0;

   // m91_87 = W*in
   wire signed [9:0] m91_87;
   assign m91_87 =10'b0;

   // m91_88 = W*in
   wire signed [9:0] m91_88;
   assign m91_88 =10'b0;

   // m91_89 = W*in
   wire signed [9:0] m91_89;
   assign m91_89 =10'b0;

   // m91_90 = W*in
   wire signed [9:0] m91_90;
   assign m91_90 =10'b0;

   // m91_91 = W*in
   wire signed [9:0] m91_91;
   assign m91_91 =10'b0;

   // m91_92 = W*in
   wire signed [9:0] m91_92;
   assign m91_92 =10'b0;

   // m91_93 = W*in
   wire signed [9:0] m91_93;
   assign m91_93 ={ {4{in91[5]}} , in91[5:0] };

   // m91_94 = W*in
   wire signed [9:0] m91_94;
   assign m91_94 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_95 = W*in
   wire signed [9:0] m91_95;
   assign m91_95 ={ {4{in91[5]}} , in91[5:0] };

   // m91_96 = W*in
   wire signed [9:0] m91_96;
   assign m91_96 =10'b0;

   // m91_97 = W*in
   wire signed [9:0] m91_97;
   assign m91_97 =10'b0;

   // m91_98 = W*in
   wire signed [9:0] m91_98;
   assign m91_98 =10'b0;

   // m91_99 = W*in
   wire signed [9:0] m91_99;
   assign m91_99 =10'b0;

   // m91_100 = W*in
   wire signed [9:0] m91_100;
   assign m91_100 ={ {4{neg91[5]}} , neg91[5:0] };

   // m91_101 = W*in
   wire signed [9:0] m91_101;
   assign m91_101 =10'b0;

   // m91_102 = W*in
   wire signed [9:0] m91_102;
   assign m91_102 =10'b0;

   // m91_103 = W*in
   wire signed [9:0] m91_103;
   assign m91_103 =10'b0;

   // m91_104 = W*in
   wire signed [9:0] m91_104;
   assign m91_104 =10'b0;

   // m91_105 = W*in
   wire signed [9:0] m91_105;
   assign m91_105 =10'b0;

   // m91_106 = W*in
   wire signed [9:0] m91_106;
   assign m91_106 =10'b0;

   // m91_107 = W*in
   wire signed [9:0] m91_107;
   assign m91_107 =10'b0;

   // m91_108 = W*in
   wire signed [9:0] m91_108;
   assign m91_108 =10'b0;

   // m91_109 = W*in
   wire signed [9:0] m91_109;
   assign m91_109 =10'b0;

   // m91_110 = W*in
   wire signed [9:0] m91_110;
   assign m91_110 =10'b0;

   // m91_111 = W*in
   wire signed [9:0] m91_111;
   assign m91_111 =10'b0;

   // m91_112 = W*in
   wire signed [9:0] m91_112;
   assign m91_112 =10'b0;

   // m91_113 = W*in
   wire signed [9:0] m91_113;
   assign m91_113 =10'b0;

   // m91_114 = W*in
   wire signed [9:0] m91_114;
   assign m91_114 ={ {5{in91[5]}} , in91[5:1] };

   // m91_115 = W*in
   wire signed [9:0] m91_115;
   assign m91_115 =10'b0;

   // m91_116 = W*in
   wire signed [9:0] m91_116;
   assign m91_116 =10'b0;

   // m91_117 = W*in
   wire signed [9:0] m91_117;
   assign m91_117 =10'b0;

   // m92_1 = W*in
   wire signed [9:0] m92_1;
   assign m92_1 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_2 = W*in
   wire signed [9:0] m92_2;
   assign m92_2 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_3 = W*in
   wire signed [9:0] m92_3;
   assign m92_3 =10'b0;

   // m92_4 = W*in
   wire signed [9:0] m92_4;
   assign m92_4 =10'b0;

   // m92_5 = W*in
   wire signed [9:0] m92_5;
   assign m92_5 =10'b0;

   // m92_6 = W*in
   wire signed [9:0] m92_6;
   assign m92_6 =10'b0;

   // m92_7 = W*in
   wire signed [9:0] m92_7;
   assign m92_7 =10'b0;

   // m92_8 = W*in
   wire signed [9:0] m92_8;
   assign m92_8 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_9 = W*in
   wire signed [9:0] m92_9;
   assign m92_9 =10'b0;

   // m92_10 = W*in
   wire signed [9:0] m92_10;
   assign m92_10 ={ {4{in92[5]}} , in92[5:0] };

   // m92_11 = W*in
   wire signed [9:0] m92_11;
   assign m92_11 ={ {4{in92[5]}} , in92[5:0] };

   // m92_12 = W*in
   wire signed [9:0] m92_12;
   assign m92_12 =10'b0;

   // m92_13 = W*in
   wire signed [9:0] m92_13;
   assign m92_13 =10'b0;

   // m92_14 = W*in
   wire signed [9:0] m92_14;
   assign m92_14 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_15 = W*in
   wire signed [9:0] m92_15;
   assign m92_15 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_16 = W*in
   wire signed [9:0] m92_16;
   assign m92_16 =10'b0;

   // m92_17 = W*in
   wire signed [9:0] m92_17;
   assign m92_17 =10'b0;

   // m92_18 = W*in
   wire signed [9:0] m92_18;
   assign m92_18 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_19 = W*in
   wire signed [9:0] m92_19;
   assign m92_19 =10'b0;

   // m92_20 = W*in
   wire signed [9:0] m92_20;
   assign m92_20 =10'b0;

   // m92_21 = W*in
   wire signed [9:0] m92_21;
   assign m92_21 ={ {4{in92[5]}} , in92[5:0] };

   // m92_22 = W*in
   wire signed [9:0] m92_22;
   assign m92_22 =10'b0;

   // m92_23 = W*in
   wire signed [9:0] m92_23;
   assign m92_23 =10'b0;

   // m92_24 = W*in
   wire signed [9:0] m92_24;
   assign m92_24 =10'b0;

   // m92_25 = W*in
   wire signed [9:0] m92_25;
   assign m92_25 =10'b0;

   // m92_26 = W*in
   wire signed [9:0] m92_26;
   assign m92_26 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_27 = W*in
   wire signed [9:0] m92_27;
   assign m92_27 =10'b0;

   // m92_28 = W*in
   wire signed [9:0] m92_28;
   assign m92_28 =10'b0;

   // m92_29 = W*in
   wire signed [9:0] m92_29;
   assign m92_29 ={ {4{in92[5]}} , in92[5:0] };

   // m92_30 = W*in
   wire signed [9:0] m92_30;
   assign m92_30 =10'b0;

   // m92_31 = W*in
   wire signed [9:0] m92_31;
   assign m92_31 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_32 = W*in
   wire signed [9:0] m92_32;
   assign m92_32 =10'b0;

   // m92_33 = W*in
   wire signed [9:0] m92_33;
   assign m92_33 =10'b0;

   // m92_34 = W*in
   wire signed [9:0] m92_34;
   assign m92_34 =10'b0;

   // m92_35 = W*in
   wire signed [9:0] m92_35;
   assign m92_35 ={ {5{in92[5]}} , in92[5:1] };

   // m92_36 = W*in
   wire signed [9:0] m92_36;
   assign m92_36 =10'b0;

   // m92_37 = W*in
   wire signed [9:0] m92_37;
   assign m92_37 =10'b0;

   // m92_38 = W*in
   wire signed [9:0] m92_38;
   assign m92_38 =10'b0;

   // m92_39 = W*in
   wire signed [9:0] m92_39;
   assign m92_39 =10'b0;

   // m92_40 = W*in
   wire signed [9:0] m92_40;
   assign m92_40 =10'b0;

   // m92_41 = W*in
   wire signed [9:0] m92_41;
   assign m92_41 =10'b0;

   // m92_42 = W*in
   wire signed [9:0] m92_42;
   assign m92_42 =10'b0;

   // m92_43 = W*in
   wire signed [9:0] m92_43;
   assign m92_43 =10'b0;

   // m92_44 = W*in
   wire signed [9:0] m92_44;
   assign m92_44 =10'b0;

   // m92_45 = W*in
   wire signed [9:0] m92_45;
   assign m92_45 =10'b0;

   // m92_46 = W*in
   wire signed [9:0] m92_46;
   assign m92_46 =10'b0;

   // m92_47 = W*in
   wire signed [9:0] m92_47;
   assign m92_47 =10'b0;

   // m92_48 = W*in
   wire signed [9:0] m92_48;
   assign m92_48 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_49 = W*in
   wire signed [9:0] m92_49;
   assign m92_49 =10'b0;

   // m92_50 = W*in
   wire signed [9:0] m92_50;
   assign m92_50 ={ {3{neg92[5]}} , neg92 , {1{1'b0}} };

   // m92_51 = W*in
   wire signed [9:0] m92_51;
   assign m92_51 =10'b0;

   // m92_52 = W*in
   wire signed [9:0] m92_52;
   assign m92_52 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_53 = W*in
   wire signed [9:0] m92_53;
   assign m92_53 =10'b0;

   // m92_54 = W*in
   wire signed [9:0] m92_54;
   assign m92_54 ={ {4{in92[5]}} , in92[5:0] };

   // m92_55 = W*in
   wire signed [9:0] m92_55;
   assign m92_55 =10'b0;

   // m92_56 = W*in
   wire signed [9:0] m92_56;
   assign m92_56 =10'b0;

   // m92_57 = W*in
   wire signed [9:0] m92_57;
   assign m92_57 =10'b0;

   // m92_58 = W*in
   wire signed [9:0] m92_58;
   assign m92_58 =10'b0;

   // m92_59 = W*in
   wire signed [9:0] m92_59;
   assign m92_59 =10'b0;

   // m92_60 = W*in
   wire signed [9:0] m92_60;
   assign m92_60 =10'b0;

   // m92_61 = W*in
   wire signed [9:0] m92_61;
   assign m92_61 =10'b0;

   // m92_62 = W*in
   wire signed [9:0] m92_62;
   assign m92_62 =10'b0;

   // m92_63 = W*in
   wire signed [9:0] m92_63;
   assign m92_63 =10'b0;

   // m92_64 = W*in
   wire signed [9:0] m92_64;
   assign m92_64 =10'b0;

   // m92_65 = W*in
   wire signed [9:0] m92_65;
   assign m92_65 =10'b0;

   // m92_66 = W*in
   wire signed [9:0] m92_66;
   assign m92_66 =10'b0;

   // m92_67 = W*in
   wire signed [9:0] m92_67;
   assign m92_67 =10'b0;

   // m92_68 = W*in
   wire signed [9:0] m92_68;
   assign m92_68 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_69 = W*in
   wire signed [9:0] m92_69;
   assign m92_69 =10'b0;

   // m92_70 = W*in
   wire signed [9:0] m92_70;
   assign m92_70 ={ {4{in92[5]}} , in92[5:0] };

   // m92_71 = W*in
   wire signed [9:0] m92_71;
   assign m92_71 =10'b0;

   // m92_72 = W*in
   wire signed [9:0] m92_72;
   assign m92_72 =10'b0;

   // m92_73 = W*in
   wire signed [9:0] m92_73;
   assign m92_73 ={ {5{neg92[5]}} , neg92[5:1] };

   // m92_74 = W*in
   wire signed [9:0] m92_74;
   assign m92_74 =10'b0;

   // m92_75 = W*in
   wire signed [9:0] m92_75;
   assign m92_75 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_76 = W*in
   wire signed [9:0] m92_76;
   assign m92_76 =10'b0;

   // m92_77 = W*in
   wire signed [9:0] m92_77;
   assign m92_77 =10'b0;

   // m92_78 = W*in
   wire signed [9:0] m92_78;
   assign m92_78 ={ {5{neg92[5]}} , neg92[5:1] };

   // m92_79 = W*in
   wire signed [9:0] m92_79;
   assign m92_79 ={ {4{in92[5]}} , in92[5:0] };

   // m92_80 = W*in
   wire signed [9:0] m92_80;
   assign m92_80 =10'b0;

   // m92_81 = W*in
   wire signed [9:0] m92_81;
   assign m92_81 =10'b0;

   // m92_82 = W*in
   wire signed [9:0] m92_82;
   assign m92_82 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_83 = W*in
   wire signed [9:0] m92_83;
   assign m92_83 =10'b0;

   // m92_84 = W*in
   wire signed [9:0] m92_84;
   assign m92_84 =10'b0;

   // m92_85 = W*in
   wire signed [9:0] m92_85;
   assign m92_85 ={ {4{in92[5]}} , in92[5:0] };

   // m92_86 = W*in
   wire signed [9:0] m92_86;
   assign m92_86 ={ {4{in92[5]}} , in92[5:0] };

   // m92_87 = W*in
   wire signed [9:0] m92_87;
   assign m92_87 =10'b0;

   // m92_88 = W*in
   wire signed [9:0] m92_88;
   assign m92_88 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_89 = W*in
   wire signed [9:0] m92_89;
   assign m92_89 =10'b0;

   // m92_90 = W*in
   wire signed [9:0] m92_90;
   assign m92_90 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_91 = W*in
   wire signed [9:0] m92_91;
   assign m92_91 =10'b0;

   // m92_92 = W*in
   wire signed [9:0] m92_92;
   assign m92_92 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_93 = W*in
   wire signed [9:0] m92_93;
   assign m92_93 ={ {4{in92[5]}} , in92[5:0] };

   // m92_94 = W*in
   wire signed [9:0] m92_94;
   assign m92_94 =10'b0;

   // m92_95 = W*in
   wire signed [9:0] m92_95;
   assign m92_95 ={ {4{in92[5]}} , in92[5:0] };

   // m92_96 = W*in
   wire signed [9:0] m92_96;
   assign m92_96 =10'b0;

   // m92_97 = W*in
   wire signed [9:0] m92_97;
   assign m92_97 =10'b0;

   // m92_98 = W*in
   wire signed [9:0] m92_98;
   assign m92_98 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_99 = W*in
   wire signed [9:0] m92_99;
   assign m92_99 =10'b0;

   // m92_100 = W*in
   wire signed [9:0] m92_100;
   assign m92_100 =10'b0;

   // m92_101 = W*in
   wire signed [9:0] m92_101;
   assign m92_101 =10'b0;

   // m92_102 = W*in
   wire signed [9:0] m92_102;
   assign m92_102 =10'b0;

   // m92_103 = W*in
   wire signed [9:0] m92_103;
   assign m92_103 =10'b0;

   // m92_104 = W*in
   wire signed [9:0] m92_104;
   assign m92_104 =10'b0;

   // m92_105 = W*in
   wire signed [9:0] m92_105;
   assign m92_105 =10'b0;

   // m92_106 = W*in
   wire signed [9:0] m92_106;
   assign m92_106 =10'b0;

   // m92_107 = W*in
   wire signed [9:0] m92_107;
   assign m92_107 =10'b0;

   // m92_108 = W*in
   wire signed [9:0] m92_108;
   assign m92_108 ={ {4{in92[5]}} , in92[5:0] };

   // m92_109 = W*in
   wire signed [9:0] m92_109;
   assign m92_109 ={ {5{in92[5]}} , in92[5:1] };

   // m92_110 = W*in
   wire signed [9:0] m92_110;
   assign m92_110 =10'b0;

   // m92_111 = W*in
   wire signed [9:0] m92_111;
   assign m92_111 =10'b0;

   // m92_112 = W*in
   wire signed [9:0] m92_112;
   assign m92_112 =10'b0;

   // m92_113 = W*in
   wire signed [9:0] m92_113;
   assign m92_113 ={ {4{neg92[5]}} , neg92[5:0] };

   // m92_114 = W*in
   wire signed [9:0] m92_114;
   assign m92_114 ={ {5{in92[5]}} , in92[5:1] };

   // m92_115 = W*in
   wire signed [9:0] m92_115;
   assign m92_115 =10'b0;

   // m92_116 = W*in
   wire signed [9:0] m92_116;
   assign m92_116 =10'b0;

   // m92_117 = W*in
   wire signed [9:0] m92_117;
   assign m92_117 ={ {4{in92[5]}} , in92[5:0] };

   // m93_1 = W*in
   wire signed [9:0] m93_1;
   assign m93_1 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_2 = W*in
   wire signed [9:0] m93_2;
   assign m93_2 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_3 = W*in
   wire signed [9:0] m93_3;
   assign m93_3 =10'b0;

   // m93_4 = W*in
   wire signed [9:0] m93_4;
   assign m93_4 =10'b0;

   // m93_5 = W*in
   wire signed [9:0] m93_5;
   assign m93_5 =10'b0;

   // m93_6 = W*in
   wire signed [9:0] m93_6;
   assign m93_6 ={ {4{in93[5]}} , in93[5:0] };

   // m93_7 = W*in
   wire signed [9:0] m93_7;
   assign m93_7 =10'b0;

   // m93_8 = W*in
   wire signed [9:0] m93_8;
   assign m93_8 =10'b0;

   // m93_9 = W*in
   wire signed [9:0] m93_9;
   assign m93_9 =10'b0;

   // m93_10 = W*in
   wire signed [9:0] m93_10;
   assign m93_10 ={ {4{in93[5]}} , in93[5:0] };

   // m93_11 = W*in
   wire signed [9:0] m93_11;
   assign m93_11 =10'b0;

   // m93_12 = W*in
   wire signed [9:0] m93_12;
   assign m93_12 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_13 = W*in
   wire signed [9:0] m93_13;
   assign m93_13 =10'b0;

   // m93_14 = W*in
   wire signed [9:0] m93_14;
   assign m93_14 =10'b0;

   // m93_15 = W*in
   wire signed [9:0] m93_15;
   assign m93_15 =10'b0;

   // m93_16 = W*in
   wire signed [9:0] m93_16;
   assign m93_16 =10'b0;

   // m93_17 = W*in
   wire signed [9:0] m93_17;
   assign m93_17 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_18 = W*in
   wire signed [9:0] m93_18;
   assign m93_18 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_19 = W*in
   wire signed [9:0] m93_19;
   assign m93_19 ={ {5{neg93[5]}} , neg93[5:1] };

   // m93_20 = W*in
   wire signed [9:0] m93_20;
   assign m93_20 ={ {5{in93[5]}} , in93[5:1] };

   // m93_21 = W*in
   wire signed [9:0] m93_21;
   assign m93_21 ={ {4{in93[5]}} , in93[5:0] };

   // m93_22 = W*in
   wire signed [9:0] m93_22;
   assign m93_22 =10'b0;

   // m93_23 = W*in
   wire signed [9:0] m93_23;
   assign m93_23 =10'b0;

   // m93_24 = W*in
   wire signed [9:0] m93_24;
   assign m93_24 =10'b0;

   // m93_25 = W*in
   wire signed [9:0] m93_25;
   assign m93_25 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_26 = W*in
   wire signed [9:0] m93_26;
   assign m93_26 =10'b0;

   // m93_27 = W*in
   wire signed [9:0] m93_27;
   assign m93_27 =10'b0;

   // m93_28 = W*in
   wire signed [9:0] m93_28;
   assign m93_28 =10'b0;

   // m93_29 = W*in
   wire signed [9:0] m93_29;
   assign m93_29 ={ {5{in93[5]}} , in93[5:1] };

   // m93_30 = W*in
   wire signed [9:0] m93_30;
   assign m93_30 =10'b0;

   // m93_31 = W*in
   wire signed [9:0] m93_31;
   assign m93_31 ={ {5{neg93[5]}} , neg93[5:1] };

   // m93_32 = W*in
   wire signed [9:0] m93_32;
   assign m93_32 ={ {4{in93[5]}} , in93[5:0] };

   // m93_33 = W*in
   wire signed [9:0] m93_33;
   assign m93_33 =10'b0;

   // m93_34 = W*in
   wire signed [9:0] m93_34;
   assign m93_34 =10'b0;

   // m93_35 = W*in
   wire signed [9:0] m93_35;
   assign m93_35 =10'b0;

   // m93_36 = W*in
   wire signed [9:0] m93_36;
   assign m93_36 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_37 = W*in
   wire signed [9:0] m93_37;
   assign m93_37 ={ {5{neg93[5]}} , neg93[5:1] };

   // m93_38 = W*in
   wire signed [9:0] m93_38;
   assign m93_38 =10'b0;

   // m93_39 = W*in
   wire signed [9:0] m93_39;
   assign m93_39 =10'b0;

   // m93_40 = W*in
   wire signed [9:0] m93_40;
   assign m93_40 =10'b0;

   // m93_41 = W*in
   wire signed [9:0] m93_41;
   assign m93_41 =10'b0;

   // m93_42 = W*in
   wire signed [9:0] m93_42;
   assign m93_42 =10'b0;

   // m93_43 = W*in
   wire signed [9:0] m93_43;
   assign m93_43 =10'b0;

   // m93_44 = W*in
   wire signed [9:0] m93_44;
   assign m93_44 =10'b0;

   // m93_45 = W*in
   wire signed [9:0] m93_45;
   assign m93_45 =10'b0;

   // m93_46 = W*in
   wire signed [9:0] m93_46;
   assign m93_46 =10'b0;

   // m93_47 = W*in
   wire signed [9:0] m93_47;
   assign m93_47 =10'b0;

   // m93_48 = W*in
   wire signed [9:0] m93_48;
   assign m93_48 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_49 = W*in
   wire signed [9:0] m93_49;
   assign m93_49 =10'b0;

   // m93_50 = W*in
   wire signed [9:0] m93_50;
   assign m93_50 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_51 = W*in
   wire signed [9:0] m93_51;
   assign m93_51 =10'b0;

   // m93_52 = W*in
   wire signed [9:0] m93_52;
   assign m93_52 =10'b0;

   // m93_53 = W*in
   wire signed [9:0] m93_53;
   assign m93_53 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_54 = W*in
   wire signed [9:0] m93_54;
   assign m93_54 =10'b0;

   // m93_55 = W*in
   wire signed [9:0] m93_55;
   assign m93_55 =10'b0;

   // m93_56 = W*in
   wire signed [9:0] m93_56;
   assign m93_56 =10'b0;

   // m93_57 = W*in
   wire signed [9:0] m93_57;
   assign m93_57 =10'b0;

   // m93_58 = W*in
   wire signed [9:0] m93_58;
   assign m93_58 =10'b0;

   // m93_59 = W*in
   wire signed [9:0] m93_59;
   assign m93_59 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_60 = W*in
   wire signed [9:0] m93_60;
   assign m93_60 =10'b0;

   // m93_61 = W*in
   wire signed [9:0] m93_61;
   assign m93_61 =10'b0;

   // m93_62 = W*in
   wire signed [9:0] m93_62;
   assign m93_62 =10'b0;

   // m93_63 = W*in
   wire signed [9:0] m93_63;
   assign m93_63 =10'b0;

   // m93_64 = W*in
   wire signed [9:0] m93_64;
   assign m93_64 =10'b0;

   // m93_65 = W*in
   wire signed [9:0] m93_65;
   assign m93_65 =10'b0;

   // m93_66 = W*in
   wire signed [9:0] m93_66;
   assign m93_66 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_67 = W*in
   wire signed [9:0] m93_67;
   assign m93_67 =10'b0;

   // m93_68 = W*in
   wire signed [9:0] m93_68;
   assign m93_68 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_69 = W*in
   wire signed [9:0] m93_69;
   assign m93_69 =10'b0;

   // m93_70 = W*in
   wire signed [9:0] m93_70;
   assign m93_70 =10'b0;

   // m93_71 = W*in
   wire signed [9:0] m93_71;
   assign m93_71 =10'b0;

   // m93_72 = W*in
   wire signed [9:0] m93_72;
   assign m93_72 =10'b0;

   // m93_73 = W*in
   wire signed [9:0] m93_73;
   assign m93_73 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_74 = W*in
   wire signed [9:0] m93_74;
   assign m93_74 ={ {4{in93[5]}} , in93[5:0] };

   // m93_75 = W*in
   wire signed [9:0] m93_75;
   assign m93_75 =10'b0;

   // m93_76 = W*in
   wire signed [9:0] m93_76;
   assign m93_76 =10'b0;

   // m93_77 = W*in
   wire signed [9:0] m93_77;
   assign m93_77 =10'b0;

   // m93_78 = W*in
   wire signed [9:0] m93_78;
   assign m93_78 =10'b0;

   // m93_79 = W*in
   wire signed [9:0] m93_79;
   assign m93_79 =10'b0;

   // m93_80 = W*in
   wire signed [9:0] m93_80;
   assign m93_80 =10'b0;

   // m93_81 = W*in
   wire signed [9:0] m93_81;
   assign m93_81 =10'b0;

   // m93_82 = W*in
   wire signed [9:0] m93_82;
   assign m93_82 =10'b0;

   // m93_83 = W*in
   wire signed [9:0] m93_83;
   assign m93_83 =10'b0;

   // m93_84 = W*in
   wire signed [9:0] m93_84;
   assign m93_84 =10'b0;

   // m93_85 = W*in
   wire signed [9:0] m93_85;
   assign m93_85 =10'b0;

   // m93_86 = W*in
   wire signed [9:0] m93_86;
   assign m93_86 =10'b0;

   // m93_87 = W*in
   wire signed [9:0] m93_87;
   assign m93_87 =10'b0;

   // m93_88 = W*in
   wire signed [9:0] m93_88;
   assign m93_88 =10'b0;

   // m93_89 = W*in
   wire signed [9:0] m93_89;
   assign m93_89 ={ {4{in93[5]}} , in93[5:0] };

   // m93_90 = W*in
   wire signed [9:0] m93_90;
   assign m93_90 =10'b0;

   // m93_91 = W*in
   wire signed [9:0] m93_91;
   assign m93_91 =10'b0;

   // m93_92 = W*in
   wire signed [9:0] m93_92;
   assign m93_92 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_93 = W*in
   wire signed [9:0] m93_93;
   assign m93_93 =10'b0;

   // m93_94 = W*in
   wire signed [9:0] m93_94;
   assign m93_94 =10'b0;

   // m93_95 = W*in
   wire signed [9:0] m93_95;
   assign m93_95 =10'b0;

   // m93_96 = W*in
   wire signed [9:0] m93_96;
   assign m93_96 =10'b0;

   // m93_97 = W*in
   wire signed [9:0] m93_97;
   assign m93_97 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_98 = W*in
   wire signed [9:0] m93_98;
   assign m93_98 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_99 = W*in
   wire signed [9:0] m93_99;
   assign m93_99 =10'b0;

   // m93_100 = W*in
   wire signed [9:0] m93_100;
   assign m93_100 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_101 = W*in
   wire signed [9:0] m93_101;
   assign m93_101 =10'b0;

   // m93_102 = W*in
   wire signed [9:0] m93_102;
   assign m93_102 =10'b0;

   // m93_103 = W*in
   wire signed [9:0] m93_103;
   assign m93_103 =10'b0;

   // m93_104 = W*in
   wire signed [9:0] m93_104;
   assign m93_104 =10'b0;

   // m93_105 = W*in
   wire signed [9:0] m93_105;
   assign m93_105 =10'b0;

   // m93_106 = W*in
   wire signed [9:0] m93_106;
   assign m93_106 =10'b0;

   // m93_107 = W*in
   wire signed [9:0] m93_107;
   assign m93_107 =10'b0;

   // m93_108 = W*in
   wire signed [9:0] m93_108;
   assign m93_108 =10'b0;

   // m93_109 = W*in
   wire signed [9:0] m93_109;
   assign m93_109 =10'b0;

   // m93_110 = W*in
   wire signed [9:0] m93_110;
   assign m93_110 =10'b0;

   // m93_111 = W*in
   wire signed [9:0] m93_111;
   assign m93_111 =10'b0;

   // m93_112 = W*in
   wire signed [9:0] m93_112;
   assign m93_112 ={ {4{neg93[5]}} , neg93[5:0] };

   // m93_113 = W*in
   wire signed [9:0] m93_113;
   assign m93_113 =10'b0;

   // m93_114 = W*in
   wire signed [9:0] m93_114;
   assign m93_114 =10'b0;

   // m93_115 = W*in
   wire signed [9:0] m93_115;
   assign m93_115 =10'b0;

   // m93_116 = W*in
   wire signed [9:0] m93_116;
   assign m93_116 =10'b0;

   // m93_117 = W*in
   wire signed [9:0] m93_117;
   assign m93_117 =10'b0;

   // m94_1 = W*in
   wire signed [9:0] m94_1;
   assign m94_1 =10'b0;

   // m94_2 = W*in
   wire signed [9:0] m94_2;
   assign m94_2 =10'b0;

   // m94_3 = W*in
   wire signed [9:0] m94_3;
   assign m94_3 =10'b0;

   // m94_4 = W*in
   wire signed [9:0] m94_4;
   assign m94_4 =10'b0;

   // m94_5 = W*in
   wire signed [9:0] m94_5;
   assign m94_5 =10'b0;

   // m94_6 = W*in
   wire signed [9:0] m94_6;
   assign m94_6 ={ {4{in94[5]}} , in94[5:0] };

   // m94_7 = W*in
   wire signed [9:0] m94_7;
   assign m94_7 =10'b0;

   // m94_8 = W*in
   wire signed [9:0] m94_8;
   assign m94_8 =10'b0;

   // m94_9 = W*in
   wire signed [9:0] m94_9;
   assign m94_9 =10'b0;

   // m94_10 = W*in
   wire signed [9:0] m94_10;
   assign m94_10 =10'b0;

   // m94_11 = W*in
   wire signed [9:0] m94_11;
   assign m94_11 =10'b0;

   // m94_12 = W*in
   wire signed [9:0] m94_12;
   assign m94_12 =10'b0;

   // m94_13 = W*in
   wire signed [9:0] m94_13;
   assign m94_13 =10'b0;

   // m94_14 = W*in
   wire signed [9:0] m94_14;
   assign m94_14 =10'b0;

   // m94_15 = W*in
   wire signed [9:0] m94_15;
   assign m94_15 =10'b0;

   // m94_16 = W*in
   wire signed [9:0] m94_16;
   assign m94_16 =10'b0;

   // m94_17 = W*in
   wire signed [9:0] m94_17;
   assign m94_17 =10'b0;

   // m94_18 = W*in
   wire signed [9:0] m94_18;
   assign m94_18 =10'b0;

   // m94_19 = W*in
   wire signed [9:0] m94_19;
   assign m94_19 ={ {5{neg94[5]}} , neg94[5:1] };

   // m94_20 = W*in
   wire signed [9:0] m94_20;
   assign m94_20 =10'b0;

   // m94_21 = W*in
   wire signed [9:0] m94_21;
   assign m94_21 =10'b0;

   // m94_22 = W*in
   wire signed [9:0] m94_22;
   assign m94_22 =10'b0;

   // m94_23 = W*in
   wire signed [9:0] m94_23;
   assign m94_23 =10'b0;

   // m94_24 = W*in
   wire signed [9:0] m94_24;
   assign m94_24 =10'b0;

   // m94_25 = W*in
   wire signed [9:0] m94_25;
   assign m94_25 =10'b0;

   // m94_26 = W*in
   wire signed [9:0] m94_26;
   assign m94_26 =10'b0;

   // m94_27 = W*in
   wire signed [9:0] m94_27;
   assign m94_27 =10'b0;

   // m94_28 = W*in
   wire signed [9:0] m94_28;
   assign m94_28 =10'b0;

   // m94_29 = W*in
   wire signed [9:0] m94_29;
   assign m94_29 =10'b0;

   // m94_30 = W*in
   wire signed [9:0] m94_30;
   assign m94_30 =10'b0;

   // m94_31 = W*in
   wire signed [9:0] m94_31;
   assign m94_31 =10'b0;

   // m94_32 = W*in
   wire signed [9:0] m94_32;
   assign m94_32 =10'b0;

   // m94_33 = W*in
   wire signed [9:0] m94_33;
   assign m94_33 =10'b0;

   // m94_34 = W*in
   wire signed [9:0] m94_34;
   assign m94_34 =10'b0;

   // m94_35 = W*in
   wire signed [9:0] m94_35;
   assign m94_35 =10'b0;

   // m94_36 = W*in
   wire signed [9:0] m94_36;
   assign m94_36 ={ {5{neg94[5]}} , neg94[5:1] };

   // m94_37 = W*in
   wire signed [9:0] m94_37;
   assign m94_37 =10'b0;

   // m94_38 = W*in
   wire signed [9:0] m94_38;
   assign m94_38 =10'b0;

   // m94_39 = W*in
   wire signed [9:0] m94_39;
   assign m94_39 =10'b0;

   // m94_40 = W*in
   wire signed [9:0] m94_40;
   assign m94_40 =10'b0;

   // m94_41 = W*in
   wire signed [9:0] m94_41;
   assign m94_41 =10'b0;

   // m94_42 = W*in
   wire signed [9:0] m94_42;
   assign m94_42 =10'b0;

   // m94_43 = W*in
   wire signed [9:0] m94_43;
   assign m94_43 =10'b0;

   // m94_44 = W*in
   wire signed [9:0] m94_44;
   assign m94_44 =10'b0;

   // m94_45 = W*in
   wire signed [9:0] m94_45;
   assign m94_45 =10'b0;

   // m94_46 = W*in
   wire signed [9:0] m94_46;
   assign m94_46 =10'b0;

   // m94_47 = W*in
   wire signed [9:0] m94_47;
   assign m94_47 =10'b0;

   // m94_48 = W*in
   wire signed [9:0] m94_48;
   assign m94_48 =10'b0;

   // m94_49 = W*in
   wire signed [9:0] m94_49;
   assign m94_49 =10'b0;

   // m94_50 = W*in
   wire signed [9:0] m94_50;
   assign m94_50 =10'b0;

   // m94_51 = W*in
   wire signed [9:0] m94_51;
   assign m94_51 =10'b0;

   // m94_52 = W*in
   wire signed [9:0] m94_52;
   assign m94_52 =10'b0;

   // m94_53 = W*in
   wire signed [9:0] m94_53;
   assign m94_53 =10'b0;

   // m94_54 = W*in
   wire signed [9:0] m94_54;
   assign m94_54 =10'b0;

   // m94_55 = W*in
   wire signed [9:0] m94_55;
   assign m94_55 =10'b0;

   // m94_56 = W*in
   wire signed [9:0] m94_56;
   assign m94_56 =10'b0;

   // m94_57 = W*in
   wire signed [9:0] m94_57;
   assign m94_57 =10'b0;

   // m94_58 = W*in
   wire signed [9:0] m94_58;
   assign m94_58 =10'b0;

   // m94_59 = W*in
   wire signed [9:0] m94_59;
   assign m94_59 =10'b0;

   // m94_60 = W*in
   wire signed [9:0] m94_60;
   assign m94_60 =10'b0;

   // m94_61 = W*in
   wire signed [9:0] m94_61;
   assign m94_61 =10'b0;

   // m94_62 = W*in
   wire signed [9:0] m94_62;
   assign m94_62 =10'b0;

   // m94_63 = W*in
   wire signed [9:0] m94_63;
   assign m94_63 =10'b0;

   // m94_64 = W*in
   wire signed [9:0] m94_64;
   assign m94_64 =10'b0;

   // m94_65 = W*in
   wire signed [9:0] m94_65;
   assign m94_65 ={ {5{in94[5]}} , in94[5:1] };

   // m94_66 = W*in
   wire signed [9:0] m94_66;
   assign m94_66 ={ {4{in94[5]}} , in94[5:0] };

   // m94_67 = W*in
   wire signed [9:0] m94_67;
   assign m94_67 =10'b0;

   // m94_68 = W*in
   wire signed [9:0] m94_68;
   assign m94_68 =10'b0;

   // m94_69 = W*in
   wire signed [9:0] m94_69;
   assign m94_69 =10'b0;

   // m94_70 = W*in
   wire signed [9:0] m94_70;
   assign m94_70 =10'b0;

   // m94_71 = W*in
   wire signed [9:0] m94_71;
   assign m94_71 =10'b0;

   // m94_72 = W*in
   wire signed [9:0] m94_72;
   assign m94_72 ={ {5{neg94[5]}} , neg94[5:1] };

   // m94_73 = W*in
   wire signed [9:0] m94_73;
   assign m94_73 ={ {5{neg94[5]}} , neg94[5:1] };

   // m94_74 = W*in
   wire signed [9:0] m94_74;
   assign m94_74 =10'b0;

   // m94_75 = W*in
   wire signed [9:0] m94_75;
   assign m94_75 =10'b0;

   // m94_76 = W*in
   wire signed [9:0] m94_76;
   assign m94_76 =10'b0;

   // m94_77 = W*in
   wire signed [9:0] m94_77;
   assign m94_77 ={ {4{in94[5]}} , in94[5:0] };

   // m94_78 = W*in
   wire signed [9:0] m94_78;
   assign m94_78 =10'b0;

   // m94_79 = W*in
   wire signed [9:0] m94_79;
   assign m94_79 =10'b0;

   // m94_80 = W*in
   wire signed [9:0] m94_80;
   assign m94_80 =10'b0;

   // m94_81 = W*in
   wire signed [9:0] m94_81;
   assign m94_81 ={ {5{in94[5]}} , in94[5:1] };

   // m94_82 = W*in
   wire signed [9:0] m94_82;
   assign m94_82 =10'b0;

   // m94_83 = W*in
   wire signed [9:0] m94_83;
   assign m94_83 =10'b0;

   // m94_84 = W*in
   wire signed [9:0] m94_84;
   assign m94_84 =10'b0;

   // m94_85 = W*in
   wire signed [9:0] m94_85;
   assign m94_85 =10'b0;

   // m94_86 = W*in
   wire signed [9:0] m94_86;
   assign m94_86 =10'b0;

   // m94_87 = W*in
   wire signed [9:0] m94_87;
   assign m94_87 =10'b0;

   // m94_88 = W*in
   wire signed [9:0] m94_88;
   assign m94_88 =10'b0;

   // m94_89 = W*in
   wire signed [9:0] m94_89;
   assign m94_89 =10'b0;

   // m94_90 = W*in
   wire signed [9:0] m94_90;
   assign m94_90 =10'b0;

   // m94_91 = W*in
   wire signed [9:0] m94_91;
   assign m94_91 ={ {4{in94[5]}} , in94[5:0] };

   // m94_92 = W*in
   wire signed [9:0] m94_92;
   assign m94_92 =10'b0;

   // m94_93 = W*in
   wire signed [9:0] m94_93;
   assign m94_93 =10'b0;

   // m94_94 = W*in
   wire signed [9:0] m94_94;
   assign m94_94 =10'b0;

   // m94_95 = W*in
   wire signed [9:0] m94_95;
   assign m94_95 =10'b0;

   // m94_96 = W*in
   wire signed [9:0] m94_96;
   assign m94_96 =10'b0;

   // m94_97 = W*in
   wire signed [9:0] m94_97;
   assign m94_97 ={ {4{in94[5]}} , in94[5:0] };

   // m94_98 = W*in
   wire signed [9:0] m94_98;
   assign m94_98 =10'b0;

   // m94_99 = W*in
   wire signed [9:0] m94_99;
   assign m94_99 =10'b0;

   // m94_100 = W*in
   wire signed [9:0] m94_100;
   assign m94_100 =10'b0;

   // m94_101 = W*in
   wire signed [9:0] m94_101;
   assign m94_101 =10'b0;

   // m94_102 = W*in
   wire signed [9:0] m94_102;
   assign m94_102 =10'b0;

   // m94_103 = W*in
   wire signed [9:0] m94_103;
   assign m94_103 =10'b0;

   // m94_104 = W*in
   wire signed [9:0] m94_104;
   assign m94_104 =10'b0;

   // m94_105 = W*in
   wire signed [9:0] m94_105;
   assign m94_105 =10'b0;

   // m94_106 = W*in
   wire signed [9:0] m94_106;
   assign m94_106 =10'b0;

   // m94_107 = W*in
   wire signed [9:0] m94_107;
   assign m94_107 =10'b0;

   // m94_108 = W*in
   wire signed [9:0] m94_108;
   assign m94_108 ={ {5{in94[5]}} , in94[5:1] };

   // m94_109 = W*in
   wire signed [9:0] m94_109;
   assign m94_109 =10'b0;

   // m94_110 = W*in
   wire signed [9:0] m94_110;
   assign m94_110 =10'b0;

   // m94_111 = W*in
   wire signed [9:0] m94_111;
   assign m94_111 =10'b0;

   // m94_112 = W*in
   wire signed [9:0] m94_112;
   assign m94_112 =10'b0;

   // m94_113 = W*in
   wire signed [9:0] m94_113;
   assign m94_113 =10'b0;

   // m94_114 = W*in
   wire signed [9:0] m94_114;
   assign m94_114 =10'b0;

   // m94_115 = W*in
   wire signed [9:0] m94_115;
   assign m94_115 =10'b0;

   // m94_116 = W*in
   wire signed [9:0] m94_116;
   assign m94_116 =10'b0;

   // m94_117 = W*in
   wire signed [9:0] m94_117;
   assign m94_117 =10'b0;

   // m95_1 = W*in
   wire signed [9:0] m95_1;
   assign m95_1 =10'b0;

   // m95_2 = W*in
   wire signed [9:0] m95_2;
   assign m95_2 =10'b0;

   // m95_3 = W*in
   wire signed [9:0] m95_3;
   assign m95_3 =10'b0;

   // m95_4 = W*in
   wire signed [9:0] m95_4;
   assign m95_4 =10'b0;

   // m95_5 = W*in
   wire signed [9:0] m95_5;
   assign m95_5 =10'b0;

   // m95_6 = W*in
   wire signed [9:0] m95_6;
   assign m95_6 =10'b0;

   // m95_7 = W*in
   wire signed [9:0] m95_7;
   assign m95_7 =10'b0;

   // m95_8 = W*in
   wire signed [9:0] m95_8;
   assign m95_8 =10'b0;

   // m95_9 = W*in
   wire signed [9:0] m95_9;
   assign m95_9 =10'b0;

   // m95_10 = W*in
   wire signed [9:0] m95_10;
   assign m95_10 =10'b0;

   // m95_11 = W*in
   wire signed [9:0] m95_11;
   assign m95_11 =10'b0;

   // m95_12 = W*in
   wire signed [9:0] m95_12;
   assign m95_12 =10'b0;

   // m95_13 = W*in
   wire signed [9:0] m95_13;
   assign m95_13 =10'b0;

   // m95_14 = W*in
   wire signed [9:0] m95_14;
   assign m95_14 =10'b0;

   // m95_15 = W*in
   wire signed [9:0] m95_15;
   assign m95_15 =10'b0;

   // m95_16 = W*in
   wire signed [9:0] m95_16;
   assign m95_16 =10'b0;

   // m95_17 = W*in
   wire signed [9:0] m95_17;
   assign m95_17 =10'b0;

   // m95_18 = W*in
   wire signed [9:0] m95_18;
   assign m95_18 =10'b0;

   // m95_19 = W*in
   wire signed [9:0] m95_19;
   assign m95_19 =10'b0;

   // m95_20 = W*in
   wire signed [9:0] m95_20;
   assign m95_20 =10'b0;

   // m95_21 = W*in
   wire signed [9:0] m95_21;
   assign m95_21 =10'b0;

   // m95_22 = W*in
   wire signed [9:0] m95_22;
   assign m95_22 =10'b0;

   // m95_23 = W*in
   wire signed [9:0] m95_23;
   assign m95_23 =10'b0;

   // m95_24 = W*in
   wire signed [9:0] m95_24;
   assign m95_24 =10'b0;

   // m95_25 = W*in
   wire signed [9:0] m95_25;
   assign m95_25 =10'b0;

   // m95_26 = W*in
   wire signed [9:0] m95_26;
   assign m95_26 =10'b0;

   // m95_27 = W*in
   wire signed [9:0] m95_27;
   assign m95_27 =10'b0;

   // m95_28 = W*in
   wire signed [9:0] m95_28;
   assign m95_28 =10'b0;

   // m95_29 = W*in
   wire signed [9:0] m95_29;
   assign m95_29 =10'b0;

   // m95_30 = W*in
   wire signed [9:0] m95_30;
   assign m95_30 =10'b0;

   // m95_31 = W*in
   wire signed [9:0] m95_31;
   assign m95_31 =10'b0;

   // m95_32 = W*in
   wire signed [9:0] m95_32;
   assign m95_32 =10'b0;

   // m95_33 = W*in
   wire signed [9:0] m95_33;
   assign m95_33 =10'b0;

   // m95_34 = W*in
   wire signed [9:0] m95_34;
   assign m95_34 =10'b0;

   // m95_35 = W*in
   wire signed [9:0] m95_35;
   assign m95_35 =10'b0;

   // m95_36 = W*in
   wire signed [9:0] m95_36;
   assign m95_36 =10'b0;

   // m95_37 = W*in
   wire signed [9:0] m95_37;
   assign m95_37 =10'b0;

   // m95_38 = W*in
   wire signed [9:0] m95_38;
   assign m95_38 =10'b0;

   // m95_39 = W*in
   wire signed [9:0] m95_39;
   assign m95_39 =10'b0;

   // m95_40 = W*in
   wire signed [9:0] m95_40;
   assign m95_40 =10'b0;

   // m95_41 = W*in
   wire signed [9:0] m95_41;
   assign m95_41 =10'b0;

   // m95_42 = W*in
   wire signed [9:0] m95_42;
   assign m95_42 =10'b0;

   // m95_43 = W*in
   wire signed [9:0] m95_43;
   assign m95_43 =10'b0;

   // m95_44 = W*in
   wire signed [9:0] m95_44;
   assign m95_44 =10'b0;

   // m95_45 = W*in
   wire signed [9:0] m95_45;
   assign m95_45 =10'b0;

   // m95_46 = W*in
   wire signed [9:0] m95_46;
   assign m95_46 =10'b0;

   // m95_47 = W*in
   wire signed [9:0] m95_47;
   assign m95_47 =10'b0;

   // m95_48 = W*in
   wire signed [9:0] m95_48;
   assign m95_48 =10'b0;

   // m95_49 = W*in
   wire signed [9:0] m95_49;
   assign m95_49 =10'b0;

   // m95_50 = W*in
   wire signed [9:0] m95_50;
   assign m95_50 =10'b0;

   // m95_51 = W*in
   wire signed [9:0] m95_51;
   assign m95_51 =10'b0;

   // m95_52 = W*in
   wire signed [9:0] m95_52;
   assign m95_52 =10'b0;

   // m95_53 = W*in
   wire signed [9:0] m95_53;
   assign m95_53 =10'b0;

   // m95_54 = W*in
   wire signed [9:0] m95_54;
   assign m95_54 =10'b0;

   // m95_55 = W*in
   wire signed [9:0] m95_55;
   assign m95_55 =10'b0;

   // m95_56 = W*in
   wire signed [9:0] m95_56;
   assign m95_56 =10'b0;

   // m95_57 = W*in
   wire signed [9:0] m95_57;
   assign m95_57 =10'b0;

   // m95_58 = W*in
   wire signed [9:0] m95_58;
   assign m95_58 =10'b0;

   // m95_59 = W*in
   wire signed [9:0] m95_59;
   assign m95_59 =10'b0;

   // m95_60 = W*in
   wire signed [9:0] m95_60;
   assign m95_60 =10'b0;

   // m95_61 = W*in
   wire signed [9:0] m95_61;
   assign m95_61 =10'b0;

   // m95_62 = W*in
   wire signed [9:0] m95_62;
   assign m95_62 =10'b0;

   // m95_63 = W*in
   wire signed [9:0] m95_63;
   assign m95_63 =10'b0;

   // m95_64 = W*in
   wire signed [9:0] m95_64;
   assign m95_64 =10'b0;

   // m95_65 = W*in
   wire signed [9:0] m95_65;
   assign m95_65 =10'b0;

   // m95_66 = W*in
   wire signed [9:0] m95_66;
   assign m95_66 =10'b0;

   // m95_67 = W*in
   wire signed [9:0] m95_67;
   assign m95_67 =10'b0;

   // m95_68 = W*in
   wire signed [9:0] m95_68;
   assign m95_68 =10'b0;

   // m95_69 = W*in
   wire signed [9:0] m95_69;
   assign m95_69 =10'b0;

   // m95_70 = W*in
   wire signed [9:0] m95_70;
   assign m95_70 =10'b0;

   // m95_71 = W*in
   wire signed [9:0] m95_71;
   assign m95_71 =10'b0;

   // m95_72 = W*in
   wire signed [9:0] m95_72;
   assign m95_72 =10'b0;

   // m95_73 = W*in
   wire signed [9:0] m95_73;
   assign m95_73 =10'b0;

   // m95_74 = W*in
   wire signed [9:0] m95_74;
   assign m95_74 =10'b0;

   // m95_75 = W*in
   wire signed [9:0] m95_75;
   assign m95_75 =10'b0;

   // m95_76 = W*in
   wire signed [9:0] m95_76;
   assign m95_76 =10'b0;

   // m95_77 = W*in
   wire signed [9:0] m95_77;
   assign m95_77 =10'b0;

   // m95_78 = W*in
   wire signed [9:0] m95_78;
   assign m95_78 =10'b0;

   // m95_79 = W*in
   wire signed [9:0] m95_79;
   assign m95_79 =10'b0;

   // m95_80 = W*in
   wire signed [9:0] m95_80;
   assign m95_80 =10'b0;

   // m95_81 = W*in
   wire signed [9:0] m95_81;
   assign m95_81 =10'b0;

   // m95_82 = W*in
   wire signed [9:0] m95_82;
   assign m95_82 =10'b0;

   // m95_83 = W*in
   wire signed [9:0] m95_83;
   assign m95_83 =10'b0;

   // m95_84 = W*in
   wire signed [9:0] m95_84;
   assign m95_84 =10'b0;

   // m95_85 = W*in
   wire signed [9:0] m95_85;
   assign m95_85 =10'b0;

   // m95_86 = W*in
   wire signed [9:0] m95_86;
   assign m95_86 =10'b0;

   // m95_87 = W*in
   wire signed [9:0] m95_87;
   assign m95_87 =10'b0;

   // m95_88 = W*in
   wire signed [9:0] m95_88;
   assign m95_88 =10'b0;

   // m95_89 = W*in
   wire signed [9:0] m95_89;
   assign m95_89 =10'b0;

   // m95_90 = W*in
   wire signed [9:0] m95_90;
   assign m95_90 =10'b0;

   // m95_91 = W*in
   wire signed [9:0] m95_91;
   assign m95_91 =10'b0;

   // m95_92 = W*in
   wire signed [9:0] m95_92;
   assign m95_92 =10'b0;

   // m95_93 = W*in
   wire signed [9:0] m95_93;
   assign m95_93 =10'b0;

   // m95_94 = W*in
   wire signed [9:0] m95_94;
   assign m95_94 =10'b0;

   // m95_95 = W*in
   wire signed [9:0] m95_95;
   assign m95_95 =10'b0;

   // m95_96 = W*in
   wire signed [9:0] m95_96;
   assign m95_96 =10'b0;

   // m95_97 = W*in
   wire signed [9:0] m95_97;
   assign m95_97 =10'b0;

   // m95_98 = W*in
   wire signed [9:0] m95_98;
   assign m95_98 =10'b0;

   // m95_99 = W*in
   wire signed [9:0] m95_99;
   assign m95_99 =10'b0;

   // m95_100 = W*in
   wire signed [9:0] m95_100;
   assign m95_100 =10'b0;

   // m95_101 = W*in
   wire signed [9:0] m95_101;
   assign m95_101 =10'b0;

   // m95_102 = W*in
   wire signed [9:0] m95_102;
   assign m95_102 =10'b0;

   // m95_103 = W*in
   wire signed [9:0] m95_103;
   assign m95_103 =10'b0;

   // m95_104 = W*in
   wire signed [9:0] m95_104;
   assign m95_104 =10'b0;

   // m95_105 = W*in
   wire signed [9:0] m95_105;
   assign m95_105 =10'b0;

   // m95_106 = W*in
   wire signed [9:0] m95_106;
   assign m95_106 =10'b0;

   // m95_107 = W*in
   wire signed [9:0] m95_107;
   assign m95_107 =10'b0;

   // m95_108 = W*in
   wire signed [9:0] m95_108;
   assign m95_108 ={ {5{in95[5]}} , in95[5:1] };

   // m95_109 = W*in
   wire signed [9:0] m95_109;
   assign m95_109 =10'b0;

   // m95_110 = W*in
   wire signed [9:0] m95_110;
   assign m95_110 =10'b0;

   // m95_111 = W*in
   wire signed [9:0] m95_111;
   assign m95_111 =10'b0;

   // m95_112 = W*in
   wire signed [9:0] m95_112;
   assign m95_112 =10'b0;

   // m95_113 = W*in
   wire signed [9:0] m95_113;
   assign m95_113 =10'b0;

   // m95_114 = W*in
   wire signed [9:0] m95_114;
   assign m95_114 =10'b0;

   // m95_115 = W*in
   wire signed [9:0] m95_115;
   assign m95_115 =10'b0;

   // m95_116 = W*in
   wire signed [9:0] m95_116;
   assign m95_116 =10'b0;

   // m95_117 = W*in
   wire signed [9:0] m95_117;
   assign m95_117 =10'b0;

   // m96_1 = W*in
   wire signed [9:0] m96_1;
   assign m96_1 ={ {4{in96[5]}} , in96[5:0] };

   // m96_2 = W*in
   wire signed [9:0] m96_2;
   assign m96_2 =10'b0;

   // m96_3 = W*in
   wire signed [9:0] m96_3;
   assign m96_3 =10'b0;

   // m96_4 = W*in
   wire signed [9:0] m96_4;
   assign m96_4 =10'b0;

   // m96_5 = W*in
   wire signed [9:0] m96_5;
   assign m96_5 =10'b0;

   // m96_6 = W*in
   wire signed [9:0] m96_6;
   assign m96_6 ={ {4{neg96[5]}} , neg96[5:0] };

   // m96_7 = W*in
   wire signed [9:0] m96_7;
   assign m96_7 =10'b0;

   // m96_8 = W*in
   wire signed [9:0] m96_8;
   assign m96_8 =10'b0;

   // m96_9 = W*in
   wire signed [9:0] m96_9;
   assign m96_9 =10'b0;

   // m96_10 = W*in
   wire signed [9:0] m96_10;
   assign m96_10 =10'b0;

   // m96_11 = W*in
   wire signed [9:0] m96_11;
   assign m96_11 =10'b0;

   // m96_12 = W*in
   wire signed [9:0] m96_12;
   assign m96_12 =10'b0;

   // m96_13 = W*in
   wire signed [9:0] m96_13;
   assign m96_13 =10'b0;

   // m96_14 = W*in
   wire signed [9:0] m96_14;
   assign m96_14 =10'b0;

   // m96_15 = W*in
   wire signed [9:0] m96_15;
   assign m96_15 =10'b0;

   // m96_16 = W*in
   wire signed [9:0] m96_16;
   assign m96_16 ={ {4{in96[5]}} , in96[5:0] };

   // m96_17 = W*in
   wire signed [9:0] m96_17;
   assign m96_17 =10'b0;

   // m96_18 = W*in
   wire signed [9:0] m96_18;
   assign m96_18 ={ {5{neg96[5]}} , neg96[5:1] };

   // m96_19 = W*in
   wire signed [9:0] m96_19;
   assign m96_19 =10'b0;

   // m96_20 = W*in
   wire signed [9:0] m96_20;
   assign m96_20 ={ {4{in96[5]}} , in96[5:0] };

   // m96_21 = W*in
   wire signed [9:0] m96_21;
   assign m96_21 ={ {5{neg96[5]}} , neg96[5:1] };

   // m96_22 = W*in
   wire signed [9:0] m96_22;
   assign m96_22 =10'b0;

   // m96_23 = W*in
   wire signed [9:0] m96_23;
   assign m96_23 =10'b0;

   // m96_24 = W*in
   wire signed [9:0] m96_24;
   assign m96_24 =10'b0;

   // m96_25 = W*in
   wire signed [9:0] m96_25;
   assign m96_25 ={ {4{in96[5]}} , in96[5:0] };

   // m96_26 = W*in
   wire signed [9:0] m96_26;
   assign m96_26 =10'b0;

   // m96_27 = W*in
   wire signed [9:0] m96_27;
   assign m96_27 ={ {5{neg96[5]}} , neg96[5:1] };

   // m96_28 = W*in
   wire signed [9:0] m96_28;
   assign m96_28 =10'b0;

   // m96_29 = W*in
   wire signed [9:0] m96_29;
   assign m96_29 =10'b0;

   // m96_30 = W*in
   wire signed [9:0] m96_30;
   assign m96_30 ={ {4{in96[5]}} , in96[5:0] };

   // m96_31 = W*in
   wire signed [9:0] m96_31;
   assign m96_31 =10'b0;

   // m96_32 = W*in
   wire signed [9:0] m96_32;
   assign m96_32 =10'b0;

   // m96_33 = W*in
   wire signed [9:0] m96_33;
   assign m96_33 =10'b0;

   // m96_34 = W*in
   wire signed [9:0] m96_34;
   assign m96_34 =10'b0;

   // m96_35 = W*in
   wire signed [9:0] m96_35;
   assign m96_35 ={ {5{in96[5]}} , in96[5:1] };

   // m96_36 = W*in
   wire signed [9:0] m96_36;
   assign m96_36 =10'b0;

   // m96_37 = W*in
   wire signed [9:0] m96_37;
   assign m96_37 =10'b0;

   // m96_38 = W*in
   wire signed [9:0] m96_38;
   assign m96_38 =10'b0;

   // m96_39 = W*in
   wire signed [9:0] m96_39;
   assign m96_39 =10'b0;

   // m96_40 = W*in
   wire signed [9:0] m96_40;
   assign m96_40 =10'b0;

   // m96_41 = W*in
   wire signed [9:0] m96_41;
   assign m96_41 =10'b0;

   // m96_42 = W*in
   wire signed [9:0] m96_42;
   assign m96_42 ={ {4{in96[5]}} , in96[5:0] };

   // m96_43 = W*in
   wire signed [9:0] m96_43;
   assign m96_43 =10'b0;

   // m96_44 = W*in
   wire signed [9:0] m96_44;
   assign m96_44 =10'b0;

   // m96_45 = W*in
   wire signed [9:0] m96_45;
   assign m96_45 =10'b0;

   // m96_46 = W*in
   wire signed [9:0] m96_46;
   assign m96_46 =10'b0;

   // m96_47 = W*in
   wire signed [9:0] m96_47;
   assign m96_47 =10'b0;

   // m96_48 = W*in
   wire signed [9:0] m96_48;
   assign m96_48 =10'b0;

   // m96_49 = W*in
   wire signed [9:0] m96_49;
   assign m96_49 =10'b0;

   // m96_50 = W*in
   wire signed [9:0] m96_50;
   assign m96_50 =10'b0;

   // m96_51 = W*in
   wire signed [9:0] m96_51;
   assign m96_51 =10'b0;

   // m96_52 = W*in
   wire signed [9:0] m96_52;
   assign m96_52 =10'b0;

   // m96_53 = W*in
   wire signed [9:0] m96_53;
   assign m96_53 =10'b0;

   // m96_54 = W*in
   wire signed [9:0] m96_54;
   assign m96_54 =10'b0;

   // m96_55 = W*in
   wire signed [9:0] m96_55;
   assign m96_55 =10'b0;

   // m96_56 = W*in
   wire signed [9:0] m96_56;
   assign m96_56 ={ {4{in96[5]}} , in96[5:0] };

   // m96_57 = W*in
   wire signed [9:0] m96_57;
   assign m96_57 =10'b0;

   // m96_58 = W*in
   wire signed [9:0] m96_58;
   assign m96_58 =10'b0;

   // m96_59 = W*in
   wire signed [9:0] m96_59;
   assign m96_59 =10'b0;

   // m96_60 = W*in
   wire signed [9:0] m96_60;
   assign m96_60 =10'b0;

   // m96_61 = W*in
   wire signed [9:0] m96_61;
   assign m96_61 =10'b0;

   // m96_62 = W*in
   wire signed [9:0] m96_62;
   assign m96_62 =10'b0;

   // m96_63 = W*in
   wire signed [9:0] m96_63;
   assign m96_63 =10'b0;

   // m96_64 = W*in
   wire signed [9:0] m96_64;
   assign m96_64 =10'b0;

   // m96_65 = W*in
   wire signed [9:0] m96_65;
   assign m96_65 =10'b0;

   // m96_66 = W*in
   wire signed [9:0] m96_66;
   assign m96_66 =10'b0;

   // m96_67 = W*in
   wire signed [9:0] m96_67;
   assign m96_67 =10'b0;

   // m96_68 = W*in
   wire signed [9:0] m96_68;
   assign m96_68 =10'b0;

   // m96_69 = W*in
   wire signed [9:0] m96_69;
   assign m96_69 ={ {4{neg96[5]}} , neg96[5:0] };

   // m96_70 = W*in
   wire signed [9:0] m96_70;
   assign m96_70 =10'b0;

   // m96_71 = W*in
   wire signed [9:0] m96_71;
   assign m96_71 ={ {5{neg96[5]}} , neg96[5:1] };

   // m96_72 = W*in
   wire signed [9:0] m96_72;
   assign m96_72 =10'b0;

   // m96_73 = W*in
   wire signed [9:0] m96_73;
   assign m96_73 =10'b0;

   // m96_74 = W*in
   wire signed [9:0] m96_74;
   assign m96_74 ={ {5{neg96[5]}} , neg96[5:1] };

   // m96_75 = W*in
   wire signed [9:0] m96_75;
   assign m96_75 =10'b0;

   // m96_76 = W*in
   wire signed [9:0] m96_76;
   assign m96_76 =10'b0;

   // m96_77 = W*in
   wire signed [9:0] m96_77;
   assign m96_77 =10'b0;

   // m96_78 = W*in
   wire signed [9:0] m96_78;
   assign m96_78 =10'b0;

   // m96_79 = W*in
   wire signed [9:0] m96_79;
   assign m96_79 ={ {4{in96[5]}} , in96[5:0] };

   // m96_80 = W*in
   wire signed [9:0] m96_80;
   assign m96_80 =10'b0;

   // m96_81 = W*in
   wire signed [9:0] m96_81;
   assign m96_81 ={ {4{in96[5]}} , in96[5:0] };

   // m96_82 = W*in
   wire signed [9:0] m96_82;
   assign m96_82 ={ {5{neg96[5]}} , neg96[5:1] };

   // m96_83 = W*in
   wire signed [9:0] m96_83;
   assign m96_83 =10'b0;

   // m96_84 = W*in
   wire signed [9:0] m96_84;
   assign m96_84 =10'b0;

   // m96_85 = W*in
   wire signed [9:0] m96_85;
   assign m96_85 =10'b0;

   // m96_86 = W*in
   wire signed [9:0] m96_86;
   assign m96_86 =10'b0;

   // m96_87 = W*in
   wire signed [9:0] m96_87;
   assign m96_87 ={ {4{neg96[5]}} , neg96[5:0] };

   // m96_88 = W*in
   wire signed [9:0] m96_88;
   assign m96_88 ={ {4{neg96[5]}} , neg96[5:0] };

   // m96_89 = W*in
   wire signed [9:0] m96_89;
   assign m96_89 =10'b0;

   // m96_90 = W*in
   wire signed [9:0] m96_90;
   assign m96_90 =10'b0;

   // m96_91 = W*in
   wire signed [9:0] m96_91;
   assign m96_91 =10'b0;

   // m96_92 = W*in
   wire signed [9:0] m96_92;
   assign m96_92 =10'b0;

   // m96_93 = W*in
   wire signed [9:0] m96_93;
   assign m96_93 =10'b0;

   // m96_94 = W*in
   wire signed [9:0] m96_94;
   assign m96_94 ={ {4{in96[5]}} , in96[5:0] };

   // m96_95 = W*in
   wire signed [9:0] m96_95;
   assign m96_95 =10'b0;

   // m96_96 = W*in
   wire signed [9:0] m96_96;
   assign m96_96 =10'b0;

   // m96_97 = W*in
   wire signed [9:0] m96_97;
   assign m96_97 =10'b0;

   // m96_98 = W*in
   wire signed [9:0] m96_98;
   assign m96_98 =10'b0;

   // m96_99 = W*in
   wire signed [9:0] m96_99;
   assign m96_99 =10'b0;

   // m96_100 = W*in
   wire signed [9:0] m96_100;
   assign m96_100 ={ {4{in96[5]}} , in96[5:0] };

   // m96_101 = W*in
   wire signed [9:0] m96_101;
   assign m96_101 =10'b0;

   // m96_102 = W*in
   wire signed [9:0] m96_102;
   assign m96_102 =10'b0;

   // m96_103 = W*in
   wire signed [9:0] m96_103;
   assign m96_103 =10'b0;

   // m96_104 = W*in
   wire signed [9:0] m96_104;
   assign m96_104 =10'b0;

   // m96_105 = W*in
   wire signed [9:0] m96_105;
   assign m96_105 =10'b0;

   // m96_106 = W*in
   wire signed [9:0] m96_106;
   assign m96_106 ={ {4{in96[5]}} , in96[5:0] };

   // m96_107 = W*in
   wire signed [9:0] m96_107;
   assign m96_107 =10'b0;

   // m96_108 = W*in
   wire signed [9:0] m96_108;
   assign m96_108 ={ {5{in96[5]}} , in96[5:1] };

   // m96_109 = W*in
   wire signed [9:0] m96_109;
   assign m96_109 =10'b0;

   // m96_110 = W*in
   wire signed [9:0] m96_110;
   assign m96_110 =10'b0;

   // m96_111 = W*in
   wire signed [9:0] m96_111;
   assign m96_111 ={ {4{in96[5]}} , in96[5:0] };

   // m96_112 = W*in
   wire signed [9:0] m96_112;
   assign m96_112 =10'b0;

   // m96_113 = W*in
   wire signed [9:0] m96_113;
   assign m96_113 ={ {4{in96[5]}} , in96[5:0] };

   // m96_114 = W*in
   wire signed [9:0] m96_114;
   assign m96_114 =10'b0;

   // m96_115 = W*in
   wire signed [9:0] m96_115;
   assign m96_115 =10'b0;

   // m96_116 = W*in
   wire signed [9:0] m96_116;
   assign m96_116 ={ {4{in96[5]}} , in96[5:0] };

   // m96_117 = W*in
   wire signed [9:0] m96_117;
   assign m96_117 =10'b0;

   // m97_1 = W*in
   wire signed [9:0] m97_1;
   assign m97_1 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_2 = W*in
   wire signed [9:0] m97_2;
   assign m97_2 ={ {4{in97[5]}} , in97[5:0] };

   // m97_3 = W*in
   wire signed [9:0] m97_3;
   assign m97_3 =10'b0;

   // m97_4 = W*in
   wire signed [9:0] m97_4;
   assign m97_4 =10'b0;

   // m97_5 = W*in
   wire signed [9:0] m97_5;
   assign m97_5 =10'b0;

   // m97_6 = W*in
   wire signed [9:0] m97_6;
   assign m97_6 =10'b0;

   // m97_7 = W*in
   wire signed [9:0] m97_7;
   assign m97_7 ={ {4{in97[5]}} , in97[5:0] };

   // m97_8 = W*in
   wire signed [9:0] m97_8;
   assign m97_8 =10'b0;

   // m97_9 = W*in
   wire signed [9:0] m97_9;
   assign m97_9 =10'b0;

   // m97_10 = W*in
   wire signed [9:0] m97_10;
   assign m97_10 =10'b0;

   // m97_11 = W*in
   wire signed [9:0] m97_11;
   assign m97_11 =10'b0;

   // m97_12 = W*in
   wire signed [9:0] m97_12;
   assign m97_12 =10'b0;

   // m97_13 = W*in
   wire signed [9:0] m97_13;
   assign m97_13 ={ {4{in97[5]}} , in97[5:0] };

   // m97_14 = W*in
   wire signed [9:0] m97_14;
   assign m97_14 =10'b0;

   // m97_15 = W*in
   wire signed [9:0] m97_15;
   assign m97_15 =10'b0;

   // m97_16 = W*in
   wire signed [9:0] m97_16;
   assign m97_16 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_17 = W*in
   wire signed [9:0] m97_17;
   assign m97_17 =10'b0;

   // m97_18 = W*in
   wire signed [9:0] m97_18;
   assign m97_18 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_19 = W*in
   wire signed [9:0] m97_19;
   assign m97_19 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_20 = W*in
   wire signed [9:0] m97_20;
   assign m97_20 ={ {4{in97[5]}} , in97[5:0] };

   // m97_21 = W*in
   wire signed [9:0] m97_21;
   assign m97_21 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_22 = W*in
   wire signed [9:0] m97_22;
   assign m97_22 =10'b0;

   // m97_23 = W*in
   wire signed [9:0] m97_23;
   assign m97_23 =10'b0;

   // m97_24 = W*in
   wire signed [9:0] m97_24;
   assign m97_24 =10'b0;

   // m97_25 = W*in
   wire signed [9:0] m97_25;
   assign m97_25 =10'b0;

   // m97_26 = W*in
   wire signed [9:0] m97_26;
   assign m97_26 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_27 = W*in
   wire signed [9:0] m97_27;
   assign m97_27 =10'b0;

   // m97_28 = W*in
   wire signed [9:0] m97_28;
   assign m97_28 ={ {5{in97[5]}} , in97[5:1] };

   // m97_29 = W*in
   wire signed [9:0] m97_29;
   assign m97_29 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_30 = W*in
   wire signed [9:0] m97_30;
   assign m97_30 ={ {4{in97[5]}} , in97[5:0] };

   // m97_31 = W*in
   wire signed [9:0] m97_31;
   assign m97_31 =10'b0;

   // m97_32 = W*in
   wire signed [9:0] m97_32;
   assign m97_32 ={ {4{in97[5]}} , in97[5:0] };

   // m97_33 = W*in
   wire signed [9:0] m97_33;
   assign m97_33 ={ {4{in97[5]}} , in97[5:0] };

   // m97_34 = W*in
   wire signed [9:0] m97_34;
   assign m97_34 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_35 = W*in
   wire signed [9:0] m97_35;
   assign m97_35 =10'b0;

   // m97_36 = W*in
   wire signed [9:0] m97_36;
   assign m97_36 ={ {4{in97[5]}} , in97[5:0] };

   // m97_37 = W*in
   wire signed [9:0] m97_37;
   assign m97_37 ={ {5{in97[5]}} , in97[5:1] };

   // m97_38 = W*in
   wire signed [9:0] m97_38;
   assign m97_38 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_39 = W*in
   wire signed [9:0] m97_39;
   assign m97_39 =10'b0;

   // m97_40 = W*in
   wire signed [9:0] m97_40;
   assign m97_40 =10'b0;

   // m97_41 = W*in
   wire signed [9:0] m97_41;
   assign m97_41 ={ {4{in97[5]}} , in97[5:0] };

   // m97_42 = W*in
   wire signed [9:0] m97_42;
   assign m97_42 =10'b0;

   // m97_43 = W*in
   wire signed [9:0] m97_43;
   assign m97_43 =10'b0;

   // m97_44 = W*in
   wire signed [9:0] m97_44;
   assign m97_44 =10'b0;

   // m97_45 = W*in
   wire signed [9:0] m97_45;
   assign m97_45 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_46 = W*in
   wire signed [9:0] m97_46;
   assign m97_46 =10'b0;

   // m97_47 = W*in
   wire signed [9:0] m97_47;
   assign m97_47 =10'b0;

   // m97_48 = W*in
   wire signed [9:0] m97_48;
   assign m97_48 =10'b0;

   // m97_49 = W*in
   wire signed [9:0] m97_49;
   assign m97_49 =10'b0;

   // m97_50 = W*in
   wire signed [9:0] m97_50;
   assign m97_50 =10'b0;

   // m97_51 = W*in
   wire signed [9:0] m97_51;
   assign m97_51 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_52 = W*in
   wire signed [9:0] m97_52;
   assign m97_52 ={ {4{in97[5]}} , in97[5:0] };

   // m97_53 = W*in
   wire signed [9:0] m97_53;
   assign m97_53 =10'b0;

   // m97_54 = W*in
   wire signed [9:0] m97_54;
   assign m97_54 =10'b0;

   // m97_55 = W*in
   wire signed [9:0] m97_55;
   assign m97_55 =10'b0;

   // m97_56 = W*in
   wire signed [9:0] m97_56;
   assign m97_56 ={ {3{in97[5]}} , in97 , {1{1'b0}} };

   // m97_57 = W*in
   wire signed [9:0] m97_57;
   assign m97_57 =10'b0;

   // m97_58 = W*in
   wire signed [9:0] m97_58;
   assign m97_58 =10'b0;

   // m97_59 = W*in
   wire signed [9:0] m97_59;
   assign m97_59 ={ {4{in97[5]}} , in97[5:0] };

   // m97_60 = W*in
   wire signed [9:0] m97_60;
   assign m97_60 =10'b0;

   // m97_61 = W*in
   wire signed [9:0] m97_61;
   assign m97_61 ={ {4{in97[5]}} , in97[5:0] };

   // m97_62 = W*in
   wire signed [9:0] m97_62;
   assign m97_62 =10'b0;

   // m97_63 = W*in
   wire signed [9:0] m97_63;
   assign m97_63 =10'b0;

   // m97_64 = W*in
   wire signed [9:0] m97_64;
   assign m97_64 =10'b0;

   // m97_65 = W*in
   wire signed [9:0] m97_65;
   assign m97_65 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_66 = W*in
   wire signed [9:0] m97_66;
   assign m97_66 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_67 = W*in
   wire signed [9:0] m97_67;
   assign m97_67 =10'b0;

   // m97_68 = W*in
   wire signed [9:0] m97_68;
   assign m97_68 =10'b0;

   // m97_69 = W*in
   wire signed [9:0] m97_69;
   assign m97_69 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_70 = W*in
   wire signed [9:0] m97_70;
   assign m97_70 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_71 = W*in
   wire signed [9:0] m97_71;
   assign m97_71 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_72 = W*in
   wire signed [9:0] m97_72;
   assign m97_72 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_73 = W*in
   wire signed [9:0] m97_73;
   assign m97_73 ={ {4{in97[5]}} , in97[5:0] };

   // m97_74 = W*in
   wire signed [9:0] m97_74;
   assign m97_74 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_75 = W*in
   wire signed [9:0] m97_75;
   assign m97_75 =10'b0;

   // m97_76 = W*in
   wire signed [9:0] m97_76;
   assign m97_76 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_77 = W*in
   wire signed [9:0] m97_77;
   assign m97_77 =10'b0;

   // m97_78 = W*in
   wire signed [9:0] m97_78;
   assign m97_78 ={ {5{in97[5]}} , in97[5:1] };

   // m97_79 = W*in
   wire signed [9:0] m97_79;
   assign m97_79 =10'b0;

   // m97_80 = W*in
   wire signed [9:0] m97_80;
   assign m97_80 =10'b0;

   // m97_81 = W*in
   wire signed [9:0] m97_81;
   assign m97_81 ={ {5{in97[5]}} , in97[5:1] };

   // m97_82 = W*in
   wire signed [9:0] m97_82;
   assign m97_82 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_83 = W*in
   wire signed [9:0] m97_83;
   assign m97_83 ={ {4{in97[5]}} , in97[5:0] };

   // m97_84 = W*in
   wire signed [9:0] m97_84;
   assign m97_84 =10'b0;

   // m97_85 = W*in
   wire signed [9:0] m97_85;
   assign m97_85 ={ {4{in97[5]}} , in97[5:0] };

   // m97_86 = W*in
   wire signed [9:0] m97_86;
   assign m97_86 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_87 = W*in
   wire signed [9:0] m97_87;
   assign m97_87 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_88 = W*in
   wire signed [9:0] m97_88;
   assign m97_88 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_89 = W*in
   wire signed [9:0] m97_89;
   assign m97_89 =10'b0;

   // m97_90 = W*in
   wire signed [9:0] m97_90;
   assign m97_90 =10'b0;

   // m97_91 = W*in
   wire signed [9:0] m97_91;
   assign m97_91 =10'b0;

   // m97_92 = W*in
   wire signed [9:0] m97_92;
   assign m97_92 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_93 = W*in
   wire signed [9:0] m97_93;
   assign m97_93 =10'b0;

   // m97_94 = W*in
   wire signed [9:0] m97_94;
   assign m97_94 =10'b0;

   // m97_95 = W*in
   wire signed [9:0] m97_95;
   assign m97_95 =10'b0;

   // m97_96 = W*in
   wire signed [9:0] m97_96;
   assign m97_96 =10'b0;

   // m97_97 = W*in
   wire signed [9:0] m97_97;
   assign m97_97 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_98 = W*in
   wire signed [9:0] m97_98;
   assign m97_98 ={ {4{in97[5]}} , in97[5:0] };

   // m97_99 = W*in
   wire signed [9:0] m97_99;
   assign m97_99 ={ {3{neg97[5]}} , neg97 , {1{1'b0}} };

   // m97_100 = W*in
   wire signed [9:0] m97_100;
   assign m97_100 =10'b0;

   // m97_101 = W*in
   wire signed [9:0] m97_101;
   assign m97_101 ={ {4{neg97[5]}} , neg97[5:0] };

   // m97_102 = W*in
   wire signed [9:0] m97_102;
   assign m97_102 ={ {4{in97[5]}} , in97[5:0] };

   // m97_103 = W*in
   wire signed [9:0] m97_103;
   assign m97_103 =10'b0;

   // m97_104 = W*in
   wire signed [9:0] m97_104;
   assign m97_104 =10'b0;

   // m97_105 = W*in
   wire signed [9:0] m97_105;
   assign m97_105 =10'b0;

   // m97_106 = W*in
   wire signed [9:0] m97_106;
   assign m97_106 ={ {4{in97[5]}} , in97[5:0] };

   // m97_107 = W*in
   wire signed [9:0] m97_107;
   assign m97_107 =10'b0;

   // m97_108 = W*in
   wire signed [9:0] m97_108;
   assign m97_108 =10'b0;

   // m97_109 = W*in
   wire signed [9:0] m97_109;
   assign m97_109 =10'b0;

   // m97_110 = W*in
   wire signed [9:0] m97_110;
   assign m97_110 =10'b0;

   // m97_111 = W*in
   wire signed [9:0] m97_111;
   assign m97_111 ={ {4{in97[5]}} , in97[5:0] };

   // m97_112 = W*in
   wire signed [9:0] m97_112;
   assign m97_112 =10'b0;

   // m97_113 = W*in
   wire signed [9:0] m97_113;
   assign m97_113 ={ {4{in97[5]}} , in97[5:0] };

   // m97_114 = W*in
   wire signed [9:0] m97_114;
   assign m97_114 ={ {5{neg97[5]}} , neg97[5:1] };

   // m97_115 = W*in
   wire signed [9:0] m97_115;
   assign m97_115 ={ {4{in97[5]}} , in97[5:0] };

   // m97_116 = W*in
   wire signed [9:0] m97_116;
   assign m97_116 ={ {4{in97[5]}} , in97[5:0] };

   // m97_117 = W*in
   wire signed [9:0] m97_117;
   assign m97_117 =10'b0;

   // m98_1 = W*in
   wire signed [9:0] m98_1;
   assign m98_1 ={ {4{in98[5]}} , in98[5:0] };

   // m98_2 = W*in
   wire signed [9:0] m98_2;
   assign m98_2 =10'b0;

   // m98_3 = W*in
   wire signed [9:0] m98_3;
   assign m98_3 =10'b0;

   // m98_4 = W*in
   wire signed [9:0] m98_4;
   assign m98_4 =10'b0;

   // m98_5 = W*in
   wire signed [9:0] m98_5;
   assign m98_5 ={ {4{in98[5]}} , in98[5:0] };

   // m98_6 = W*in
   wire signed [9:0] m98_6;
   assign m98_6 =10'b0;

   // m98_7 = W*in
   wire signed [9:0] m98_7;
   assign m98_7 ={ {4{in98[5]}} , in98[5:0] };

   // m98_8 = W*in
   wire signed [9:0] m98_8;
   assign m98_8 =10'b0;

   // m98_9 = W*in
   wire signed [9:0] m98_9;
   assign m98_9 =10'b0;

   // m98_10 = W*in
   wire signed [9:0] m98_10;
   assign m98_10 =10'b0;

   // m98_11 = W*in
   wire signed [9:0] m98_11;
   assign m98_11 =10'b0;

   // m98_12 = W*in
   wire signed [9:0] m98_12;
   assign m98_12 ={ {4{neg98[5]}} , neg98[5:0] };

   // m98_13 = W*in
   wire signed [9:0] m98_13;
   assign m98_13 ={ {4{in98[5]}} , in98[5:0] };

   // m98_14 = W*in
   wire signed [9:0] m98_14;
   assign m98_14 =10'b0;

   // m98_15 = W*in
   wire signed [9:0] m98_15;
   assign m98_15 =10'b0;

   // m98_16 = W*in
   wire signed [9:0] m98_16;
   assign m98_16 ={ {4{in98[5]}} , in98[5:0] };

   // m98_17 = W*in
   wire signed [9:0] m98_17;
   assign m98_17 =10'b0;

   // m98_18 = W*in
   wire signed [9:0] m98_18;
   assign m98_18 =10'b0;

   // m98_19 = W*in
   wire signed [9:0] m98_19;
   assign m98_19 =10'b0;

   // m98_20 = W*in
   wire signed [9:0] m98_20;
   assign m98_20 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_21 = W*in
   wire signed [9:0] m98_21;
   assign m98_21 =10'b0;

   // m98_22 = W*in
   wire signed [9:0] m98_22;
   assign m98_22 =10'b0;

   // m98_23 = W*in
   wire signed [9:0] m98_23;
   assign m98_23 =10'b0;

   // m98_24 = W*in
   wire signed [9:0] m98_24;
   assign m98_24 =10'b0;

   // m98_25 = W*in
   wire signed [9:0] m98_25;
   assign m98_25 ={ {4{in98[5]}} , in98[5:0] };

   // m98_26 = W*in
   wire signed [9:0] m98_26;
   assign m98_26 =10'b0;

   // m98_27 = W*in
   wire signed [9:0] m98_27;
   assign m98_27 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_28 = W*in
   wire signed [9:0] m98_28;
   assign m98_28 =10'b0;

   // m98_29 = W*in
   wire signed [9:0] m98_29;
   assign m98_29 =10'b0;

   // m98_30 = W*in
   wire signed [9:0] m98_30;
   assign m98_30 =10'b0;

   // m98_31 = W*in
   wire signed [9:0] m98_31;
   assign m98_31 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_32 = W*in
   wire signed [9:0] m98_32;
   assign m98_32 =10'b0;

   // m98_33 = W*in
   wire signed [9:0] m98_33;
   assign m98_33 ={ {4{in98[5]}} , in98[5:0] };

   // m98_34 = W*in
   wire signed [9:0] m98_34;
   assign m98_34 =10'b0;

   // m98_35 = W*in
   wire signed [9:0] m98_35;
   assign m98_35 =10'b0;

   // m98_36 = W*in
   wire signed [9:0] m98_36;
   assign m98_36 ={ {5{in98[5]}} , in98[5:1] };

   // m98_37 = W*in
   wire signed [9:0] m98_37;
   assign m98_37 =10'b0;

   // m98_38 = W*in
   wire signed [9:0] m98_38;
   assign m98_38 =10'b0;

   // m98_39 = W*in
   wire signed [9:0] m98_39;
   assign m98_39 =10'b0;

   // m98_40 = W*in
   wire signed [9:0] m98_40;
   assign m98_40 =10'b0;

   // m98_41 = W*in
   wire signed [9:0] m98_41;
   assign m98_41 =10'b0;

   // m98_42 = W*in
   wire signed [9:0] m98_42;
   assign m98_42 =10'b0;

   // m98_43 = W*in
   wire signed [9:0] m98_43;
   assign m98_43 =10'b0;

   // m98_44 = W*in
   wire signed [9:0] m98_44;
   assign m98_44 =10'b0;

   // m98_45 = W*in
   wire signed [9:0] m98_45;
   assign m98_45 ={ {4{in98[5]}} , in98[5:0] };

   // m98_46 = W*in
   wire signed [9:0] m98_46;
   assign m98_46 =10'b0;

   // m98_47 = W*in
   wire signed [9:0] m98_47;
   assign m98_47 =10'b0;

   // m98_48 = W*in
   wire signed [9:0] m98_48;
   assign m98_48 =10'b0;

   // m98_49 = W*in
   wire signed [9:0] m98_49;
   assign m98_49 =10'b0;

   // m98_50 = W*in
   wire signed [9:0] m98_50;
   assign m98_50 =10'b0;

   // m98_51 = W*in
   wire signed [9:0] m98_51;
   assign m98_51 =10'b0;

   // m98_52 = W*in
   wire signed [9:0] m98_52;
   assign m98_52 =10'b0;

   // m98_53 = W*in
   wire signed [9:0] m98_53;
   assign m98_53 =10'b0;

   // m98_54 = W*in
   wire signed [9:0] m98_54;
   assign m98_54 =10'b0;

   // m98_55 = W*in
   wire signed [9:0] m98_55;
   assign m98_55 =10'b0;

   // m98_56 = W*in
   wire signed [9:0] m98_56;
   assign m98_56 ={ {4{in98[5]}} , in98[5:0] };

   // m98_57 = W*in
   wire signed [9:0] m98_57;
   assign m98_57 =10'b0;

   // m98_58 = W*in
   wire signed [9:0] m98_58;
   assign m98_58 =10'b0;

   // m98_59 = W*in
   wire signed [9:0] m98_59;
   assign m98_59 ={ {4{in98[5]}} , in98[5:0] };

   // m98_60 = W*in
   wire signed [9:0] m98_60;
   assign m98_60 =10'b0;

   // m98_61 = W*in
   wire signed [9:0] m98_61;
   assign m98_61 =10'b0;

   // m98_62 = W*in
   wire signed [9:0] m98_62;
   assign m98_62 =10'b0;

   // m98_63 = W*in
   wire signed [9:0] m98_63;
   assign m98_63 =10'b0;

   // m98_64 = W*in
   wire signed [9:0] m98_64;
   assign m98_64 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_65 = W*in
   wire signed [9:0] m98_65;
   assign m98_65 =10'b0;

   // m98_66 = W*in
   wire signed [9:0] m98_66;
   assign m98_66 =10'b0;

   // m98_67 = W*in
   wire signed [9:0] m98_67;
   assign m98_67 =10'b0;

   // m98_68 = W*in
   wire signed [9:0] m98_68;
   assign m98_68 =10'b0;

   // m98_69 = W*in
   wire signed [9:0] m98_69;
   assign m98_69 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_70 = W*in
   wire signed [9:0] m98_70;
   assign m98_70 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_71 = W*in
   wire signed [9:0] m98_71;
   assign m98_71 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_72 = W*in
   wire signed [9:0] m98_72;
   assign m98_72 =10'b0;

   // m98_73 = W*in
   wire signed [9:0] m98_73;
   assign m98_73 ={ {5{in98[5]}} , in98[5:1] };

   // m98_74 = W*in
   wire signed [9:0] m98_74;
   assign m98_74 =10'b0;

   // m98_75 = W*in
   wire signed [9:0] m98_75;
   assign m98_75 ={ {5{in98[5]}} , in98[5:1] };

   // m98_76 = W*in
   wire signed [9:0] m98_76;
   assign m98_76 =10'b0;

   // m98_77 = W*in
   wire signed [9:0] m98_77;
   assign m98_77 =10'b0;

   // m98_78 = W*in
   wire signed [9:0] m98_78;
   assign m98_78 ={ {4{in98[5]}} , in98[5:0] };

   // m98_79 = W*in
   wire signed [9:0] m98_79;
   assign m98_79 =10'b0;

   // m98_80 = W*in
   wire signed [9:0] m98_80;
   assign m98_80 =10'b0;

   // m98_81 = W*in
   wire signed [9:0] m98_81;
   assign m98_81 ={ {5{in98[5]}} , in98[5:1] };

   // m98_82 = W*in
   wire signed [9:0] m98_82;
   assign m98_82 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_83 = W*in
   wire signed [9:0] m98_83;
   assign m98_83 =10'b0;

   // m98_84 = W*in
   wire signed [9:0] m98_84;
   assign m98_84 =10'b0;

   // m98_85 = W*in
   wire signed [9:0] m98_85;
   assign m98_85 =10'b0;

   // m98_86 = W*in
   wire signed [9:0] m98_86;
   assign m98_86 =10'b0;

   // m98_87 = W*in
   wire signed [9:0] m98_87;
   assign m98_87 =10'b0;

   // m98_88 = W*in
   wire signed [9:0] m98_88;
   assign m98_88 ={ {4{neg98[5]}} , neg98[5:0] };

   // m98_89 = W*in
   wire signed [9:0] m98_89;
   assign m98_89 =10'b0;

   // m98_90 = W*in
   wire signed [9:0] m98_90;
   assign m98_90 =10'b0;

   // m98_91 = W*in
   wire signed [9:0] m98_91;
   assign m98_91 =10'b0;

   // m98_92 = W*in
   wire signed [9:0] m98_92;
   assign m98_92 =10'b0;

   // m98_93 = W*in
   wire signed [9:0] m98_93;
   assign m98_93 =10'b0;

   // m98_94 = W*in
   wire signed [9:0] m98_94;
   assign m98_94 =10'b0;

   // m98_95 = W*in
   wire signed [9:0] m98_95;
   assign m98_95 =10'b0;

   // m98_96 = W*in
   wire signed [9:0] m98_96;
   assign m98_96 =10'b0;

   // m98_97 = W*in
   wire signed [9:0] m98_97;
   assign m98_97 =10'b0;

   // m98_98 = W*in
   wire signed [9:0] m98_98;
   assign m98_98 =10'b0;

   // m98_99 = W*in
   wire signed [9:0] m98_99;
   assign m98_99 =10'b0;

   // m98_100 = W*in
   wire signed [9:0] m98_100;
   assign m98_100 =10'b0;

   // m98_101 = W*in
   wire signed [9:0] m98_101;
   assign m98_101 =10'b0;

   // m98_102 = W*in
   wire signed [9:0] m98_102;
   assign m98_102 ={ {4{in98[5]}} , in98[5:0] };

   // m98_103 = W*in
   wire signed [9:0] m98_103;
   assign m98_103 =10'b0;

   // m98_104 = W*in
   wire signed [9:0] m98_104;
   assign m98_104 =10'b0;

   // m98_105 = W*in
   wire signed [9:0] m98_105;
   assign m98_105 =10'b0;

   // m98_106 = W*in
   wire signed [9:0] m98_106;
   assign m98_106 =10'b0;

   // m98_107 = W*in
   wire signed [9:0] m98_107;
   assign m98_107 =10'b0;

   // m98_108 = W*in
   wire signed [9:0] m98_108;
   assign m98_108 ={ {5{neg98[5]}} , neg98[5:1] };

   // m98_109 = W*in
   wire signed [9:0] m98_109;
   assign m98_109 =10'b0;

   // m98_110 = W*in
   wire signed [9:0] m98_110;
   assign m98_110 =10'b0;

   // m98_111 = W*in
   wire signed [9:0] m98_111;
   assign m98_111 =10'b0;

   // m98_112 = W*in
   wire signed [9:0] m98_112;
   assign m98_112 =10'b0;

   // m98_113 = W*in
   wire signed [9:0] m98_113;
   assign m98_113 =10'b0;

   // m98_114 = W*in
   wire signed [9:0] m98_114;
   assign m98_114 =10'b0;

   // m98_115 = W*in
   wire signed [9:0] m98_115;
   assign m98_115 =10'b0;

   // m98_116 = W*in
   wire signed [9:0] m98_116;
   assign m98_116 =10'b0;

   // m98_117 = W*in
   wire signed [9:0] m98_117;
   assign m98_117 =10'b0;

   // m99_1 = W*in
   wire signed [9:0] m99_1;
   assign m99_1 ={ {4{in99[5]}} , in99[5:0] };

   // m99_2 = W*in
   wire signed [9:0] m99_2;
   assign m99_2 =10'b0;

   // m99_3 = W*in
   wire signed [9:0] m99_3;
   assign m99_3 =10'b0;

   // m99_4 = W*in
   wire signed [9:0] m99_4;
   assign m99_4 =10'b0;

   // m99_5 = W*in
   wire signed [9:0] m99_5;
   assign m99_5 =10'b0;

   // m99_6 = W*in
   wire signed [9:0] m99_6;
   assign m99_6 =10'b0;

   // m99_7 = W*in
   wire signed [9:0] m99_7;
   assign m99_7 ={ {4{in99[5]}} , in99[5:0] };

   // m99_8 = W*in
   wire signed [9:0] m99_8;
   assign m99_8 =10'b0;

   // m99_9 = W*in
   wire signed [9:0] m99_9;
   assign m99_9 =10'b0;

   // m99_10 = W*in
   wire signed [9:0] m99_10;
   assign m99_10 =10'b0;

   // m99_11 = W*in
   wire signed [9:0] m99_11;
   assign m99_11 =10'b0;

   // m99_12 = W*in
   wire signed [9:0] m99_12;
   assign m99_12 =10'b0;

   // m99_13 = W*in
   wire signed [9:0] m99_13;
   assign m99_13 =10'b0;

   // m99_14 = W*in
   wire signed [9:0] m99_14;
   assign m99_14 =10'b0;

   // m99_15 = W*in
   wire signed [9:0] m99_15;
   assign m99_15 =10'b0;

   // m99_16 = W*in
   wire signed [9:0] m99_16;
   assign m99_16 =10'b0;

   // m99_17 = W*in
   wire signed [9:0] m99_17;
   assign m99_17 =10'b0;

   // m99_18 = W*in
   wire signed [9:0] m99_18;
   assign m99_18 =10'b0;

   // m99_19 = W*in
   wire signed [9:0] m99_19;
   assign m99_19 =10'b0;

   // m99_20 = W*in
   wire signed [9:0] m99_20;
   assign m99_20 =10'b0;

   // m99_21 = W*in
   wire signed [9:0] m99_21;
   assign m99_21 =10'b0;

   // m99_22 = W*in
   wire signed [9:0] m99_22;
   assign m99_22 ={ {5{in99[5]}} , in99[5:1] };

   // m99_23 = W*in
   wire signed [9:0] m99_23;
   assign m99_23 =10'b0;

   // m99_24 = W*in
   wire signed [9:0] m99_24;
   assign m99_24 =10'b0;

   // m99_25 = W*in
   wire signed [9:0] m99_25;
   assign m99_25 =10'b0;

   // m99_26 = W*in
   wire signed [9:0] m99_26;
   assign m99_26 =10'b0;

   // m99_27 = W*in
   wire signed [9:0] m99_27;
   assign m99_27 =10'b0;

   // m99_28 = W*in
   wire signed [9:0] m99_28;
   assign m99_28 ={ {5{in99[5]}} , in99[5:1] };

   // m99_29 = W*in
   wire signed [9:0] m99_29;
   assign m99_29 =10'b0;

   // m99_30 = W*in
   wire signed [9:0] m99_30;
   assign m99_30 =10'b0;

   // m99_31 = W*in
   wire signed [9:0] m99_31;
   assign m99_31 ={ {5{neg99[5]}} , neg99[5:1] };

   // m99_32 = W*in
   wire signed [9:0] m99_32;
   assign m99_32 =10'b0;

   // m99_33 = W*in
   wire signed [9:0] m99_33;
   assign m99_33 ={ {4{in99[5]}} , in99[5:0] };

   // m99_34 = W*in
   wire signed [9:0] m99_34;
   assign m99_34 =10'b0;

   // m99_35 = W*in
   wire signed [9:0] m99_35;
   assign m99_35 =10'b0;

   // m99_36 = W*in
   wire signed [9:0] m99_36;
   assign m99_36 =10'b0;

   // m99_37 = W*in
   wire signed [9:0] m99_37;
   assign m99_37 =10'b0;

   // m99_38 = W*in
   wire signed [9:0] m99_38;
   assign m99_38 =10'b0;

   // m99_39 = W*in
   wire signed [9:0] m99_39;
   assign m99_39 =10'b0;

   // m99_40 = W*in
   wire signed [9:0] m99_40;
   assign m99_40 =10'b0;

   // m99_41 = W*in
   wire signed [9:0] m99_41;
   assign m99_41 =10'b0;

   // m99_42 = W*in
   wire signed [9:0] m99_42;
   assign m99_42 =10'b0;

   // m99_43 = W*in
   wire signed [9:0] m99_43;
   assign m99_43 =10'b0;

   // m99_44 = W*in
   wire signed [9:0] m99_44;
   assign m99_44 =10'b0;

   // m99_45 = W*in
   wire signed [9:0] m99_45;
   assign m99_45 ={ {4{in99[5]}} , in99[5:0] };

   // m99_46 = W*in
   wire signed [9:0] m99_46;
   assign m99_46 =10'b0;

   // m99_47 = W*in
   wire signed [9:0] m99_47;
   assign m99_47 =10'b0;

   // m99_48 = W*in
   wire signed [9:0] m99_48;
   assign m99_48 =10'b0;

   // m99_49 = W*in
   wire signed [9:0] m99_49;
   assign m99_49 =10'b0;

   // m99_50 = W*in
   wire signed [9:0] m99_50;
   assign m99_50 =10'b0;

   // m99_51 = W*in
   wire signed [9:0] m99_51;
   assign m99_51 ={ {4{in99[5]}} , in99[5:0] };

   // m99_52 = W*in
   wire signed [9:0] m99_52;
   assign m99_52 =10'b0;

   // m99_53 = W*in
   wire signed [9:0] m99_53;
   assign m99_53 =10'b0;

   // m99_54 = W*in
   wire signed [9:0] m99_54;
   assign m99_54 =10'b0;

   // m99_55 = W*in
   wire signed [9:0] m99_55;
   assign m99_55 =10'b0;

   // m99_56 = W*in
   wire signed [9:0] m99_56;
   assign m99_56 ={ {4{in99[5]}} , in99[5:0] };

   // m99_57 = W*in
   wire signed [9:0] m99_57;
   assign m99_57 =10'b0;

   // m99_58 = W*in
   wire signed [9:0] m99_58;
   assign m99_58 =10'b0;

   // m99_59 = W*in
   wire signed [9:0] m99_59;
   assign m99_59 =10'b0;

   // m99_60 = W*in
   wire signed [9:0] m99_60;
   assign m99_60 =10'b0;

   // m99_61 = W*in
   wire signed [9:0] m99_61;
   assign m99_61 =10'b0;

   // m99_62 = W*in
   wire signed [9:0] m99_62;
   assign m99_62 =10'b0;

   // m99_63 = W*in
   wire signed [9:0] m99_63;
   assign m99_63 =10'b0;

   // m99_64 = W*in
   wire signed [9:0] m99_64;
   assign m99_64 =10'b0;

   // m99_65 = W*in
   wire signed [9:0] m99_65;
   assign m99_65 ={ {5{neg99[5]}} , neg99[5:1] };

   // m99_66 = W*in
   wire signed [9:0] m99_66;
   assign m99_66 ={ {4{neg99[5]}} , neg99[5:0] };

   // m99_67 = W*in
   wire signed [9:0] m99_67;
   assign m99_67 =10'b0;

   // m99_68 = W*in
   wire signed [9:0] m99_68;
   assign m99_68 =10'b0;

   // m99_69 = W*in
   wire signed [9:0] m99_69;
   assign m99_69 =10'b0;

   // m99_70 = W*in
   wire signed [9:0] m99_70;
   assign m99_70 ={ {5{neg99[5]}} , neg99[5:1] };

   // m99_71 = W*in
   wire signed [9:0] m99_71;
   assign m99_71 =10'b0;

   // m99_72 = W*in
   wire signed [9:0] m99_72;
   assign m99_72 =10'b0;

   // m99_73 = W*in
   wire signed [9:0] m99_73;
   assign m99_73 =10'b0;

   // m99_74 = W*in
   wire signed [9:0] m99_74;
   assign m99_74 ={ {4{neg99[5]}} , neg99[5:0] };

   // m99_75 = W*in
   wire signed [9:0] m99_75;
   assign m99_75 =10'b0;

   // m99_76 = W*in
   wire signed [9:0] m99_76;
   assign m99_76 =10'b0;

   // m99_77 = W*in
   wire signed [9:0] m99_77;
   assign m99_77 =10'b0;

   // m99_78 = W*in
   wire signed [9:0] m99_78;
   assign m99_78 ={ {5{in99[5]}} , in99[5:1] };

   // m99_79 = W*in
   wire signed [9:0] m99_79;
   assign m99_79 =10'b0;

   // m99_80 = W*in
   wire signed [9:0] m99_80;
   assign m99_80 =10'b0;

   // m99_81 = W*in
   wire signed [9:0] m99_81;
   assign m99_81 =10'b0;

   // m99_82 = W*in
   wire signed [9:0] m99_82;
   assign m99_82 =10'b0;

   // m99_83 = W*in
   wire signed [9:0] m99_83;
   assign m99_83 ={ {5{in99[5]}} , in99[5:1] };

   // m99_84 = W*in
   wire signed [9:0] m99_84;
   assign m99_84 =10'b0;

   // m99_85 = W*in
   wire signed [9:0] m99_85;
   assign m99_85 =10'b0;

   // m99_86 = W*in
   wire signed [9:0] m99_86;
   assign m99_86 =10'b0;

   // m99_87 = W*in
   wire signed [9:0] m99_87;
   assign m99_87 =10'b0;

   // m99_88 = W*in
   wire signed [9:0] m99_88;
   assign m99_88 =10'b0;

   // m99_89 = W*in
   wire signed [9:0] m99_89;
   assign m99_89 =10'b0;

   // m99_90 = W*in
   wire signed [9:0] m99_90;
   assign m99_90 =10'b0;

   // m99_91 = W*in
   wire signed [9:0] m99_91;
   assign m99_91 =10'b0;

   // m99_92 = W*in
   wire signed [9:0] m99_92;
   assign m99_92 =10'b0;

   // m99_93 = W*in
   wire signed [9:0] m99_93;
   assign m99_93 =10'b0;

   // m99_94 = W*in
   wire signed [9:0] m99_94;
   assign m99_94 =10'b0;

   // m99_95 = W*in
   wire signed [9:0] m99_95;
   assign m99_95 =10'b0;

   // m99_96 = W*in
   wire signed [9:0] m99_96;
   assign m99_96 =10'b0;

   // m99_97 = W*in
   wire signed [9:0] m99_97;
   assign m99_97 =10'b0;

   // m99_98 = W*in
   wire signed [9:0] m99_98;
   assign m99_98 =10'b0;

   // m99_99 = W*in
   wire signed [9:0] m99_99;
   assign m99_99 =10'b0;

   // m99_100 = W*in
   wire signed [9:0] m99_100;
   assign m99_100 =10'b0;

   // m99_101 = W*in
   wire signed [9:0] m99_101;
   assign m99_101 =10'b0;

   // m99_102 = W*in
   wire signed [9:0] m99_102;
   assign m99_102 =10'b0;

   // m99_103 = W*in
   wire signed [9:0] m99_103;
   assign m99_103 =10'b0;

   // m99_104 = W*in
   wire signed [9:0] m99_104;
   assign m99_104 =10'b0;

   // m99_105 = W*in
   wire signed [9:0] m99_105;
   assign m99_105 =10'b0;

   // m99_106 = W*in
   wire signed [9:0] m99_106;
   assign m99_106 =10'b0;

   // m99_107 = W*in
   wire signed [9:0] m99_107;
   assign m99_107 =10'b0;

   // m99_108 = W*in
   wire signed [9:0] m99_108;
   assign m99_108 ={ {5{neg99[5]}} , neg99[5:1] };

   // m99_109 = W*in
   wire signed [9:0] m99_109;
   assign m99_109 =10'b0;

   // m99_110 = W*in
   wire signed [9:0] m99_110;
   assign m99_110 =10'b0;

   // m99_111 = W*in
   wire signed [9:0] m99_111;
   assign m99_111 =10'b0;

   // m99_112 = W*in
   wire signed [9:0] m99_112;
   assign m99_112 =10'b0;

   // m99_113 = W*in
   wire signed [9:0] m99_113;
   assign m99_113 ={ {4{in99[5]}} , in99[5:0] };

   // m99_114 = W*in
   wire signed [9:0] m99_114;
   assign m99_114 =10'b0;

   // m99_115 = W*in
   wire signed [9:0] m99_115;
   assign m99_115 =10'b0;

   // m99_116 = W*in
   wire signed [9:0] m99_116;
   assign m99_116 ={ {4{neg99[5]}} , neg99[5:0] };

   // m99_117 = W*in
   wire signed [9:0] m99_117;
   assign m99_117 =10'b0;

   // m100_1 = W*in
   wire signed [9:0] m100_1;
   assign m100_1 ={ {4{in100[5]}} , in100[5:0] };

   // m100_2 = W*in
   wire signed [9:0] m100_2;
   assign m100_2 =10'b0;

   // m100_3 = W*in
   wire signed [9:0] m100_3;
   assign m100_3 =10'b0;

   // m100_4 = W*in
   wire signed [9:0] m100_4;
   assign m100_4 =10'b0;

   // m100_5 = W*in
   wire signed [9:0] m100_5;
   assign m100_5 =10'b0;

   // m100_6 = W*in
   wire signed [9:0] m100_6;
   assign m100_6 =10'b0;

   // m100_7 = W*in
   wire signed [9:0] m100_7;
   assign m100_7 =10'b0;

   // m100_8 = W*in
   wire signed [9:0] m100_8;
   assign m100_8 =10'b0;

   // m100_9 = W*in
   wire signed [9:0] m100_9;
   assign m100_9 =10'b0;

   // m100_10 = W*in
   wire signed [9:0] m100_10;
   assign m100_10 =10'b0;

   // m100_11 = W*in
   wire signed [9:0] m100_11;
   assign m100_11 =10'b0;

   // m100_12 = W*in
   wire signed [9:0] m100_12;
   assign m100_12 =10'b0;

   // m100_13 = W*in
   wire signed [9:0] m100_13;
   assign m100_13 =10'b0;

   // m100_14 = W*in
   wire signed [9:0] m100_14;
   assign m100_14 =10'b0;

   // m100_15 = W*in
   wire signed [9:0] m100_15;
   assign m100_15 =10'b0;

   // m100_16 = W*in
   wire signed [9:0] m100_16;
   assign m100_16 =10'b0;

   // m100_17 = W*in
   wire signed [9:0] m100_17;
   assign m100_17 =10'b0;

   // m100_18 = W*in
   wire signed [9:0] m100_18;
   assign m100_18 =10'b0;

   // m100_19 = W*in
   wire signed [9:0] m100_19;
   assign m100_19 =10'b0;

   // m100_20 = W*in
   wire signed [9:0] m100_20;
   assign m100_20 ={ {5{in100[5]}} , in100[5:1] };

   // m100_21 = W*in
   wire signed [9:0] m100_21;
   assign m100_21 =10'b0;

   // m100_22 = W*in
   wire signed [9:0] m100_22;
   assign m100_22 ={ {5{in100[5]}} , in100[5:1] };

   // m100_23 = W*in
   wire signed [9:0] m100_23;
   assign m100_23 =10'b0;

   // m100_24 = W*in
   wire signed [9:0] m100_24;
   assign m100_24 =10'b0;

   // m100_25 = W*in
   wire signed [9:0] m100_25;
   assign m100_25 =10'b0;

   // m100_26 = W*in
   wire signed [9:0] m100_26;
   assign m100_26 =10'b0;

   // m100_27 = W*in
   wire signed [9:0] m100_27;
   assign m100_27 =10'b0;

   // m100_28 = W*in
   wire signed [9:0] m100_28;
   assign m100_28 =10'b0;

   // m100_29 = W*in
   wire signed [9:0] m100_29;
   assign m100_29 =10'b0;

   // m100_30 = W*in
   wire signed [9:0] m100_30;
   assign m100_30 ={ {5{in100[5]}} , in100[5:1] };

   // m100_31 = W*in
   wire signed [9:0] m100_31;
   assign m100_31 =10'b0;

   // m100_32 = W*in
   wire signed [9:0] m100_32;
   assign m100_32 =10'b0;

   // m100_33 = W*in
   wire signed [9:0] m100_33;
   assign m100_33 =10'b0;

   // m100_34 = W*in
   wire signed [9:0] m100_34;
   assign m100_34 =10'b0;

   // m100_35 = W*in
   wire signed [9:0] m100_35;
   assign m100_35 ={ {5{in100[5]}} , in100[5:1] };

   // m100_36 = W*in
   wire signed [9:0] m100_36;
   assign m100_36 =10'b0;

   // m100_37 = W*in
   wire signed [9:0] m100_37;
   assign m100_37 =10'b0;

   // m100_38 = W*in
   wire signed [9:0] m100_38;
   assign m100_38 =10'b0;

   // m100_39 = W*in
   wire signed [9:0] m100_39;
   assign m100_39 =10'b0;

   // m100_40 = W*in
   wire signed [9:0] m100_40;
   assign m100_40 =10'b0;

   // m100_41 = W*in
   wire signed [9:0] m100_41;
   assign m100_41 =10'b0;

   // m100_42 = W*in
   wire signed [9:0] m100_42;
   assign m100_42 =10'b0;

   // m100_43 = W*in
   wire signed [9:0] m100_43;
   assign m100_43 =10'b0;

   // m100_44 = W*in
   wire signed [9:0] m100_44;
   assign m100_44 =10'b0;

   // m100_45 = W*in
   wire signed [9:0] m100_45;
   assign m100_45 =10'b0;

   // m100_46 = W*in
   wire signed [9:0] m100_46;
   assign m100_46 =10'b0;

   // m100_47 = W*in
   wire signed [9:0] m100_47;
   assign m100_47 =10'b0;

   // m100_48 = W*in
   wire signed [9:0] m100_48;
   assign m100_48 =10'b0;

   // m100_49 = W*in
   wire signed [9:0] m100_49;
   assign m100_49 =10'b0;

   // m100_50 = W*in
   wire signed [9:0] m100_50;
   assign m100_50 =10'b0;

   // m100_51 = W*in
   wire signed [9:0] m100_51;
   assign m100_51 =10'b0;

   // m100_52 = W*in
   wire signed [9:0] m100_52;
   assign m100_52 =10'b0;

   // m100_53 = W*in
   wire signed [9:0] m100_53;
   assign m100_53 =10'b0;

   // m100_54 = W*in
   wire signed [9:0] m100_54;
   assign m100_54 =10'b0;

   // m100_55 = W*in
   wire signed [9:0] m100_55;
   assign m100_55 =10'b0;

   // m100_56 = W*in
   wire signed [9:0] m100_56;
   assign m100_56 =10'b0;

   // m100_57 = W*in
   wire signed [9:0] m100_57;
   assign m100_57 =10'b0;

   // m100_58 = W*in
   wire signed [9:0] m100_58;
   assign m100_58 =10'b0;

   // m100_59 = W*in
   wire signed [9:0] m100_59;
   assign m100_59 =10'b0;

   // m100_60 = W*in
   wire signed [9:0] m100_60;
   assign m100_60 =10'b0;

   // m100_61 = W*in
   wire signed [9:0] m100_61;
   assign m100_61 =10'b0;

   // m100_62 = W*in
   wire signed [9:0] m100_62;
   assign m100_62 =10'b0;

   // m100_63 = W*in
   wire signed [9:0] m100_63;
   assign m100_63 =10'b0;

   // m100_64 = W*in
   wire signed [9:0] m100_64;
   assign m100_64 ={ {5{in100[5]}} , in100[5:1] };

   // m100_65 = W*in
   wire signed [9:0] m100_65;
   assign m100_65 =10'b0;

   // m100_66 = W*in
   wire signed [9:0] m100_66;
   assign m100_66 =10'b0;

   // m100_67 = W*in
   wire signed [9:0] m100_67;
   assign m100_67 =10'b0;

   // m100_68 = W*in
   wire signed [9:0] m100_68;
   assign m100_68 =10'b0;

   // m100_69 = W*in
   wire signed [9:0] m100_69;
   assign m100_69 =10'b0;

   // m100_70 = W*in
   wire signed [9:0] m100_70;
   assign m100_70 =10'b0;

   // m100_71 = W*in
   wire signed [9:0] m100_71;
   assign m100_71 =10'b0;

   // m100_72 = W*in
   wire signed [9:0] m100_72;
   assign m100_72 =10'b0;

   // m100_73 = W*in
   wire signed [9:0] m100_73;
   assign m100_73 =10'b0;

   // m100_74 = W*in
   wire signed [9:0] m100_74;
   assign m100_74 =10'b0;

   // m100_75 = W*in
   wire signed [9:0] m100_75;
   assign m100_75 =10'b0;

   // m100_76 = W*in
   wire signed [9:0] m100_76;
   assign m100_76 =10'b0;

   // m100_77 = W*in
   wire signed [9:0] m100_77;
   assign m100_77 =10'b0;

   // m100_78 = W*in
   wire signed [9:0] m100_78;
   assign m100_78 =10'b0;

   // m100_79 = W*in
   wire signed [9:0] m100_79;
   assign m100_79 =10'b0;

   // m100_80 = W*in
   wire signed [9:0] m100_80;
   assign m100_80 =10'b0;

   // m100_81 = W*in
   wire signed [9:0] m100_81;
   assign m100_81 ={ {5{in100[5]}} , in100[5:1] };

   // m100_82 = W*in
   wire signed [9:0] m100_82;
   assign m100_82 =10'b0;

   // m100_83 = W*in
   wire signed [9:0] m100_83;
   assign m100_83 ={ {5{in100[5]}} , in100[5:1] };

   // m100_84 = W*in
   wire signed [9:0] m100_84;
   assign m100_84 =10'b0;

   // m100_85 = W*in
   wire signed [9:0] m100_85;
   assign m100_85 =10'b0;

   // m100_86 = W*in
   wire signed [9:0] m100_86;
   assign m100_86 =10'b0;

   // m100_87 = W*in
   wire signed [9:0] m100_87;
   assign m100_87 =10'b0;

   // m100_88 = W*in
   wire signed [9:0] m100_88;
   assign m100_88 =10'b0;

   // m100_89 = W*in
   wire signed [9:0] m100_89;
   assign m100_89 =10'b0;

   // m100_90 = W*in
   wire signed [9:0] m100_90;
   assign m100_90 =10'b0;

   // m100_91 = W*in
   wire signed [9:0] m100_91;
   assign m100_91 =10'b0;

   // m100_92 = W*in
   wire signed [9:0] m100_92;
   assign m100_92 =10'b0;

   // m100_93 = W*in
   wire signed [9:0] m100_93;
   assign m100_93 =10'b0;

   // m100_94 = W*in
   wire signed [9:0] m100_94;
   assign m100_94 =10'b0;

   // m100_95 = W*in
   wire signed [9:0] m100_95;
   assign m100_95 =10'b0;

   // m100_96 = W*in
   wire signed [9:0] m100_96;
   assign m100_96 =10'b0;

   // m100_97 = W*in
   wire signed [9:0] m100_97;
   assign m100_97 =10'b0;

   // m100_98 = W*in
   wire signed [9:0] m100_98;
   assign m100_98 =10'b0;

   // m100_99 = W*in
   wire signed [9:0] m100_99;
   assign m100_99 =10'b0;

   // m100_100 = W*in
   wire signed [9:0] m100_100;
   assign m100_100 =10'b0;

   // m100_101 = W*in
   wire signed [9:0] m100_101;
   assign m100_101 =10'b0;

   // m100_102 = W*in
   wire signed [9:0] m100_102;
   assign m100_102 =10'b0;

   // m100_103 = W*in
   wire signed [9:0] m100_103;
   assign m100_103 =10'b0;

   // m100_104 = W*in
   wire signed [9:0] m100_104;
   assign m100_104 =10'b0;

   // m100_105 = W*in
   wire signed [9:0] m100_105;
   assign m100_105 =10'b0;

   // m100_106 = W*in
   wire signed [9:0] m100_106;
   assign m100_106 =10'b0;

   // m100_107 = W*in
   wire signed [9:0] m100_107;
   assign m100_107 =10'b0;

   // m100_108 = W*in
   wire signed [9:0] m100_108;
   assign m100_108 ={ {5{in100[5]}} , in100[5:1] };

   // m100_109 = W*in
   wire signed [9:0] m100_109;
   assign m100_109 ={ {4{in100[5]}} , in100[5:0] };

   // m100_110 = W*in
   wire signed [9:0] m100_110;
   assign m100_110 =10'b0;

   // m100_111 = W*in
   wire signed [9:0] m100_111;
   assign m100_111 =10'b0;

   // m100_112 = W*in
   wire signed [9:0] m100_112;
   assign m100_112 =10'b0;

   // m100_113 = W*in
   wire signed [9:0] m100_113;
   assign m100_113 =10'b0;

   // m100_114 = W*in
   wire signed [9:0] m100_114;
   assign m100_114 =10'b0;

   // m100_115 = W*in
   wire signed [9:0] m100_115;
   assign m100_115 =10'b0;

   // m100_116 = W*in
   wire signed [9:0] m100_116;
   assign m100_116 =10'b0;

   // m100_117 = W*in
   wire signed [9:0] m100_117;
   assign m100_117 =10'b0;

   // m101_1 = W*in
   wire signed [9:0] m101_1;
   assign m101_1 =10'b0;

   // m101_2 = W*in
   wire signed [9:0] m101_2;
   assign m101_2 =10'b0;

   // m101_3 = W*in
   wire signed [9:0] m101_3;
   assign m101_3 =10'b0;

   // m101_4 = W*in
   wire signed [9:0] m101_4;
   assign m101_4 =10'b0;

   // m101_5 = W*in
   wire signed [9:0] m101_5;
   assign m101_5 =10'b0;

   // m101_6 = W*in
   wire signed [9:0] m101_6;
   assign m101_6 =10'b0;

   // m101_7 = W*in
   wire signed [9:0] m101_7;
   assign m101_7 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_8 = W*in
   wire signed [9:0] m101_8;
   assign m101_8 =10'b0;

   // m101_9 = W*in
   wire signed [9:0] m101_9;
   assign m101_9 =10'b0;

   // m101_10 = W*in
   wire signed [9:0] m101_10;
   assign m101_10 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_11 = W*in
   wire signed [9:0] m101_11;
   assign m101_11 =10'b0;

   // m101_12 = W*in
   wire signed [9:0] m101_12;
   assign m101_12 =10'b0;

   // m101_13 = W*in
   wire signed [9:0] m101_13;
   assign m101_13 =10'b0;

   // m101_14 = W*in
   wire signed [9:0] m101_14;
   assign m101_14 =10'b0;

   // m101_15 = W*in
   wire signed [9:0] m101_15;
   assign m101_15 =10'b0;

   // m101_16 = W*in
   wire signed [9:0] m101_16;
   assign m101_16 ={ {4{in101[5]}} , in101[5:0] };

   // m101_17 = W*in
   wire signed [9:0] m101_17;
   assign m101_17 ={ {5{neg101[5]}} , neg101[5:1] };

   // m101_18 = W*in
   wire signed [9:0] m101_18;
   assign m101_18 ={ {5{in101[5]}} , in101[5:1] };

   // m101_19 = W*in
   wire signed [9:0] m101_19;
   assign m101_19 =10'b0;

   // m101_20 = W*in
   wire signed [9:0] m101_20;
   assign m101_20 =10'b0;

   // m101_21 = W*in
   wire signed [9:0] m101_21;
   assign m101_21 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_22 = W*in
   wire signed [9:0] m101_22;
   assign m101_22 =10'b0;

   // m101_23 = W*in
   wire signed [9:0] m101_23;
   assign m101_23 =10'b0;

   // m101_24 = W*in
   wire signed [9:0] m101_24;
   assign m101_24 =10'b0;

   // m101_25 = W*in
   wire signed [9:0] m101_25;
   assign m101_25 =10'b0;

   // m101_26 = W*in
   wire signed [9:0] m101_26;
   assign m101_26 =10'b0;

   // m101_27 = W*in
   wire signed [9:0] m101_27;
   assign m101_27 =10'b0;

   // m101_28 = W*in
   wire signed [9:0] m101_28;
   assign m101_28 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_29 = W*in
   wire signed [9:0] m101_29;
   assign m101_29 =10'b0;

   // m101_30 = W*in
   wire signed [9:0] m101_30;
   assign m101_30 ={ {4{in101[5]}} , in101[5:0] };

   // m101_31 = W*in
   wire signed [9:0] m101_31;
   assign m101_31 =10'b0;

   // m101_32 = W*in
   wire signed [9:0] m101_32;
   assign m101_32 =10'b0;

   // m101_33 = W*in
   wire signed [9:0] m101_33;
   assign m101_33 =10'b0;

   // m101_34 = W*in
   wire signed [9:0] m101_34;
   assign m101_34 =10'b0;

   // m101_35 = W*in
   wire signed [9:0] m101_35;
   assign m101_35 ={ {4{in101[5]}} , in101[5:0] };

   // m101_36 = W*in
   wire signed [9:0] m101_36;
   assign m101_36 =10'b0;

   // m101_37 = W*in
   wire signed [9:0] m101_37;
   assign m101_37 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_38 = W*in
   wire signed [9:0] m101_38;
   assign m101_38 =10'b0;

   // m101_39 = W*in
   wire signed [9:0] m101_39;
   assign m101_39 =10'b0;

   // m101_40 = W*in
   wire signed [9:0] m101_40;
   assign m101_40 =10'b0;

   // m101_41 = W*in
   wire signed [9:0] m101_41;
   assign m101_41 =10'b0;

   // m101_42 = W*in
   wire signed [9:0] m101_42;
   assign m101_42 ={ {4{in101[5]}} , in101[5:0] };

   // m101_43 = W*in
   wire signed [9:0] m101_43;
   assign m101_43 =10'b0;

   // m101_44 = W*in
   wire signed [9:0] m101_44;
   assign m101_44 =10'b0;

   // m101_45 = W*in
   wire signed [9:0] m101_45;
   assign m101_45 =10'b0;

   // m101_46 = W*in
   wire signed [9:0] m101_46;
   assign m101_46 =10'b0;

   // m101_47 = W*in
   wire signed [9:0] m101_47;
   assign m101_47 =10'b0;

   // m101_48 = W*in
   wire signed [9:0] m101_48;
   assign m101_48 =10'b0;

   // m101_49 = W*in
   wire signed [9:0] m101_49;
   assign m101_49 =10'b0;

   // m101_50 = W*in
   wire signed [9:0] m101_50;
   assign m101_50 ={ {4{in101[5]}} , in101[5:0] };

   // m101_51 = W*in
   wire signed [9:0] m101_51;
   assign m101_51 =10'b0;

   // m101_52 = W*in
   wire signed [9:0] m101_52;
   assign m101_52 =10'b0;

   // m101_53 = W*in
   wire signed [9:0] m101_53;
   assign m101_53 =10'b0;

   // m101_54 = W*in
   wire signed [9:0] m101_54;
   assign m101_54 =10'b0;

   // m101_55 = W*in
   wire signed [9:0] m101_55;
   assign m101_55 =10'b0;

   // m101_56 = W*in
   wire signed [9:0] m101_56;
   assign m101_56 ={ {4{in101[5]}} , in101[5:0] };

   // m101_57 = W*in
   wire signed [9:0] m101_57;
   assign m101_57 =10'b0;

   // m101_58 = W*in
   wire signed [9:0] m101_58;
   assign m101_58 =10'b0;

   // m101_59 = W*in
   wire signed [9:0] m101_59;
   assign m101_59 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_60 = W*in
   wire signed [9:0] m101_60;
   assign m101_60 =10'b0;

   // m101_61 = W*in
   wire signed [9:0] m101_61;
   assign m101_61 =10'b0;

   // m101_62 = W*in
   wire signed [9:0] m101_62;
   assign m101_62 =10'b0;

   // m101_63 = W*in
   wire signed [9:0] m101_63;
   assign m101_63 =10'b0;

   // m101_64 = W*in
   wire signed [9:0] m101_64;
   assign m101_64 ={ {4{in101[5]}} , in101[5:0] };

   // m101_65 = W*in
   wire signed [9:0] m101_65;
   assign m101_65 ={ {5{neg101[5]}} , neg101[5:1] };

   // m101_66 = W*in
   wire signed [9:0] m101_66;
   assign m101_66 =10'b0;

   // m101_67 = W*in
   wire signed [9:0] m101_67;
   assign m101_67 =10'b0;

   // m101_68 = W*in
   wire signed [9:0] m101_68;
   assign m101_68 =10'b0;

   // m101_69 = W*in
   wire signed [9:0] m101_69;
   assign m101_69 =10'b0;

   // m101_70 = W*in
   wire signed [9:0] m101_70;
   assign m101_70 ={ {5{neg101[5]}} , neg101[5:1] };

   // m101_71 = W*in
   wire signed [9:0] m101_71;
   assign m101_71 ={ {5{neg101[5]}} , neg101[5:1] };

   // m101_72 = W*in
   wire signed [9:0] m101_72;
   assign m101_72 ={ {5{neg101[5]}} , neg101[5:1] };

   // m101_73 = W*in
   wire signed [9:0] m101_73;
   assign m101_73 =10'b0;

   // m101_74 = W*in
   wire signed [9:0] m101_74;
   assign m101_74 =10'b0;

   // m101_75 = W*in
   wire signed [9:0] m101_75;
   assign m101_75 =10'b0;

   // m101_76 = W*in
   wire signed [9:0] m101_76;
   assign m101_76 =10'b0;

   // m101_77 = W*in
   wire signed [9:0] m101_77;
   assign m101_77 =10'b0;

   // m101_78 = W*in
   wire signed [9:0] m101_78;
   assign m101_78 =10'b0;

   // m101_79 = W*in
   wire signed [9:0] m101_79;
   assign m101_79 =10'b0;

   // m101_80 = W*in
   wire signed [9:0] m101_80;
   assign m101_80 =10'b0;

   // m101_81 = W*in
   wire signed [9:0] m101_81;
   assign m101_81 ={ {4{in101[5]}} , in101[5:0] };

   // m101_82 = W*in
   wire signed [9:0] m101_82;
   assign m101_82 =10'b0;

   // m101_83 = W*in
   wire signed [9:0] m101_83;
   assign m101_83 =10'b0;

   // m101_84 = W*in
   wire signed [9:0] m101_84;
   assign m101_84 =10'b0;

   // m101_85 = W*in
   wire signed [9:0] m101_85;
   assign m101_85 =10'b0;

   // m101_86 = W*in
   wire signed [9:0] m101_86;
   assign m101_86 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_87 = W*in
   wire signed [9:0] m101_87;
   assign m101_87 =10'b0;

   // m101_88 = W*in
   wire signed [9:0] m101_88;
   assign m101_88 =10'b0;

   // m101_89 = W*in
   wire signed [9:0] m101_89;
   assign m101_89 =10'b0;

   // m101_90 = W*in
   wire signed [9:0] m101_90;
   assign m101_90 =10'b0;

   // m101_91 = W*in
   wire signed [9:0] m101_91;
   assign m101_91 =10'b0;

   // m101_92 = W*in
   wire signed [9:0] m101_92;
   assign m101_92 =10'b0;

   // m101_93 = W*in
   wire signed [9:0] m101_93;
   assign m101_93 =10'b0;

   // m101_94 = W*in
   wire signed [9:0] m101_94;
   assign m101_94 ={ {4{in101[5]}} , in101[5:0] };

   // m101_95 = W*in
   wire signed [9:0] m101_95;
   assign m101_95 =10'b0;

   // m101_96 = W*in
   wire signed [9:0] m101_96;
   assign m101_96 =10'b0;

   // m101_97 = W*in
   wire signed [9:0] m101_97;
   assign m101_97 =10'b0;

   // m101_98 = W*in
   wire signed [9:0] m101_98;
   assign m101_98 =10'b0;

   // m101_99 = W*in
   wire signed [9:0] m101_99;
   assign m101_99 =10'b0;

   // m101_100 = W*in
   wire signed [9:0] m101_100;
   assign m101_100 =10'b0;

   // m101_101 = W*in
   wire signed [9:0] m101_101;
   assign m101_101 =10'b0;

   // m101_102 = W*in
   wire signed [9:0] m101_102;
   assign m101_102 ={ {4{in101[5]}} , in101[5:0] };

   // m101_103 = W*in
   wire signed [9:0] m101_103;
   assign m101_103 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_104 = W*in
   wire signed [9:0] m101_104;
   assign m101_104 ={ {4{neg101[5]}} , neg101[5:0] };

   // m101_105 = W*in
   wire signed [9:0] m101_105;
   assign m101_105 =10'b0;

   // m101_106 = W*in
   wire signed [9:0] m101_106;
   assign m101_106 ={ {4{in101[5]}} , in101[5:0] };

   // m101_107 = W*in
   wire signed [9:0] m101_107;
   assign m101_107 =10'b0;

   // m101_108 = W*in
   wire signed [9:0] m101_108;
   assign m101_108 =10'b0;

   // m101_109 = W*in
   wire signed [9:0] m101_109;
   assign m101_109 =10'b0;

   // m101_110 = W*in
   wire signed [9:0] m101_110;
   assign m101_110 =10'b0;

   // m101_111 = W*in
   wire signed [9:0] m101_111;
   assign m101_111 =10'b0;

   // m101_112 = W*in
   wire signed [9:0] m101_112;
   assign m101_112 =10'b0;

   // m101_113 = W*in
   wire signed [9:0] m101_113;
   assign m101_113 ={ {5{in101[5]}} , in101[5:1] };

   // m101_114 = W*in
   wire signed [9:0] m101_114;
   assign m101_114 =10'b0;

   // m101_115 = W*in
   wire signed [9:0] m101_115;
   assign m101_115 ={ {4{in101[5]}} , in101[5:0] };

   // m101_116 = W*in
   wire signed [9:0] m101_116;
   assign m101_116 =10'b0;

   // m101_117 = W*in
   wire signed [9:0] m101_117;
   assign m101_117 =10'b0;

   // m102_1 = W*in
   wire signed [9:0] m102_1;
   assign m102_1 ={ {4{in102[5]}} , in102[5:0] };

   // m102_2 = W*in
   wire signed [9:0] m102_2;
   assign m102_2 ={ {4{in102[5]}} , in102[5:0] };

   // m102_3 = W*in
   wire signed [9:0] m102_3;
   assign m102_3 =10'b0;

   // m102_4 = W*in
   wire signed [9:0] m102_4;
   assign m102_4 =10'b0;

   // m102_5 = W*in
   wire signed [9:0] m102_5;
   assign m102_5 ={ {4{in102[5]}} , in102[5:0] };

   // m102_6 = W*in
   wire signed [9:0] m102_6;
   assign m102_6 =10'b0;

   // m102_7 = W*in
   wire signed [9:0] m102_7;
   assign m102_7 =10'b0;

   // m102_8 = W*in
   wire signed [9:0] m102_8;
   assign m102_8 =10'b0;

   // m102_9 = W*in
   wire signed [9:0] m102_9;
   assign m102_9 =10'b0;

   // m102_10 = W*in
   wire signed [9:0] m102_10;
   assign m102_10 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_11 = W*in
   wire signed [9:0] m102_11;
   assign m102_11 =10'b0;

   // m102_12 = W*in
   wire signed [9:0] m102_12;
   assign m102_12 ={ {5{neg102[5]}} , neg102[5:1] };

   // m102_13 = W*in
   wire signed [9:0] m102_13;
   assign m102_13 =10'b0;

   // m102_14 = W*in
   wire signed [9:0] m102_14;
   assign m102_14 =10'b0;

   // m102_15 = W*in
   wire signed [9:0] m102_15;
   assign m102_15 =10'b0;

   // m102_16 = W*in
   wire signed [9:0] m102_16;
   assign m102_16 ={ {4{in102[5]}} , in102[5:0] };

   // m102_17 = W*in
   wire signed [9:0] m102_17;
   assign m102_17 =10'b0;

   // m102_18 = W*in
   wire signed [9:0] m102_18;
   assign m102_18 ={ {5{neg102[5]}} , neg102[5:1] };

   // m102_19 = W*in
   wire signed [9:0] m102_19;
   assign m102_19 =10'b0;

   // m102_20 = W*in
   wire signed [9:0] m102_20;
   assign m102_20 ={ {4{in102[5]}} , in102[5:0] };

   // m102_21 = W*in
   wire signed [9:0] m102_21;
   assign m102_21 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_22 = W*in
   wire signed [9:0] m102_22;
   assign m102_22 ={ {5{in102[5]}} , in102[5:1] };

   // m102_23 = W*in
   wire signed [9:0] m102_23;
   assign m102_23 =10'b0;

   // m102_24 = W*in
   wire signed [9:0] m102_24;
   assign m102_24 =10'b0;

   // m102_25 = W*in
   wire signed [9:0] m102_25;
   assign m102_25 =10'b0;

   // m102_26 = W*in
   wire signed [9:0] m102_26;
   assign m102_26 =10'b0;

   // m102_27 = W*in
   wire signed [9:0] m102_27;
   assign m102_27 ={ {5{in102[5]}} , in102[5:1] };

   // m102_28 = W*in
   wire signed [9:0] m102_28;
   assign m102_28 =10'b0;

   // m102_29 = W*in
   wire signed [9:0] m102_29;
   assign m102_29 ={ {5{neg102[5]}} , neg102[5:1] };

   // m102_30 = W*in
   wire signed [9:0] m102_30;
   assign m102_30 =10'b0;

   // m102_31 = W*in
   wire signed [9:0] m102_31;
   assign m102_31 =10'b0;

   // m102_32 = W*in
   wire signed [9:0] m102_32;
   assign m102_32 =10'b0;

   // m102_33 = W*in
   wire signed [9:0] m102_33;
   assign m102_33 ={ {5{in102[5]}} , in102[5:1] };

   // m102_34 = W*in
   wire signed [9:0] m102_34;
   assign m102_34 =10'b0;

   // m102_35 = W*in
   wire signed [9:0] m102_35;
   assign m102_35 ={ {5{in102[5]}} , in102[5:1] };

   // m102_36 = W*in
   wire signed [9:0] m102_36;
   assign m102_36 =10'b0;

   // m102_37 = W*in
   wire signed [9:0] m102_37;
   assign m102_37 =10'b0;

   // m102_38 = W*in
   wire signed [9:0] m102_38;
   assign m102_38 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_39 = W*in
   wire signed [9:0] m102_39;
   assign m102_39 =10'b0;

   // m102_40 = W*in
   wire signed [9:0] m102_40;
   assign m102_40 =10'b0;

   // m102_41 = W*in
   wire signed [9:0] m102_41;
   assign m102_41 ={ {4{in102[5]}} , in102[5:0] };

   // m102_42 = W*in
   wire signed [9:0] m102_42;
   assign m102_42 =10'b0;

   // m102_43 = W*in
   wire signed [9:0] m102_43;
   assign m102_43 =10'b0;

   // m102_44 = W*in
   wire signed [9:0] m102_44;
   assign m102_44 =10'b0;

   // m102_45 = W*in
   wire signed [9:0] m102_45;
   assign m102_45 =10'b0;

   // m102_46 = W*in
   wire signed [9:0] m102_46;
   assign m102_46 =10'b0;

   // m102_47 = W*in
   wire signed [9:0] m102_47;
   assign m102_47 =10'b0;

   // m102_48 = W*in
   wire signed [9:0] m102_48;
   assign m102_48 =10'b0;

   // m102_49 = W*in
   wire signed [9:0] m102_49;
   assign m102_49 =10'b0;

   // m102_50 = W*in
   wire signed [9:0] m102_50;
   assign m102_50 =10'b0;

   // m102_51 = W*in
   wire signed [9:0] m102_51;
   assign m102_51 ={ {4{in102[5]}} , in102[5:0] };

   // m102_52 = W*in
   wire signed [9:0] m102_52;
   assign m102_52 ={ {4{in102[5]}} , in102[5:0] };

   // m102_53 = W*in
   wire signed [9:0] m102_53;
   assign m102_53 =10'b0;

   // m102_54 = W*in
   wire signed [9:0] m102_54;
   assign m102_54 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_55 = W*in
   wire signed [9:0] m102_55;
   assign m102_55 =10'b0;

   // m102_56 = W*in
   wire signed [9:0] m102_56;
   assign m102_56 =10'b0;

   // m102_57 = W*in
   wire signed [9:0] m102_57;
   assign m102_57 =10'b0;

   // m102_58 = W*in
   wire signed [9:0] m102_58;
   assign m102_58 =10'b0;

   // m102_59 = W*in
   wire signed [9:0] m102_59;
   assign m102_59 =10'b0;

   // m102_60 = W*in
   wire signed [9:0] m102_60;
   assign m102_60 =10'b0;

   // m102_61 = W*in
   wire signed [9:0] m102_61;
   assign m102_61 =10'b0;

   // m102_62 = W*in
   wire signed [9:0] m102_62;
   assign m102_62 ={ {4{in102[5]}} , in102[5:0] };

   // m102_63 = W*in
   wire signed [9:0] m102_63;
   assign m102_63 =10'b0;

   // m102_64 = W*in
   wire signed [9:0] m102_64;
   assign m102_64 =10'b0;

   // m102_65 = W*in
   wire signed [9:0] m102_65;
   assign m102_65 =10'b0;

   // m102_66 = W*in
   wire signed [9:0] m102_66;
   assign m102_66 =10'b0;

   // m102_67 = W*in
   wire signed [9:0] m102_67;
   assign m102_67 =10'b0;

   // m102_68 = W*in
   wire signed [9:0] m102_68;
   assign m102_68 =10'b0;

   // m102_69 = W*in
   wire signed [9:0] m102_69;
   assign m102_69 ={ {5{neg102[5]}} , neg102[5:1] };

   // m102_70 = W*in
   wire signed [9:0] m102_70;
   assign m102_70 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_71 = W*in
   wire signed [9:0] m102_71;
   assign m102_71 =10'b0;

   // m102_72 = W*in
   wire signed [9:0] m102_72;
   assign m102_72 ={ {5{neg102[5]}} , neg102[5:1] };

   // m102_73 = W*in
   wire signed [9:0] m102_73;
   assign m102_73 =10'b0;

   // m102_74 = W*in
   wire signed [9:0] m102_74;
   assign m102_74 ={ {5{neg102[5]}} , neg102[5:1] };

   // m102_75 = W*in
   wire signed [9:0] m102_75;
   assign m102_75 ={ {4{in102[5]}} , in102[5:0] };

   // m102_76 = W*in
   wire signed [9:0] m102_76;
   assign m102_76 =10'b0;

   // m102_77 = W*in
   wire signed [9:0] m102_77;
   assign m102_77 =10'b0;

   // m102_78 = W*in
   wire signed [9:0] m102_78;
   assign m102_78 =10'b0;

   // m102_79 = W*in
   wire signed [9:0] m102_79;
   assign m102_79 =10'b0;

   // m102_80 = W*in
   wire signed [9:0] m102_80;
   assign m102_80 =10'b0;

   // m102_81 = W*in
   wire signed [9:0] m102_81;
   assign m102_81 ={ {4{in102[5]}} , in102[5:0] };

   // m102_82 = W*in
   wire signed [9:0] m102_82;
   assign m102_82 =10'b0;

   // m102_83 = W*in
   wire signed [9:0] m102_83;
   assign m102_83 =10'b0;

   // m102_84 = W*in
   wire signed [9:0] m102_84;
   assign m102_84 =10'b0;

   // m102_85 = W*in
   wire signed [9:0] m102_85;
   assign m102_85 =10'b0;

   // m102_86 = W*in
   wire signed [9:0] m102_86;
   assign m102_86 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_87 = W*in
   wire signed [9:0] m102_87;
   assign m102_87 =10'b0;

   // m102_88 = W*in
   wire signed [9:0] m102_88;
   assign m102_88 =10'b0;

   // m102_89 = W*in
   wire signed [9:0] m102_89;
   assign m102_89 =10'b0;

   // m102_90 = W*in
   wire signed [9:0] m102_90;
   assign m102_90 =10'b0;

   // m102_91 = W*in
   wire signed [9:0] m102_91;
   assign m102_91 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_92 = W*in
   wire signed [9:0] m102_92;
   assign m102_92 =10'b0;

   // m102_93 = W*in
   wire signed [9:0] m102_93;
   assign m102_93 =10'b0;

   // m102_94 = W*in
   wire signed [9:0] m102_94;
   assign m102_94 =10'b0;

   // m102_95 = W*in
   wire signed [9:0] m102_95;
   assign m102_95 =10'b0;

   // m102_96 = W*in
   wire signed [9:0] m102_96;
   assign m102_96 =10'b0;

   // m102_97 = W*in
   wire signed [9:0] m102_97;
   assign m102_97 =10'b0;

   // m102_98 = W*in
   wire signed [9:0] m102_98;
   assign m102_98 ={ {4{in102[5]}} , in102[5:0] };

   // m102_99 = W*in
   wire signed [9:0] m102_99;
   assign m102_99 ={ {4{neg102[5]}} , neg102[5:0] };

   // m102_100 = W*in
   wire signed [9:0] m102_100;
   assign m102_100 =10'b0;

   // m102_101 = W*in
   wire signed [9:0] m102_101;
   assign m102_101 =10'b0;

   // m102_102 = W*in
   wire signed [9:0] m102_102;
   assign m102_102 =10'b0;

   // m102_103 = W*in
   wire signed [9:0] m102_103;
   assign m102_103 =10'b0;

   // m102_104 = W*in
   wire signed [9:0] m102_104;
   assign m102_104 =10'b0;

   // m102_105 = W*in
   wire signed [9:0] m102_105;
   assign m102_105 =10'b0;

   // m102_106 = W*in
   wire signed [9:0] m102_106;
   assign m102_106 ={ {4{in102[5]}} , in102[5:0] };

   // m102_107 = W*in
   wire signed [9:0] m102_107;
   assign m102_107 =10'b0;

   // m102_108 = W*in
   wire signed [9:0] m102_108;
   assign m102_108 ={ {4{in102[5]}} , in102[5:0] };

   // m102_109 = W*in
   wire signed [9:0] m102_109;
   assign m102_109 =10'b0;

   // m102_110 = W*in
   wire signed [9:0] m102_110;
   assign m102_110 =10'b0;

   // m102_111 = W*in
   wire signed [9:0] m102_111;
   assign m102_111 =10'b0;

   // m102_112 = W*in
   wire signed [9:0] m102_112;
   assign m102_112 =10'b0;

   // m102_113 = W*in
   wire signed [9:0] m102_113;
   assign m102_113 =10'b0;

   // m102_114 = W*in
   wire signed [9:0] m102_114;
   assign m102_114 =10'b0;

   // m102_115 = W*in
   wire signed [9:0] m102_115;
   assign m102_115 ={ {4{in102[5]}} , in102[5:0] };

   // m102_116 = W*in
   wire signed [9:0] m102_116;
   assign m102_116 ={ {4{in102[5]}} , in102[5:0] };

   // m102_117 = W*in
   wire signed [9:0] m102_117;
   assign m102_117 ={ {4{in102[5]}} , in102[5:0] };

   // m103_1 = W*in
   wire signed [9:0] m103_1;
   assign m103_1 ={ {4{in103[5]}} , in103[5:0] };

   // m103_2 = W*in
   wire signed [9:0] m103_2;
   assign m103_2 =10'b0;

   // m103_3 = W*in
   wire signed [9:0] m103_3;
   assign m103_3 =10'b0;

   // m103_4 = W*in
   wire signed [9:0] m103_4;
   assign m103_4 =10'b0;

   // m103_5 = W*in
   wire signed [9:0] m103_5;
   assign m103_5 =10'b0;

   // m103_6 = W*in
   wire signed [9:0] m103_6;
   assign m103_6 =10'b0;

   // m103_7 = W*in
   wire signed [9:0] m103_7;
   assign m103_7 =10'b0;

   // m103_8 = W*in
   wire signed [9:0] m103_8;
   assign m103_8 =10'b0;

   // m103_9 = W*in
   wire signed [9:0] m103_9;
   assign m103_9 =10'b0;

   // m103_10 = W*in
   wire signed [9:0] m103_10;
   assign m103_10 =10'b0;

   // m103_11 = W*in
   wire signed [9:0] m103_11;
   assign m103_11 =10'b0;

   // m103_12 = W*in
   wire signed [9:0] m103_12;
   assign m103_12 =10'b0;

   // m103_13 = W*in
   wire signed [9:0] m103_13;
   assign m103_13 ={ {4{in103[5]}} , in103[5:0] };

   // m103_14 = W*in
   wire signed [9:0] m103_14;
   assign m103_14 =10'b0;

   // m103_15 = W*in
   wire signed [9:0] m103_15;
   assign m103_15 =10'b0;

   // m103_16 = W*in
   wire signed [9:0] m103_16;
   assign m103_16 =10'b0;

   // m103_17 = W*in
   wire signed [9:0] m103_17;
   assign m103_17 ={ {4{in103[5]}} , in103[5:0] };

   // m103_18 = W*in
   wire signed [9:0] m103_18;
   assign m103_18 =10'b0;

   // m103_19 = W*in
   wire signed [9:0] m103_19;
   assign m103_19 =10'b0;

   // m103_20 = W*in
   wire signed [9:0] m103_20;
   assign m103_20 =10'b0;

   // m103_21 = W*in
   wire signed [9:0] m103_21;
   assign m103_21 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_22 = W*in
   wire signed [9:0] m103_22;
   assign m103_22 ={ {5{in103[5]}} , in103[5:1] };

   // m103_23 = W*in
   wire signed [9:0] m103_23;
   assign m103_23 =10'b0;

   // m103_24 = W*in
   wire signed [9:0] m103_24;
   assign m103_24 =10'b0;

   // m103_25 = W*in
   wire signed [9:0] m103_25;
   assign m103_25 ={ {4{in103[5]}} , in103[5:0] };

   // m103_26 = W*in
   wire signed [9:0] m103_26;
   assign m103_26 =10'b0;

   // m103_27 = W*in
   wire signed [9:0] m103_27;
   assign m103_27 =10'b0;

   // m103_28 = W*in
   wire signed [9:0] m103_28;
   assign m103_28 =10'b0;

   // m103_29 = W*in
   wire signed [9:0] m103_29;
   assign m103_29 =10'b0;

   // m103_30 = W*in
   wire signed [9:0] m103_30;
   assign m103_30 =10'b0;

   // m103_31 = W*in
   wire signed [9:0] m103_31;
   assign m103_31 =10'b0;

   // m103_32 = W*in
   wire signed [9:0] m103_32;
   assign m103_32 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_33 = W*in
   wire signed [9:0] m103_33;
   assign m103_33 ={ {4{in103[5]}} , in103[5:0] };

   // m103_34 = W*in
   wire signed [9:0] m103_34;
   assign m103_34 =10'b0;

   // m103_35 = W*in
   wire signed [9:0] m103_35;
   assign m103_35 =10'b0;

   // m103_36 = W*in
   wire signed [9:0] m103_36;
   assign m103_36 ={ {4{in103[5]}} , in103[5:0] };

   // m103_37 = W*in
   wire signed [9:0] m103_37;
   assign m103_37 =10'b0;

   // m103_38 = W*in
   wire signed [9:0] m103_38;
   assign m103_38 =10'b0;

   // m103_39 = W*in
   wire signed [9:0] m103_39;
   assign m103_39 =10'b0;

   // m103_40 = W*in
   wire signed [9:0] m103_40;
   assign m103_40 =10'b0;

   // m103_41 = W*in
   wire signed [9:0] m103_41;
   assign m103_41 =10'b0;

   // m103_42 = W*in
   wire signed [9:0] m103_42;
   assign m103_42 =10'b0;

   // m103_43 = W*in
   wire signed [9:0] m103_43;
   assign m103_43 =10'b0;

   // m103_44 = W*in
   wire signed [9:0] m103_44;
   assign m103_44 =10'b0;

   // m103_45 = W*in
   wire signed [9:0] m103_45;
   assign m103_45 =10'b0;

   // m103_46 = W*in
   wire signed [9:0] m103_46;
   assign m103_46 =10'b0;

   // m103_47 = W*in
   wire signed [9:0] m103_47;
   assign m103_47 =10'b0;

   // m103_48 = W*in
   wire signed [9:0] m103_48;
   assign m103_48 =10'b0;

   // m103_49 = W*in
   wire signed [9:0] m103_49;
   assign m103_49 =10'b0;

   // m103_50 = W*in
   wire signed [9:0] m103_50;
   assign m103_50 =10'b0;

   // m103_51 = W*in
   wire signed [9:0] m103_51;
   assign m103_51 =10'b0;

   // m103_52 = W*in
   wire signed [9:0] m103_52;
   assign m103_52 =10'b0;

   // m103_53 = W*in
   wire signed [9:0] m103_53;
   assign m103_53 =10'b0;

   // m103_54 = W*in
   wire signed [9:0] m103_54;
   assign m103_54 =10'b0;

   // m103_55 = W*in
   wire signed [9:0] m103_55;
   assign m103_55 =10'b0;

   // m103_56 = W*in
   wire signed [9:0] m103_56;
   assign m103_56 =10'b0;

   // m103_57 = W*in
   wire signed [9:0] m103_57;
   assign m103_57 =10'b0;

   // m103_58 = W*in
   wire signed [9:0] m103_58;
   assign m103_58 =10'b0;

   // m103_59 = W*in
   wire signed [9:0] m103_59;
   assign m103_59 ={ {4{in103[5]}} , in103[5:0] };

   // m103_60 = W*in
   wire signed [9:0] m103_60;
   assign m103_60 =10'b0;

   // m103_61 = W*in
   wire signed [9:0] m103_61;
   assign m103_61 =10'b0;

   // m103_62 = W*in
   wire signed [9:0] m103_62;
   assign m103_62 =10'b0;

   // m103_63 = W*in
   wire signed [9:0] m103_63;
   assign m103_63 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_64 = W*in
   wire signed [9:0] m103_64;
   assign m103_64 ={ {5{neg103[5]}} , neg103[5:1] };

   // m103_65 = W*in
   wire signed [9:0] m103_65;
   assign m103_65 =10'b0;

   // m103_66 = W*in
   wire signed [9:0] m103_66;
   assign m103_66 =10'b0;

   // m103_67 = W*in
   wire signed [9:0] m103_67;
   assign m103_67 =10'b0;

   // m103_68 = W*in
   wire signed [9:0] m103_68;
   assign m103_68 =10'b0;

   // m103_69 = W*in
   wire signed [9:0] m103_69;
   assign m103_69 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_70 = W*in
   wire signed [9:0] m103_70;
   assign m103_70 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_71 = W*in
   wire signed [9:0] m103_71;
   assign m103_71 ={ {5{neg103[5]}} , neg103[5:1] };

   // m103_72 = W*in
   wire signed [9:0] m103_72;
   assign m103_72 ={ {5{neg103[5]}} , neg103[5:1] };

   // m103_73 = W*in
   wire signed [9:0] m103_73;
   assign m103_73 =10'b0;

   // m103_74 = W*in
   wire signed [9:0] m103_74;
   assign m103_74 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_75 = W*in
   wire signed [9:0] m103_75;
   assign m103_75 ={ {5{in103[5]}} , in103[5:1] };

   // m103_76 = W*in
   wire signed [9:0] m103_76;
   assign m103_76 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_77 = W*in
   wire signed [9:0] m103_77;
   assign m103_77 =10'b0;

   // m103_78 = W*in
   wire signed [9:0] m103_78;
   assign m103_78 ={ {4{in103[5]}} , in103[5:0] };

   // m103_79 = W*in
   wire signed [9:0] m103_79;
   assign m103_79 =10'b0;

   // m103_80 = W*in
   wire signed [9:0] m103_80;
   assign m103_80 =10'b0;

   // m103_81 = W*in
   wire signed [9:0] m103_81;
   assign m103_81 =10'b0;

   // m103_82 = W*in
   wire signed [9:0] m103_82;
   assign m103_82 ={ {5{neg103[5]}} , neg103[5:1] };

   // m103_83 = W*in
   wire signed [9:0] m103_83;
   assign m103_83 =10'b0;

   // m103_84 = W*in
   wire signed [9:0] m103_84;
   assign m103_84 =10'b0;

   // m103_85 = W*in
   wire signed [9:0] m103_85;
   assign m103_85 =10'b0;

   // m103_86 = W*in
   wire signed [9:0] m103_86;
   assign m103_86 =10'b0;

   // m103_87 = W*in
   wire signed [9:0] m103_87;
   assign m103_87 =10'b0;

   // m103_88 = W*in
   wire signed [9:0] m103_88;
   assign m103_88 =10'b0;

   // m103_89 = W*in
   wire signed [9:0] m103_89;
   assign m103_89 =10'b0;

   // m103_90 = W*in
   wire signed [9:0] m103_90;
   assign m103_90 =10'b0;

   // m103_91 = W*in
   wire signed [9:0] m103_91;
   assign m103_91 =10'b0;

   // m103_92 = W*in
   wire signed [9:0] m103_92;
   assign m103_92 =10'b0;

   // m103_93 = W*in
   wire signed [9:0] m103_93;
   assign m103_93 =10'b0;

   // m103_94 = W*in
   wire signed [9:0] m103_94;
   assign m103_94 =10'b0;

   // m103_95 = W*in
   wire signed [9:0] m103_95;
   assign m103_95 =10'b0;

   // m103_96 = W*in
   wire signed [9:0] m103_96;
   assign m103_96 =10'b0;

   // m103_97 = W*in
   wire signed [9:0] m103_97;
   assign m103_97 =10'b0;

   // m103_98 = W*in
   wire signed [9:0] m103_98;
   assign m103_98 =10'b0;

   // m103_99 = W*in
   wire signed [9:0] m103_99;
   assign m103_99 ={ {4{neg103[5]}} , neg103[5:0] };

   // m103_100 = W*in
   wire signed [9:0] m103_100;
   assign m103_100 =10'b0;

   // m103_101 = W*in
   wire signed [9:0] m103_101;
   assign m103_101 =10'b0;

   // m103_102 = W*in
   wire signed [9:0] m103_102;
   assign m103_102 =10'b0;

   // m103_103 = W*in
   wire signed [9:0] m103_103;
   assign m103_103 =10'b0;

   // m103_104 = W*in
   wire signed [9:0] m103_104;
   assign m103_104 =10'b0;

   // m103_105 = W*in
   wire signed [9:0] m103_105;
   assign m103_105 =10'b0;

   // m103_106 = W*in
   wire signed [9:0] m103_106;
   assign m103_106 =10'b0;

   // m103_107 = W*in
   wire signed [9:0] m103_107;
   assign m103_107 =10'b0;

   // m103_108 = W*in
   wire signed [9:0] m103_108;
   assign m103_108 =10'b0;

   // m103_109 = W*in
   wire signed [9:0] m103_109;
   assign m103_109 =10'b0;

   // m103_110 = W*in
   wire signed [9:0] m103_110;
   assign m103_110 =10'b0;

   // m103_111 = W*in
   wire signed [9:0] m103_111;
   assign m103_111 =10'b0;

   // m103_112 = W*in
   wire signed [9:0] m103_112;
   assign m103_112 =10'b0;

   // m103_113 = W*in
   wire signed [9:0] m103_113;
   assign m103_113 =10'b0;

   // m103_114 = W*in
   wire signed [9:0] m103_114;
   assign m103_114 =10'b0;

   // m103_115 = W*in
   wire signed [9:0] m103_115;
   assign m103_115 =10'b0;

   // m103_116 = W*in
   wire signed [9:0] m103_116;
   assign m103_116 =10'b0;

   // m103_117 = W*in
   wire signed [9:0] m103_117;
   assign m103_117 =10'b0;

   // m104_1 = W*in
   wire signed [9:0] m104_1;
   assign m104_1 =10'b0;

   // m104_2 = W*in
   wire signed [9:0] m104_2;
   assign m104_2 =10'b0;

   // m104_3 = W*in
   wire signed [9:0] m104_3;
   assign m104_3 =10'b0;

   // m104_4 = W*in
   wire signed [9:0] m104_4;
   assign m104_4 =10'b0;

   // m104_5 = W*in
   wire signed [9:0] m104_5;
   assign m104_5 =10'b0;

   // m104_6 = W*in
   wire signed [9:0] m104_6;
   assign m104_6 =10'b0;

   // m104_7 = W*in
   wire signed [9:0] m104_7;
   assign m104_7 =10'b0;

   // m104_8 = W*in
   wire signed [9:0] m104_8;
   assign m104_8 =10'b0;

   // m104_9 = W*in
   wire signed [9:0] m104_9;
   assign m104_9 =10'b0;

   // m104_10 = W*in
   wire signed [9:0] m104_10;
   assign m104_10 =10'b0;

   // m104_11 = W*in
   wire signed [9:0] m104_11;
   assign m104_11 =10'b0;

   // m104_12 = W*in
   wire signed [9:0] m104_12;
   assign m104_12 =10'b0;

   // m104_13 = W*in
   wire signed [9:0] m104_13;
   assign m104_13 ={ {4{in104[5]}} , in104[5:0] };

   // m104_14 = W*in
   wire signed [9:0] m104_14;
   assign m104_14 =10'b0;

   // m104_15 = W*in
   wire signed [9:0] m104_15;
   assign m104_15 =10'b0;

   // m104_16 = W*in
   wire signed [9:0] m104_16;
   assign m104_16 =10'b0;

   // m104_17 = W*in
   wire signed [9:0] m104_17;
   assign m104_17 =10'b0;

   // m104_18 = W*in
   wire signed [9:0] m104_18;
   assign m104_18 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_19 = W*in
   wire signed [9:0] m104_19;
   assign m104_19 =10'b0;

   // m104_20 = W*in
   wire signed [9:0] m104_20;
   assign m104_20 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_21 = W*in
   wire signed [9:0] m104_21;
   assign m104_21 =10'b0;

   // m104_22 = W*in
   wire signed [9:0] m104_22;
   assign m104_22 =10'b0;

   // m104_23 = W*in
   wire signed [9:0] m104_23;
   assign m104_23 =10'b0;

   // m104_24 = W*in
   wire signed [9:0] m104_24;
   assign m104_24 =10'b0;

   // m104_25 = W*in
   wire signed [9:0] m104_25;
   assign m104_25 =10'b0;

   // m104_26 = W*in
   wire signed [9:0] m104_26;
   assign m104_26 =10'b0;

   // m104_27 = W*in
   wire signed [9:0] m104_27;
   assign m104_27 =10'b0;

   // m104_28 = W*in
   wire signed [9:0] m104_28;
   assign m104_28 =10'b0;

   // m104_29 = W*in
   wire signed [9:0] m104_29;
   assign m104_29 =10'b0;

   // m104_30 = W*in
   wire signed [9:0] m104_30;
   assign m104_30 ={ {4{neg104[5]}} , neg104[5:0] };

   // m104_31 = W*in
   wire signed [9:0] m104_31;
   assign m104_31 =10'b0;

   // m104_32 = W*in
   wire signed [9:0] m104_32;
   assign m104_32 =10'b0;

   // m104_33 = W*in
   wire signed [9:0] m104_33;
   assign m104_33 =10'b0;

   // m104_34 = W*in
   wire signed [9:0] m104_34;
   assign m104_34 =10'b0;

   // m104_35 = W*in
   wire signed [9:0] m104_35;
   assign m104_35 =10'b0;

   // m104_36 = W*in
   wire signed [9:0] m104_36;
   assign m104_36 ={ {4{in104[5]}} , in104[5:0] };

   // m104_37 = W*in
   wire signed [9:0] m104_37;
   assign m104_37 =10'b0;

   // m104_38 = W*in
   wire signed [9:0] m104_38;
   assign m104_38 =10'b0;

   // m104_39 = W*in
   wire signed [9:0] m104_39;
   assign m104_39 =10'b0;

   // m104_40 = W*in
   wire signed [9:0] m104_40;
   assign m104_40 =10'b0;

   // m104_41 = W*in
   wire signed [9:0] m104_41;
   assign m104_41 =10'b0;

   // m104_42 = W*in
   wire signed [9:0] m104_42;
   assign m104_42 =10'b0;

   // m104_43 = W*in
   wire signed [9:0] m104_43;
   assign m104_43 =10'b0;

   // m104_44 = W*in
   wire signed [9:0] m104_44;
   assign m104_44 =10'b0;

   // m104_45 = W*in
   wire signed [9:0] m104_45;
   assign m104_45 =10'b0;

   // m104_46 = W*in
   wire signed [9:0] m104_46;
   assign m104_46 =10'b0;

   // m104_47 = W*in
   wire signed [9:0] m104_47;
   assign m104_47 =10'b0;

   // m104_48 = W*in
   wire signed [9:0] m104_48;
   assign m104_48 =10'b0;

   // m104_49 = W*in
   wire signed [9:0] m104_49;
   assign m104_49 =10'b0;

   // m104_50 = W*in
   wire signed [9:0] m104_50;
   assign m104_50 =10'b0;

   // m104_51 = W*in
   wire signed [9:0] m104_51;
   assign m104_51 =10'b0;

   // m104_52 = W*in
   wire signed [9:0] m104_52;
   assign m104_52 =10'b0;

   // m104_53 = W*in
   wire signed [9:0] m104_53;
   assign m104_53 =10'b0;

   // m104_54 = W*in
   wire signed [9:0] m104_54;
   assign m104_54 =10'b0;

   // m104_55 = W*in
   wire signed [9:0] m104_55;
   assign m104_55 =10'b0;

   // m104_56 = W*in
   wire signed [9:0] m104_56;
   assign m104_56 ={ {4{in104[5]}} , in104[5:0] };

   // m104_57 = W*in
   wire signed [9:0] m104_57;
   assign m104_57 =10'b0;

   // m104_58 = W*in
   wire signed [9:0] m104_58;
   assign m104_58 =10'b0;

   // m104_59 = W*in
   wire signed [9:0] m104_59;
   assign m104_59 =10'b0;

   // m104_60 = W*in
   wire signed [9:0] m104_60;
   assign m104_60 =10'b0;

   // m104_61 = W*in
   wire signed [9:0] m104_61;
   assign m104_61 =10'b0;

   // m104_62 = W*in
   wire signed [9:0] m104_62;
   assign m104_62 =10'b0;

   // m104_63 = W*in
   wire signed [9:0] m104_63;
   assign m104_63 =10'b0;

   // m104_64 = W*in
   wire signed [9:0] m104_64;
   assign m104_64 =10'b0;

   // m104_65 = W*in
   wire signed [9:0] m104_65;
   assign m104_65 =10'b0;

   // m104_66 = W*in
   wire signed [9:0] m104_66;
   assign m104_66 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_67 = W*in
   wire signed [9:0] m104_67;
   assign m104_67 =10'b0;

   // m104_68 = W*in
   wire signed [9:0] m104_68;
   assign m104_68 =10'b0;

   // m104_69 = W*in
   wire signed [9:0] m104_69;
   assign m104_69 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_70 = W*in
   wire signed [9:0] m104_70;
   assign m104_70 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_71 = W*in
   wire signed [9:0] m104_71;
   assign m104_71 =10'b0;

   // m104_72 = W*in
   wire signed [9:0] m104_72;
   assign m104_72 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_73 = W*in
   wire signed [9:0] m104_73;
   assign m104_73 =10'b0;

   // m104_74 = W*in
   wire signed [9:0] m104_74;
   assign m104_74 ={ {4{neg104[5]}} , neg104[5:0] };

   // m104_75 = W*in
   wire signed [9:0] m104_75;
   assign m104_75 =10'b0;

   // m104_76 = W*in
   wire signed [9:0] m104_76;
   assign m104_76 =10'b0;

   // m104_77 = W*in
   wire signed [9:0] m104_77;
   assign m104_77 =10'b0;

   // m104_78 = W*in
   wire signed [9:0] m104_78;
   assign m104_78 ={ {4{in104[5]}} , in104[5:0] };

   // m104_79 = W*in
   wire signed [9:0] m104_79;
   assign m104_79 =10'b0;

   // m104_80 = W*in
   wire signed [9:0] m104_80;
   assign m104_80 =10'b0;

   // m104_81 = W*in
   wire signed [9:0] m104_81;
   assign m104_81 ={ {5{neg104[5]}} , neg104[5:1] };

   // m104_82 = W*in
   wire signed [9:0] m104_82;
   assign m104_82 =10'b0;

   // m104_83 = W*in
   wire signed [9:0] m104_83;
   assign m104_83 =10'b0;

   // m104_84 = W*in
   wire signed [9:0] m104_84;
   assign m104_84 =10'b0;

   // m104_85 = W*in
   wire signed [9:0] m104_85;
   assign m104_85 =10'b0;

   // m104_86 = W*in
   wire signed [9:0] m104_86;
   assign m104_86 =10'b0;

   // m104_87 = W*in
   wire signed [9:0] m104_87;
   assign m104_87 =10'b0;

   // m104_88 = W*in
   wire signed [9:0] m104_88;
   assign m104_88 ={ {4{neg104[5]}} , neg104[5:0] };

   // m104_89 = W*in
   wire signed [9:0] m104_89;
   assign m104_89 =10'b0;

   // m104_90 = W*in
   wire signed [9:0] m104_90;
   assign m104_90 =10'b0;

   // m104_91 = W*in
   wire signed [9:0] m104_91;
   assign m104_91 =10'b0;

   // m104_92 = W*in
   wire signed [9:0] m104_92;
   assign m104_92 =10'b0;

   // m104_93 = W*in
   wire signed [9:0] m104_93;
   assign m104_93 =10'b0;

   // m104_94 = W*in
   wire signed [9:0] m104_94;
   assign m104_94 =10'b0;

   // m104_95 = W*in
   wire signed [9:0] m104_95;
   assign m104_95 =10'b0;

   // m104_96 = W*in
   wire signed [9:0] m104_96;
   assign m104_96 =10'b0;

   // m104_97 = W*in
   wire signed [9:0] m104_97;
   assign m104_97 =10'b0;

   // m104_98 = W*in
   wire signed [9:0] m104_98;
   assign m104_98 =10'b0;

   // m104_99 = W*in
   wire signed [9:0] m104_99;
   assign m104_99 =10'b0;

   // m104_100 = W*in
   wire signed [9:0] m104_100;
   assign m104_100 =10'b0;

   // m104_101 = W*in
   wire signed [9:0] m104_101;
   assign m104_101 =10'b0;

   // m104_102 = W*in
   wire signed [9:0] m104_102;
   assign m104_102 =10'b0;

   // m104_103 = W*in
   wire signed [9:0] m104_103;
   assign m104_103 =10'b0;

   // m104_104 = W*in
   wire signed [9:0] m104_104;
   assign m104_104 =10'b0;

   // m104_105 = W*in
   wire signed [9:0] m104_105;
   assign m104_105 =10'b0;

   // m104_106 = W*in
   wire signed [9:0] m104_106;
   assign m104_106 =10'b0;

   // m104_107 = W*in
   wire signed [9:0] m104_107;
   assign m104_107 =10'b0;

   // m104_108 = W*in
   wire signed [9:0] m104_108;
   assign m104_108 ={ {4{neg104[5]}} , neg104[5:0] };

   // m104_109 = W*in
   wire signed [9:0] m104_109;
   assign m104_109 ={ {4{neg104[5]}} , neg104[5:0] };

   // m104_110 = W*in
   wire signed [9:0] m104_110;
   assign m104_110 =10'b0;

   // m104_111 = W*in
   wire signed [9:0] m104_111;
   assign m104_111 =10'b0;

   // m104_112 = W*in
   wire signed [9:0] m104_112;
   assign m104_112 =10'b0;

   // m104_113 = W*in
   wire signed [9:0] m104_113;
   assign m104_113 =10'b0;

   // m104_114 = W*in
   wire signed [9:0] m104_114;
   assign m104_114 =10'b0;

   // m104_115 = W*in
   wire signed [9:0] m104_115;
   assign m104_115 =10'b0;

   // m104_116 = W*in
   wire signed [9:0] m104_116;
   assign m104_116 =10'b0;

   // m104_117 = W*in
   wire signed [9:0] m104_117;
   assign m104_117 =10'b0;

   // m105_1 = W*in
   wire signed [9:0] m105_1;
   assign m105_1 =10'b0;

   // m105_2 = W*in
   wire signed [9:0] m105_2;
   assign m105_2 =10'b0;

   // m105_3 = W*in
   wire signed [9:0] m105_3;
   assign m105_3 =10'b0;

   // m105_4 = W*in
   wire signed [9:0] m105_4;
   assign m105_4 =10'b0;

   // m105_5 = W*in
   wire signed [9:0] m105_5;
   assign m105_5 =10'b0;

   // m105_6 = W*in
   wire signed [9:0] m105_6;
   assign m105_6 =10'b0;

   // m105_7 = W*in
   wire signed [9:0] m105_7;
   assign m105_7 =10'b0;

   // m105_8 = W*in
   wire signed [9:0] m105_8;
   assign m105_8 =10'b0;

   // m105_9 = W*in
   wire signed [9:0] m105_9;
   assign m105_9 =10'b0;

   // m105_10 = W*in
   wire signed [9:0] m105_10;
   assign m105_10 =10'b0;

   // m105_11 = W*in
   wire signed [9:0] m105_11;
   assign m105_11 =10'b0;

   // m105_12 = W*in
   wire signed [9:0] m105_12;
   assign m105_12 =10'b0;

   // m105_13 = W*in
   wire signed [9:0] m105_13;
   assign m105_13 =10'b0;

   // m105_14 = W*in
   wire signed [9:0] m105_14;
   assign m105_14 =10'b0;

   // m105_15 = W*in
   wire signed [9:0] m105_15;
   assign m105_15 =10'b0;

   // m105_16 = W*in
   wire signed [9:0] m105_16;
   assign m105_16 =10'b0;

   // m105_17 = W*in
   wire signed [9:0] m105_17;
   assign m105_17 =10'b0;

   // m105_18 = W*in
   wire signed [9:0] m105_18;
   assign m105_18 ={ {5{in105[5]}} , in105[5:1] };

   // m105_19 = W*in
   wire signed [9:0] m105_19;
   assign m105_19 ={ {5{neg105[5]}} , neg105[5:1] };

   // m105_20 = W*in
   wire signed [9:0] m105_20;
   assign m105_20 ={ {4{in105[5]}} , in105[5:0] };

   // m105_21 = W*in
   wire signed [9:0] m105_21;
   assign m105_21 ={ {5{neg105[5]}} , neg105[5:1] };

   // m105_22 = W*in
   wire signed [9:0] m105_22;
   assign m105_22 =10'b0;

   // m105_23 = W*in
   wire signed [9:0] m105_23;
   assign m105_23 =10'b0;

   // m105_24 = W*in
   wire signed [9:0] m105_24;
   assign m105_24 =10'b0;

   // m105_25 = W*in
   wire signed [9:0] m105_25;
   assign m105_25 =10'b0;

   // m105_26 = W*in
   wire signed [9:0] m105_26;
   assign m105_26 =10'b0;

   // m105_27 = W*in
   wire signed [9:0] m105_27;
   assign m105_27 =10'b0;

   // m105_28 = W*in
   wire signed [9:0] m105_28;
   assign m105_28 =10'b0;

   // m105_29 = W*in
   wire signed [9:0] m105_29;
   assign m105_29 ={ {5{neg105[5]}} , neg105[5:1] };

   // m105_30 = W*in
   wire signed [9:0] m105_30;
   assign m105_30 ={ {4{in105[5]}} , in105[5:0] };

   // m105_31 = W*in
   wire signed [9:0] m105_31;
   assign m105_31 =10'b0;

   // m105_32 = W*in
   wire signed [9:0] m105_32;
   assign m105_32 =10'b0;

   // m105_33 = W*in
   wire signed [9:0] m105_33;
   assign m105_33 =10'b0;

   // m105_34 = W*in
   wire signed [9:0] m105_34;
   assign m105_34 =10'b0;

   // m105_35 = W*in
   wire signed [9:0] m105_35;
   assign m105_35 =10'b0;

   // m105_36 = W*in
   wire signed [9:0] m105_36;
   assign m105_36 =10'b0;

   // m105_37 = W*in
   wire signed [9:0] m105_37;
   assign m105_37 =10'b0;

   // m105_38 = W*in
   wire signed [9:0] m105_38;
   assign m105_38 =10'b0;

   // m105_39 = W*in
   wire signed [9:0] m105_39;
   assign m105_39 =10'b0;

   // m105_40 = W*in
   wire signed [9:0] m105_40;
   assign m105_40 =10'b0;

   // m105_41 = W*in
   wire signed [9:0] m105_41;
   assign m105_41 =10'b0;

   // m105_42 = W*in
   wire signed [9:0] m105_42;
   assign m105_42 =10'b0;

   // m105_43 = W*in
   wire signed [9:0] m105_43;
   assign m105_43 =10'b0;

   // m105_44 = W*in
   wire signed [9:0] m105_44;
   assign m105_44 =10'b0;

   // m105_45 = W*in
   wire signed [9:0] m105_45;
   assign m105_45 =10'b0;

   // m105_46 = W*in
   wire signed [9:0] m105_46;
   assign m105_46 =10'b0;

   // m105_47 = W*in
   wire signed [9:0] m105_47;
   assign m105_47 =10'b0;

   // m105_48 = W*in
   wire signed [9:0] m105_48;
   assign m105_48 ={ {4{in105[5]}} , in105[5:0] };

   // m105_49 = W*in
   wire signed [9:0] m105_49;
   assign m105_49 =10'b0;

   // m105_50 = W*in
   wire signed [9:0] m105_50;
   assign m105_50 ={ {4{in105[5]}} , in105[5:0] };

   // m105_51 = W*in
   wire signed [9:0] m105_51;
   assign m105_51 =10'b0;

   // m105_52 = W*in
   wire signed [9:0] m105_52;
   assign m105_52 =10'b0;

   // m105_53 = W*in
   wire signed [9:0] m105_53;
   assign m105_53 =10'b0;

   // m105_54 = W*in
   wire signed [9:0] m105_54;
   assign m105_54 =10'b0;

   // m105_55 = W*in
   wire signed [9:0] m105_55;
   assign m105_55 =10'b0;

   // m105_56 = W*in
   wire signed [9:0] m105_56;
   assign m105_56 =10'b0;

   // m105_57 = W*in
   wire signed [9:0] m105_57;
   assign m105_57 =10'b0;

   // m105_58 = W*in
   wire signed [9:0] m105_58;
   assign m105_58 =10'b0;

   // m105_59 = W*in
   wire signed [9:0] m105_59;
   assign m105_59 =10'b0;

   // m105_60 = W*in
   wire signed [9:0] m105_60;
   assign m105_60 ={ {4{neg105[5]}} , neg105[5:0] };

   // m105_61 = W*in
   wire signed [9:0] m105_61;
   assign m105_61 =10'b0;

   // m105_62 = W*in
   wire signed [9:0] m105_62;
   assign m105_62 =10'b0;

   // m105_63 = W*in
   wire signed [9:0] m105_63;
   assign m105_63 =10'b0;

   // m105_64 = W*in
   wire signed [9:0] m105_64;
   assign m105_64 =10'b0;

   // m105_65 = W*in
   wire signed [9:0] m105_65;
   assign m105_65 ={ {5{neg105[5]}} , neg105[5:1] };

   // m105_66 = W*in
   wire signed [9:0] m105_66;
   assign m105_66 =10'b0;

   // m105_67 = W*in
   wire signed [9:0] m105_67;
   assign m105_67 =10'b0;

   // m105_68 = W*in
   wire signed [9:0] m105_68;
   assign m105_68 =10'b0;

   // m105_69 = W*in
   wire signed [9:0] m105_69;
   assign m105_69 =10'b0;

   // m105_70 = W*in
   wire signed [9:0] m105_70;
   assign m105_70 ={ {5{neg105[5]}} , neg105[5:1] };

   // m105_71 = W*in
   wire signed [9:0] m105_71;
   assign m105_71 =10'b0;

   // m105_72 = W*in
   wire signed [9:0] m105_72;
   assign m105_72 ={ {5{in105[5]}} , in105[5:1] };

   // m105_73 = W*in
   wire signed [9:0] m105_73;
   assign m105_73 =10'b0;

   // m105_74 = W*in
   wire signed [9:0] m105_74;
   assign m105_74 ={ {5{in105[5]}} , in105[5:1] };

   // m105_75 = W*in
   wire signed [9:0] m105_75;
   assign m105_75 =10'b0;

   // m105_76 = W*in
   wire signed [9:0] m105_76;
   assign m105_76 =10'b0;

   // m105_77 = W*in
   wire signed [9:0] m105_77;
   assign m105_77 =10'b0;

   // m105_78 = W*in
   wire signed [9:0] m105_78;
   assign m105_78 =10'b0;

   // m105_79 = W*in
   wire signed [9:0] m105_79;
   assign m105_79 =10'b0;

   // m105_80 = W*in
   wire signed [9:0] m105_80;
   assign m105_80 =10'b0;

   // m105_81 = W*in
   wire signed [9:0] m105_81;
   assign m105_81 =10'b0;

   // m105_82 = W*in
   wire signed [9:0] m105_82;
   assign m105_82 =10'b0;

   // m105_83 = W*in
   wire signed [9:0] m105_83;
   assign m105_83 =10'b0;

   // m105_84 = W*in
   wire signed [9:0] m105_84;
   assign m105_84 =10'b0;

   // m105_85 = W*in
   wire signed [9:0] m105_85;
   assign m105_85 =10'b0;

   // m105_86 = W*in
   wire signed [9:0] m105_86;
   assign m105_86 =10'b0;

   // m105_87 = W*in
   wire signed [9:0] m105_87;
   assign m105_87 =10'b0;

   // m105_88 = W*in
   wire signed [9:0] m105_88;
   assign m105_88 =10'b0;

   // m105_89 = W*in
   wire signed [9:0] m105_89;
   assign m105_89 =10'b0;

   // m105_90 = W*in
   wire signed [9:0] m105_90;
   assign m105_90 =10'b0;

   // m105_91 = W*in
   wire signed [9:0] m105_91;
   assign m105_91 =10'b0;

   // m105_92 = W*in
   wire signed [9:0] m105_92;
   assign m105_92 ={ {4{in105[5]}} , in105[5:0] };

   // m105_93 = W*in
   wire signed [9:0] m105_93;
   assign m105_93 =10'b0;

   // m105_94 = W*in
   wire signed [9:0] m105_94;
   assign m105_94 =10'b0;

   // m105_95 = W*in
   wire signed [9:0] m105_95;
   assign m105_95 =10'b0;

   // m105_96 = W*in
   wire signed [9:0] m105_96;
   assign m105_96 =10'b0;

   // m105_97 = W*in
   wire signed [9:0] m105_97;
   assign m105_97 =10'b0;

   // m105_98 = W*in
   wire signed [9:0] m105_98;
   assign m105_98 =10'b0;

   // m105_99 = W*in
   wire signed [9:0] m105_99;
   assign m105_99 =10'b0;

   // m105_100 = W*in
   wire signed [9:0] m105_100;
   assign m105_100 =10'b0;

   // m105_101 = W*in
   wire signed [9:0] m105_101;
   assign m105_101 =10'b0;

   // m105_102 = W*in
   wire signed [9:0] m105_102;
   assign m105_102 =10'b0;

   // m105_103 = W*in
   wire signed [9:0] m105_103;
   assign m105_103 =10'b0;

   // m105_104 = W*in
   wire signed [9:0] m105_104;
   assign m105_104 =10'b0;

   // m105_105 = W*in
   wire signed [9:0] m105_105;
   assign m105_105 =10'b0;

   // m105_106 = W*in
   wire signed [9:0] m105_106;
   assign m105_106 =10'b0;

   // m105_107 = W*in
   wire signed [9:0] m105_107;
   assign m105_107 =10'b0;

   // m105_108 = W*in
   wire signed [9:0] m105_108;
   assign m105_108 =10'b0;

   // m105_109 = W*in
   wire signed [9:0] m105_109;
   assign m105_109 =10'b0;

   // m105_110 = W*in
   wire signed [9:0] m105_110;
   assign m105_110 =10'b0;

   // m105_111 = W*in
   wire signed [9:0] m105_111;
   assign m105_111 =10'b0;

   // m105_112 = W*in
   wire signed [9:0] m105_112;
   assign m105_112 =10'b0;

   // m105_113 = W*in
   wire signed [9:0] m105_113;
   assign m105_113 ={ {4{in105[5]}} , in105[5:0] };

   // m105_114 = W*in
   wire signed [9:0] m105_114;
   assign m105_114 =10'b0;

   // m105_115 = W*in
   wire signed [9:0] m105_115;
   assign m105_115 =10'b0;

   // m105_116 = W*in
   wire signed [9:0] m105_116;
   assign m105_116 =10'b0;

   // m105_117 = W*in
   wire signed [9:0] m105_117;
   assign m105_117 =10'b0;

   // m106_1 = W*in
   wire signed [9:0] m106_1;
   assign m106_1 =10'b0;

   // m106_2 = W*in
   wire signed [9:0] m106_2;
   assign m106_2 =10'b0;

   // m106_3 = W*in
   wire signed [9:0] m106_3;
   assign m106_3 =10'b0;

   // m106_4 = W*in
   wire signed [9:0] m106_4;
   assign m106_4 =10'b0;

   // m106_5 = W*in
   wire signed [9:0] m106_5;
   assign m106_5 =10'b0;

   // m106_6 = W*in
   wire signed [9:0] m106_6;
   assign m106_6 =10'b0;

   // m106_7 = W*in
   wire signed [9:0] m106_7;
   assign m106_7 =10'b0;

   // m106_8 = W*in
   wire signed [9:0] m106_8;
   assign m106_8 =10'b0;

   // m106_9 = W*in
   wire signed [9:0] m106_9;
   assign m106_9 =10'b0;

   // m106_10 = W*in
   wire signed [9:0] m106_10;
   assign m106_10 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_11 = W*in
   wire signed [9:0] m106_11;
   assign m106_11 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_12 = W*in
   wire signed [9:0] m106_12;
   assign m106_12 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_13 = W*in
   wire signed [9:0] m106_13;
   assign m106_13 =10'b0;

   // m106_14 = W*in
   wire signed [9:0] m106_14;
   assign m106_14 =10'b0;

   // m106_15 = W*in
   wire signed [9:0] m106_15;
   assign m106_15 ={ {4{in106[5]}} , in106[5:0] };

   // m106_16 = W*in
   wire signed [9:0] m106_16;
   assign m106_16 =10'b0;

   // m106_17 = W*in
   wire signed [9:0] m106_17;
   assign m106_17 =10'b0;

   // m106_18 = W*in
   wire signed [9:0] m106_18;
   assign m106_18 =10'b0;

   // m106_19 = W*in
   wire signed [9:0] m106_19;
   assign m106_19 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_20 = W*in
   wire signed [9:0] m106_20;
   assign m106_20 ={ {5{in106[5]}} , in106[5:1] };

   // m106_21 = W*in
   wire signed [9:0] m106_21;
   assign m106_21 ={ {5{neg106[5]}} , neg106[5:1] };

   // m106_22 = W*in
   wire signed [9:0] m106_22;
   assign m106_22 ={ {4{in106[5]}} , in106[5:0] };

   // m106_23 = W*in
   wire signed [9:0] m106_23;
   assign m106_23 ={ {4{in106[5]}} , in106[5:0] };

   // m106_24 = W*in
   wire signed [9:0] m106_24;
   assign m106_24 ={ {4{in106[5]}} , in106[5:0] };

   // m106_25 = W*in
   wire signed [9:0] m106_25;
   assign m106_25 =10'b0;

   // m106_26 = W*in
   wire signed [9:0] m106_26;
   assign m106_26 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_27 = W*in
   wire signed [9:0] m106_27;
   assign m106_27 =10'b0;

   // m106_28 = W*in
   wire signed [9:0] m106_28;
   assign m106_28 =10'b0;

   // m106_29 = W*in
   wire signed [9:0] m106_29;
   assign m106_29 ={ {5{neg106[5]}} , neg106[5:1] };

   // m106_30 = W*in
   wire signed [9:0] m106_30;
   assign m106_30 =10'b0;

   // m106_31 = W*in
   wire signed [9:0] m106_31;
   assign m106_31 =10'b0;

   // m106_32 = W*in
   wire signed [9:0] m106_32;
   assign m106_32 =10'b0;

   // m106_33 = W*in
   wire signed [9:0] m106_33;
   assign m106_33 =10'b0;

   // m106_34 = W*in
   wire signed [9:0] m106_34;
   assign m106_34 ={ {4{in106[5]}} , in106[5:0] };

   // m106_35 = W*in
   wire signed [9:0] m106_35;
   assign m106_35 =10'b0;

   // m106_36 = W*in
   wire signed [9:0] m106_36;
   assign m106_36 =10'b0;

   // m106_37 = W*in
   wire signed [9:0] m106_37;
   assign m106_37 =10'b0;

   // m106_38 = W*in
   wire signed [9:0] m106_38;
   assign m106_38 =10'b0;

   // m106_39 = W*in
   wire signed [9:0] m106_39;
   assign m106_39 =10'b0;

   // m106_40 = W*in
   wire signed [9:0] m106_40;
   assign m106_40 =10'b0;

   // m106_41 = W*in
   wire signed [9:0] m106_41;
   assign m106_41 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_42 = W*in
   wire signed [9:0] m106_42;
   assign m106_42 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_43 = W*in
   wire signed [9:0] m106_43;
   assign m106_43 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_44 = W*in
   wire signed [9:0] m106_44;
   assign m106_44 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_45 = W*in
   wire signed [9:0] m106_45;
   assign m106_45 =10'b0;

   // m106_46 = W*in
   wire signed [9:0] m106_46;
   assign m106_46 =10'b0;

   // m106_47 = W*in
   wire signed [9:0] m106_47;
   assign m106_47 ={ {4{in106[5]}} , in106[5:0] };

   // m106_48 = W*in
   wire signed [9:0] m106_48;
   assign m106_48 =10'b0;

   // m106_49 = W*in
   wire signed [9:0] m106_49;
   assign m106_49 =10'b0;

   // m106_50 = W*in
   wire signed [9:0] m106_50;
   assign m106_50 ={ {4{in106[5]}} , in106[5:0] };

   // m106_51 = W*in
   wire signed [9:0] m106_51;
   assign m106_51 ={ {4{in106[5]}} , in106[5:0] };

   // m106_52 = W*in
   wire signed [9:0] m106_52;
   assign m106_52 =10'b0;

   // m106_53 = W*in
   wire signed [9:0] m106_53;
   assign m106_53 =10'b0;

   // m106_54 = W*in
   wire signed [9:0] m106_54;
   assign m106_54 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_55 = W*in
   wire signed [9:0] m106_55;
   assign m106_55 =10'b0;

   // m106_56 = W*in
   wire signed [9:0] m106_56;
   assign m106_56 =10'b0;

   // m106_57 = W*in
   wire signed [9:0] m106_57;
   assign m106_57 =10'b0;

   // m106_58 = W*in
   wire signed [9:0] m106_58;
   assign m106_58 =10'b0;

   // m106_59 = W*in
   wire signed [9:0] m106_59;
   assign m106_59 =10'b0;

   // m106_60 = W*in
   wire signed [9:0] m106_60;
   assign m106_60 ={ {4{in106[5]}} , in106[5:0] };

   // m106_61 = W*in
   wire signed [9:0] m106_61;
   assign m106_61 =10'b0;

   // m106_62 = W*in
   wire signed [9:0] m106_62;
   assign m106_62 =10'b0;

   // m106_63 = W*in
   wire signed [9:0] m106_63;
   assign m106_63 =10'b0;

   // m106_64 = W*in
   wire signed [9:0] m106_64;
   assign m106_64 =10'b0;

   // m106_65 = W*in
   wire signed [9:0] m106_65;
   assign m106_65 =10'b0;

   // m106_66 = W*in
   wire signed [9:0] m106_66;
   assign m106_66 ={ {5{neg106[5]}} , neg106[5:1] };

   // m106_67 = W*in
   wire signed [9:0] m106_67;
   assign m106_67 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_68 = W*in
   wire signed [9:0] m106_68;
   assign m106_68 =10'b0;

   // m106_69 = W*in
   wire signed [9:0] m106_69;
   assign m106_69 =10'b0;

   // m106_70 = W*in
   wire signed [9:0] m106_70;
   assign m106_70 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_71 = W*in
   wire signed [9:0] m106_71;
   assign m106_71 =10'b0;

   // m106_72 = W*in
   wire signed [9:0] m106_72;
   assign m106_72 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_73 = W*in
   wire signed [9:0] m106_73;
   assign m106_73 ={ {4{in106[5]}} , in106[5:0] };

   // m106_74 = W*in
   wire signed [9:0] m106_74;
   assign m106_74 =10'b0;

   // m106_75 = W*in
   wire signed [9:0] m106_75;
   assign m106_75 ={ {5{in106[5]}} , in106[5:1] };

   // m106_76 = W*in
   wire signed [9:0] m106_76;
   assign m106_76 =10'b0;

   // m106_77 = W*in
   wire signed [9:0] m106_77;
   assign m106_77 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_78 = W*in
   wire signed [9:0] m106_78;
   assign m106_78 =10'b0;

   // m106_79 = W*in
   wire signed [9:0] m106_79;
   assign m106_79 =10'b0;

   // m106_80 = W*in
   wire signed [9:0] m106_80;
   assign m106_80 =10'b0;

   // m106_81 = W*in
   wire signed [9:0] m106_81;
   assign m106_81 =10'b0;

   // m106_82 = W*in
   wire signed [9:0] m106_82;
   assign m106_82 ={ {5{in106[5]}} , in106[5:1] };

   // m106_83 = W*in
   wire signed [9:0] m106_83;
   assign m106_83 =10'b0;

   // m106_84 = W*in
   wire signed [9:0] m106_84;
   assign m106_84 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_85 = W*in
   wire signed [9:0] m106_85;
   assign m106_85 =10'b0;

   // m106_86 = W*in
   wire signed [9:0] m106_86;
   assign m106_86 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_87 = W*in
   wire signed [9:0] m106_87;
   assign m106_87 ={ {4{in106[5]}} , in106[5:0] };

   // m106_88 = W*in
   wire signed [9:0] m106_88;
   assign m106_88 =10'b0;

   // m106_89 = W*in
   wire signed [9:0] m106_89;
   assign m106_89 =10'b0;

   // m106_90 = W*in
   wire signed [9:0] m106_90;
   assign m106_90 ={ {4{in106[5]}} , in106[5:0] };

   // m106_91 = W*in
   wire signed [9:0] m106_91;
   assign m106_91 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_92 = W*in
   wire signed [9:0] m106_92;
   assign m106_92 =10'b0;

   // m106_93 = W*in
   wire signed [9:0] m106_93;
   assign m106_93 =10'b0;

   // m106_94 = W*in
   wire signed [9:0] m106_94;
   assign m106_94 =10'b0;

   // m106_95 = W*in
   wire signed [9:0] m106_95;
   assign m106_95 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_96 = W*in
   wire signed [9:0] m106_96;
   assign m106_96 =10'b0;

   // m106_97 = W*in
   wire signed [9:0] m106_97;
   assign m106_97 ={ {3{neg106[5]}} , neg106 , {1{1'b0}} };

   // m106_98 = W*in
   wire signed [9:0] m106_98;
   assign m106_98 =10'b0;

   // m106_99 = W*in
   wire signed [9:0] m106_99;
   assign m106_99 =10'b0;

   // m106_100 = W*in
   wire signed [9:0] m106_100;
   assign m106_100 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_101 = W*in
   wire signed [9:0] m106_101;
   assign m106_101 =10'b0;

   // m106_102 = W*in
   wire signed [9:0] m106_102;
   assign m106_102 =10'b0;

   // m106_103 = W*in
   wire signed [9:0] m106_103;
   assign m106_103 =10'b0;

   // m106_104 = W*in
   wire signed [9:0] m106_104;
   assign m106_104 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_105 = W*in
   wire signed [9:0] m106_105;
   assign m106_105 =10'b0;

   // m106_106 = W*in
   wire signed [9:0] m106_106;
   assign m106_106 =10'b0;

   // m106_107 = W*in
   wire signed [9:0] m106_107;
   assign m106_107 =10'b0;

   // m106_108 = W*in
   wire signed [9:0] m106_108;
   assign m106_108 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_109 = W*in
   wire signed [9:0] m106_109;
   assign m106_109 ={ {3{in106[5]}} , in106 , {1{1'b0}} };

   // m106_110 = W*in
   wire signed [9:0] m106_110;
   assign m106_110 =10'b0;

   // m106_111 = W*in
   wire signed [9:0] m106_111;
   assign m106_111 =10'b0;

   // m106_112 = W*in
   wire signed [9:0] m106_112;
   assign m106_112 ={ {4{neg106[5]}} , neg106[5:0] };

   // m106_113 = W*in
   wire signed [9:0] m106_113;
   assign m106_113 =10'b0;

   // m106_114 = W*in
   wire signed [9:0] m106_114;
   assign m106_114 ={ {4{in106[5]}} , in106[5:0] };

   // m106_115 = W*in
   wire signed [9:0] m106_115;
   assign m106_115 =10'b0;

   // m106_116 = W*in
   wire signed [9:0] m106_116;
   assign m106_116 =10'b0;

   // m106_117 = W*in
   wire signed [9:0] m106_117;
   assign m106_117 ={ {4{in106[5]}} , in106[5:0] };

   // m107_1 = W*in
   wire signed [9:0] m107_1;
   assign m107_1 ={ {4{in107[5]}} , in107[5:0] };

   // m107_2 = W*in
   wire signed [9:0] m107_2;
   assign m107_2 =10'b0;

   // m107_3 = W*in
   wire signed [9:0] m107_3;
   assign m107_3 =10'b0;

   // m107_4 = W*in
   wire signed [9:0] m107_4;
   assign m107_4 ={ {5{in107[5]}} , in107[5:1] };

   // m107_5 = W*in
   wire signed [9:0] m107_5;
   assign m107_5 =10'b0;

   // m107_6 = W*in
   wire signed [9:0] m107_6;
   assign m107_6 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_7 = W*in
   wire signed [9:0] m107_7;
   assign m107_7 =10'b0;

   // m107_8 = W*in
   wire signed [9:0] m107_8;
   assign m107_8 =10'b0;

   // m107_9 = W*in
   wire signed [9:0] m107_9;
   assign m107_9 =10'b0;

   // m107_10 = W*in
   wire signed [9:0] m107_10;
   assign m107_10 =10'b0;

   // m107_11 = W*in
   wire signed [9:0] m107_11;
   assign m107_11 =10'b0;

   // m107_12 = W*in
   wire signed [9:0] m107_12;
   assign m107_12 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_13 = W*in
   wire signed [9:0] m107_13;
   assign m107_13 =10'b0;

   // m107_14 = W*in
   wire signed [9:0] m107_14;
   assign m107_14 =10'b0;

   // m107_15 = W*in
   wire signed [9:0] m107_15;
   assign m107_15 =10'b0;

   // m107_16 = W*in
   wire signed [9:0] m107_16;
   assign m107_16 =10'b0;

   // m107_17 = W*in
   wire signed [9:0] m107_17;
   assign m107_17 ={ {5{in107[5]}} , in107[5:1] };

   // m107_18 = W*in
   wire signed [9:0] m107_18;
   assign m107_18 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_19 = W*in
   wire signed [9:0] m107_19;
   assign m107_19 ={ {5{neg107[5]}} , neg107[5:1] };

   // m107_20 = W*in
   wire signed [9:0] m107_20;
   assign m107_20 ={ {5{in107[5]}} , in107[5:1] };

   // m107_21 = W*in
   wire signed [9:0] m107_21;
   assign m107_21 ={ {5{neg107[5]}} , neg107[5:1] };

   // m107_22 = W*in
   wire signed [9:0] m107_22;
   assign m107_22 ={ {5{in107[5]}} , in107[5:1] };

   // m107_23 = W*in
   wire signed [9:0] m107_23;
   assign m107_23 =10'b0;

   // m107_24 = W*in
   wire signed [9:0] m107_24;
   assign m107_24 ={ {5{in107[5]}} , in107[5:1] };

   // m107_25 = W*in
   wire signed [9:0] m107_25;
   assign m107_25 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_26 = W*in
   wire signed [9:0] m107_26;
   assign m107_26 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_27 = W*in
   wire signed [9:0] m107_27;
   assign m107_27 ={ {5{in107[5]}} , in107[5:1] };

   // m107_28 = W*in
   wire signed [9:0] m107_28;
   assign m107_28 ={ {5{neg107[5]}} , neg107[5:1] };

   // m107_29 = W*in
   wire signed [9:0] m107_29;
   assign m107_29 =10'b0;

   // m107_30 = W*in
   wire signed [9:0] m107_30;
   assign m107_30 =10'b0;

   // m107_31 = W*in
   wire signed [9:0] m107_31;
   assign m107_31 =10'b0;

   // m107_32 = W*in
   wire signed [9:0] m107_32;
   assign m107_32 =10'b0;

   // m107_33 = W*in
   wire signed [9:0] m107_33;
   assign m107_33 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_34 = W*in
   wire signed [9:0] m107_34;
   assign m107_34 =10'b0;

   // m107_35 = W*in
   wire signed [9:0] m107_35;
   assign m107_35 =10'b0;

   // m107_36 = W*in
   wire signed [9:0] m107_36;
   assign m107_36 ={ {5{neg107[5]}} , neg107[5:1] };

   // m107_37 = W*in
   wire signed [9:0] m107_37;
   assign m107_37 ={ {5{in107[5]}} , in107[5:1] };

   // m107_38 = W*in
   wire signed [9:0] m107_38;
   assign m107_38 =10'b0;

   // m107_39 = W*in
   wire signed [9:0] m107_39;
   assign m107_39 =10'b0;

   // m107_40 = W*in
   wire signed [9:0] m107_40;
   assign m107_40 =10'b0;

   // m107_41 = W*in
   wire signed [9:0] m107_41;
   assign m107_41 ={ {4{in107[5]}} , in107[5:0] };

   // m107_42 = W*in
   wire signed [9:0] m107_42;
   assign m107_42 =10'b0;

   // m107_43 = W*in
   wire signed [9:0] m107_43;
   assign m107_43 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_44 = W*in
   wire signed [9:0] m107_44;
   assign m107_44 =10'b0;

   // m107_45 = W*in
   wire signed [9:0] m107_45;
   assign m107_45 ={ {4{in107[5]}} , in107[5:0] };

   // m107_46 = W*in
   wire signed [9:0] m107_46;
   assign m107_46 =10'b0;

   // m107_47 = W*in
   wire signed [9:0] m107_47;
   assign m107_47 =10'b0;

   // m107_48 = W*in
   wire signed [9:0] m107_48;
   assign m107_48 =10'b0;

   // m107_49 = W*in
   wire signed [9:0] m107_49;
   assign m107_49 =10'b0;

   // m107_50 = W*in
   wire signed [9:0] m107_50;
   assign m107_50 =10'b0;

   // m107_51 = W*in
   wire signed [9:0] m107_51;
   assign m107_51 =10'b0;

   // m107_52 = W*in
   wire signed [9:0] m107_52;
   assign m107_52 ={ {4{in107[5]}} , in107[5:0] };

   // m107_53 = W*in
   wire signed [9:0] m107_53;
   assign m107_53 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_54 = W*in
   wire signed [9:0] m107_54;
   assign m107_54 =10'b0;

   // m107_55 = W*in
   wire signed [9:0] m107_55;
   assign m107_55 =10'b0;

   // m107_56 = W*in
   wire signed [9:0] m107_56;
   assign m107_56 =10'b0;

   // m107_57 = W*in
   wire signed [9:0] m107_57;
   assign m107_57 =10'b0;

   // m107_58 = W*in
   wire signed [9:0] m107_58;
   assign m107_58 =10'b0;

   // m107_59 = W*in
   wire signed [9:0] m107_59;
   assign m107_59 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_60 = W*in
   wire signed [9:0] m107_60;
   assign m107_60 ={ {4{in107[5]}} , in107[5:0] };

   // m107_61 = W*in
   wire signed [9:0] m107_61;
   assign m107_61 =10'b0;

   // m107_62 = W*in
   wire signed [9:0] m107_62;
   assign m107_62 ={ {4{in107[5]}} , in107[5:0] };

   // m107_63 = W*in
   wire signed [9:0] m107_63;
   assign m107_63 =10'b0;

   // m107_64 = W*in
   wire signed [9:0] m107_64;
   assign m107_64 =10'b0;

   // m107_65 = W*in
   wire signed [9:0] m107_65;
   assign m107_65 ={ {5{in107[5]}} , in107[5:1] };

   // m107_66 = W*in
   wire signed [9:0] m107_66;
   assign m107_66 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_67 = W*in
   wire signed [9:0] m107_67;
   assign m107_67 =10'b0;

   // m107_68 = W*in
   wire signed [9:0] m107_68;
   assign m107_68 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_69 = W*in
   wire signed [9:0] m107_69;
   assign m107_69 ={ {4{in107[5]}} , in107[5:0] };

   // m107_70 = W*in
   wire signed [9:0] m107_70;
   assign m107_70 =10'b0;

   // m107_71 = W*in
   wire signed [9:0] m107_71;
   assign m107_71 =10'b0;

   // m107_72 = W*in
   wire signed [9:0] m107_72;
   assign m107_72 =10'b0;

   // m107_73 = W*in
   wire signed [9:0] m107_73;
   assign m107_73 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_74 = W*in
   wire signed [9:0] m107_74;
   assign m107_74 ={ {5{neg107[5]}} , neg107[5:1] };

   // m107_75 = W*in
   wire signed [9:0] m107_75;
   assign m107_75 =10'b0;

   // m107_76 = W*in
   wire signed [9:0] m107_76;
   assign m107_76 ={ {3{in107[5]}} , in107 , {1{1'b0}} };

   // m107_77 = W*in
   wire signed [9:0] m107_77;
   assign m107_77 =10'b0;

   // m107_78 = W*in
   wire signed [9:0] m107_78;
   assign m107_78 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_79 = W*in
   wire signed [9:0] m107_79;
   assign m107_79 =10'b0;

   // m107_80 = W*in
   wire signed [9:0] m107_80;
   assign m107_80 =10'b0;

   // m107_81 = W*in
   wire signed [9:0] m107_81;
   assign m107_81 =10'b0;

   // m107_82 = W*in
   wire signed [9:0] m107_82;
   assign m107_82 ={ {4{in107[5]}} , in107[5:0] };

   // m107_83 = W*in
   wire signed [9:0] m107_83;
   assign m107_83 ={ {4{in107[5]}} , in107[5:0] };

   // m107_84 = W*in
   wire signed [9:0] m107_84;
   assign m107_84 =10'b0;

   // m107_85 = W*in
   wire signed [9:0] m107_85;
   assign m107_85 ={ {4{in107[5]}} , in107[5:0] };

   // m107_86 = W*in
   wire signed [9:0] m107_86;
   assign m107_86 =10'b0;

   // m107_87 = W*in
   wire signed [9:0] m107_87;
   assign m107_87 =10'b0;

   // m107_88 = W*in
   wire signed [9:0] m107_88;
   assign m107_88 =10'b0;

   // m107_89 = W*in
   wire signed [9:0] m107_89;
   assign m107_89 =10'b0;

   // m107_90 = W*in
   wire signed [9:0] m107_90;
   assign m107_90 =10'b0;

   // m107_91 = W*in
   wire signed [9:0] m107_91;
   assign m107_91 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_92 = W*in
   wire signed [9:0] m107_92;
   assign m107_92 =10'b0;

   // m107_93 = W*in
   wire signed [9:0] m107_93;
   assign m107_93 =10'b0;

   // m107_94 = W*in
   wire signed [9:0] m107_94;
   assign m107_94 =10'b0;

   // m107_95 = W*in
   wire signed [9:0] m107_95;
   assign m107_95 ={ {4{in107[5]}} , in107[5:0] };

   // m107_96 = W*in
   wire signed [9:0] m107_96;
   assign m107_96 =10'b0;

   // m107_97 = W*in
   wire signed [9:0] m107_97;
   assign m107_97 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_98 = W*in
   wire signed [9:0] m107_98;
   assign m107_98 ={ {4{in107[5]}} , in107[5:0] };

   // m107_99 = W*in
   wire signed [9:0] m107_99;
   assign m107_99 =10'b0;

   // m107_100 = W*in
   wire signed [9:0] m107_100;
   assign m107_100 =10'b0;

   // m107_101 = W*in
   wire signed [9:0] m107_101;
   assign m107_101 =10'b0;

   // m107_102 = W*in
   wire signed [9:0] m107_102;
   assign m107_102 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_103 = W*in
   wire signed [9:0] m107_103;
   assign m107_103 =10'b0;

   // m107_104 = W*in
   wire signed [9:0] m107_104;
   assign m107_104 =10'b0;

   // m107_105 = W*in
   wire signed [9:0] m107_105;
   assign m107_105 =10'b0;

   // m107_106 = W*in
   wire signed [9:0] m107_106;
   assign m107_106 ={ {4{neg107[5]}} , neg107[5:0] };

   // m107_107 = W*in
   wire signed [9:0] m107_107;
   assign m107_107 =10'b0;

   // m107_108 = W*in
   wire signed [9:0] m107_108;
   assign m107_108 ={ {4{in107[5]}} , in107[5:0] };

   // m107_109 = W*in
   wire signed [9:0] m107_109;
   assign m107_109 ={ {4{in107[5]}} , in107[5:0] };

   // m107_110 = W*in
   wire signed [9:0] m107_110;
   assign m107_110 =10'b0;

   // m107_111 = W*in
   wire signed [9:0] m107_111;
   assign m107_111 =10'b0;

   // m107_112 = W*in
   wire signed [9:0] m107_112;
   assign m107_112 =10'b0;

   // m107_113 = W*in
   wire signed [9:0] m107_113;
   assign m107_113 =10'b0;

   // m107_114 = W*in
   wire signed [9:0] m107_114;
   assign m107_114 ={ {5{in107[5]}} , in107[5:1] };

   // m107_115 = W*in
   wire signed [9:0] m107_115;
   assign m107_115 ={ {4{in107[5]}} , in107[5:0] };

   // m107_116 = W*in
   wire signed [9:0] m107_116;
   assign m107_116 ={ {4{in107[5]}} , in107[5:0] };

   // m107_117 = W*in
   wire signed [9:0] m107_117;
   assign m107_117 =10'b0;

   // m108_1 = W*in
   wire signed [9:0] m108_1;
   assign m108_1 =10'b0;

   // m108_2 = W*in
   wire signed [9:0] m108_2;
   assign m108_2 =10'b0;

   // m108_3 = W*in
   wire signed [9:0] m108_3;
   assign m108_3 =10'b0;

   // m108_4 = W*in
   wire signed [9:0] m108_4;
   assign m108_4 ={ {4{in108[5]}} , in108[5:0] };

   // m108_5 = W*in
   wire signed [9:0] m108_5;
   assign m108_5 =10'b0;

   // m108_6 = W*in
   wire signed [9:0] m108_6;
   assign m108_6 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_7 = W*in
   wire signed [9:0] m108_7;
   assign m108_7 =10'b0;

   // m108_8 = W*in
   wire signed [9:0] m108_8;
   assign m108_8 =10'b0;

   // m108_9 = W*in
   wire signed [9:0] m108_9;
   assign m108_9 =10'b0;

   // m108_10 = W*in
   wire signed [9:0] m108_10;
   assign m108_10 =10'b0;

   // m108_11 = W*in
   wire signed [9:0] m108_11;
   assign m108_11 =10'b0;

   // m108_12 = W*in
   wire signed [9:0] m108_12;
   assign m108_12 =10'b0;

   // m108_13 = W*in
   wire signed [9:0] m108_13;
   assign m108_13 =10'b0;

   // m108_14 = W*in
   wire signed [9:0] m108_14;
   assign m108_14 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_15 = W*in
   wire signed [9:0] m108_15;
   assign m108_15 =10'b0;

   // m108_16 = W*in
   wire signed [9:0] m108_16;
   assign m108_16 =10'b0;

   // m108_17 = W*in
   wire signed [9:0] m108_17;
   assign m108_17 ={ {5{in108[5]}} , in108[5:1] };

   // m108_18 = W*in
   wire signed [9:0] m108_18;
   assign m108_18 =10'b0;

   // m108_19 = W*in
   wire signed [9:0] m108_19;
   assign m108_19 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_20 = W*in
   wire signed [9:0] m108_20;
   assign m108_20 =10'b0;

   // m108_21 = W*in
   wire signed [9:0] m108_21;
   assign m108_21 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_22 = W*in
   wire signed [9:0] m108_22;
   assign m108_22 ={ {4{in108[5]}} , in108[5:0] };

   // m108_23 = W*in
   wire signed [9:0] m108_23;
   assign m108_23 ={ {4{in108[5]}} , in108[5:0] };

   // m108_24 = W*in
   wire signed [9:0] m108_24;
   assign m108_24 ={ {4{in108[5]}} , in108[5:0] };

   // m108_25 = W*in
   wire signed [9:0] m108_25;
   assign m108_25 =10'b0;

   // m108_26 = W*in
   wire signed [9:0] m108_26;
   assign m108_26 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_27 = W*in
   wire signed [9:0] m108_27;
   assign m108_27 ={ {4{in108[5]}} , in108[5:0] };

   // m108_28 = W*in
   wire signed [9:0] m108_28;
   assign m108_28 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_29 = W*in
   wire signed [9:0] m108_29;
   assign m108_29 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_30 = W*in
   wire signed [9:0] m108_30;
   assign m108_30 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_31 = W*in
   wire signed [9:0] m108_31;
   assign m108_31 =10'b0;

   // m108_32 = W*in
   wire signed [9:0] m108_32;
   assign m108_32 =10'b0;

   // m108_33 = W*in
   wire signed [9:0] m108_33;
   assign m108_33 =10'b0;

   // m108_34 = W*in
   wire signed [9:0] m108_34;
   assign m108_34 =10'b0;

   // m108_35 = W*in
   wire signed [9:0] m108_35;
   assign m108_35 =10'b0;

   // m108_36 = W*in
   wire signed [9:0] m108_36;
   assign m108_36 =10'b0;

   // m108_37 = W*in
   wire signed [9:0] m108_37;
   assign m108_37 =10'b0;

   // m108_38 = W*in
   wire signed [9:0] m108_38;
   assign m108_38 =10'b0;

   // m108_39 = W*in
   wire signed [9:0] m108_39;
   assign m108_39 ={ {4{in108[5]}} , in108[5:0] };

   // m108_40 = W*in
   wire signed [9:0] m108_40;
   assign m108_40 =10'b0;

   // m108_41 = W*in
   wire signed [9:0] m108_41;
   assign m108_41 =10'b0;

   // m108_42 = W*in
   wire signed [9:0] m108_42;
   assign m108_42 =10'b0;

   // m108_43 = W*in
   wire signed [9:0] m108_43;
   assign m108_43 =10'b0;

   // m108_44 = W*in
   wire signed [9:0] m108_44;
   assign m108_44 =10'b0;

   // m108_45 = W*in
   wire signed [9:0] m108_45;
   assign m108_45 =10'b0;

   // m108_46 = W*in
   wire signed [9:0] m108_46;
   assign m108_46 ={ {4{in108[5]}} , in108[5:0] };

   // m108_47 = W*in
   wire signed [9:0] m108_47;
   assign m108_47 =10'b0;

   // m108_48 = W*in
   wire signed [9:0] m108_48;
   assign m108_48 =10'b0;

   // m108_49 = W*in
   wire signed [9:0] m108_49;
   assign m108_49 =10'b0;

   // m108_50 = W*in
   wire signed [9:0] m108_50;
   assign m108_50 =10'b0;

   // m108_51 = W*in
   wire signed [9:0] m108_51;
   assign m108_51 =10'b0;

   // m108_52 = W*in
   wire signed [9:0] m108_52;
   assign m108_52 =10'b0;

   // m108_53 = W*in
   wire signed [9:0] m108_53;
   assign m108_53 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_54 = W*in
   wire signed [9:0] m108_54;
   assign m108_54 =10'b0;

   // m108_55 = W*in
   wire signed [9:0] m108_55;
   assign m108_55 =10'b0;

   // m108_56 = W*in
   wire signed [9:0] m108_56;
   assign m108_56 =10'b0;

   // m108_57 = W*in
   wire signed [9:0] m108_57;
   assign m108_57 =10'b0;

   // m108_58 = W*in
   wire signed [9:0] m108_58;
   assign m108_58 =10'b0;

   // m108_59 = W*in
   wire signed [9:0] m108_59;
   assign m108_59 =10'b0;

   // m108_60 = W*in
   wire signed [9:0] m108_60;
   assign m108_60 =10'b0;

   // m108_61 = W*in
   wire signed [9:0] m108_61;
   assign m108_61 =10'b0;

   // m108_62 = W*in
   wire signed [9:0] m108_62;
   assign m108_62 =10'b0;

   // m108_63 = W*in
   wire signed [9:0] m108_63;
   assign m108_63 =10'b0;

   // m108_64 = W*in
   wire signed [9:0] m108_64;
   assign m108_64 =10'b0;

   // m108_65 = W*in
   wire signed [9:0] m108_65;
   assign m108_65 =10'b0;

   // m108_66 = W*in
   wire signed [9:0] m108_66;
   assign m108_66 ={ {5{in108[5]}} , in108[5:1] };

   // m108_67 = W*in
   wire signed [9:0] m108_67;
   assign m108_67 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_68 = W*in
   wire signed [9:0] m108_68;
   assign m108_68 =10'b0;

   // m108_69 = W*in
   wire signed [9:0] m108_69;
   assign m108_69 =10'b0;

   // m108_70 = W*in
   wire signed [9:0] m108_70;
   assign m108_70 =10'b0;

   // m108_71 = W*in
   wire signed [9:0] m108_71;
   assign m108_71 ={ {5{in108[5]}} , in108[5:1] };

   // m108_72 = W*in
   wire signed [9:0] m108_72;
   assign m108_72 =10'b0;

   // m108_73 = W*in
   wire signed [9:0] m108_73;
   assign m108_73 =10'b0;

   // m108_74 = W*in
   wire signed [9:0] m108_74;
   assign m108_74 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_75 = W*in
   wire signed [9:0] m108_75;
   assign m108_75 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_76 = W*in
   wire signed [9:0] m108_76;
   assign m108_76 =10'b0;

   // m108_77 = W*in
   wire signed [9:0] m108_77;
   assign m108_77 =10'b0;

   // m108_78 = W*in
   wire signed [9:0] m108_78;
   assign m108_78 ={ {5{neg108[5]}} , neg108[5:1] };

   // m108_79 = W*in
   wire signed [9:0] m108_79;
   assign m108_79 =10'b0;

   // m108_80 = W*in
   wire signed [9:0] m108_80;
   assign m108_80 ={ {4{in108[5]}} , in108[5:0] };

   // m108_81 = W*in
   wire signed [9:0] m108_81;
   assign m108_81 ={ {5{in108[5]}} , in108[5:1] };

   // m108_82 = W*in
   wire signed [9:0] m108_82;
   assign m108_82 =10'b0;

   // m108_83 = W*in
   wire signed [9:0] m108_83;
   assign m108_83 ={ {4{in108[5]}} , in108[5:0] };

   // m108_84 = W*in
   wire signed [9:0] m108_84;
   assign m108_84 =10'b0;

   // m108_85 = W*in
   wire signed [9:0] m108_85;
   assign m108_85 =10'b0;

   // m108_86 = W*in
   wire signed [9:0] m108_86;
   assign m108_86 =10'b0;

   // m108_87 = W*in
   wire signed [9:0] m108_87;
   assign m108_87 =10'b0;

   // m108_88 = W*in
   wire signed [9:0] m108_88;
   assign m108_88 =10'b0;

   // m108_89 = W*in
   wire signed [9:0] m108_89;
   assign m108_89 =10'b0;

   // m108_90 = W*in
   wire signed [9:0] m108_90;
   assign m108_90 =10'b0;

   // m108_91 = W*in
   wire signed [9:0] m108_91;
   assign m108_91 =10'b0;

   // m108_92 = W*in
   wire signed [9:0] m108_92;
   assign m108_92 =10'b0;

   // m108_93 = W*in
   wire signed [9:0] m108_93;
   assign m108_93 =10'b0;

   // m108_94 = W*in
   wire signed [9:0] m108_94;
   assign m108_94 =10'b0;

   // m108_95 = W*in
   wire signed [9:0] m108_95;
   assign m108_95 =10'b0;

   // m108_96 = W*in
   wire signed [9:0] m108_96;
   assign m108_96 =10'b0;

   // m108_97 = W*in
   wire signed [9:0] m108_97;
   assign m108_97 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_98 = W*in
   wire signed [9:0] m108_98;
   assign m108_98 =10'b0;

   // m108_99 = W*in
   wire signed [9:0] m108_99;
   assign m108_99 =10'b0;

   // m108_100 = W*in
   wire signed [9:0] m108_100;
   assign m108_100 =10'b0;

   // m108_101 = W*in
   wire signed [9:0] m108_101;
   assign m108_101 =10'b0;

   // m108_102 = W*in
   wire signed [9:0] m108_102;
   assign m108_102 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_103 = W*in
   wire signed [9:0] m108_103;
   assign m108_103 =10'b0;

   // m108_104 = W*in
   wire signed [9:0] m108_104;
   assign m108_104 ={ {4{in108[5]}} , in108[5:0] };

   // m108_105 = W*in
   wire signed [9:0] m108_105;
   assign m108_105 =10'b0;

   // m108_106 = W*in
   wire signed [9:0] m108_106;
   assign m108_106 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_107 = W*in
   wire signed [9:0] m108_107;
   assign m108_107 ={ {4{in108[5]}} , in108[5:0] };

   // m108_108 = W*in
   wire signed [9:0] m108_108;
   assign m108_108 =10'b0;

   // m108_109 = W*in
   wire signed [9:0] m108_109;
   assign m108_109 ={ {5{in108[5]}} , in108[5:1] };

   // m108_110 = W*in
   wire signed [9:0] m108_110;
   assign m108_110 =10'b0;

   // m108_111 = W*in
   wire signed [9:0] m108_111;
   assign m108_111 ={ {4{neg108[5]}} , neg108[5:0] };

   // m108_112 = W*in
   wire signed [9:0] m108_112;
   assign m108_112 =10'b0;

   // m108_113 = W*in
   wire signed [9:0] m108_113;
   assign m108_113 =10'b0;

   // m108_114 = W*in
   wire signed [9:0] m108_114;
   assign m108_114 ={ {5{in108[5]}} , in108[5:1] };

   // m108_115 = W*in
   wire signed [9:0] m108_115;
   assign m108_115 =10'b0;

   // m108_116 = W*in
   wire signed [9:0] m108_116;
   assign m108_116 =10'b0;

   // m108_117 = W*in
   wire signed [9:0] m108_117;
   assign m108_117 =10'b0;

   // m109_1 = W*in
   wire signed [9:0] m109_1;
   assign m109_1 =10'b0;

   // m109_2 = W*in
   wire signed [9:0] m109_2;
   assign m109_2 =10'b0;

   // m109_3 = W*in
   wire signed [9:0] m109_3;
   assign m109_3 =10'b0;

   // m109_4 = W*in
   wire signed [9:0] m109_4;
   assign m109_4 =10'b0;

   // m109_5 = W*in
   wire signed [9:0] m109_5;
   assign m109_5 =10'b0;

   // m109_6 = W*in
   wire signed [9:0] m109_6;
   assign m109_6 =10'b0;

   // m109_7 = W*in
   wire signed [9:0] m109_7;
   assign m109_7 =10'b0;

   // m109_8 = W*in
   wire signed [9:0] m109_8;
   assign m109_8 =10'b0;

   // m109_9 = W*in
   wire signed [9:0] m109_9;
   assign m109_9 =10'b0;

   // m109_10 = W*in
   wire signed [9:0] m109_10;
   assign m109_10 =10'b0;

   // m109_11 = W*in
   wire signed [9:0] m109_11;
   assign m109_11 =10'b0;

   // m109_12 = W*in
   wire signed [9:0] m109_12;
   assign m109_12 =10'b0;

   // m109_13 = W*in
   wire signed [9:0] m109_13;
   assign m109_13 =10'b0;

   // m109_14 = W*in
   wire signed [9:0] m109_14;
   assign m109_14 =10'b0;

   // m109_15 = W*in
   wire signed [9:0] m109_15;
   assign m109_15 =10'b0;

   // m109_16 = W*in
   wire signed [9:0] m109_16;
   assign m109_16 =10'b0;

   // m109_17 = W*in
   wire signed [9:0] m109_17;
   assign m109_17 ={ {5{in109[5]}} , in109[5:1] };

   // m109_18 = W*in
   wire signed [9:0] m109_18;
   assign m109_18 =10'b0;

   // m109_19 = W*in
   wire signed [9:0] m109_19;
   assign m109_19 =10'b0;

   // m109_20 = W*in
   wire signed [9:0] m109_20;
   assign m109_20 =10'b0;

   // m109_21 = W*in
   wire signed [9:0] m109_21;
   assign m109_21 =10'b0;

   // m109_22 = W*in
   wire signed [9:0] m109_22;
   assign m109_22 =10'b0;

   // m109_23 = W*in
   wire signed [9:0] m109_23;
   assign m109_23 =10'b0;

   // m109_24 = W*in
   wire signed [9:0] m109_24;
   assign m109_24 =10'b0;

   // m109_25 = W*in
   wire signed [9:0] m109_25;
   assign m109_25 =10'b0;

   // m109_26 = W*in
   wire signed [9:0] m109_26;
   assign m109_26 =10'b0;

   // m109_27 = W*in
   wire signed [9:0] m109_27;
   assign m109_27 ={ {5{in109[5]}} , in109[5:1] };

   // m109_28 = W*in
   wire signed [9:0] m109_28;
   assign m109_28 =10'b0;

   // m109_29 = W*in
   wire signed [9:0] m109_29;
   assign m109_29 =10'b0;

   // m109_30 = W*in
   wire signed [9:0] m109_30;
   assign m109_30 ={ {5{neg109[5]}} , neg109[5:1] };

   // m109_31 = W*in
   wire signed [9:0] m109_31;
   assign m109_31 =10'b0;

   // m109_32 = W*in
   wire signed [9:0] m109_32;
   assign m109_32 =10'b0;

   // m109_33 = W*in
   wire signed [9:0] m109_33;
   assign m109_33 =10'b0;

   // m109_34 = W*in
   wire signed [9:0] m109_34;
   assign m109_34 =10'b0;

   // m109_35 = W*in
   wire signed [9:0] m109_35;
   assign m109_35 =10'b0;

   // m109_36 = W*in
   wire signed [9:0] m109_36;
   assign m109_36 ={ {5{in109[5]}} , in109[5:1] };

   // m109_37 = W*in
   wire signed [9:0] m109_37;
   assign m109_37 =10'b0;

   // m109_38 = W*in
   wire signed [9:0] m109_38;
   assign m109_38 =10'b0;

   // m109_39 = W*in
   wire signed [9:0] m109_39;
   assign m109_39 =10'b0;

   // m109_40 = W*in
   wire signed [9:0] m109_40;
   assign m109_40 =10'b0;

   // m109_41 = W*in
   wire signed [9:0] m109_41;
   assign m109_41 =10'b0;

   // m109_42 = W*in
   wire signed [9:0] m109_42;
   assign m109_42 ={ {4{neg109[5]}} , neg109[5:0] };

   // m109_43 = W*in
   wire signed [9:0] m109_43;
   assign m109_43 =10'b0;

   // m109_44 = W*in
   wire signed [9:0] m109_44;
   assign m109_44 =10'b0;

   // m109_45 = W*in
   wire signed [9:0] m109_45;
   assign m109_45 =10'b0;

   // m109_46 = W*in
   wire signed [9:0] m109_46;
   assign m109_46 =10'b0;

   // m109_47 = W*in
   wire signed [9:0] m109_47;
   assign m109_47 =10'b0;

   // m109_48 = W*in
   wire signed [9:0] m109_48;
   assign m109_48 ={ {4{in109[5]}} , in109[5:0] };

   // m109_49 = W*in
   wire signed [9:0] m109_49;
   assign m109_49 =10'b0;

   // m109_50 = W*in
   wire signed [9:0] m109_50;
   assign m109_50 ={ {4{in109[5]}} , in109[5:0] };

   // m109_51 = W*in
   wire signed [9:0] m109_51;
   assign m109_51 =10'b0;

   // m109_52 = W*in
   wire signed [9:0] m109_52;
   assign m109_52 =10'b0;

   // m109_53 = W*in
   wire signed [9:0] m109_53;
   assign m109_53 =10'b0;

   // m109_54 = W*in
   wire signed [9:0] m109_54;
   assign m109_54 =10'b0;

   // m109_55 = W*in
   wire signed [9:0] m109_55;
   assign m109_55 =10'b0;

   // m109_56 = W*in
   wire signed [9:0] m109_56;
   assign m109_56 =10'b0;

   // m109_57 = W*in
   wire signed [9:0] m109_57;
   assign m109_57 =10'b0;

   // m109_58 = W*in
   wire signed [9:0] m109_58;
   assign m109_58 =10'b0;

   // m109_59 = W*in
   wire signed [9:0] m109_59;
   assign m109_59 =10'b0;

   // m109_60 = W*in
   wire signed [9:0] m109_60;
   assign m109_60 =10'b0;

   // m109_61 = W*in
   wire signed [9:0] m109_61;
   assign m109_61 =10'b0;

   // m109_62 = W*in
   wire signed [9:0] m109_62;
   assign m109_62 =10'b0;

   // m109_63 = W*in
   wire signed [9:0] m109_63;
   assign m109_63 =10'b0;

   // m109_64 = W*in
   wire signed [9:0] m109_64;
   assign m109_64 ={ {5{neg109[5]}} , neg109[5:1] };

   // m109_65 = W*in
   wire signed [9:0] m109_65;
   assign m109_65 =10'b0;

   // m109_66 = W*in
   wire signed [9:0] m109_66;
   assign m109_66 =10'b0;

   // m109_67 = W*in
   wire signed [9:0] m109_67;
   assign m109_67 =10'b0;

   // m109_68 = W*in
   wire signed [9:0] m109_68;
   assign m109_68 =10'b0;

   // m109_69 = W*in
   wire signed [9:0] m109_69;
   assign m109_69 =10'b0;

   // m109_70 = W*in
   wire signed [9:0] m109_70;
   assign m109_70 =10'b0;

   // m109_71 = W*in
   wire signed [9:0] m109_71;
   assign m109_71 ={ {5{in109[5]}} , in109[5:1] };

   // m109_72 = W*in
   wire signed [9:0] m109_72;
   assign m109_72 =10'b0;

   // m109_73 = W*in
   wire signed [9:0] m109_73;
   assign m109_73 ={ {4{in109[5]}} , in109[5:0] };

   // m109_74 = W*in
   wire signed [9:0] m109_74;
   assign m109_74 =10'b0;

   // m109_75 = W*in
   wire signed [9:0] m109_75;
   assign m109_75 ={ {5{neg109[5]}} , neg109[5:1] };

   // m109_76 = W*in
   wire signed [9:0] m109_76;
   assign m109_76 =10'b0;

   // m109_77 = W*in
   wire signed [9:0] m109_77;
   assign m109_77 =10'b0;

   // m109_78 = W*in
   wire signed [9:0] m109_78;
   assign m109_78 =10'b0;

   // m109_79 = W*in
   wire signed [9:0] m109_79;
   assign m109_79 =10'b0;

   // m109_80 = W*in
   wire signed [9:0] m109_80;
   assign m109_80 =10'b0;

   // m109_81 = W*in
   wire signed [9:0] m109_81;
   assign m109_81 ={ {5{neg109[5]}} , neg109[5:1] };

   // m109_82 = W*in
   wire signed [9:0] m109_82;
   assign m109_82 =10'b0;

   // m109_83 = W*in
   wire signed [9:0] m109_83;
   assign m109_83 =10'b0;

   // m109_84 = W*in
   wire signed [9:0] m109_84;
   assign m109_84 =10'b0;

   // m109_85 = W*in
   wire signed [9:0] m109_85;
   assign m109_85 =10'b0;

   // m109_86 = W*in
   wire signed [9:0] m109_86;
   assign m109_86 =10'b0;

   // m109_87 = W*in
   wire signed [9:0] m109_87;
   assign m109_87 =10'b0;

   // m109_88 = W*in
   wire signed [9:0] m109_88;
   assign m109_88 =10'b0;

   // m109_89 = W*in
   wire signed [9:0] m109_89;
   assign m109_89 =10'b0;

   // m109_90 = W*in
   wire signed [9:0] m109_90;
   assign m109_90 =10'b0;

   // m109_91 = W*in
   wire signed [9:0] m109_91;
   assign m109_91 =10'b0;

   // m109_92 = W*in
   wire signed [9:0] m109_92;
   assign m109_92 =10'b0;

   // m109_93 = W*in
   wire signed [9:0] m109_93;
   assign m109_93 =10'b0;

   // m109_94 = W*in
   wire signed [9:0] m109_94;
   assign m109_94 =10'b0;

   // m109_95 = W*in
   wire signed [9:0] m109_95;
   assign m109_95 =10'b0;

   // m109_96 = W*in
   wire signed [9:0] m109_96;
   assign m109_96 =10'b0;

   // m109_97 = W*in
   wire signed [9:0] m109_97;
   assign m109_97 =10'b0;

   // m109_98 = W*in
   wire signed [9:0] m109_98;
   assign m109_98 =10'b0;

   // m109_99 = W*in
   wire signed [9:0] m109_99;
   assign m109_99 =10'b0;

   // m109_100 = W*in
   wire signed [9:0] m109_100;
   assign m109_100 =10'b0;

   // m109_101 = W*in
   wire signed [9:0] m109_101;
   assign m109_101 =10'b0;

   // m109_102 = W*in
   wire signed [9:0] m109_102;
   assign m109_102 =10'b0;

   // m109_103 = W*in
   wire signed [9:0] m109_103;
   assign m109_103 =10'b0;

   // m109_104 = W*in
   wire signed [9:0] m109_104;
   assign m109_104 =10'b0;

   // m109_105 = W*in
   wire signed [9:0] m109_105;
   assign m109_105 =10'b0;

   // m109_106 = W*in
   wire signed [9:0] m109_106;
   assign m109_106 =10'b0;

   // m109_107 = W*in
   wire signed [9:0] m109_107;
   assign m109_107 =10'b0;

   // m109_108 = W*in
   wire signed [9:0] m109_108;
   assign m109_108 =10'b0;

   // m109_109 = W*in
   wire signed [9:0] m109_109;
   assign m109_109 =10'b0;

   // m109_110 = W*in
   wire signed [9:0] m109_110;
   assign m109_110 =10'b0;

   // m109_111 = W*in
   wire signed [9:0] m109_111;
   assign m109_111 =10'b0;

   // m109_112 = W*in
   wire signed [9:0] m109_112;
   assign m109_112 =10'b0;

   // m109_113 = W*in
   wire signed [9:0] m109_113;
   assign m109_113 =10'b0;

   // m109_114 = W*in
   wire signed [9:0] m109_114;
   assign m109_114 =10'b0;

   // m109_115 = W*in
   wire signed [9:0] m109_115;
   assign m109_115 =10'b0;

   // m109_116 = W*in
   wire signed [9:0] m109_116;
   assign m109_116 =10'b0;

   // m109_117 = W*in
   wire signed [9:0] m109_117;
   assign m109_117 ={ {5{in109[5]}} , in109[5:1] };

   // m110_1 = W*in
   wire signed [9:0] m110_1;
   assign m110_1 =10'b0;

   // m110_2 = W*in
   wire signed [9:0] m110_2;
   assign m110_2 =10'b0;

   // m110_3 = W*in
   wire signed [9:0] m110_3;
   assign m110_3 =10'b0;

   // m110_4 = W*in
   wire signed [9:0] m110_4;
   assign m110_4 =10'b0;

   // m110_5 = W*in
   wire signed [9:0] m110_5;
   assign m110_5 =10'b0;

   // m110_6 = W*in
   wire signed [9:0] m110_6;
   assign m110_6 =10'b0;

   // m110_7 = W*in
   wire signed [9:0] m110_7;
   assign m110_7 =10'b0;

   // m110_8 = W*in
   wire signed [9:0] m110_8;
   assign m110_8 =10'b0;

   // m110_9 = W*in
   wire signed [9:0] m110_9;
   assign m110_9 =10'b0;

   // m110_10 = W*in
   wire signed [9:0] m110_10;
   assign m110_10 =10'b0;

   // m110_11 = W*in
   wire signed [9:0] m110_11;
   assign m110_11 =10'b0;

   // m110_12 = W*in
   wire signed [9:0] m110_12;
   assign m110_12 =10'b0;

   // m110_13 = W*in
   wire signed [9:0] m110_13;
   assign m110_13 =10'b0;

   // m110_14 = W*in
   wire signed [9:0] m110_14;
   assign m110_14 =10'b0;

   // m110_15 = W*in
   wire signed [9:0] m110_15;
   assign m110_15 =10'b0;

   // m110_16 = W*in
   wire signed [9:0] m110_16;
   assign m110_16 =10'b0;

   // m110_17 = W*in
   wire signed [9:0] m110_17;
   assign m110_17 ={ {5{neg110[5]}} , neg110[5:1] };

   // m110_18 = W*in
   wire signed [9:0] m110_18;
   assign m110_18 =10'b0;

   // m110_19 = W*in
   wire signed [9:0] m110_19;
   assign m110_19 =10'b0;

   // m110_20 = W*in
   wire signed [9:0] m110_20;
   assign m110_20 =10'b0;

   // m110_21 = W*in
   wire signed [9:0] m110_21;
   assign m110_21 ={ {5{in110[5]}} , in110[5:1] };

   // m110_22 = W*in
   wire signed [9:0] m110_22;
   assign m110_22 =10'b0;

   // m110_23 = W*in
   wire signed [9:0] m110_23;
   assign m110_23 =10'b0;

   // m110_24 = W*in
   wire signed [9:0] m110_24;
   assign m110_24 =10'b0;

   // m110_25 = W*in
   wire signed [9:0] m110_25;
   assign m110_25 =10'b0;

   // m110_26 = W*in
   wire signed [9:0] m110_26;
   assign m110_26 =10'b0;

   // m110_27 = W*in
   wire signed [9:0] m110_27;
   assign m110_27 =10'b0;

   // m110_28 = W*in
   wire signed [9:0] m110_28;
   assign m110_28 =10'b0;

   // m110_29 = W*in
   wire signed [9:0] m110_29;
   assign m110_29 =10'b0;

   // m110_30 = W*in
   wire signed [9:0] m110_30;
   assign m110_30 =10'b0;

   // m110_31 = W*in
   wire signed [9:0] m110_31;
   assign m110_31 =10'b0;

   // m110_32 = W*in
   wire signed [9:0] m110_32;
   assign m110_32 =10'b0;

   // m110_33 = W*in
   wire signed [9:0] m110_33;
   assign m110_33 =10'b0;

   // m110_34 = W*in
   wire signed [9:0] m110_34;
   assign m110_34 =10'b0;

   // m110_35 = W*in
   wire signed [9:0] m110_35;
   assign m110_35 ={ {5{in110[5]}} , in110[5:1] };

   // m110_36 = W*in
   wire signed [9:0] m110_36;
   assign m110_36 =10'b0;

   // m110_37 = W*in
   wire signed [9:0] m110_37;
   assign m110_37 =10'b0;

   // m110_38 = W*in
   wire signed [9:0] m110_38;
   assign m110_38 =10'b0;

   // m110_39 = W*in
   wire signed [9:0] m110_39;
   assign m110_39 =10'b0;

   // m110_40 = W*in
   wire signed [9:0] m110_40;
   assign m110_40 =10'b0;

   // m110_41 = W*in
   wire signed [9:0] m110_41;
   assign m110_41 =10'b0;

   // m110_42 = W*in
   wire signed [9:0] m110_42;
   assign m110_42 =10'b0;

   // m110_43 = W*in
   wire signed [9:0] m110_43;
   assign m110_43 =10'b0;

   // m110_44 = W*in
   wire signed [9:0] m110_44;
   assign m110_44 =10'b0;

   // m110_45 = W*in
   wire signed [9:0] m110_45;
   assign m110_45 =10'b0;

   // m110_46 = W*in
   wire signed [9:0] m110_46;
   assign m110_46 =10'b0;

   // m110_47 = W*in
   wire signed [9:0] m110_47;
   assign m110_47 =10'b0;

   // m110_48 = W*in
   wire signed [9:0] m110_48;
   assign m110_48 =10'b0;

   // m110_49 = W*in
   wire signed [9:0] m110_49;
   assign m110_49 =10'b0;

   // m110_50 = W*in
   wire signed [9:0] m110_50;
   assign m110_50 =10'b0;

   // m110_51 = W*in
   wire signed [9:0] m110_51;
   assign m110_51 =10'b0;

   // m110_52 = W*in
   wire signed [9:0] m110_52;
   assign m110_52 =10'b0;

   // m110_53 = W*in
   wire signed [9:0] m110_53;
   assign m110_53 =10'b0;

   // m110_54 = W*in
   wire signed [9:0] m110_54;
   assign m110_54 =10'b0;

   // m110_55 = W*in
   wire signed [9:0] m110_55;
   assign m110_55 =10'b0;

   // m110_56 = W*in
   wire signed [9:0] m110_56;
   assign m110_56 =10'b0;

   // m110_57 = W*in
   wire signed [9:0] m110_57;
   assign m110_57 =10'b0;

   // m110_58 = W*in
   wire signed [9:0] m110_58;
   assign m110_58 =10'b0;

   // m110_59 = W*in
   wire signed [9:0] m110_59;
   assign m110_59 =10'b0;

   // m110_60 = W*in
   wire signed [9:0] m110_60;
   assign m110_60 =10'b0;

   // m110_61 = W*in
   wire signed [9:0] m110_61;
   assign m110_61 =10'b0;

   // m110_62 = W*in
   wire signed [9:0] m110_62;
   assign m110_62 =10'b0;

   // m110_63 = W*in
   wire signed [9:0] m110_63;
   assign m110_63 =10'b0;

   // m110_64 = W*in
   wire signed [9:0] m110_64;
   assign m110_64 =10'b0;

   // m110_65 = W*in
   wire signed [9:0] m110_65;
   assign m110_65 =10'b0;

   // m110_66 = W*in
   wire signed [9:0] m110_66;
   assign m110_66 =10'b0;

   // m110_67 = W*in
   wire signed [9:0] m110_67;
   assign m110_67 =10'b0;

   // m110_68 = W*in
   wire signed [9:0] m110_68;
   assign m110_68 =10'b0;

   // m110_69 = W*in
   wire signed [9:0] m110_69;
   assign m110_69 ={ {5{in110[5]}} , in110[5:1] };

   // m110_70 = W*in
   wire signed [9:0] m110_70;
   assign m110_70 =10'b0;

   // m110_71 = W*in
   wire signed [9:0] m110_71;
   assign m110_71 =10'b0;

   // m110_72 = W*in
   wire signed [9:0] m110_72;
   assign m110_72 =10'b0;

   // m110_73 = W*in
   wire signed [9:0] m110_73;
   assign m110_73 =10'b0;

   // m110_74 = W*in
   wire signed [9:0] m110_74;
   assign m110_74 =10'b0;

   // m110_75 = W*in
   wire signed [9:0] m110_75;
   assign m110_75 =10'b0;

   // m110_76 = W*in
   wire signed [9:0] m110_76;
   assign m110_76 =10'b0;

   // m110_77 = W*in
   wire signed [9:0] m110_77;
   assign m110_77 =10'b0;

   // m110_78 = W*in
   wire signed [9:0] m110_78;
   assign m110_78 =10'b0;

   // m110_79 = W*in
   wire signed [9:0] m110_79;
   assign m110_79 =10'b0;

   // m110_80 = W*in
   wire signed [9:0] m110_80;
   assign m110_80 =10'b0;

   // m110_81 = W*in
   wire signed [9:0] m110_81;
   assign m110_81 =10'b0;

   // m110_82 = W*in
   wire signed [9:0] m110_82;
   assign m110_82 ={ {5{in110[5]}} , in110[5:1] };

   // m110_83 = W*in
   wire signed [9:0] m110_83;
   assign m110_83 =10'b0;

   // m110_84 = W*in
   wire signed [9:0] m110_84;
   assign m110_84 =10'b0;

   // m110_85 = W*in
   wire signed [9:0] m110_85;
   assign m110_85 =10'b0;

   // m110_86 = W*in
   wire signed [9:0] m110_86;
   assign m110_86 =10'b0;

   // m110_87 = W*in
   wire signed [9:0] m110_87;
   assign m110_87 =10'b0;

   // m110_88 = W*in
   wire signed [9:0] m110_88;
   assign m110_88 =10'b0;

   // m110_89 = W*in
   wire signed [9:0] m110_89;
   assign m110_89 =10'b0;

   // m110_90 = W*in
   wire signed [9:0] m110_90;
   assign m110_90 =10'b0;

   // m110_91 = W*in
   wire signed [9:0] m110_91;
   assign m110_91 =10'b0;

   // m110_92 = W*in
   wire signed [9:0] m110_92;
   assign m110_92 =10'b0;

   // m110_93 = W*in
   wire signed [9:0] m110_93;
   assign m110_93 =10'b0;

   // m110_94 = W*in
   wire signed [9:0] m110_94;
   assign m110_94 =10'b0;

   // m110_95 = W*in
   wire signed [9:0] m110_95;
   assign m110_95 =10'b0;

   // m110_96 = W*in
   wire signed [9:0] m110_96;
   assign m110_96 =10'b0;

   // m110_97 = W*in
   wire signed [9:0] m110_97;
   assign m110_97 =10'b0;

   // m110_98 = W*in
   wire signed [9:0] m110_98;
   assign m110_98 =10'b0;

   // m110_99 = W*in
   wire signed [9:0] m110_99;
   assign m110_99 ={ {4{in110[5]}} , in110[5:0] };

   // m110_100 = W*in
   wire signed [9:0] m110_100;
   assign m110_100 =10'b0;

   // m110_101 = W*in
   wire signed [9:0] m110_101;
   assign m110_101 =10'b0;

   // m110_102 = W*in
   wire signed [9:0] m110_102;
   assign m110_102 =10'b0;

   // m110_103 = W*in
   wire signed [9:0] m110_103;
   assign m110_103 =10'b0;

   // m110_104 = W*in
   wire signed [9:0] m110_104;
   assign m110_104 =10'b0;

   // m110_105 = W*in
   wire signed [9:0] m110_105;
   assign m110_105 =10'b0;

   // m110_106 = W*in
   wire signed [9:0] m110_106;
   assign m110_106 =10'b0;

   // m110_107 = W*in
   wire signed [9:0] m110_107;
   assign m110_107 =10'b0;

   // m110_108 = W*in
   wire signed [9:0] m110_108;
   assign m110_108 ={ {5{in110[5]}} , in110[5:1] };

   // m110_109 = W*in
   wire signed [9:0] m110_109;
   assign m110_109 =10'b0;

   // m110_110 = W*in
   wire signed [9:0] m110_110;
   assign m110_110 =10'b0;

   // m110_111 = W*in
   wire signed [9:0] m110_111;
   assign m110_111 =10'b0;

   // m110_112 = W*in
   wire signed [9:0] m110_112;
   assign m110_112 =10'b0;

   // m110_113 = W*in
   wire signed [9:0] m110_113;
   assign m110_113 =10'b0;

   // m110_114 = W*in
   wire signed [9:0] m110_114;
   assign m110_114 =10'b0;

   // m110_115 = W*in
   wire signed [9:0] m110_115;
   assign m110_115 =10'b0;

   // m110_116 = W*in
   wire signed [9:0] m110_116;
   assign m110_116 =10'b0;

   // m110_117 = W*in
   wire signed [9:0] m110_117;
   assign m110_117 =10'b0;

   // m111_1 = W*in
   wire signed [9:0] m111_1;
   assign m111_1 =10'b0;

   // m111_2 = W*in
   wire signed [9:0] m111_2;
   assign m111_2 =10'b0;

   // m111_3 = W*in
   wire signed [9:0] m111_3;
   assign m111_3 =10'b0;

   // m111_4 = W*in
   wire signed [9:0] m111_4;
   assign m111_4 ={ {4{in111[5]}} , in111[5:0] };

   // m111_5 = W*in
   wire signed [9:0] m111_5;
   assign m111_5 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_6 = W*in
   wire signed [9:0] m111_6;
   assign m111_6 =10'b0;

   // m111_7 = W*in
   wire signed [9:0] m111_7;
   assign m111_7 =10'b0;

   // m111_8 = W*in
   wire signed [9:0] m111_8;
   assign m111_8 =10'b0;

   // m111_9 = W*in
   wire signed [9:0] m111_9;
   assign m111_9 =10'b0;

   // m111_10 = W*in
   wire signed [9:0] m111_10;
   assign m111_10 =10'b0;

   // m111_11 = W*in
   wire signed [9:0] m111_11;
   assign m111_11 =10'b0;

   // m111_12 = W*in
   wire signed [9:0] m111_12;
   assign m111_12 =10'b0;

   // m111_13 = W*in
   wire signed [9:0] m111_13;
   assign m111_13 =10'b0;

   // m111_14 = W*in
   wire signed [9:0] m111_14;
   assign m111_14 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_15 = W*in
   wire signed [9:0] m111_15;
   assign m111_15 =10'b0;

   // m111_16 = W*in
   wire signed [9:0] m111_16;
   assign m111_16 =10'b0;

   // m111_17 = W*in
   wire signed [9:0] m111_17;
   assign m111_17 ={ {4{in111[5]}} , in111[5:0] };

   // m111_18 = W*in
   wire signed [9:0] m111_18;
   assign m111_18 =10'b0;

   // m111_19 = W*in
   wire signed [9:0] m111_19;
   assign m111_19 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_20 = W*in
   wire signed [9:0] m111_20;
   assign m111_20 ={ {4{in111[5]}} , in111[5:0] };

   // m111_21 = W*in
   wire signed [9:0] m111_21;
   assign m111_21 ={ {5{neg111[5]}} , neg111[5:1] };

   // m111_22 = W*in
   wire signed [9:0] m111_22;
   assign m111_22 ={ {5{in111[5]}} , in111[5:1] };

   // m111_23 = W*in
   wire signed [9:0] m111_23;
   assign m111_23 =10'b0;

   // m111_24 = W*in
   wire signed [9:0] m111_24;
   assign m111_24 =10'b0;

   // m111_25 = W*in
   wire signed [9:0] m111_25;
   assign m111_25 =10'b0;

   // m111_26 = W*in
   wire signed [9:0] m111_26;
   assign m111_26 ={ {5{neg111[5]}} , neg111[5:1] };

   // m111_27 = W*in
   wire signed [9:0] m111_27;
   assign m111_27 =10'b0;

   // m111_28 = W*in
   wire signed [9:0] m111_28;
   assign m111_28 ={ {5{neg111[5]}} , neg111[5:1] };

   // m111_29 = W*in
   wire signed [9:0] m111_29;
   assign m111_29 ={ {5{neg111[5]}} , neg111[5:1] };

   // m111_30 = W*in
   wire signed [9:0] m111_30;
   assign m111_30 =10'b0;

   // m111_31 = W*in
   wire signed [9:0] m111_31;
   assign m111_31 =10'b0;

   // m111_32 = W*in
   wire signed [9:0] m111_32;
   assign m111_32 =10'b0;

   // m111_33 = W*in
   wire signed [9:0] m111_33;
   assign m111_33 =10'b0;

   // m111_34 = W*in
   wire signed [9:0] m111_34;
   assign m111_34 =10'b0;

   // m111_35 = W*in
   wire signed [9:0] m111_35;
   assign m111_35 ={ {5{in111[5]}} , in111[5:1] };

   // m111_36 = W*in
   wire signed [9:0] m111_36;
   assign m111_36 =10'b0;

   // m111_37 = W*in
   wire signed [9:0] m111_37;
   assign m111_37 =10'b0;

   // m111_38 = W*in
   wire signed [9:0] m111_38;
   assign m111_38 =10'b0;

   // m111_39 = W*in
   wire signed [9:0] m111_39;
   assign m111_39 =10'b0;

   // m111_40 = W*in
   wire signed [9:0] m111_40;
   assign m111_40 =10'b0;

   // m111_41 = W*in
   wire signed [9:0] m111_41;
   assign m111_41 =10'b0;

   // m111_42 = W*in
   wire signed [9:0] m111_42;
   assign m111_42 =10'b0;

   // m111_43 = W*in
   wire signed [9:0] m111_43;
   assign m111_43 =10'b0;

   // m111_44 = W*in
   wire signed [9:0] m111_44;
   assign m111_44 =10'b0;

   // m111_45 = W*in
   wire signed [9:0] m111_45;
   assign m111_45 =10'b0;

   // m111_46 = W*in
   wire signed [9:0] m111_46;
   assign m111_46 =10'b0;

   // m111_47 = W*in
   wire signed [9:0] m111_47;
   assign m111_47 =10'b0;

   // m111_48 = W*in
   wire signed [9:0] m111_48;
   assign m111_48 =10'b0;

   // m111_49 = W*in
   wire signed [9:0] m111_49;
   assign m111_49 =10'b0;

   // m111_50 = W*in
   wire signed [9:0] m111_50;
   assign m111_50 =10'b0;

   // m111_51 = W*in
   wire signed [9:0] m111_51;
   assign m111_51 =10'b0;

   // m111_52 = W*in
   wire signed [9:0] m111_52;
   assign m111_52 =10'b0;

   // m111_53 = W*in
   wire signed [9:0] m111_53;
   assign m111_53 =10'b0;

   // m111_54 = W*in
   wire signed [9:0] m111_54;
   assign m111_54 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_55 = W*in
   wire signed [9:0] m111_55;
   assign m111_55 =10'b0;

   // m111_56 = W*in
   wire signed [9:0] m111_56;
   assign m111_56 =10'b0;

   // m111_57 = W*in
   wire signed [9:0] m111_57;
   assign m111_57 =10'b0;

   // m111_58 = W*in
   wire signed [9:0] m111_58;
   assign m111_58 =10'b0;

   // m111_59 = W*in
   wire signed [9:0] m111_59;
   assign m111_59 =10'b0;

   // m111_60 = W*in
   wire signed [9:0] m111_60;
   assign m111_60 =10'b0;

   // m111_61 = W*in
   wire signed [9:0] m111_61;
   assign m111_61 =10'b0;

   // m111_62 = W*in
   wire signed [9:0] m111_62;
   assign m111_62 =10'b0;

   // m111_63 = W*in
   wire signed [9:0] m111_63;
   assign m111_63 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_64 = W*in
   wire signed [9:0] m111_64;
   assign m111_64 ={ {4{in111[5]}} , in111[5:0] };

   // m111_65 = W*in
   wire signed [9:0] m111_65;
   assign m111_65 =10'b0;

   // m111_66 = W*in
   wire signed [9:0] m111_66;
   assign m111_66 =10'b0;

   // m111_67 = W*in
   wire signed [9:0] m111_67;
   assign m111_67 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_68 = W*in
   wire signed [9:0] m111_68;
   assign m111_68 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_69 = W*in
   wire signed [9:0] m111_69;
   assign m111_69 =10'b0;

   // m111_70 = W*in
   wire signed [9:0] m111_70;
   assign m111_70 =10'b0;

   // m111_71 = W*in
   wire signed [9:0] m111_71;
   assign m111_71 =10'b0;

   // m111_72 = W*in
   wire signed [9:0] m111_72;
   assign m111_72 ={ {5{in111[5]}} , in111[5:1] };

   // m111_73 = W*in
   wire signed [9:0] m111_73;
   assign m111_73 =10'b0;

   // m111_74 = W*in
   wire signed [9:0] m111_74;
   assign m111_74 ={ {5{in111[5]}} , in111[5:1] };

   // m111_75 = W*in
   wire signed [9:0] m111_75;
   assign m111_75 ={ {5{in111[5]}} , in111[5:1] };

   // m111_76 = W*in
   wire signed [9:0] m111_76;
   assign m111_76 =10'b0;

   // m111_77 = W*in
   wire signed [9:0] m111_77;
   assign m111_77 ={ {4{in111[5]}} , in111[5:0] };

   // m111_78 = W*in
   wire signed [9:0] m111_78;
   assign m111_78 ={ {5{neg111[5]}} , neg111[5:1] };

   // m111_79 = W*in
   wire signed [9:0] m111_79;
   assign m111_79 =10'b0;

   // m111_80 = W*in
   wire signed [9:0] m111_80;
   assign m111_80 =10'b0;

   // m111_81 = W*in
   wire signed [9:0] m111_81;
   assign m111_81 ={ {4{in111[5]}} , in111[5:0] };

   // m111_82 = W*in
   wire signed [9:0] m111_82;
   assign m111_82 =10'b0;

   // m111_83 = W*in
   wire signed [9:0] m111_83;
   assign m111_83 ={ {5{in111[5]}} , in111[5:1] };

   // m111_84 = W*in
   wire signed [9:0] m111_84;
   assign m111_84 =10'b0;

   // m111_85 = W*in
   wire signed [9:0] m111_85;
   assign m111_85 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_86 = W*in
   wire signed [9:0] m111_86;
   assign m111_86 =10'b0;

   // m111_87 = W*in
   wire signed [9:0] m111_87;
   assign m111_87 =10'b0;

   // m111_88 = W*in
   wire signed [9:0] m111_88;
   assign m111_88 =10'b0;

   // m111_89 = W*in
   wire signed [9:0] m111_89;
   assign m111_89 =10'b0;

   // m111_90 = W*in
   wire signed [9:0] m111_90;
   assign m111_90 =10'b0;

   // m111_91 = W*in
   wire signed [9:0] m111_91;
   assign m111_91 =10'b0;

   // m111_92 = W*in
   wire signed [9:0] m111_92;
   assign m111_92 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_93 = W*in
   wire signed [9:0] m111_93;
   assign m111_93 ={ {4{neg111[5]}} , neg111[5:0] };

   // m111_94 = W*in
   wire signed [9:0] m111_94;
   assign m111_94 =10'b0;

   // m111_95 = W*in
   wire signed [9:0] m111_95;
   assign m111_95 =10'b0;

   // m111_96 = W*in
   wire signed [9:0] m111_96;
   assign m111_96 =10'b0;

   // m111_97 = W*in
   wire signed [9:0] m111_97;
   assign m111_97 =10'b0;

   // m111_98 = W*in
   wire signed [9:0] m111_98;
   assign m111_98 =10'b0;

   // m111_99 = W*in
   wire signed [9:0] m111_99;
   assign m111_99 =10'b0;

   // m111_100 = W*in
   wire signed [9:0] m111_100;
   assign m111_100 =10'b0;

   // m111_101 = W*in
   wire signed [9:0] m111_101;
   assign m111_101 =10'b0;

   // m111_102 = W*in
   wire signed [9:0] m111_102;
   assign m111_102 =10'b0;

   // m111_103 = W*in
   wire signed [9:0] m111_103;
   assign m111_103 =10'b0;

   // m111_104 = W*in
   wire signed [9:0] m111_104;
   assign m111_104 =10'b0;

   // m111_105 = W*in
   wire signed [9:0] m111_105;
   assign m111_105 =10'b0;

   // m111_106 = W*in
   wire signed [9:0] m111_106;
   assign m111_106 =10'b0;

   // m111_107 = W*in
   wire signed [9:0] m111_107;
   assign m111_107 ={ {4{in111[5]}} , in111[5:0] };

   // m111_108 = W*in
   wire signed [9:0] m111_108;
   assign m111_108 ={ {5{in111[5]}} , in111[5:1] };

   // m111_109 = W*in
   wire signed [9:0] m111_109;
   assign m111_109 ={ {5{in111[5]}} , in111[5:1] };

   // m111_110 = W*in
   wire signed [9:0] m111_110;
   assign m111_110 =10'b0;

   // m111_111 = W*in
   wire signed [9:0] m111_111;
   assign m111_111 =10'b0;

   // m111_112 = W*in
   wire signed [9:0] m111_112;
   assign m111_112 =10'b0;

   // m111_113 = W*in
   wire signed [9:0] m111_113;
   assign m111_113 =10'b0;

   // m111_114 = W*in
   wire signed [9:0] m111_114;
   assign m111_114 ={ {5{in111[5]}} , in111[5:1] };

   // m111_115 = W*in
   wire signed [9:0] m111_115;
   assign m111_115 =10'b0;

   // m111_116 = W*in
   wire signed [9:0] m111_116;
   assign m111_116 =10'b0;

   // m111_117 = W*in
   wire signed [9:0] m111_117;
   assign m111_117 =10'b0;

   // m112_1 = W*in
   wire signed [9:0] m112_1;
   assign m112_1 =10'b0;

   // m112_2 = W*in
   wire signed [9:0] m112_2;
   assign m112_2 =10'b0;

   // m112_3 = W*in
   wire signed [9:0] m112_3;
   assign m112_3 =10'b0;

   // m112_4 = W*in
   wire signed [9:0] m112_4;
   assign m112_4 ={ {4{in112[5]}} , in112[5:0] };

   // m112_5 = W*in
   wire signed [9:0] m112_5;
   assign m112_5 =10'b0;

   // m112_6 = W*in
   wire signed [9:0] m112_6;
   assign m112_6 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_7 = W*in
   wire signed [9:0] m112_7;
   assign m112_7 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_8 = W*in
   wire signed [9:0] m112_8;
   assign m112_8 =10'b0;

   // m112_9 = W*in
   wire signed [9:0] m112_9;
   assign m112_9 =10'b0;

   // m112_10 = W*in
   wire signed [9:0] m112_10;
   assign m112_10 =10'b0;

   // m112_11 = W*in
   wire signed [9:0] m112_11;
   assign m112_11 ={ {4{in112[5]}} , in112[5:0] };

   // m112_12 = W*in
   wire signed [9:0] m112_12;
   assign m112_12 =10'b0;

   // m112_13 = W*in
   wire signed [9:0] m112_13;
   assign m112_13 =10'b0;

   // m112_14 = W*in
   wire signed [9:0] m112_14;
   assign m112_14 =10'b0;

   // m112_15 = W*in
   wire signed [9:0] m112_15;
   assign m112_15 =10'b0;

   // m112_16 = W*in
   wire signed [9:0] m112_16;
   assign m112_16 ={ {4{in112[5]}} , in112[5:0] };

   // m112_17 = W*in
   wire signed [9:0] m112_17;
   assign m112_17 =10'b0;

   // m112_18 = W*in
   wire signed [9:0] m112_18;
   assign m112_18 =10'b0;

   // m112_19 = W*in
   wire signed [9:0] m112_19;
   assign m112_19 =10'b0;

   // m112_20 = W*in
   wire signed [9:0] m112_20;
   assign m112_20 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_21 = W*in
   wire signed [9:0] m112_21;
   assign m112_21 =10'b0;

   // m112_22 = W*in
   wire signed [9:0] m112_22;
   assign m112_22 =10'b0;

   // m112_23 = W*in
   wire signed [9:0] m112_23;
   assign m112_23 =10'b0;

   // m112_24 = W*in
   wire signed [9:0] m112_24;
   assign m112_24 =10'b0;

   // m112_25 = W*in
   wire signed [9:0] m112_25;
   assign m112_25 =10'b0;

   // m112_26 = W*in
   wire signed [9:0] m112_26;
   assign m112_26 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_27 = W*in
   wire signed [9:0] m112_27;
   assign m112_27 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_28 = W*in
   wire signed [9:0] m112_28;
   assign m112_28 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_29 = W*in
   wire signed [9:0] m112_29;
   assign m112_29 =10'b0;

   // m112_30 = W*in
   wire signed [9:0] m112_30;
   assign m112_30 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_31 = W*in
   wire signed [9:0] m112_31;
   assign m112_31 =10'b0;

   // m112_32 = W*in
   wire signed [9:0] m112_32;
   assign m112_32 =10'b0;

   // m112_33 = W*in
   wire signed [9:0] m112_33;
   assign m112_33 =10'b0;

   // m112_34 = W*in
   wire signed [9:0] m112_34;
   assign m112_34 =10'b0;

   // m112_35 = W*in
   wire signed [9:0] m112_35;
   assign m112_35 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_36 = W*in
   wire signed [9:0] m112_36;
   assign m112_36 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_37 = W*in
   wire signed [9:0] m112_37;
   assign m112_37 ={ {4{in112[5]}} , in112[5:0] };

   // m112_38 = W*in
   wire signed [9:0] m112_38;
   assign m112_38 =10'b0;

   // m112_39 = W*in
   wire signed [9:0] m112_39;
   assign m112_39 =10'b0;

   // m112_40 = W*in
   wire signed [9:0] m112_40;
   assign m112_40 =10'b0;

   // m112_41 = W*in
   wire signed [9:0] m112_41;
   assign m112_41 =10'b0;

   // m112_42 = W*in
   wire signed [9:0] m112_42;
   assign m112_42 =10'b0;

   // m112_43 = W*in
   wire signed [9:0] m112_43;
   assign m112_43 =10'b0;

   // m112_44 = W*in
   wire signed [9:0] m112_44;
   assign m112_44 =10'b0;

   // m112_45 = W*in
   wire signed [9:0] m112_45;
   assign m112_45 =10'b0;

   // m112_46 = W*in
   wire signed [9:0] m112_46;
   assign m112_46 =10'b0;

   // m112_47 = W*in
   wire signed [9:0] m112_47;
   assign m112_47 =10'b0;

   // m112_48 = W*in
   wire signed [9:0] m112_48;
   assign m112_48 =10'b0;

   // m112_49 = W*in
   wire signed [9:0] m112_49;
   assign m112_49 =10'b0;

   // m112_50 = W*in
   wire signed [9:0] m112_50;
   assign m112_50 =10'b0;

   // m112_51 = W*in
   wire signed [9:0] m112_51;
   assign m112_51 =10'b0;

   // m112_52 = W*in
   wire signed [9:0] m112_52;
   assign m112_52 =10'b0;

   // m112_53 = W*in
   wire signed [9:0] m112_53;
   assign m112_53 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_54 = W*in
   wire signed [9:0] m112_54;
   assign m112_54 =10'b0;

   // m112_55 = W*in
   wire signed [9:0] m112_55;
   assign m112_55 =10'b0;

   // m112_56 = W*in
   wire signed [9:0] m112_56;
   assign m112_56 =10'b0;

   // m112_57 = W*in
   wire signed [9:0] m112_57;
   assign m112_57 =10'b0;

   // m112_58 = W*in
   wire signed [9:0] m112_58;
   assign m112_58 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_59 = W*in
   wire signed [9:0] m112_59;
   assign m112_59 =10'b0;

   // m112_60 = W*in
   wire signed [9:0] m112_60;
   assign m112_60 =10'b0;

   // m112_61 = W*in
   wire signed [9:0] m112_61;
   assign m112_61 ={ {4{in112[5]}} , in112[5:0] };

   // m112_62 = W*in
   wire signed [9:0] m112_62;
   assign m112_62 ={ {4{in112[5]}} , in112[5:0] };

   // m112_63 = W*in
   wire signed [9:0] m112_63;
   assign m112_63 =10'b0;

   // m112_64 = W*in
   wire signed [9:0] m112_64;
   assign m112_64 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_65 = W*in
   wire signed [9:0] m112_65;
   assign m112_65 =10'b0;

   // m112_66 = W*in
   wire signed [9:0] m112_66;
   assign m112_66 =10'b0;

   // m112_67 = W*in
   wire signed [9:0] m112_67;
   assign m112_67 =10'b0;

   // m112_68 = W*in
   wire signed [9:0] m112_68;
   assign m112_68 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_69 = W*in
   wire signed [9:0] m112_69;
   assign m112_69 ={ {5{in112[5]}} , in112[5:1] };

   // m112_70 = W*in
   wire signed [9:0] m112_70;
   assign m112_70 =10'b0;

   // m112_71 = W*in
   wire signed [9:0] m112_71;
   assign m112_71 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_72 = W*in
   wire signed [9:0] m112_72;
   assign m112_72 =10'b0;

   // m112_73 = W*in
   wire signed [9:0] m112_73;
   assign m112_73 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_74 = W*in
   wire signed [9:0] m112_74;
   assign m112_74 =10'b0;

   // m112_75 = W*in
   wire signed [9:0] m112_75;
   assign m112_75 =10'b0;

   // m112_76 = W*in
   wire signed [9:0] m112_76;
   assign m112_76 =10'b0;

   // m112_77 = W*in
   wire signed [9:0] m112_77;
   assign m112_77 ={ {4{in112[5]}} , in112[5:0] };

   // m112_78 = W*in
   wire signed [9:0] m112_78;
   assign m112_78 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_79 = W*in
   wire signed [9:0] m112_79;
   assign m112_79 =10'b0;

   // m112_80 = W*in
   wire signed [9:0] m112_80;
   assign m112_80 =10'b0;

   // m112_81 = W*in
   wire signed [9:0] m112_81;
   assign m112_81 =10'b0;

   // m112_82 = W*in
   wire signed [9:0] m112_82;
   assign m112_82 ={ {4{in112[5]}} , in112[5:0] };

   // m112_83 = W*in
   wire signed [9:0] m112_83;
   assign m112_83 ={ {4{in112[5]}} , in112[5:0] };

   // m112_84 = W*in
   wire signed [9:0] m112_84;
   assign m112_84 =10'b0;

   // m112_85 = W*in
   wire signed [9:0] m112_85;
   assign m112_85 ={ {4{in112[5]}} , in112[5:0] };

   // m112_86 = W*in
   wire signed [9:0] m112_86;
   assign m112_86 =10'b0;

   // m112_87 = W*in
   wire signed [9:0] m112_87;
   assign m112_87 =10'b0;

   // m112_88 = W*in
   wire signed [9:0] m112_88;
   assign m112_88 =10'b0;

   // m112_89 = W*in
   wire signed [9:0] m112_89;
   assign m112_89 =10'b0;

   // m112_90 = W*in
   wire signed [9:0] m112_90;
   assign m112_90 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_91 = W*in
   wire signed [9:0] m112_91;
   assign m112_91 =10'b0;

   // m112_92 = W*in
   wire signed [9:0] m112_92;
   assign m112_92 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_93 = W*in
   wire signed [9:0] m112_93;
   assign m112_93 =10'b0;

   // m112_94 = W*in
   wire signed [9:0] m112_94;
   assign m112_94 =10'b0;

   // m112_95 = W*in
   wire signed [9:0] m112_95;
   assign m112_95 ={ {4{in112[5]}} , in112[5:0] };

   // m112_96 = W*in
   wire signed [9:0] m112_96;
   assign m112_96 =10'b0;

   // m112_97 = W*in
   wire signed [9:0] m112_97;
   assign m112_97 =10'b0;

   // m112_98 = W*in
   wire signed [9:0] m112_98;
   assign m112_98 ={ {4{in112[5]}} , in112[5:0] };

   // m112_99 = W*in
   wire signed [9:0] m112_99;
   assign m112_99 =10'b0;

   // m112_100 = W*in
   wire signed [9:0] m112_100;
   assign m112_100 =10'b0;

   // m112_101 = W*in
   wire signed [9:0] m112_101;
   assign m112_101 =10'b0;

   // m112_102 = W*in
   wire signed [9:0] m112_102;
   assign m112_102 =10'b0;

   // m112_103 = W*in
   wire signed [9:0] m112_103;
   assign m112_103 =10'b0;

   // m112_104 = W*in
   wire signed [9:0] m112_104;
   assign m112_104 =10'b0;

   // m112_105 = W*in
   wire signed [9:0] m112_105;
   assign m112_105 =10'b0;

   // m112_106 = W*in
   wire signed [9:0] m112_106;
   assign m112_106 ={ {4{neg112[5]}} , neg112[5:0] };

   // m112_107 = W*in
   wire signed [9:0] m112_107;
   assign m112_107 =10'b0;

   // m112_108 = W*in
   wire signed [9:0] m112_108;
   assign m112_108 =10'b0;

   // m112_109 = W*in
   wire signed [9:0] m112_109;
   assign m112_109 =10'b0;

   // m112_110 = W*in
   wire signed [9:0] m112_110;
   assign m112_110 =10'b0;

   // m112_111 = W*in
   wire signed [9:0] m112_111;
   assign m112_111 =10'b0;

   // m112_112 = W*in
   wire signed [9:0] m112_112;
   assign m112_112 =10'b0;

   // m112_113 = W*in
   wire signed [9:0] m112_113;
   assign m112_113 =10'b0;

   // m112_114 = W*in
   wire signed [9:0] m112_114;
   assign m112_114 ={ {5{neg112[5]}} , neg112[5:1] };

   // m112_115 = W*in
   wire signed [9:0] m112_115;
   assign m112_115 =10'b0;

   // m112_116 = W*in
   wire signed [9:0] m112_116;
   assign m112_116 =10'b0;

   // m112_117 = W*in
   wire signed [9:0] m112_117;
   assign m112_117 ={ {4{neg112[5]}} , neg112[5:0] };

   // m113_1 = W*in
   wire signed [9:0] m113_1;
   assign m113_1 ={ {4{neg113[5]}} , neg113[5:0] };

   // m113_2 = W*in
   wire signed [9:0] m113_2;
   assign m113_2 =10'b0;

   // m113_3 = W*in
   wire signed [9:0] m113_3;
   assign m113_3 =10'b0;

   // m113_4 = W*in
   wire signed [9:0] m113_4;
   assign m113_4 =10'b0;

   // m113_5 = W*in
   wire signed [9:0] m113_5;
   assign m113_5 =10'b0;

   // m113_6 = W*in
   wire signed [9:0] m113_6;
   assign m113_6 =10'b0;

   // m113_7 = W*in
   wire signed [9:0] m113_7;
   assign m113_7 =10'b0;

   // m113_8 = W*in
   wire signed [9:0] m113_8;
   assign m113_8 =10'b0;

   // m113_9 = W*in
   wire signed [9:0] m113_9;
   assign m113_9 =10'b0;

   // m113_10 = W*in
   wire signed [9:0] m113_10;
   assign m113_10 =10'b0;

   // m113_11 = W*in
   wire signed [9:0] m113_11;
   assign m113_11 =10'b0;

   // m113_12 = W*in
   wire signed [9:0] m113_12;
   assign m113_12 =10'b0;

   // m113_13 = W*in
   wire signed [9:0] m113_13;
   assign m113_13 =10'b0;

   // m113_14 = W*in
   wire signed [9:0] m113_14;
   assign m113_14 =10'b0;

   // m113_15 = W*in
   wire signed [9:0] m113_15;
   assign m113_15 =10'b0;

   // m113_16 = W*in
   wire signed [9:0] m113_16;
   assign m113_16 =10'b0;

   // m113_17 = W*in
   wire signed [9:0] m113_17;
   assign m113_17 =10'b0;

   // m113_18 = W*in
   wire signed [9:0] m113_18;
   assign m113_18 ={ {5{neg113[5]}} , neg113[5:1] };

   // m113_19 = W*in
   wire signed [9:0] m113_19;
   assign m113_19 ={ {5{neg113[5]}} , neg113[5:1] };

   // m113_20 = W*in
   wire signed [9:0] m113_20;
   assign m113_20 ={ {5{in113[5]}} , in113[5:1] };

   // m113_21 = W*in
   wire signed [9:0] m113_21;
   assign m113_21 ={ {5{in113[5]}} , in113[5:1] };

   // m113_22 = W*in
   wire signed [9:0] m113_22;
   assign m113_22 =10'b0;

   // m113_23 = W*in
   wire signed [9:0] m113_23;
   assign m113_23 ={ {4{in113[5]}} , in113[5:0] };

   // m113_24 = W*in
   wire signed [9:0] m113_24;
   assign m113_24 =10'b0;

   // m113_25 = W*in
   wire signed [9:0] m113_25;
   assign m113_25 ={ {4{neg113[5]}} , neg113[5:0] };

   // m113_26 = W*in
   wire signed [9:0] m113_26;
   assign m113_26 =10'b0;

   // m113_27 = W*in
   wire signed [9:0] m113_27;
   assign m113_27 ={ {5{in113[5]}} , in113[5:1] };

   // m113_28 = W*in
   wire signed [9:0] m113_28;
   assign m113_28 ={ {4{neg113[5]}} , neg113[5:0] };

   // m113_29 = W*in
   wire signed [9:0] m113_29;
   assign m113_29 =10'b0;

   // m113_30 = W*in
   wire signed [9:0] m113_30;
   assign m113_30 ={ {5{neg113[5]}} , neg113[5:1] };

   // m113_31 = W*in
   wire signed [9:0] m113_31;
   assign m113_31 =10'b0;

   // m113_32 = W*in
   wire signed [9:0] m113_32;
   assign m113_32 =10'b0;

   // m113_33 = W*in
   wire signed [9:0] m113_33;
   assign m113_33 =10'b0;

   // m113_34 = W*in
   wire signed [9:0] m113_34;
   assign m113_34 ={ {4{in113[5]}} , in113[5:0] };

   // m113_35 = W*in
   wire signed [9:0] m113_35;
   assign m113_35 =10'b0;

   // m113_36 = W*in
   wire signed [9:0] m113_36;
   assign m113_36 =10'b0;

   // m113_37 = W*in
   wire signed [9:0] m113_37;
   assign m113_37 =10'b0;

   // m113_38 = W*in
   wire signed [9:0] m113_38;
   assign m113_38 =10'b0;

   // m113_39 = W*in
   wire signed [9:0] m113_39;
   assign m113_39 =10'b0;

   // m113_40 = W*in
   wire signed [9:0] m113_40;
   assign m113_40 =10'b0;

   // m113_41 = W*in
   wire signed [9:0] m113_41;
   assign m113_41 =10'b0;

   // m113_42 = W*in
   wire signed [9:0] m113_42;
   assign m113_42 =10'b0;

   // m113_43 = W*in
   wire signed [9:0] m113_43;
   assign m113_43 =10'b0;

   // m113_44 = W*in
   wire signed [9:0] m113_44;
   assign m113_44 =10'b0;

   // m113_45 = W*in
   wire signed [9:0] m113_45;
   assign m113_45 =10'b0;

   // m113_46 = W*in
   wire signed [9:0] m113_46;
   assign m113_46 =10'b0;

   // m113_47 = W*in
   wire signed [9:0] m113_47;
   assign m113_47 =10'b0;

   // m113_48 = W*in
   wire signed [9:0] m113_48;
   assign m113_48 =10'b0;

   // m113_49 = W*in
   wire signed [9:0] m113_49;
   assign m113_49 =10'b0;

   // m113_50 = W*in
   wire signed [9:0] m113_50;
   assign m113_50 =10'b0;

   // m113_51 = W*in
   wire signed [9:0] m113_51;
   assign m113_51 =10'b0;

   // m113_52 = W*in
   wire signed [9:0] m113_52;
   assign m113_52 =10'b0;

   // m113_53 = W*in
   wire signed [9:0] m113_53;
   assign m113_53 =10'b0;

   // m113_54 = W*in
   wire signed [9:0] m113_54;
   assign m113_54 =10'b0;

   // m113_55 = W*in
   wire signed [9:0] m113_55;
   assign m113_55 =10'b0;

   // m113_56 = W*in
   wire signed [9:0] m113_56;
   assign m113_56 =10'b0;

   // m113_57 = W*in
   wire signed [9:0] m113_57;
   assign m113_57 =10'b0;

   // m113_58 = W*in
   wire signed [9:0] m113_58;
   assign m113_58 =10'b0;

   // m113_59 = W*in
   wire signed [9:0] m113_59;
   assign m113_59 =10'b0;

   // m113_60 = W*in
   wire signed [9:0] m113_60;
   assign m113_60 =10'b0;

   // m113_61 = W*in
   wire signed [9:0] m113_61;
   assign m113_61 =10'b0;

   // m113_62 = W*in
   wire signed [9:0] m113_62;
   assign m113_62 =10'b0;

   // m113_63 = W*in
   wire signed [9:0] m113_63;
   assign m113_63 =10'b0;

   // m113_64 = W*in
   wire signed [9:0] m113_64;
   assign m113_64 =10'b0;

   // m113_65 = W*in
   wire signed [9:0] m113_65;
   assign m113_65 =10'b0;

   // m113_66 = W*in
   wire signed [9:0] m113_66;
   assign m113_66 =10'b0;

   // m113_67 = W*in
   wire signed [9:0] m113_67;
   assign m113_67 =10'b0;

   // m113_68 = W*in
   wire signed [9:0] m113_68;
   assign m113_68 =10'b0;

   // m113_69 = W*in
   wire signed [9:0] m113_69;
   assign m113_69 ={ {5{in113[5]}} , in113[5:1] };

   // m113_70 = W*in
   wire signed [9:0] m113_70;
   assign m113_70 ={ {5{in113[5]}} , in113[5:1] };

   // m113_71 = W*in
   wire signed [9:0] m113_71;
   assign m113_71 =10'b0;

   // m113_72 = W*in
   wire signed [9:0] m113_72;
   assign m113_72 ={ {5{in113[5]}} , in113[5:1] };

   // m113_73 = W*in
   wire signed [9:0] m113_73;
   assign m113_73 =10'b0;

   // m113_74 = W*in
   wire signed [9:0] m113_74;
   assign m113_74 =10'b0;

   // m113_75 = W*in
   wire signed [9:0] m113_75;
   assign m113_75 ={ {5{neg113[5]}} , neg113[5:1] };

   // m113_76 = W*in
   wire signed [9:0] m113_76;
   assign m113_76 ={ {4{in113[5]}} , in113[5:0] };

   // m113_77 = W*in
   wire signed [9:0] m113_77;
   assign m113_77 =10'b0;

   // m113_78 = W*in
   wire signed [9:0] m113_78;
   assign m113_78 ={ {4{neg113[5]}} , neg113[5:0] };

   // m113_79 = W*in
   wire signed [9:0] m113_79;
   assign m113_79 =10'b0;

   // m113_80 = W*in
   wire signed [9:0] m113_80;
   assign m113_80 =10'b0;

   // m113_81 = W*in
   wire signed [9:0] m113_81;
   assign m113_81 =10'b0;

   // m113_82 = W*in
   wire signed [9:0] m113_82;
   assign m113_82 ={ {5{in113[5]}} , in113[5:1] };

   // m113_83 = W*in
   wire signed [9:0] m113_83;
   assign m113_83 ={ {5{neg113[5]}} , neg113[5:1] };

   // m113_84 = W*in
   wire signed [9:0] m113_84;
   assign m113_84 =10'b0;

   // m113_85 = W*in
   wire signed [9:0] m113_85;
   assign m113_85 =10'b0;

   // m113_86 = W*in
   wire signed [9:0] m113_86;
   assign m113_86 =10'b0;

   // m113_87 = W*in
   wire signed [9:0] m113_87;
   assign m113_87 =10'b0;

   // m113_88 = W*in
   wire signed [9:0] m113_88;
   assign m113_88 =10'b0;

   // m113_89 = W*in
   wire signed [9:0] m113_89;
   assign m113_89 =10'b0;

   // m113_90 = W*in
   wire signed [9:0] m113_90;
   assign m113_90 =10'b0;

   // m113_91 = W*in
   wire signed [9:0] m113_91;
   assign m113_91 =10'b0;

   // m113_92 = W*in
   wire signed [9:0] m113_92;
   assign m113_92 =10'b0;

   // m113_93 = W*in
   wire signed [9:0] m113_93;
   assign m113_93 =10'b0;

   // m113_94 = W*in
   wire signed [9:0] m113_94;
   assign m113_94 =10'b0;

   // m113_95 = W*in
   wire signed [9:0] m113_95;
   assign m113_95 =10'b0;

   // m113_96 = W*in
   wire signed [9:0] m113_96;
   assign m113_96 =10'b0;

   // m113_97 = W*in
   wire signed [9:0] m113_97;
   assign m113_97 =10'b0;

   // m113_98 = W*in
   wire signed [9:0] m113_98;
   assign m113_98 =10'b0;

   // m113_99 = W*in
   wire signed [9:0] m113_99;
   assign m113_99 ={ {4{in113[5]}} , in113[5:0] };

   // m113_100 = W*in
   wire signed [9:0] m113_100;
   assign m113_100 =10'b0;

   // m113_101 = W*in
   wire signed [9:0] m113_101;
   assign m113_101 =10'b0;

   // m113_102 = W*in
   wire signed [9:0] m113_102;
   assign m113_102 =10'b0;

   // m113_103 = W*in
   wire signed [9:0] m113_103;
   assign m113_103 =10'b0;

   // m113_104 = W*in
   wire signed [9:0] m113_104;
   assign m113_104 =10'b0;

   // m113_105 = W*in
   wire signed [9:0] m113_105;
   assign m113_105 =10'b0;

   // m113_106 = W*in
   wire signed [9:0] m113_106;
   assign m113_106 =10'b0;

   // m113_107 = W*in
   wire signed [9:0] m113_107;
   assign m113_107 =10'b0;

   // m113_108 = W*in
   wire signed [9:0] m113_108;
   assign m113_108 =10'b0;

   // m113_109 = W*in
   wire signed [9:0] m113_109;
   assign m113_109 ={ {4{in113[5]}} , in113[5:0] };

   // m113_110 = W*in
   wire signed [9:0] m113_110;
   assign m113_110 =10'b0;

   // m113_111 = W*in
   wire signed [9:0] m113_111;
   assign m113_111 =10'b0;

   // m113_112 = W*in
   wire signed [9:0] m113_112;
   assign m113_112 ={ {4{neg113[5]}} , neg113[5:0] };

   // m113_113 = W*in
   wire signed [9:0] m113_113;
   assign m113_113 =10'b0;

   // m113_114 = W*in
   wire signed [9:0] m113_114;
   assign m113_114 ={ {4{in113[5]}} , in113[5:0] };

   // m113_115 = W*in
   wire signed [9:0] m113_115;
   assign m113_115 =10'b0;

   // m113_116 = W*in
   wire signed [9:0] m113_116;
   assign m113_116 =10'b0;

   // m113_117 = W*in
   wire signed [9:0] m113_117;
   assign m113_117 =10'b0;

   // m114_1 = W*in
   wire signed [9:0] m114_1;
   assign m114_1 =10'b0;

   // m114_2 = W*in
   wire signed [9:0] m114_2;
   assign m114_2 =10'b0;

   // m114_3 = W*in
   wire signed [9:0] m114_3;
   assign m114_3 =10'b0;

   // m114_4 = W*in
   wire signed [9:0] m114_4;
   assign m114_4 =10'b0;

   // m114_5 = W*in
   wire signed [9:0] m114_5;
   assign m114_5 =10'b0;

   // m114_6 = W*in
   wire signed [9:0] m114_6;
   assign m114_6 =10'b0;

   // m114_7 = W*in
   wire signed [9:0] m114_7;
   assign m114_7 =10'b0;

   // m114_8 = W*in
   wire signed [9:0] m114_8;
   assign m114_8 =10'b0;

   // m114_9 = W*in
   wire signed [9:0] m114_9;
   assign m114_9 =10'b0;

   // m114_10 = W*in
   wire signed [9:0] m114_10;
   assign m114_10 =10'b0;

   // m114_11 = W*in
   wire signed [9:0] m114_11;
   assign m114_11 =10'b0;

   // m114_12 = W*in
   wire signed [9:0] m114_12;
   assign m114_12 =10'b0;

   // m114_13 = W*in
   wire signed [9:0] m114_13;
   assign m114_13 =10'b0;

   // m114_14 = W*in
   wire signed [9:0] m114_14;
   assign m114_14 =10'b0;

   // m114_15 = W*in
   wire signed [9:0] m114_15;
   assign m114_15 =10'b0;

   // m114_16 = W*in
   wire signed [9:0] m114_16;
   assign m114_16 =10'b0;

   // m114_17 = W*in
   wire signed [9:0] m114_17;
   assign m114_17 =10'b0;

   // m114_18 = W*in
   wire signed [9:0] m114_18;
   assign m114_18 ={ {5{in114[5]}} , in114[5:1] };

   // m114_19 = W*in
   wire signed [9:0] m114_19;
   assign m114_19 =10'b0;

   // m114_20 = W*in
   wire signed [9:0] m114_20;
   assign m114_20 =10'b0;

   // m114_21 = W*in
   wire signed [9:0] m114_21;
   assign m114_21 =10'b0;

   // m114_22 = W*in
   wire signed [9:0] m114_22;
   assign m114_22 =10'b0;

   // m114_23 = W*in
   wire signed [9:0] m114_23;
   assign m114_23 =10'b0;

   // m114_24 = W*in
   wire signed [9:0] m114_24;
   assign m114_24 =10'b0;

   // m114_25 = W*in
   wire signed [9:0] m114_25;
   assign m114_25 =10'b0;

   // m114_26 = W*in
   wire signed [9:0] m114_26;
   assign m114_26 =10'b0;

   // m114_27 = W*in
   wire signed [9:0] m114_27;
   assign m114_27 =10'b0;

   // m114_28 = W*in
   wire signed [9:0] m114_28;
   assign m114_28 =10'b0;

   // m114_29 = W*in
   wire signed [9:0] m114_29;
   assign m114_29 ={ {5{in114[5]}} , in114[5:1] };

   // m114_30 = W*in
   wire signed [9:0] m114_30;
   assign m114_30 =10'b0;

   // m114_31 = W*in
   wire signed [9:0] m114_31;
   assign m114_31 =10'b0;

   // m114_32 = W*in
   wire signed [9:0] m114_32;
   assign m114_32 =10'b0;

   // m114_33 = W*in
   wire signed [9:0] m114_33;
   assign m114_33 =10'b0;

   // m114_34 = W*in
   wire signed [9:0] m114_34;
   assign m114_34 =10'b0;

   // m114_35 = W*in
   wire signed [9:0] m114_35;
   assign m114_35 =10'b0;

   // m114_36 = W*in
   wire signed [9:0] m114_36;
   assign m114_36 =10'b0;

   // m114_37 = W*in
   wire signed [9:0] m114_37;
   assign m114_37 =10'b0;

   // m114_38 = W*in
   wire signed [9:0] m114_38;
   assign m114_38 =10'b0;

   // m114_39 = W*in
   wire signed [9:0] m114_39;
   assign m114_39 =10'b0;

   // m114_40 = W*in
   wire signed [9:0] m114_40;
   assign m114_40 =10'b0;

   // m114_41 = W*in
   wire signed [9:0] m114_41;
   assign m114_41 =10'b0;

   // m114_42 = W*in
   wire signed [9:0] m114_42;
   assign m114_42 =10'b0;

   // m114_43 = W*in
   wire signed [9:0] m114_43;
   assign m114_43 =10'b0;

   // m114_44 = W*in
   wire signed [9:0] m114_44;
   assign m114_44 =10'b0;

   // m114_45 = W*in
   wire signed [9:0] m114_45;
   assign m114_45 =10'b0;

   // m114_46 = W*in
   wire signed [9:0] m114_46;
   assign m114_46 =10'b0;

   // m114_47 = W*in
   wire signed [9:0] m114_47;
   assign m114_47 =10'b0;

   // m114_48 = W*in
   wire signed [9:0] m114_48;
   assign m114_48 =10'b0;

   // m114_49 = W*in
   wire signed [9:0] m114_49;
   assign m114_49 =10'b0;

   // m114_50 = W*in
   wire signed [9:0] m114_50;
   assign m114_50 =10'b0;

   // m114_51 = W*in
   wire signed [9:0] m114_51;
   assign m114_51 =10'b0;

   // m114_52 = W*in
   wire signed [9:0] m114_52;
   assign m114_52 =10'b0;

   // m114_53 = W*in
   wire signed [9:0] m114_53;
   assign m114_53 =10'b0;

   // m114_54 = W*in
   wire signed [9:0] m114_54;
   assign m114_54 =10'b0;

   // m114_55 = W*in
   wire signed [9:0] m114_55;
   assign m114_55 =10'b0;

   // m114_56 = W*in
   wire signed [9:0] m114_56;
   assign m114_56 =10'b0;

   // m114_57 = W*in
   wire signed [9:0] m114_57;
   assign m114_57 =10'b0;

   // m114_58 = W*in
   wire signed [9:0] m114_58;
   assign m114_58 =10'b0;

   // m114_59 = W*in
   wire signed [9:0] m114_59;
   assign m114_59 =10'b0;

   // m114_60 = W*in
   wire signed [9:0] m114_60;
   assign m114_60 =10'b0;

   // m114_61 = W*in
   wire signed [9:0] m114_61;
   assign m114_61 =10'b0;

   // m114_62 = W*in
   wire signed [9:0] m114_62;
   assign m114_62 =10'b0;

   // m114_63 = W*in
   wire signed [9:0] m114_63;
   assign m114_63 =10'b0;

   // m114_64 = W*in
   wire signed [9:0] m114_64;
   assign m114_64 ={ {5{neg114[5]}} , neg114[5:1] };

   // m114_65 = W*in
   wire signed [9:0] m114_65;
   assign m114_65 =10'b0;

   // m114_66 = W*in
   wire signed [9:0] m114_66;
   assign m114_66 =10'b0;

   // m114_67 = W*in
   wire signed [9:0] m114_67;
   assign m114_67 =10'b0;

   // m114_68 = W*in
   wire signed [9:0] m114_68;
   assign m114_68 =10'b0;

   // m114_69 = W*in
   wire signed [9:0] m114_69;
   assign m114_69 =10'b0;

   // m114_70 = W*in
   wire signed [9:0] m114_70;
   assign m114_70 =10'b0;

   // m114_71 = W*in
   wire signed [9:0] m114_71;
   assign m114_71 =10'b0;

   // m114_72 = W*in
   wire signed [9:0] m114_72;
   assign m114_72 =10'b0;

   // m114_73 = W*in
   wire signed [9:0] m114_73;
   assign m114_73 =10'b0;

   // m114_74 = W*in
   wire signed [9:0] m114_74;
   assign m114_74 =10'b0;

   // m114_75 = W*in
   wire signed [9:0] m114_75;
   assign m114_75 =10'b0;

   // m114_76 = W*in
   wire signed [9:0] m114_76;
   assign m114_76 =10'b0;

   // m114_77 = W*in
   wire signed [9:0] m114_77;
   assign m114_77 =10'b0;

   // m114_78 = W*in
   wire signed [9:0] m114_78;
   assign m114_78 =10'b0;

   // m114_79 = W*in
   wire signed [9:0] m114_79;
   assign m114_79 =10'b0;

   // m114_80 = W*in
   wire signed [9:0] m114_80;
   assign m114_80 =10'b0;

   // m114_81 = W*in
   wire signed [9:0] m114_81;
   assign m114_81 =10'b0;

   // m114_82 = W*in
   wire signed [9:0] m114_82;
   assign m114_82 ={ {5{in114[5]}} , in114[5:1] };

   // m114_83 = W*in
   wire signed [9:0] m114_83;
   assign m114_83 =10'b0;

   // m114_84 = W*in
   wire signed [9:0] m114_84;
   assign m114_84 =10'b0;

   // m114_85 = W*in
   wire signed [9:0] m114_85;
   assign m114_85 =10'b0;

   // m114_86 = W*in
   wire signed [9:0] m114_86;
   assign m114_86 =10'b0;

   // m114_87 = W*in
   wire signed [9:0] m114_87;
   assign m114_87 =10'b0;

   // m114_88 = W*in
   wire signed [9:0] m114_88;
   assign m114_88 =10'b0;

   // m114_89 = W*in
   wire signed [9:0] m114_89;
   assign m114_89 =10'b0;

   // m114_90 = W*in
   wire signed [9:0] m114_90;
   assign m114_90 =10'b0;

   // m114_91 = W*in
   wire signed [9:0] m114_91;
   assign m114_91 =10'b0;

   // m114_92 = W*in
   wire signed [9:0] m114_92;
   assign m114_92 =10'b0;

   // m114_93 = W*in
   wire signed [9:0] m114_93;
   assign m114_93 =10'b0;

   // m114_94 = W*in
   wire signed [9:0] m114_94;
   assign m114_94 =10'b0;

   // m114_95 = W*in
   wire signed [9:0] m114_95;
   assign m114_95 =10'b0;

   // m114_96 = W*in
   wire signed [9:0] m114_96;
   assign m114_96 =10'b0;

   // m114_97 = W*in
   wire signed [9:0] m114_97;
   assign m114_97 =10'b0;

   // m114_98 = W*in
   wire signed [9:0] m114_98;
   assign m114_98 =10'b0;

   // m114_99 = W*in
   wire signed [9:0] m114_99;
   assign m114_99 =10'b0;

   // m114_100 = W*in
   wire signed [9:0] m114_100;
   assign m114_100 =10'b0;

   // m114_101 = W*in
   wire signed [9:0] m114_101;
   assign m114_101 =10'b0;

   // m114_102 = W*in
   wire signed [9:0] m114_102;
   assign m114_102 =10'b0;

   // m114_103 = W*in
   wire signed [9:0] m114_103;
   assign m114_103 =10'b0;

   // m114_104 = W*in
   wire signed [9:0] m114_104;
   assign m114_104 =10'b0;

   // m114_105 = W*in
   wire signed [9:0] m114_105;
   assign m114_105 =10'b0;

   // m114_106 = W*in
   wire signed [9:0] m114_106;
   assign m114_106 =10'b0;

   // m114_107 = W*in
   wire signed [9:0] m114_107;
   assign m114_107 =10'b0;

   // m114_108 = W*in
   wire signed [9:0] m114_108;
   assign m114_108 =10'b0;

   // m114_109 = W*in
   wire signed [9:0] m114_109;
   assign m114_109 =10'b0;

   // m114_110 = W*in
   wire signed [9:0] m114_110;
   assign m114_110 =10'b0;

   // m114_111 = W*in
   wire signed [9:0] m114_111;
   assign m114_111 =10'b0;

   // m114_112 = W*in
   wire signed [9:0] m114_112;
   assign m114_112 =10'b0;

   // m114_113 = W*in
   wire signed [9:0] m114_113;
   assign m114_113 =10'b0;

   // m114_114 = W*in
   wire signed [9:0] m114_114;
   assign m114_114 =10'b0;

   // m114_115 = W*in
   wire signed [9:0] m114_115;
   assign m114_115 =10'b0;

   // m114_116 = W*in
   wire signed [9:0] m114_116;
   assign m114_116 =10'b0;

   // m114_117 = W*in
   wire signed [9:0] m114_117;
   assign m114_117 =10'b0;

   // m115_1 = W*in
   wire signed [9:0] m115_1;
   assign m115_1 =10'b0;

   // m115_2 = W*in
   wire signed [9:0] m115_2;
   assign m115_2 =10'b0;

   // m115_3 = W*in
   wire signed [9:0] m115_3;
   assign m115_3 =10'b0;

   // m115_4 = W*in
   wire signed [9:0] m115_4;
   assign m115_4 =10'b0;

   // m115_5 = W*in
   wire signed [9:0] m115_5;
   assign m115_5 =10'b0;

   // m115_6 = W*in
   wire signed [9:0] m115_6;
   assign m115_6 =10'b0;

   // m115_7 = W*in
   wire signed [9:0] m115_7;
   assign m115_7 =10'b0;

   // m115_8 = W*in
   wire signed [9:0] m115_8;
   assign m115_8 =10'b0;

   // m115_9 = W*in
   wire signed [9:0] m115_9;
   assign m115_9 =10'b0;

   // m115_10 = W*in
   wire signed [9:0] m115_10;
   assign m115_10 =10'b0;

   // m115_11 = W*in
   wire signed [9:0] m115_11;
   assign m115_11 =10'b0;

   // m115_12 = W*in
   wire signed [9:0] m115_12;
   assign m115_12 =10'b0;

   // m115_13 = W*in
   wire signed [9:0] m115_13;
   assign m115_13 =10'b0;

   // m115_14 = W*in
   wire signed [9:0] m115_14;
   assign m115_14 =10'b0;

   // m115_15 = W*in
   wire signed [9:0] m115_15;
   assign m115_15 =10'b0;

   // m115_16 = W*in
   wire signed [9:0] m115_16;
   assign m115_16 =10'b0;

   // m115_17 = W*in
   wire signed [9:0] m115_17;
   assign m115_17 =10'b0;

   // m115_18 = W*in
   wire signed [9:0] m115_18;
   assign m115_18 =10'b0;

   // m115_19 = W*in
   wire signed [9:0] m115_19;
   assign m115_19 =10'b0;

   // m115_20 = W*in
   wire signed [9:0] m115_20;
   assign m115_20 =10'b0;

   // m115_21 = W*in
   wire signed [9:0] m115_21;
   assign m115_21 =10'b0;

   // m115_22 = W*in
   wire signed [9:0] m115_22;
   assign m115_22 =10'b0;

   // m115_23 = W*in
   wire signed [9:0] m115_23;
   assign m115_23 =10'b0;

   // m115_24 = W*in
   wire signed [9:0] m115_24;
   assign m115_24 =10'b0;

   // m115_25 = W*in
   wire signed [9:0] m115_25;
   assign m115_25 =10'b0;

   // m115_26 = W*in
   wire signed [9:0] m115_26;
   assign m115_26 =10'b0;

   // m115_27 = W*in
   wire signed [9:0] m115_27;
   assign m115_27 =10'b0;

   // m115_28 = W*in
   wire signed [9:0] m115_28;
   assign m115_28 =10'b0;

   // m115_29 = W*in
   wire signed [9:0] m115_29;
   assign m115_29 =10'b0;

   // m115_30 = W*in
   wire signed [9:0] m115_30;
   assign m115_30 =10'b0;

   // m115_31 = W*in
   wire signed [9:0] m115_31;
   assign m115_31 ={ {5{in115[5]}} , in115[5:1] };

   // m115_32 = W*in
   wire signed [9:0] m115_32;
   assign m115_32 =10'b0;

   // m115_33 = W*in
   wire signed [9:0] m115_33;
   assign m115_33 =10'b0;

   // m115_34 = W*in
   wire signed [9:0] m115_34;
   assign m115_34 =10'b0;

   // m115_35 = W*in
   wire signed [9:0] m115_35;
   assign m115_35 =10'b0;

   // m115_36 = W*in
   wire signed [9:0] m115_36;
   assign m115_36 =10'b0;

   // m115_37 = W*in
   wire signed [9:0] m115_37;
   assign m115_37 =10'b0;

   // m115_38 = W*in
   wire signed [9:0] m115_38;
   assign m115_38 =10'b0;

   // m115_39 = W*in
   wire signed [9:0] m115_39;
   assign m115_39 =10'b0;

   // m115_40 = W*in
   wire signed [9:0] m115_40;
   assign m115_40 =10'b0;

   // m115_41 = W*in
   wire signed [9:0] m115_41;
   assign m115_41 =10'b0;

   // m115_42 = W*in
   wire signed [9:0] m115_42;
   assign m115_42 =10'b0;

   // m115_43 = W*in
   wire signed [9:0] m115_43;
   assign m115_43 =10'b0;

   // m115_44 = W*in
   wire signed [9:0] m115_44;
   assign m115_44 =10'b0;

   // m115_45 = W*in
   wire signed [9:0] m115_45;
   assign m115_45 =10'b0;

   // m115_46 = W*in
   wire signed [9:0] m115_46;
   assign m115_46 =10'b0;

   // m115_47 = W*in
   wire signed [9:0] m115_47;
   assign m115_47 =10'b0;

   // m115_48 = W*in
   wire signed [9:0] m115_48;
   assign m115_48 =10'b0;

   // m115_49 = W*in
   wire signed [9:0] m115_49;
   assign m115_49 =10'b0;

   // m115_50 = W*in
   wire signed [9:0] m115_50;
   assign m115_50 =10'b0;

   // m115_51 = W*in
   wire signed [9:0] m115_51;
   assign m115_51 =10'b0;

   // m115_52 = W*in
   wire signed [9:0] m115_52;
   assign m115_52 =10'b0;

   // m115_53 = W*in
   wire signed [9:0] m115_53;
   assign m115_53 =10'b0;

   // m115_54 = W*in
   wire signed [9:0] m115_54;
   assign m115_54 =10'b0;

   // m115_55 = W*in
   wire signed [9:0] m115_55;
   assign m115_55 =10'b0;

   // m115_56 = W*in
   wire signed [9:0] m115_56;
   assign m115_56 =10'b0;

   // m115_57 = W*in
   wire signed [9:0] m115_57;
   assign m115_57 =10'b0;

   // m115_58 = W*in
   wire signed [9:0] m115_58;
   assign m115_58 =10'b0;

   // m115_59 = W*in
   wire signed [9:0] m115_59;
   assign m115_59 =10'b0;

   // m115_60 = W*in
   wire signed [9:0] m115_60;
   assign m115_60 =10'b0;

   // m115_61 = W*in
   wire signed [9:0] m115_61;
   assign m115_61 =10'b0;

   // m115_62 = W*in
   wire signed [9:0] m115_62;
   assign m115_62 =10'b0;

   // m115_63 = W*in
   wire signed [9:0] m115_63;
   assign m115_63 =10'b0;

   // m115_64 = W*in
   wire signed [9:0] m115_64;
   assign m115_64 =10'b0;

   // m115_65 = W*in
   wire signed [9:0] m115_65;
   assign m115_65 =10'b0;

   // m115_66 = W*in
   wire signed [9:0] m115_66;
   assign m115_66 =10'b0;

   // m115_67 = W*in
   wire signed [9:0] m115_67;
   assign m115_67 =10'b0;

   // m115_68 = W*in
   wire signed [9:0] m115_68;
   assign m115_68 =10'b0;

   // m115_69 = W*in
   wire signed [9:0] m115_69;
   assign m115_69 =10'b0;

   // m115_70 = W*in
   wire signed [9:0] m115_70;
   assign m115_70 =10'b0;

   // m115_71 = W*in
   wire signed [9:0] m115_71;
   assign m115_71 =10'b0;

   // m115_72 = W*in
   wire signed [9:0] m115_72;
   assign m115_72 ={ {5{in115[5]}} , in115[5:1] };

   // m115_73 = W*in
   wire signed [9:0] m115_73;
   assign m115_73 =10'b0;

   // m115_74 = W*in
   wire signed [9:0] m115_74;
   assign m115_74 =10'b0;

   // m115_75 = W*in
   wire signed [9:0] m115_75;
   assign m115_75 =10'b0;

   // m115_76 = W*in
   wire signed [9:0] m115_76;
   assign m115_76 =10'b0;

   // m115_77 = W*in
   wire signed [9:0] m115_77;
   assign m115_77 =10'b0;

   // m115_78 = W*in
   wire signed [9:0] m115_78;
   assign m115_78 =10'b0;

   // m115_79 = W*in
   wire signed [9:0] m115_79;
   assign m115_79 =10'b0;

   // m115_80 = W*in
   wire signed [9:0] m115_80;
   assign m115_80 =10'b0;

   // m115_81 = W*in
   wire signed [9:0] m115_81;
   assign m115_81 =10'b0;

   // m115_82 = W*in
   wire signed [9:0] m115_82;
   assign m115_82 =10'b0;

   // m115_83 = W*in
   wire signed [9:0] m115_83;
   assign m115_83 =10'b0;

   // m115_84 = W*in
   wire signed [9:0] m115_84;
   assign m115_84 =10'b0;

   // m115_85 = W*in
   wire signed [9:0] m115_85;
   assign m115_85 =10'b0;

   // m115_86 = W*in
   wire signed [9:0] m115_86;
   assign m115_86 =10'b0;

   // m115_87 = W*in
   wire signed [9:0] m115_87;
   assign m115_87 =10'b0;

   // m115_88 = W*in
   wire signed [9:0] m115_88;
   assign m115_88 =10'b0;

   // m115_89 = W*in
   wire signed [9:0] m115_89;
   assign m115_89 =10'b0;

   // m115_90 = W*in
   wire signed [9:0] m115_90;
   assign m115_90 =10'b0;

   // m115_91 = W*in
   wire signed [9:0] m115_91;
   assign m115_91 =10'b0;

   // m115_92 = W*in
   wire signed [9:0] m115_92;
   assign m115_92 =10'b0;

   // m115_93 = W*in
   wire signed [9:0] m115_93;
   assign m115_93 =10'b0;

   // m115_94 = W*in
   wire signed [9:0] m115_94;
   assign m115_94 =10'b0;

   // m115_95 = W*in
   wire signed [9:0] m115_95;
   assign m115_95 =10'b0;

   // m115_96 = W*in
   wire signed [9:0] m115_96;
   assign m115_96 =10'b0;

   // m115_97 = W*in
   wire signed [9:0] m115_97;
   assign m115_97 =10'b0;

   // m115_98 = W*in
   wire signed [9:0] m115_98;
   assign m115_98 =10'b0;

   // m115_99 = W*in
   wire signed [9:0] m115_99;
   assign m115_99 =10'b0;

   // m115_100 = W*in
   wire signed [9:0] m115_100;
   assign m115_100 =10'b0;

   // m115_101 = W*in
   wire signed [9:0] m115_101;
   assign m115_101 =10'b0;

   // m115_102 = W*in
   wire signed [9:0] m115_102;
   assign m115_102 =10'b0;

   // m115_103 = W*in
   wire signed [9:0] m115_103;
   assign m115_103 =10'b0;

   // m115_104 = W*in
   wire signed [9:0] m115_104;
   assign m115_104 =10'b0;

   // m115_105 = W*in
   wire signed [9:0] m115_105;
   assign m115_105 =10'b0;

   // m115_106 = W*in
   wire signed [9:0] m115_106;
   assign m115_106 =10'b0;

   // m115_107 = W*in
   wire signed [9:0] m115_107;
   assign m115_107 =10'b0;

   // m115_108 = W*in
   wire signed [9:0] m115_108;
   assign m115_108 =10'b0;

   // m115_109 = W*in
   wire signed [9:0] m115_109;
   assign m115_109 =10'b0;

   // m115_110 = W*in
   wire signed [9:0] m115_110;
   assign m115_110 =10'b0;

   // m115_111 = W*in
   wire signed [9:0] m115_111;
   assign m115_111 =10'b0;

   // m115_112 = W*in
   wire signed [9:0] m115_112;
   assign m115_112 =10'b0;

   // m115_113 = W*in
   wire signed [9:0] m115_113;
   assign m115_113 =10'b0;

   // m115_114 = W*in
   wire signed [9:0] m115_114;
   assign m115_114 =10'b0;

   // m115_115 = W*in
   wire signed [9:0] m115_115;
   assign m115_115 =10'b0;

   // m115_116 = W*in
   wire signed [9:0] m115_116;
   assign m115_116 =10'b0;

   // m115_117 = W*in
   wire signed [9:0] m115_117;
   assign m115_117 =10'b0;

   // m116_1 = W*in
   wire signed [9:0] m116_1;
   assign m116_1 ={ {4{in116[5]}} , in116[5:0] };

   // m116_2 = W*in
   wire signed [9:0] m116_2;
   assign m116_2 ={ {4{in116[5]}} , in116[5:0] };

   // m116_3 = W*in
   wire signed [9:0] m116_3;
   assign m116_3 =10'b0;

   // m116_4 = W*in
   wire signed [9:0] m116_4;
   assign m116_4 =10'b0;

   // m116_5 = W*in
   wire signed [9:0] m116_5;
   assign m116_5 =10'b0;

   // m116_6 = W*in
   wire signed [9:0] m116_6;
   assign m116_6 ={ {4{neg116[5]}} , neg116[5:0] };

   // m116_7 = W*in
   wire signed [9:0] m116_7;
   assign m116_7 =10'b0;

   // m116_8 = W*in
   wire signed [9:0] m116_8;
   assign m116_8 ={ {4{in116[5]}} , in116[5:0] };

   // m116_9 = W*in
   wire signed [9:0] m116_9;
   assign m116_9 =10'b0;

   // m116_10 = W*in
   wire signed [9:0] m116_10;
   assign m116_10 =10'b0;

   // m116_11 = W*in
   wire signed [9:0] m116_11;
   assign m116_11 =10'b0;

   // m116_12 = W*in
   wire signed [9:0] m116_12;
   assign m116_12 =10'b0;

   // m116_13 = W*in
   wire signed [9:0] m116_13;
   assign m116_13 =10'b0;

   // m116_14 = W*in
   wire signed [9:0] m116_14;
   assign m116_14 =10'b0;

   // m116_15 = W*in
   wire signed [9:0] m116_15;
   assign m116_15 ={ {4{in116[5]}} , in116[5:0] };

   // m116_16 = W*in
   wire signed [9:0] m116_16;
   assign m116_16 ={ {4{in116[5]}} , in116[5:0] };

   // m116_17 = W*in
   wire signed [9:0] m116_17;
   assign m116_17 ={ {5{in116[5]}} , in116[5:1] };

   // m116_18 = W*in
   wire signed [9:0] m116_18;
   assign m116_18 =10'b0;

   // m116_19 = W*in
   wire signed [9:0] m116_19;
   assign m116_19 =10'b0;

   // m116_20 = W*in
   wire signed [9:0] m116_20;
   assign m116_20 =10'b0;

   // m116_21 = W*in
   wire signed [9:0] m116_21;
   assign m116_21 ={ {5{neg116[5]}} , neg116[5:1] };

   // m116_22 = W*in
   wire signed [9:0] m116_22;
   assign m116_22 =10'b0;

   // m116_23 = W*in
   wire signed [9:0] m116_23;
   assign m116_23 =10'b0;

   // m116_24 = W*in
   wire signed [9:0] m116_24;
   assign m116_24 =10'b0;

   // m116_25 = W*in
   wire signed [9:0] m116_25;
   assign m116_25 =10'b0;

   // m116_26 = W*in
   wire signed [9:0] m116_26;
   assign m116_26 =10'b0;

   // m116_27 = W*in
   wire signed [9:0] m116_27;
   assign m116_27 ={ {5{in116[5]}} , in116[5:1] };

   // m116_28 = W*in
   wire signed [9:0] m116_28;
   assign m116_28 =10'b0;

   // m116_29 = W*in
   wire signed [9:0] m116_29;
   assign m116_29 ={ {5{neg116[5]}} , neg116[5:1] };

   // m116_30 = W*in
   wire signed [9:0] m116_30;
   assign m116_30 =10'b0;

   // m116_31 = W*in
   wire signed [9:0] m116_31;
   assign m116_31 ={ {5{in116[5]}} , in116[5:1] };

   // m116_32 = W*in
   wire signed [9:0] m116_32;
   assign m116_32 =10'b0;

   // m116_33 = W*in
   wire signed [9:0] m116_33;
   assign m116_33 =10'b0;

   // m116_34 = W*in
   wire signed [9:0] m116_34;
   assign m116_34 ={ {4{in116[5]}} , in116[5:0] };

   // m116_35 = W*in
   wire signed [9:0] m116_35;
   assign m116_35 =10'b0;

   // m116_36 = W*in
   wire signed [9:0] m116_36;
   assign m116_36 =10'b0;

   // m116_37 = W*in
   wire signed [9:0] m116_37;
   assign m116_37 =10'b0;

   // m116_38 = W*in
   wire signed [9:0] m116_38;
   assign m116_38 ={ {4{neg116[5]}} , neg116[5:0] };

   // m116_39 = W*in
   wire signed [9:0] m116_39;
   assign m116_39 =10'b0;

   // m116_40 = W*in
   wire signed [9:0] m116_40;
   assign m116_40 =10'b0;

   // m116_41 = W*in
   wire signed [9:0] m116_41;
   assign m116_41 =10'b0;

   // m116_42 = W*in
   wire signed [9:0] m116_42;
   assign m116_42 =10'b0;

   // m116_43 = W*in
   wire signed [9:0] m116_43;
   assign m116_43 =10'b0;

   // m116_44 = W*in
   wire signed [9:0] m116_44;
   assign m116_44 =10'b0;

   // m116_45 = W*in
   wire signed [9:0] m116_45;
   assign m116_45 =10'b0;

   // m116_46 = W*in
   wire signed [9:0] m116_46;
   assign m116_46 =10'b0;

   // m116_47 = W*in
   wire signed [9:0] m116_47;
   assign m116_47 =10'b0;

   // m116_48 = W*in
   wire signed [9:0] m116_48;
   assign m116_48 =10'b0;

   // m116_49 = W*in
   wire signed [9:0] m116_49;
   assign m116_49 =10'b0;

   // m116_50 = W*in
   wire signed [9:0] m116_50;
   assign m116_50 ={ {4{in116[5]}} , in116[5:0] };

   // m116_51 = W*in
   wire signed [9:0] m116_51;
   assign m116_51 ={ {4{in116[5]}} , in116[5:0] };

   // m116_52 = W*in
   wire signed [9:0] m116_52;
   assign m116_52 ={ {4{in116[5]}} , in116[5:0] };

   // m116_53 = W*in
   wire signed [9:0] m116_53;
   assign m116_53 =10'b0;

   // m116_54 = W*in
   wire signed [9:0] m116_54;
   assign m116_54 =10'b0;

   // m116_55 = W*in
   wire signed [9:0] m116_55;
   assign m116_55 =10'b0;

   // m116_56 = W*in
   wire signed [9:0] m116_56;
   assign m116_56 ={ {4{in116[5]}} , in116[5:0] };

   // m116_57 = W*in
   wire signed [9:0] m116_57;
   assign m116_57 =10'b0;

   // m116_58 = W*in
   wire signed [9:0] m116_58;
   assign m116_58 =10'b0;

   // m116_59 = W*in
   wire signed [9:0] m116_59;
   assign m116_59 =10'b0;

   // m116_60 = W*in
   wire signed [9:0] m116_60;
   assign m116_60 =10'b0;

   // m116_61 = W*in
   wire signed [9:0] m116_61;
   assign m116_61 =10'b0;

   // m116_62 = W*in
   wire signed [9:0] m116_62;
   assign m116_62 =10'b0;

   // m116_63 = W*in
   wire signed [9:0] m116_63;
   assign m116_63 =10'b0;

   // m116_64 = W*in
   wire signed [9:0] m116_64;
   assign m116_64 ={ {5{neg116[5]}} , neg116[5:1] };

   // m116_65 = W*in
   wire signed [9:0] m116_65;
   assign m116_65 ={ {4{neg116[5]}} , neg116[5:0] };

   // m116_66 = W*in
   wire signed [9:0] m116_66;
   assign m116_66 =10'b0;

   // m116_67 = W*in
   wire signed [9:0] m116_67;
   assign m116_67 =10'b0;

   // m116_68 = W*in
   wire signed [9:0] m116_68;
   assign m116_68 ={ {4{in116[5]}} , in116[5:0] };

   // m116_69 = W*in
   wire signed [9:0] m116_69;
   assign m116_69 ={ {5{neg116[5]}} , neg116[5:1] };

   // m116_70 = W*in
   wire signed [9:0] m116_70;
   assign m116_70 ={ {4{neg116[5]}} , neg116[5:0] };

   // m116_71 = W*in
   wire signed [9:0] m116_71;
   assign m116_71 =10'b0;

   // m116_72 = W*in
   wire signed [9:0] m116_72;
   assign m116_72 =10'b0;

   // m116_73 = W*in
   wire signed [9:0] m116_73;
   assign m116_73 =10'b0;

   // m116_74 = W*in
   wire signed [9:0] m116_74;
   assign m116_74 =10'b0;

   // m116_75 = W*in
   wire signed [9:0] m116_75;
   assign m116_75 ={ {5{in116[5]}} , in116[5:1] };

   // m116_76 = W*in
   wire signed [9:0] m116_76;
   assign m116_76 =10'b0;

   // m116_77 = W*in
   wire signed [9:0] m116_77;
   assign m116_77 =10'b0;

   // m116_78 = W*in
   wire signed [9:0] m116_78;
   assign m116_78 =10'b0;

   // m116_79 = W*in
   wire signed [9:0] m116_79;
   assign m116_79 =10'b0;

   // m116_80 = W*in
   wire signed [9:0] m116_80;
   assign m116_80 =10'b0;

   // m116_81 = W*in
   wire signed [9:0] m116_81;
   assign m116_81 =10'b0;

   // m116_82 = W*in
   wire signed [9:0] m116_82;
   assign m116_82 =10'b0;

   // m116_83 = W*in
   wire signed [9:0] m116_83;
   assign m116_83 =10'b0;

   // m116_84 = W*in
   wire signed [9:0] m116_84;
   assign m116_84 =10'b0;

   // m116_85 = W*in
   wire signed [9:0] m116_85;
   assign m116_85 =10'b0;

   // m116_86 = W*in
   wire signed [9:0] m116_86;
   assign m116_86 =10'b0;

   // m116_87 = W*in
   wire signed [9:0] m116_87;
   assign m116_87 =10'b0;

   // m116_88 = W*in
   wire signed [9:0] m116_88;
   assign m116_88 ={ {4{in116[5]}} , in116[5:0] };

   // m116_89 = W*in
   wire signed [9:0] m116_89;
   assign m116_89 =10'b0;

   // m116_90 = W*in
   wire signed [9:0] m116_90;
   assign m116_90 ={ {4{in116[5]}} , in116[5:0] };

   // m116_91 = W*in
   wire signed [9:0] m116_91;
   assign m116_91 =10'b0;

   // m116_92 = W*in
   wire signed [9:0] m116_92;
   assign m116_92 =10'b0;

   // m116_93 = W*in
   wire signed [9:0] m116_93;
   assign m116_93 =10'b0;

   // m116_94 = W*in
   wire signed [9:0] m116_94;
   assign m116_94 =10'b0;

   // m116_95 = W*in
   wire signed [9:0] m116_95;
   assign m116_95 =10'b0;

   // m116_96 = W*in
   wire signed [9:0] m116_96;
   assign m116_96 =10'b0;

   // m116_97 = W*in
   wire signed [9:0] m116_97;
   assign m116_97 =10'b0;

   // m116_98 = W*in
   wire signed [9:0] m116_98;
   assign m116_98 ={ {4{in116[5]}} , in116[5:0] };

   // m116_99 = W*in
   wire signed [9:0] m116_99;
   assign m116_99 ={ {4{neg116[5]}} , neg116[5:0] };

   // m116_100 = W*in
   wire signed [9:0] m116_100;
   assign m116_100 =10'b0;

   // m116_101 = W*in
   wire signed [9:0] m116_101;
   assign m116_101 =10'b0;

   // m116_102 = W*in
   wire signed [9:0] m116_102;
   assign m116_102 =10'b0;

   // m116_103 = W*in
   wire signed [9:0] m116_103;
   assign m116_103 =10'b0;

   // m116_104 = W*in
   wire signed [9:0] m116_104;
   assign m116_104 =10'b0;

   // m116_105 = W*in
   wire signed [9:0] m116_105;
   assign m116_105 ={ {4{in116[5]}} , in116[5:0] };

   // m116_106 = W*in
   wire signed [9:0] m116_106;
   assign m116_106 =10'b0;

   // m116_107 = W*in
   wire signed [9:0] m116_107;
   assign m116_107 ={ {4{in116[5]}} , in116[5:0] };

   // m116_108 = W*in
   wire signed [9:0] m116_108;
   assign m116_108 ={ {5{neg116[5]}} , neg116[5:1] };

   // m116_109 = W*in
   wire signed [9:0] m116_109;
   assign m116_109 ={ {5{neg116[5]}} , neg116[5:1] };

   // m116_110 = W*in
   wire signed [9:0] m116_110;
   assign m116_110 ={ {4{neg116[5]}} , neg116[5:0] };

   // m116_111 = W*in
   wire signed [9:0] m116_111;
   assign m116_111 =10'b0;

   // m116_112 = W*in
   wire signed [9:0] m116_112;
   assign m116_112 =10'b0;

   // m116_113 = W*in
   wire signed [9:0] m116_113;
   assign m116_113 ={ {4{in116[5]}} , in116[5:0] };

   // m116_114 = W*in
   wire signed [9:0] m116_114;
   assign m116_114 =10'b0;

   // m116_115 = W*in
   wire signed [9:0] m116_115;
   assign m116_115 =10'b0;

   // m116_116 = W*in
   wire signed [9:0] m116_116;
   assign m116_116 =10'b0;

   // m116_117 = W*in
   wire signed [9:0] m116_117;
   assign m116_117 =10'b0;

   // m117_1 = W*in
   wire signed [9:0] m117_1;
   assign m117_1 =10'b0;

   // m117_2 = W*in
   wire signed [9:0] m117_2;
   assign m117_2 =10'b0;

   // m117_3 = W*in
   wire signed [9:0] m117_3;
   assign m117_3 =10'b0;

   // m117_4 = W*in
   wire signed [9:0] m117_4;
   assign m117_4 =10'b0;

   // m117_5 = W*in
   wire signed [9:0] m117_5;
   assign m117_5 =10'b0;

   // m117_6 = W*in
   wire signed [9:0] m117_6;
   assign m117_6 ={ {4{in117[5]}} , in117[5:0] };

   // m117_7 = W*in
   wire signed [9:0] m117_7;
   assign m117_7 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_8 = W*in
   wire signed [9:0] m117_8;
   assign m117_8 =10'b0;

   // m117_9 = W*in
   wire signed [9:0] m117_9;
   assign m117_9 =10'b0;

   // m117_10 = W*in
   wire signed [9:0] m117_10;
   assign m117_10 =10'b0;

   // m117_11 = W*in
   wire signed [9:0] m117_11;
   assign m117_11 =10'b0;

   // m117_12 = W*in
   wire signed [9:0] m117_12;
   assign m117_12 =10'b0;

   // m117_13 = W*in
   wire signed [9:0] m117_13;
   assign m117_13 =10'b0;

   // m117_14 = W*in
   wire signed [9:0] m117_14;
   assign m117_14 =10'b0;

   // m117_15 = W*in
   wire signed [9:0] m117_15;
   assign m117_15 ={ {4{in117[5]}} , in117[5:0] };

   // m117_16 = W*in
   wire signed [9:0] m117_16;
   assign m117_16 =10'b0;

   // m117_17 = W*in
   wire signed [9:0] m117_17;
   assign m117_17 =10'b0;

   // m117_18 = W*in
   wire signed [9:0] m117_18;
   assign m117_18 =10'b0;

   // m117_19 = W*in
   wire signed [9:0] m117_19;
   assign m117_19 =10'b0;

   // m117_20 = W*in
   wire signed [9:0] m117_20;
   assign m117_20 =10'b0;

   // m117_21 = W*in
   wire signed [9:0] m117_21;
   assign m117_21 =10'b0;

   // m117_22 = W*in
   wire signed [9:0] m117_22;
   assign m117_22 =10'b0;

   // m117_23 = W*in
   wire signed [9:0] m117_23;
   assign m117_23 =10'b0;

   // m117_24 = W*in
   wire signed [9:0] m117_24;
   assign m117_24 =10'b0;

   // m117_25 = W*in
   wire signed [9:0] m117_25;
   assign m117_25 =10'b0;

   // m117_26 = W*in
   wire signed [9:0] m117_26;
   assign m117_26 =10'b0;

   // m117_27 = W*in
   wire signed [9:0] m117_27;
   assign m117_27 =10'b0;

   // m117_28 = W*in
   wire signed [9:0] m117_28;
   assign m117_28 =10'b0;

   // m117_29 = W*in
   wire signed [9:0] m117_29;
   assign m117_29 ={ {4{in117[5]}} , in117[5:0] };

   // m117_30 = W*in
   wire signed [9:0] m117_30;
   assign m117_30 =10'b0;

   // m117_31 = W*in
   wire signed [9:0] m117_31;
   assign m117_31 =10'b0;

   // m117_32 = W*in
   wire signed [9:0] m117_32;
   assign m117_32 =10'b0;

   // m117_33 = W*in
   wire signed [9:0] m117_33;
   assign m117_33 =10'b0;

   // m117_34 = W*in
   wire signed [9:0] m117_34;
   assign m117_34 =10'b0;

   // m117_35 = W*in
   wire signed [9:0] m117_35;
   assign m117_35 =10'b0;

   // m117_36 = W*in
   wire signed [9:0] m117_36;
   assign m117_36 =10'b0;

   // m117_37 = W*in
   wire signed [9:0] m117_37;
   assign m117_37 =10'b0;

   // m117_38 = W*in
   wire signed [9:0] m117_38;
   assign m117_38 =10'b0;

   // m117_39 = W*in
   wire signed [9:0] m117_39;
   assign m117_39 =10'b0;

   // m117_40 = W*in
   wire signed [9:0] m117_40;
   assign m117_40 =10'b0;

   // m117_41 = W*in
   wire signed [9:0] m117_41;
   assign m117_41 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_42 = W*in
   wire signed [9:0] m117_42;
   assign m117_42 =10'b0;

   // m117_43 = W*in
   wire signed [9:0] m117_43;
   assign m117_43 =10'b0;

   // m117_44 = W*in
   wire signed [9:0] m117_44;
   assign m117_44 =10'b0;

   // m117_45 = W*in
   wire signed [9:0] m117_45;
   assign m117_45 =10'b0;

   // m117_46 = W*in
   wire signed [9:0] m117_46;
   assign m117_46 =10'b0;

   // m117_47 = W*in
   wire signed [9:0] m117_47;
   assign m117_47 =10'b0;

   // m117_48 = W*in
   wire signed [9:0] m117_48;
   assign m117_48 =10'b0;

   // m117_49 = W*in
   wire signed [9:0] m117_49;
   assign m117_49 =10'b0;

   // m117_50 = W*in
   wire signed [9:0] m117_50;
   assign m117_50 =10'b0;

   // m117_51 = W*in
   wire signed [9:0] m117_51;
   assign m117_51 =10'b0;

   // m117_52 = W*in
   wire signed [9:0] m117_52;
   assign m117_52 =10'b0;

   // m117_53 = W*in
   wire signed [9:0] m117_53;
   assign m117_53 =10'b0;

   // m117_54 = W*in
   wire signed [9:0] m117_54;
   assign m117_54 =10'b0;

   // m117_55 = W*in
   wire signed [9:0] m117_55;
   assign m117_55 =10'b0;

   // m117_56 = W*in
   wire signed [9:0] m117_56;
   assign m117_56 =10'b0;

   // m117_57 = W*in
   wire signed [9:0] m117_57;
   assign m117_57 =10'b0;

   // m117_58 = W*in
   wire signed [9:0] m117_58;
   assign m117_58 =10'b0;

   // m117_59 = W*in
   wire signed [9:0] m117_59;
   assign m117_59 =10'b0;

   // m117_60 = W*in
   wire signed [9:0] m117_60;
   assign m117_60 =10'b0;

   // m117_61 = W*in
   wire signed [9:0] m117_61;
   assign m117_61 =10'b0;

   // m117_62 = W*in
   wire signed [9:0] m117_62;
   assign m117_62 =10'b0;

   // m117_63 = W*in
   wire signed [9:0] m117_63;
   assign m117_63 =10'b0;

   // m117_64 = W*in
   wire signed [9:0] m117_64;
   assign m117_64 ={ {5{neg117[5]}} , neg117[5:1] };

   // m117_65 = W*in
   wire signed [9:0] m117_65;
   assign m117_65 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_66 = W*in
   wire signed [9:0] m117_66;
   assign m117_66 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_67 = W*in
   wire signed [9:0] m117_67;
   assign m117_67 =10'b0;

   // m117_68 = W*in
   wire signed [9:0] m117_68;
   assign m117_68 ={ {4{in117[5]}} , in117[5:0] };

   // m117_69 = W*in
   wire signed [9:0] m117_69;
   assign m117_69 ={ {5{in117[5]}} , in117[5:1] };

   // m117_70 = W*in
   wire signed [9:0] m117_70;
   assign m117_70 =10'b0;

   // m117_71 = W*in
   wire signed [9:0] m117_71;
   assign m117_71 =10'b0;

   // m117_72 = W*in
   wire signed [9:0] m117_72;
   assign m117_72 ={ {5{in117[5]}} , in117[5:1] };

   // m117_73 = W*in
   wire signed [9:0] m117_73;
   assign m117_73 ={ {5{neg117[5]}} , neg117[5:1] };

   // m117_74 = W*in
   wire signed [9:0] m117_74;
   assign m117_74 =10'b0;

   // m117_75 = W*in
   wire signed [9:0] m117_75;
   assign m117_75 =10'b0;

   // m117_76 = W*in
   wire signed [9:0] m117_76;
   assign m117_76 ={ {4{in117[5]}} , in117[5:0] };

   // m117_77 = W*in
   wire signed [9:0] m117_77;
   assign m117_77 =10'b0;

   // m117_78 = W*in
   wire signed [9:0] m117_78;
   assign m117_78 =10'b0;

   // m117_79 = W*in
   wire signed [9:0] m117_79;
   assign m117_79 =10'b0;

   // m117_80 = W*in
   wire signed [9:0] m117_80;
   assign m117_80 =10'b0;

   // m117_81 = W*in
   wire signed [9:0] m117_81;
   assign m117_81 =10'b0;

   // m117_82 = W*in
   wire signed [9:0] m117_82;
   assign m117_82 =10'b0;

   // m117_83 = W*in
   wire signed [9:0] m117_83;
   assign m117_83 =10'b0;

   // m117_84 = W*in
   wire signed [9:0] m117_84;
   assign m117_84 =10'b0;

   // m117_85 = W*in
   wire signed [9:0] m117_85;
   assign m117_85 =10'b0;

   // m117_86 = W*in
   wire signed [9:0] m117_86;
   assign m117_86 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_87 = W*in
   wire signed [9:0] m117_87;
   assign m117_87 =10'b0;

   // m117_88 = W*in
   wire signed [9:0] m117_88;
   assign m117_88 ={ {4{in117[5]}} , in117[5:0] };

   // m117_89 = W*in
   wire signed [9:0] m117_89;
   assign m117_89 =10'b0;

   // m117_90 = W*in
   wire signed [9:0] m117_90;
   assign m117_90 ={ {4{in117[5]}} , in117[5:0] };

   // m117_91 = W*in
   wire signed [9:0] m117_91;
   assign m117_91 =10'b0;

   // m117_92 = W*in
   wire signed [9:0] m117_92;
   assign m117_92 ={ {4{in117[5]}} , in117[5:0] };

   // m117_93 = W*in
   wire signed [9:0] m117_93;
   assign m117_93 =10'b0;

   // m117_94 = W*in
   wire signed [9:0] m117_94;
   assign m117_94 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_95 = W*in
   wire signed [9:0] m117_95;
   assign m117_95 =10'b0;

   // m117_96 = W*in
   wire signed [9:0] m117_96;
   assign m117_96 =10'b0;

   // m117_97 = W*in
   wire signed [9:0] m117_97;
   assign m117_97 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_98 = W*in
   wire signed [9:0] m117_98;
   assign m117_98 ={ {4{in117[5]}} , in117[5:0] };

   // m117_99 = W*in
   wire signed [9:0] m117_99;
   assign m117_99 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_100 = W*in
   wire signed [9:0] m117_100;
   assign m117_100 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_101 = W*in
   wire signed [9:0] m117_101;
   assign m117_101 =10'b0;

   // m117_102 = W*in
   wire signed [9:0] m117_102;
   assign m117_102 =10'b0;

   // m117_103 = W*in
   wire signed [9:0] m117_103;
   assign m117_103 =10'b0;

   // m117_104 = W*in
   wire signed [9:0] m117_104;
   assign m117_104 =10'b0;

   // m117_105 = W*in
   wire signed [9:0] m117_105;
   assign m117_105 =10'b0;

   // m117_106 = W*in
   wire signed [9:0] m117_106;
   assign m117_106 =10'b0;

   // m117_107 = W*in
   wire signed [9:0] m117_107;
   assign m117_107 =10'b0;

   // m117_108 = W*in
   wire signed [9:0] m117_108;
   assign m117_108 ={ {5{neg117[5]}} , neg117[5:1] };

   // m117_109 = W*in
   wire signed [9:0] m117_109;
   assign m117_109 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_110 = W*in
   wire signed [9:0] m117_110;
   assign m117_110 =10'b0;

   // m117_111 = W*in
   wire signed [9:0] m117_111;
   assign m117_111 =10'b0;

   // m117_112 = W*in
   wire signed [9:0] m117_112;
   assign m117_112 =10'b0;

   // m117_113 = W*in
   wire signed [9:0] m117_113;
   assign m117_113 ={ {5{neg117[5]}} , neg117[5:1] };

   // m117_114 = W*in
   wire signed [9:0] m117_114;
   assign m117_114 ={ {5{neg117[5]}} , neg117[5:1] };

   // m117_115 = W*in
   wire signed [9:0] m117_115;
   assign m117_115 =10'b0;

   // m117_116 = W*in
   wire signed [9:0] m117_116;
   assign m117_116 ={ {4{neg117[5]}} , neg117[5:0] };

   // m117_117 = W*in
   wire signed [9:0] m117_117;
   assign m117_117 =10'b0;

   // m118_1 = W*in
   wire signed [9:0] m118_1;
   assign m118_1 =10'b0;

   // m118_2 = W*in
   wire signed [9:0] m118_2;
   assign m118_2 =10'b0;

   // m118_3 = W*in
   wire signed [9:0] m118_3;
   assign m118_3 =10'b0;

   // m118_4 = W*in
   wire signed [9:0] m118_4;
   assign m118_4 =10'b0;

   // m118_5 = W*in
   wire signed [9:0] m118_5;
   assign m118_5 =10'b0;

   // m118_6 = W*in
   wire signed [9:0] m118_6;
   assign m118_6 =10'b0;

   // m118_7 = W*in
   wire signed [9:0] m118_7;
   assign m118_7 ={ {4{in118[5]}} , in118[5:0] };

   // m118_8 = W*in
   wire signed [9:0] m118_8;
   assign m118_8 =10'b0;

   // m118_9 = W*in
   wire signed [9:0] m118_9;
   assign m118_9 =10'b0;

   // m118_10 = W*in
   wire signed [9:0] m118_10;
   assign m118_10 =10'b0;

   // m118_11 = W*in
   wire signed [9:0] m118_11;
   assign m118_11 =10'b0;

   // m118_12 = W*in
   wire signed [9:0] m118_12;
   assign m118_12 =10'b0;

   // m118_13 = W*in
   wire signed [9:0] m118_13;
   assign m118_13 =10'b0;

   // m118_14 = W*in
   wire signed [9:0] m118_14;
   assign m118_14 =10'b0;

   // m118_15 = W*in
   wire signed [9:0] m118_15;
   assign m118_15 =10'b0;

   // m118_16 = W*in
   wire signed [9:0] m118_16;
   assign m118_16 =10'b0;

   // m118_17 = W*in
   wire signed [9:0] m118_17;
   assign m118_17 =10'b0;

   // m118_18 = W*in
   wire signed [9:0] m118_18;
   assign m118_18 =10'b0;

   // m118_19 = W*in
   wire signed [9:0] m118_19;
   assign m118_19 ={ {5{neg118[5]}} , neg118[5:1] };

   // m118_20 = W*in
   wire signed [9:0] m118_20;
   assign m118_20 ={ {5{neg118[5]}} , neg118[5:1] };

   // m118_21 = W*in
   wire signed [9:0] m118_21;
   assign m118_21 ={ {5{in118[5]}} , in118[5:1] };

   // m118_22 = W*in
   wire signed [9:0] m118_22;
   assign m118_22 =10'b0;

   // m118_23 = W*in
   wire signed [9:0] m118_23;
   assign m118_23 ={ {5{in118[5]}} , in118[5:1] };

   // m118_24 = W*in
   wire signed [9:0] m118_24;
   assign m118_24 =10'b0;

   // m118_25 = W*in
   wire signed [9:0] m118_25;
   assign m118_25 =10'b0;

   // m118_26 = W*in
   wire signed [9:0] m118_26;
   assign m118_26 =10'b0;

   // m118_27 = W*in
   wire signed [9:0] m118_27;
   assign m118_27 =10'b0;

   // m118_28 = W*in
   wire signed [9:0] m118_28;
   assign m118_28 =10'b0;

   // m118_29 = W*in
   wire signed [9:0] m118_29;
   assign m118_29 ={ {5{in118[5]}} , in118[5:1] };

   // m118_30 = W*in
   wire signed [9:0] m118_30;
   assign m118_30 =10'b0;

   // m118_31 = W*in
   wire signed [9:0] m118_31;
   assign m118_31 =10'b0;

   // m118_32 = W*in
   wire signed [9:0] m118_32;
   assign m118_32 =10'b0;

   // m118_33 = W*in
   wire signed [9:0] m118_33;
   assign m118_33 =10'b0;

   // m118_34 = W*in
   wire signed [9:0] m118_34;
   assign m118_34 =10'b0;

   // m118_35 = W*in
   wire signed [9:0] m118_35;
   assign m118_35 =10'b0;

   // m118_36 = W*in
   wire signed [9:0] m118_36;
   assign m118_36 =10'b0;

   // m118_37 = W*in
   wire signed [9:0] m118_37;
   assign m118_37 =10'b0;

   // m118_38 = W*in
   wire signed [9:0] m118_38;
   assign m118_38 =10'b0;

   // m118_39 = W*in
   wire signed [9:0] m118_39;
   assign m118_39 =10'b0;

   // m118_40 = W*in
   wire signed [9:0] m118_40;
   assign m118_40 =10'b0;

   // m118_41 = W*in
   wire signed [9:0] m118_41;
   assign m118_41 =10'b0;

   // m118_42 = W*in
   wire signed [9:0] m118_42;
   assign m118_42 =10'b0;

   // m118_43 = W*in
   wire signed [9:0] m118_43;
   assign m118_43 =10'b0;

   // m118_44 = W*in
   wire signed [9:0] m118_44;
   assign m118_44 =10'b0;

   // m118_45 = W*in
   wire signed [9:0] m118_45;
   assign m118_45 =10'b0;

   // m118_46 = W*in
   wire signed [9:0] m118_46;
   assign m118_46 =10'b0;

   // m118_47 = W*in
   wire signed [9:0] m118_47;
   assign m118_47 =10'b0;

   // m118_48 = W*in
   wire signed [9:0] m118_48;
   assign m118_48 ={ {4{neg118[5]}} , neg118[5:0] };

   // m118_49 = W*in
   wire signed [9:0] m118_49;
   assign m118_49 =10'b0;

   // m118_50 = W*in
   wire signed [9:0] m118_50;
   assign m118_50 =10'b0;

   // m118_51 = W*in
   wire signed [9:0] m118_51;
   assign m118_51 =10'b0;

   // m118_52 = W*in
   wire signed [9:0] m118_52;
   assign m118_52 =10'b0;

   // m118_53 = W*in
   wire signed [9:0] m118_53;
   assign m118_53 =10'b0;

   // m118_54 = W*in
   wire signed [9:0] m118_54;
   assign m118_54 =10'b0;

   // m118_55 = W*in
   wire signed [9:0] m118_55;
   assign m118_55 =10'b0;

   // m118_56 = W*in
   wire signed [9:0] m118_56;
   assign m118_56 =10'b0;

   // m118_57 = W*in
   wire signed [9:0] m118_57;
   assign m118_57 =10'b0;

   // m118_58 = W*in
   wire signed [9:0] m118_58;
   assign m118_58 =10'b0;

   // m118_59 = W*in
   wire signed [9:0] m118_59;
   assign m118_59 =10'b0;

   // m118_60 = W*in
   wire signed [9:0] m118_60;
   assign m118_60 =10'b0;

   // m118_61 = W*in
   wire signed [9:0] m118_61;
   assign m118_61 =10'b0;

   // m118_62 = W*in
   wire signed [9:0] m118_62;
   assign m118_62 =10'b0;

   // m118_63 = W*in
   wire signed [9:0] m118_63;
   assign m118_63 =10'b0;

   // m118_64 = W*in
   wire signed [9:0] m118_64;
   assign m118_64 =10'b0;

   // m118_65 = W*in
   wire signed [9:0] m118_65;
   assign m118_65 ={ {5{neg118[5]}} , neg118[5:1] };

   // m118_66 = W*in
   wire signed [9:0] m118_66;
   assign m118_66 ={ {5{neg118[5]}} , neg118[5:1] };

   // m118_67 = W*in
   wire signed [9:0] m118_67;
   assign m118_67 =10'b0;

   // m118_68 = W*in
   wire signed [9:0] m118_68;
   assign m118_68 =10'b0;

   // m118_69 = W*in
   wire signed [9:0] m118_69;
   assign m118_69 =10'b0;

   // m118_70 = W*in
   wire signed [9:0] m118_70;
   assign m118_70 =10'b0;

   // m118_71 = W*in
   wire signed [9:0] m118_71;
   assign m118_71 =10'b0;

   // m118_72 = W*in
   wire signed [9:0] m118_72;
   assign m118_72 =10'b0;

   // m118_73 = W*in
   wire signed [9:0] m118_73;
   assign m118_73 =10'b0;

   // m118_74 = W*in
   wire signed [9:0] m118_74;
   assign m118_74 ={ {4{neg118[5]}} , neg118[5:0] };

   // m118_75 = W*in
   wire signed [9:0] m118_75;
   assign m118_75 =10'b0;

   // m118_76 = W*in
   wire signed [9:0] m118_76;
   assign m118_76 ={ {4{in118[5]}} , in118[5:0] };

   // m118_77 = W*in
   wire signed [9:0] m118_77;
   assign m118_77 =10'b0;

   // m118_78 = W*in
   wire signed [9:0] m118_78;
   assign m118_78 ={ {4{neg118[5]}} , neg118[5:0] };

   // m118_79 = W*in
   wire signed [9:0] m118_79;
   assign m118_79 =10'b0;

   // m118_80 = W*in
   wire signed [9:0] m118_80;
   assign m118_80 =10'b0;

   // m118_81 = W*in
   wire signed [9:0] m118_81;
   assign m118_81 =10'b0;

   // m118_82 = W*in
   wire signed [9:0] m118_82;
   assign m118_82 =10'b0;

   // m118_83 = W*in
   wire signed [9:0] m118_83;
   assign m118_83 =10'b0;

   // m118_84 = W*in
   wire signed [9:0] m118_84;
   assign m118_84 =10'b0;

   // m118_85 = W*in
   wire signed [9:0] m118_85;
   assign m118_85 =10'b0;

   // m118_86 = W*in
   wire signed [9:0] m118_86;
   assign m118_86 =10'b0;

   // m118_87 = W*in
   wire signed [9:0] m118_87;
   assign m118_87 =10'b0;

   // m118_88 = W*in
   wire signed [9:0] m118_88;
   assign m118_88 =10'b0;

   // m118_89 = W*in
   wire signed [9:0] m118_89;
   assign m118_89 =10'b0;

   // m118_90 = W*in
   wire signed [9:0] m118_90;
   assign m118_90 =10'b0;

   // m118_91 = W*in
   wire signed [9:0] m118_91;
   assign m118_91 =10'b0;

   // m118_92 = W*in
   wire signed [9:0] m118_92;
   assign m118_92 =10'b0;

   // m118_93 = W*in
   wire signed [9:0] m118_93;
   assign m118_93 =10'b0;

   // m118_94 = W*in
   wire signed [9:0] m118_94;
   assign m118_94 =10'b0;

   // m118_95 = W*in
   wire signed [9:0] m118_95;
   assign m118_95 =10'b0;

   // m118_96 = W*in
   wire signed [9:0] m118_96;
   assign m118_96 =10'b0;

   // m118_97 = W*in
   wire signed [9:0] m118_97;
   assign m118_97 =10'b0;

   // m118_98 = W*in
   wire signed [9:0] m118_98;
   assign m118_98 =10'b0;

   // m118_99 = W*in
   wire signed [9:0] m118_99;
   assign m118_99 =10'b0;

   // m118_100 = W*in
   wire signed [9:0] m118_100;
   assign m118_100 =10'b0;

   // m118_101 = W*in
   wire signed [9:0] m118_101;
   assign m118_101 =10'b0;

   // m118_102 = W*in
   wire signed [9:0] m118_102;
   assign m118_102 =10'b0;

   // m118_103 = W*in
   wire signed [9:0] m118_103;
   assign m118_103 =10'b0;

   // m118_104 = W*in
   wire signed [9:0] m118_104;
   assign m118_104 =10'b0;

   // m118_105 = W*in
   wire signed [9:0] m118_105;
   assign m118_105 =10'b0;

   // m118_106 = W*in
   wire signed [9:0] m118_106;
   assign m118_106 =10'b0;

   // m118_107 = W*in
   wire signed [9:0] m118_107;
   assign m118_107 =10'b0;

   // m118_108 = W*in
   wire signed [9:0] m118_108;
   assign m118_108 ={ {5{neg118[5]}} , neg118[5:1] };

   // m118_109 = W*in
   wire signed [9:0] m118_109;
   assign m118_109 =10'b0;

   // m118_110 = W*in
   wire signed [9:0] m118_110;
   assign m118_110 =10'b0;

   // m118_111 = W*in
   wire signed [9:0] m118_111;
   assign m118_111 =10'b0;

   // m118_112 = W*in
   wire signed [9:0] m118_112;
   assign m118_112 =10'b0;

   // m118_113 = W*in
   wire signed [9:0] m118_113;
   assign m118_113 =10'b0;

   // m118_114 = W*in
   wire signed [9:0] m118_114;
   assign m118_114 =10'b0;

   // m118_115 = W*in
   wire signed [9:0] m118_115;
   assign m118_115 =10'b0;

   // m118_116 = W*in
   wire signed [9:0] m118_116;
   assign m118_116 =10'b0;

   // m118_117 = W*in
   wire signed [9:0] m118_117;
   assign m118_117 =10'b0;

   // m119_1 = W*in
   wire signed [9:0] m119_1;
   assign m119_1 =10'b0;

   // m119_2 = W*in
   wire signed [9:0] m119_2;
   assign m119_2 =10'b0;

   // m119_3 = W*in
   wire signed [9:0] m119_3;
   assign m119_3 =10'b0;

   // m119_4 = W*in
   wire signed [9:0] m119_4;
   assign m119_4 =10'b0;

   // m119_5 = W*in
   wire signed [9:0] m119_5;
   assign m119_5 =10'b0;

   // m119_6 = W*in
   wire signed [9:0] m119_6;
   assign m119_6 =10'b0;

   // m119_7 = W*in
   wire signed [9:0] m119_7;
   assign m119_7 =10'b0;

   // m119_8 = W*in
   wire signed [9:0] m119_8;
   assign m119_8 =10'b0;

   // m119_9 = W*in
   wire signed [9:0] m119_9;
   assign m119_9 =10'b0;

   // m119_10 = W*in
   wire signed [9:0] m119_10;
   assign m119_10 =10'b0;

   // m119_11 = W*in
   wire signed [9:0] m119_11;
   assign m119_11 =10'b0;

   // m119_12 = W*in
   wire signed [9:0] m119_12;
   assign m119_12 =10'b0;

   // m119_13 = W*in
   wire signed [9:0] m119_13;
   assign m119_13 =10'b0;

   // m119_14 = W*in
   wire signed [9:0] m119_14;
   assign m119_14 =10'b0;

   // m119_15 = W*in
   wire signed [9:0] m119_15;
   assign m119_15 =10'b0;

   // m119_16 = W*in
   wire signed [9:0] m119_16;
   assign m119_16 =10'b0;

   // m119_17 = W*in
   wire signed [9:0] m119_17;
   assign m119_17 =10'b0;

   // m119_18 = W*in
   wire signed [9:0] m119_18;
   assign m119_18 =10'b0;

   // m119_19 = W*in
   wire signed [9:0] m119_19;
   assign m119_19 =10'b0;

   // m119_20 = W*in
   wire signed [9:0] m119_20;
   assign m119_20 =10'b0;

   // m119_21 = W*in
   wire signed [9:0] m119_21;
   assign m119_21 ={ {5{in119[5]}} , in119[5:1] };

   // m119_22 = W*in
   wire signed [9:0] m119_22;
   assign m119_22 =10'b0;

   // m119_23 = W*in
   wire signed [9:0] m119_23;
   assign m119_23 =10'b0;

   // m119_24 = W*in
   wire signed [9:0] m119_24;
   assign m119_24 =10'b0;

   // m119_25 = W*in
   wire signed [9:0] m119_25;
   assign m119_25 =10'b0;

   // m119_26 = W*in
   wire signed [9:0] m119_26;
   assign m119_26 =10'b0;

   // m119_27 = W*in
   wire signed [9:0] m119_27;
   assign m119_27 ={ {5{neg119[5]}} , neg119[5:1] };

   // m119_28 = W*in
   wire signed [9:0] m119_28;
   assign m119_28 ={ {5{neg119[5]}} , neg119[5:1] };

   // m119_29 = W*in
   wire signed [9:0] m119_29;
   assign m119_29 ={ {5{in119[5]}} , in119[5:1] };

   // m119_30 = W*in
   wire signed [9:0] m119_30;
   assign m119_30 =10'b0;

   // m119_31 = W*in
   wire signed [9:0] m119_31;
   assign m119_31 =10'b0;

   // m119_32 = W*in
   wire signed [9:0] m119_32;
   assign m119_32 =10'b0;

   // m119_33 = W*in
   wire signed [9:0] m119_33;
   assign m119_33 =10'b0;

   // m119_34 = W*in
   wire signed [9:0] m119_34;
   assign m119_34 =10'b0;

   // m119_35 = W*in
   wire signed [9:0] m119_35;
   assign m119_35 =10'b0;

   // m119_36 = W*in
   wire signed [9:0] m119_36;
   assign m119_36 =10'b0;

   // m119_37 = W*in
   wire signed [9:0] m119_37;
   assign m119_37 =10'b0;

   // m119_38 = W*in
   wire signed [9:0] m119_38;
   assign m119_38 =10'b0;

   // m119_39 = W*in
   wire signed [9:0] m119_39;
   assign m119_39 =10'b0;

   // m119_40 = W*in
   wire signed [9:0] m119_40;
   assign m119_40 =10'b0;

   // m119_41 = W*in
   wire signed [9:0] m119_41;
   assign m119_41 =10'b0;

   // m119_42 = W*in
   wire signed [9:0] m119_42;
   assign m119_42 =10'b0;

   // m119_43 = W*in
   wire signed [9:0] m119_43;
   assign m119_43 =10'b0;

   // m119_44 = W*in
   wire signed [9:0] m119_44;
   assign m119_44 =10'b0;

   // m119_45 = W*in
   wire signed [9:0] m119_45;
   assign m119_45 =10'b0;

   // m119_46 = W*in
   wire signed [9:0] m119_46;
   assign m119_46 =10'b0;

   // m119_47 = W*in
   wire signed [9:0] m119_47;
   assign m119_47 =10'b0;

   // m119_48 = W*in
   wire signed [9:0] m119_48;
   assign m119_48 =10'b0;

   // m119_49 = W*in
   wire signed [9:0] m119_49;
   assign m119_49 =10'b0;

   // m119_50 = W*in
   wire signed [9:0] m119_50;
   assign m119_50 =10'b0;

   // m119_51 = W*in
   wire signed [9:0] m119_51;
   assign m119_51 =10'b0;

   // m119_52 = W*in
   wire signed [9:0] m119_52;
   assign m119_52 =10'b0;

   // m119_53 = W*in
   wire signed [9:0] m119_53;
   assign m119_53 =10'b0;

   // m119_54 = W*in
   wire signed [9:0] m119_54;
   assign m119_54 =10'b0;

   // m119_55 = W*in
   wire signed [9:0] m119_55;
   assign m119_55 =10'b0;

   // m119_56 = W*in
   wire signed [9:0] m119_56;
   assign m119_56 =10'b0;

   // m119_57 = W*in
   wire signed [9:0] m119_57;
   assign m119_57 =10'b0;

   // m119_58 = W*in
   wire signed [9:0] m119_58;
   assign m119_58 =10'b0;

   // m119_59 = W*in
   wire signed [9:0] m119_59;
   assign m119_59 =10'b0;

   // m119_60 = W*in
   wire signed [9:0] m119_60;
   assign m119_60 =10'b0;

   // m119_61 = W*in
   wire signed [9:0] m119_61;
   assign m119_61 =10'b0;

   // m119_62 = W*in
   wire signed [9:0] m119_62;
   assign m119_62 =10'b0;

   // m119_63 = W*in
   wire signed [9:0] m119_63;
   assign m119_63 =10'b0;

   // m119_64 = W*in
   wire signed [9:0] m119_64;
   assign m119_64 =10'b0;

   // m119_65 = W*in
   wire signed [9:0] m119_65;
   assign m119_65 =10'b0;

   // m119_66 = W*in
   wire signed [9:0] m119_66;
   assign m119_66 =10'b0;

   // m119_67 = W*in
   wire signed [9:0] m119_67;
   assign m119_67 =10'b0;

   // m119_68 = W*in
   wire signed [9:0] m119_68;
   assign m119_68 =10'b0;

   // m119_69 = W*in
   wire signed [9:0] m119_69;
   assign m119_69 =10'b0;

   // m119_70 = W*in
   wire signed [9:0] m119_70;
   assign m119_70 ={ {5{in119[5]}} , in119[5:1] };

   // m119_71 = W*in
   wire signed [9:0] m119_71;
   assign m119_71 =10'b0;

   // m119_72 = W*in
   wire signed [9:0] m119_72;
   assign m119_72 =10'b0;

   // m119_73 = W*in
   wire signed [9:0] m119_73;
   assign m119_73 =10'b0;

   // m119_74 = W*in
   wire signed [9:0] m119_74;
   assign m119_74 =10'b0;

   // m119_75 = W*in
   wire signed [9:0] m119_75;
   assign m119_75 =10'b0;

   // m119_76 = W*in
   wire signed [9:0] m119_76;
   assign m119_76 =10'b0;

   // m119_77 = W*in
   wire signed [9:0] m119_77;
   assign m119_77 =10'b0;

   // m119_78 = W*in
   wire signed [9:0] m119_78;
   assign m119_78 =10'b0;

   // m119_79 = W*in
   wire signed [9:0] m119_79;
   assign m119_79 =10'b0;

   // m119_80 = W*in
   wire signed [9:0] m119_80;
   assign m119_80 =10'b0;

   // m119_81 = W*in
   wire signed [9:0] m119_81;
   assign m119_81 =10'b0;

   // m119_82 = W*in
   wire signed [9:0] m119_82;
   assign m119_82 ={ {5{in119[5]}} , in119[5:1] };

   // m119_83 = W*in
   wire signed [9:0] m119_83;
   assign m119_83 =10'b0;

   // m119_84 = W*in
   wire signed [9:0] m119_84;
   assign m119_84 =10'b0;

   // m119_85 = W*in
   wire signed [9:0] m119_85;
   assign m119_85 =10'b0;

   // m119_86 = W*in
   wire signed [9:0] m119_86;
   assign m119_86 =10'b0;

   // m119_87 = W*in
   wire signed [9:0] m119_87;
   assign m119_87 =10'b0;

   // m119_88 = W*in
   wire signed [9:0] m119_88;
   assign m119_88 =10'b0;

   // m119_89 = W*in
   wire signed [9:0] m119_89;
   assign m119_89 =10'b0;

   // m119_90 = W*in
   wire signed [9:0] m119_90;
   assign m119_90 =10'b0;

   // m119_91 = W*in
   wire signed [9:0] m119_91;
   assign m119_91 =10'b0;

   // m119_92 = W*in
   wire signed [9:0] m119_92;
   assign m119_92 =10'b0;

   // m119_93 = W*in
   wire signed [9:0] m119_93;
   assign m119_93 =10'b0;

   // m119_94 = W*in
   wire signed [9:0] m119_94;
   assign m119_94 =10'b0;

   // m119_95 = W*in
   wire signed [9:0] m119_95;
   assign m119_95 =10'b0;

   // m119_96 = W*in
   wire signed [9:0] m119_96;
   assign m119_96 =10'b0;

   // m119_97 = W*in
   wire signed [9:0] m119_97;
   assign m119_97 =10'b0;

   // m119_98 = W*in
   wire signed [9:0] m119_98;
   assign m119_98 =10'b0;

   // m119_99 = W*in
   wire signed [9:0] m119_99;
   assign m119_99 =10'b0;

   // m119_100 = W*in
   wire signed [9:0] m119_100;
   assign m119_100 =10'b0;

   // m119_101 = W*in
   wire signed [9:0] m119_101;
   assign m119_101 =10'b0;

   // m119_102 = W*in
   wire signed [9:0] m119_102;
   assign m119_102 =10'b0;

   // m119_103 = W*in
   wire signed [9:0] m119_103;
   assign m119_103 =10'b0;

   // m119_104 = W*in
   wire signed [9:0] m119_104;
   assign m119_104 =10'b0;

   // m119_105 = W*in
   wire signed [9:0] m119_105;
   assign m119_105 =10'b0;

   // m119_106 = W*in
   wire signed [9:0] m119_106;
   assign m119_106 =10'b0;

   // m119_107 = W*in
   wire signed [9:0] m119_107;
   assign m119_107 =10'b0;

   // m119_108 = W*in
   wire signed [9:0] m119_108;
   assign m119_108 =10'b0;

   // m119_109 = W*in
   wire signed [9:0] m119_109;
   assign m119_109 =10'b0;

   // m119_110 = W*in
   wire signed [9:0] m119_110;
   assign m119_110 =10'b0;

   // m119_111 = W*in
   wire signed [9:0] m119_111;
   assign m119_111 =10'b0;

   // m119_112 = W*in
   wire signed [9:0] m119_112;
   assign m119_112 =10'b0;

   // m119_113 = W*in
   wire signed [9:0] m119_113;
   assign m119_113 =10'b0;

   // m119_114 = W*in
   wire signed [9:0] m119_114;
   assign m119_114 =10'b0;

   // m119_115 = W*in
   wire signed [9:0] m119_115;
   assign m119_115 =10'b0;

   // m119_116 = W*in
   wire signed [9:0] m119_116;
   assign m119_116 =10'b0;

   // m119_117 = W*in
   wire signed [9:0] m119_117;
   assign m119_117 =10'b0;

   // m120_1 = W*in
   wire signed [9:0] m120_1;
   assign m120_1 =10'b0;

   // m120_2 = W*in
   wire signed [9:0] m120_2;
   assign m120_2 =10'b0;

   // m120_3 = W*in
   wire signed [9:0] m120_3;
   assign m120_3 =10'b0;

   // m120_4 = W*in
   wire signed [9:0] m120_4;
   assign m120_4 =10'b0;

   // m120_5 = W*in
   wire signed [9:0] m120_5;
   assign m120_5 =10'b0;

   // m120_6 = W*in
   wire signed [9:0] m120_6;
   assign m120_6 =10'b0;

   // m120_7 = W*in
   wire signed [9:0] m120_7;
   assign m120_7 =10'b0;

   // m120_8 = W*in
   wire signed [9:0] m120_8;
   assign m120_8 =10'b0;

   // m120_9 = W*in
   wire signed [9:0] m120_9;
   assign m120_9 =10'b0;

   // m120_10 = W*in
   wire signed [9:0] m120_10;
   assign m120_10 =10'b0;

   // m120_11 = W*in
   wire signed [9:0] m120_11;
   assign m120_11 =10'b0;

   // m120_12 = W*in
   wire signed [9:0] m120_12;
   assign m120_12 =10'b0;

   // m120_13 = W*in
   wire signed [9:0] m120_13;
   assign m120_13 =10'b0;

   // m120_14 = W*in
   wire signed [9:0] m120_14;
   assign m120_14 =10'b0;

   // m120_15 = W*in
   wire signed [9:0] m120_15;
   assign m120_15 =10'b0;

   // m120_16 = W*in
   wire signed [9:0] m120_16;
   assign m120_16 =10'b0;

   // m120_17 = W*in
   wire signed [9:0] m120_17;
   assign m120_17 =10'b0;

   // m120_18 = W*in
   wire signed [9:0] m120_18;
   assign m120_18 ={ {5{in120[5]}} , in120[5:1] };

   // m120_19 = W*in
   wire signed [9:0] m120_19;
   assign m120_19 ={ {5{in120[5]}} , in120[5:1] };

   // m120_20 = W*in
   wire signed [9:0] m120_20;
   assign m120_20 =10'b0;

   // m120_21 = W*in
   wire signed [9:0] m120_21;
   assign m120_21 ={ {5{in120[5]}} , in120[5:1] };

   // m120_22 = W*in
   wire signed [9:0] m120_22;
   assign m120_22 ={ {5{neg120[5]}} , neg120[5:1] };

   // m120_23 = W*in
   wire signed [9:0] m120_23;
   assign m120_23 ={ {5{neg120[5]}} , neg120[5:1] };

   // m120_24 = W*in
   wire signed [9:0] m120_24;
   assign m120_24 =10'b0;

   // m120_25 = W*in
   wire signed [9:0] m120_25;
   assign m120_25 =10'b0;

   // m120_26 = W*in
   wire signed [9:0] m120_26;
   assign m120_26 ={ {5{in120[5]}} , in120[5:1] };

   // m120_27 = W*in
   wire signed [9:0] m120_27;
   assign m120_27 =10'b0;

   // m120_28 = W*in
   wire signed [9:0] m120_28;
   assign m120_28 =10'b0;

   // m120_29 = W*in
   wire signed [9:0] m120_29;
   assign m120_29 =10'b0;

   // m120_30 = W*in
   wire signed [9:0] m120_30;
   assign m120_30 =10'b0;

   // m120_31 = W*in
   wire signed [9:0] m120_31;
   assign m120_31 =10'b0;

   // m120_32 = W*in
   wire signed [9:0] m120_32;
   assign m120_32 =10'b0;

   // m120_33 = W*in
   wire signed [9:0] m120_33;
   assign m120_33 =10'b0;

   // m120_34 = W*in
   wire signed [9:0] m120_34;
   assign m120_34 =10'b0;

   // m120_35 = W*in
   wire signed [9:0] m120_35;
   assign m120_35 =10'b0;

   // m120_36 = W*in
   wire signed [9:0] m120_36;
   assign m120_36 ={ {5{neg120[5]}} , neg120[5:1] };

   // m120_37 = W*in
   wire signed [9:0] m120_37;
   assign m120_37 ={ {4{neg120[5]}} , neg120[5:0] };

   // m120_38 = W*in
   wire signed [9:0] m120_38;
   assign m120_38 =10'b0;

   // m120_39 = W*in
   wire signed [9:0] m120_39;
   assign m120_39 =10'b0;

   // m120_40 = W*in
   wire signed [9:0] m120_40;
   assign m120_40 =10'b0;

   // m120_41 = W*in
   wire signed [9:0] m120_41;
   assign m120_41 =10'b0;

   // m120_42 = W*in
   wire signed [9:0] m120_42;
   assign m120_42 =10'b0;

   // m120_43 = W*in
   wire signed [9:0] m120_43;
   assign m120_43 =10'b0;

   // m120_44 = W*in
   wire signed [9:0] m120_44;
   assign m120_44 =10'b0;

   // m120_45 = W*in
   wire signed [9:0] m120_45;
   assign m120_45 =10'b0;

   // m120_46 = W*in
   wire signed [9:0] m120_46;
   assign m120_46 =10'b0;

   // m120_47 = W*in
   wire signed [9:0] m120_47;
   assign m120_47 =10'b0;

   // m120_48 = W*in
   wire signed [9:0] m120_48;
   assign m120_48 =10'b0;

   // m120_49 = W*in
   wire signed [9:0] m120_49;
   assign m120_49 =10'b0;

   // m120_50 = W*in
   wire signed [9:0] m120_50;
   assign m120_50 =10'b0;

   // m120_51 = W*in
   wire signed [9:0] m120_51;
   assign m120_51 =10'b0;

   // m120_52 = W*in
   wire signed [9:0] m120_52;
   assign m120_52 =10'b0;

   // m120_53 = W*in
   wire signed [9:0] m120_53;
   assign m120_53 =10'b0;

   // m120_54 = W*in
   wire signed [9:0] m120_54;
   assign m120_54 =10'b0;

   // m120_55 = W*in
   wire signed [9:0] m120_55;
   assign m120_55 =10'b0;

   // m120_56 = W*in
   wire signed [9:0] m120_56;
   assign m120_56 =10'b0;

   // m120_57 = W*in
   wire signed [9:0] m120_57;
   assign m120_57 =10'b0;

   // m120_58 = W*in
   wire signed [9:0] m120_58;
   assign m120_58 =10'b0;

   // m120_59 = W*in
   wire signed [9:0] m120_59;
   assign m120_59 =10'b0;

   // m120_60 = W*in
   wire signed [9:0] m120_60;
   assign m120_60 =10'b0;

   // m120_61 = W*in
   wire signed [9:0] m120_61;
   assign m120_61 =10'b0;

   // m120_62 = W*in
   wire signed [9:0] m120_62;
   assign m120_62 =10'b0;

   // m120_63 = W*in
   wire signed [9:0] m120_63;
   assign m120_63 =10'b0;

   // m120_64 = W*in
   wire signed [9:0] m120_64;
   assign m120_64 =10'b0;

   // m120_65 = W*in
   wire signed [9:0] m120_65;
   assign m120_65 =10'b0;

   // m120_66 = W*in
   wire signed [9:0] m120_66;
   assign m120_66 =10'b0;

   // m120_67 = W*in
   wire signed [9:0] m120_67;
   assign m120_67 =10'b0;

   // m120_68 = W*in
   wire signed [9:0] m120_68;
   assign m120_68 =10'b0;

   // m120_69 = W*in
   wire signed [9:0] m120_69;
   assign m120_69 =10'b0;

   // m120_70 = W*in
   wire signed [9:0] m120_70;
   assign m120_70 =10'b0;

   // m120_71 = W*in
   wire signed [9:0] m120_71;
   assign m120_71 =10'b0;

   // m120_72 = W*in
   wire signed [9:0] m120_72;
   assign m120_72 =10'b0;

   // m120_73 = W*in
   wire signed [9:0] m120_73;
   assign m120_73 =10'b0;

   // m120_74 = W*in
   wire signed [9:0] m120_74;
   assign m120_74 =10'b0;

   // m120_75 = W*in
   wire signed [9:0] m120_75;
   assign m120_75 =10'b0;

   // m120_76 = W*in
   wire signed [9:0] m120_76;
   assign m120_76 =10'b0;

   // m120_77 = W*in
   wire signed [9:0] m120_77;
   assign m120_77 =10'b0;

   // m120_78 = W*in
   wire signed [9:0] m120_78;
   assign m120_78 =10'b0;

   // m120_79 = W*in
   wire signed [9:0] m120_79;
   assign m120_79 =10'b0;

   // m120_80 = W*in
   wire signed [9:0] m120_80;
   assign m120_80 =10'b0;

   // m120_81 = W*in
   wire signed [9:0] m120_81;
   assign m120_81 =10'b0;

   // m120_82 = W*in
   wire signed [9:0] m120_82;
   assign m120_82 ={ {5{neg120[5]}} , neg120[5:1] };

   // m120_83 = W*in
   wire signed [9:0] m120_83;
   assign m120_83 ={ {5{neg120[5]}} , neg120[5:1] };

   // m120_84 = W*in
   wire signed [9:0] m120_84;
   assign m120_84 =10'b0;

   // m120_85 = W*in
   wire signed [9:0] m120_85;
   assign m120_85 =10'b0;

   // m120_86 = W*in
   wire signed [9:0] m120_86;
   assign m120_86 =10'b0;

   // m120_87 = W*in
   wire signed [9:0] m120_87;
   assign m120_87 =10'b0;

   // m120_88 = W*in
   wire signed [9:0] m120_88;
   assign m120_88 =10'b0;

   // m120_89 = W*in
   wire signed [9:0] m120_89;
   assign m120_89 =10'b0;

   // m120_90 = W*in
   wire signed [9:0] m120_90;
   assign m120_90 =10'b0;

   // m120_91 = W*in
   wire signed [9:0] m120_91;
   assign m120_91 =10'b0;

   // m120_92 = W*in
   wire signed [9:0] m120_92;
   assign m120_92 =10'b0;

   // m120_93 = W*in
   wire signed [9:0] m120_93;
   assign m120_93 =10'b0;

   // m120_94 = W*in
   wire signed [9:0] m120_94;
   assign m120_94 =10'b0;

   // m120_95 = W*in
   wire signed [9:0] m120_95;
   assign m120_95 =10'b0;

   // m120_96 = W*in
   wire signed [9:0] m120_96;
   assign m120_96 =10'b0;

   // m120_97 = W*in
   wire signed [9:0] m120_97;
   assign m120_97 =10'b0;

   // m120_98 = W*in
   wire signed [9:0] m120_98;
   assign m120_98 =10'b0;

   // m120_99 = W*in
   wire signed [9:0] m120_99;
   assign m120_99 =10'b0;

   // m120_100 = W*in
   wire signed [9:0] m120_100;
   assign m120_100 =10'b0;

   // m120_101 = W*in
   wire signed [9:0] m120_101;
   assign m120_101 =10'b0;

   // m120_102 = W*in
   wire signed [9:0] m120_102;
   assign m120_102 =10'b0;

   // m120_103 = W*in
   wire signed [9:0] m120_103;
   assign m120_103 =10'b0;

   // m120_104 = W*in
   wire signed [9:0] m120_104;
   assign m120_104 =10'b0;

   // m120_105 = W*in
   wire signed [9:0] m120_105;
   assign m120_105 =10'b0;

   // m120_106 = W*in
   wire signed [9:0] m120_106;
   assign m120_106 =10'b0;

   // m120_107 = W*in
   wire signed [9:0] m120_107;
   assign m120_107 =10'b0;

   // m120_108 = W*in
   wire signed [9:0] m120_108;
   assign m120_108 ={ {5{neg120[5]}} , neg120[5:1] };

   // m120_109 = W*in
   wire signed [9:0] m120_109;
   assign m120_109 ={ {4{neg120[5]}} , neg120[5:0] };

   // m120_110 = W*in
   wire signed [9:0] m120_110;
   assign m120_110 =10'b0;

   // m120_111 = W*in
   wire signed [9:0] m120_111;
   assign m120_111 =10'b0;

   // m120_112 = W*in
   wire signed [9:0] m120_112;
   assign m120_112 =10'b0;

   // m120_113 = W*in
   wire signed [9:0] m120_113;
   assign m120_113 =10'b0;

   // m120_114 = W*in
   wire signed [9:0] m120_114;
   assign m120_114 =10'b0;

   // m120_115 = W*in
   wire signed [9:0] m120_115;
   assign m120_115 =10'b0;

   // m120_116 = W*in
   wire signed [9:0] m120_116;
   assign m120_116 =10'b0;

   // m120_117 = W*in
   wire signed [9:0] m120_117;
   assign m120_117 =10'b0;

   // m121_1 = W*in
   wire signed [9:0] m121_1;
   assign m121_1 ={ {3{neg121[5]}} , neg121 , {1{1'b0}} };

   // m121_2 = W*in
   wire signed [9:0] m121_2;
   assign m121_2 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_3 = W*in
   wire signed [9:0] m121_3;
   assign m121_3 =10'b0;

   // m121_4 = W*in
   wire signed [9:0] m121_4;
   assign m121_4 =10'b0;

   // m121_5 = W*in
   wire signed [9:0] m121_5;
   assign m121_5 =10'b0;

   // m121_6 = W*in
   wire signed [9:0] m121_6;
   assign m121_6 =10'b0;

   // m121_7 = W*in
   wire signed [9:0] m121_7;
   assign m121_7 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_8 = W*in
   wire signed [9:0] m121_8;
   assign m121_8 =10'b0;

   // m121_9 = W*in
   wire signed [9:0] m121_9;
   assign m121_9 =10'b0;

   // m121_10 = W*in
   wire signed [9:0] m121_10;
   assign m121_10 =10'b0;

   // m121_11 = W*in
   wire signed [9:0] m121_11;
   assign m121_11 =10'b0;

   // m121_12 = W*in
   wire signed [9:0] m121_12;
   assign m121_12 =10'b0;

   // m121_13 = W*in
   wire signed [9:0] m121_13;
   assign m121_13 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_14 = W*in
   wire signed [9:0] m121_14;
   assign m121_14 =10'b0;

   // m121_15 = W*in
   wire signed [9:0] m121_15;
   assign m121_15 ={ {4{in121[5]}} , in121[5:0] };

   // m121_16 = W*in
   wire signed [9:0] m121_16;
   assign m121_16 ={ {3{neg121[5]}} , neg121 , {1{1'b0}} };

   // m121_17 = W*in
   wire signed [9:0] m121_17;
   assign m121_17 =10'b0;

   // m121_18 = W*in
   wire signed [9:0] m121_18;
   assign m121_18 ={ {5{in121[5]}} , in121[5:1] };

   // m121_19 = W*in
   wire signed [9:0] m121_19;
   assign m121_19 =10'b0;

   // m121_20 = W*in
   wire signed [9:0] m121_20;
   assign m121_20 =10'b0;

   // m121_21 = W*in
   wire signed [9:0] m121_21;
   assign m121_21 ={ {4{in121[5]}} , in121[5:0] };

   // m121_22 = W*in
   wire signed [9:0] m121_22;
   assign m121_22 =10'b0;

   // m121_23 = W*in
   wire signed [9:0] m121_23;
   assign m121_23 =10'b0;

   // m121_24 = W*in
   wire signed [9:0] m121_24;
   assign m121_24 =10'b0;

   // m121_25 = W*in
   wire signed [9:0] m121_25;
   assign m121_25 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_26 = W*in
   wire signed [9:0] m121_26;
   assign m121_26 =10'b0;

   // m121_27 = W*in
   wire signed [9:0] m121_27;
   assign m121_27 ={ {5{in121[5]}} , in121[5:1] };

   // m121_28 = W*in
   wire signed [9:0] m121_28;
   assign m121_28 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_29 = W*in
   wire signed [9:0] m121_29;
   assign m121_29 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_30 = W*in
   wire signed [9:0] m121_30;
   assign m121_30 =10'b0;

   // m121_31 = W*in
   wire signed [9:0] m121_31;
   assign m121_31 =10'b0;

   // m121_32 = W*in
   wire signed [9:0] m121_32;
   assign m121_32 =10'b0;

   // m121_33 = W*in
   wire signed [9:0] m121_33;
   assign m121_33 ={ {3{neg121[5]}} , neg121 , {1{1'b0}} };

   // m121_34 = W*in
   wire signed [9:0] m121_34;
   assign m121_34 =10'b0;

   // m121_35 = W*in
   wire signed [9:0] m121_35;
   assign m121_35 =10'b0;

   // m121_36 = W*in
   wire signed [9:0] m121_36;
   assign m121_36 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_37 = W*in
   wire signed [9:0] m121_37;
   assign m121_37 =10'b0;

   // m121_38 = W*in
   wire signed [9:0] m121_38;
   assign m121_38 ={ {3{in121[5]}} , in121 , {1{1'b0}} };

   // m121_39 = W*in
   wire signed [9:0] m121_39;
   assign m121_39 =10'b0;

   // m121_40 = W*in
   wire signed [9:0] m121_40;
   assign m121_40 =10'b0;

   // m121_41 = W*in
   wire signed [9:0] m121_41;
   assign m121_41 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_42 = W*in
   wire signed [9:0] m121_42;
   assign m121_42 =10'b0;

   // m121_43 = W*in
   wire signed [9:0] m121_43;
   assign m121_43 =10'b0;

   // m121_44 = W*in
   wire signed [9:0] m121_44;
   assign m121_44 =10'b0;

   // m121_45 = W*in
   wire signed [9:0] m121_45;
   assign m121_45 ={ {3{neg121[5]}} , neg121 , {1{1'b0}} };

   // m121_46 = W*in
   wire signed [9:0] m121_46;
   assign m121_46 =10'b0;

   // m121_47 = W*in
   wire signed [9:0] m121_47;
   assign m121_47 =10'b0;

   // m121_48 = W*in
   wire signed [9:0] m121_48;
   assign m121_48 =10'b0;

   // m121_49 = W*in
   wire signed [9:0] m121_49;
   assign m121_49 =10'b0;

   // m121_50 = W*in
   wire signed [9:0] m121_50;
   assign m121_50 =10'b0;

   // m121_51 = W*in
   wire signed [9:0] m121_51;
   assign m121_51 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_52 = W*in
   wire signed [9:0] m121_52;
   assign m121_52 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_53 = W*in
   wire signed [9:0] m121_53;
   assign m121_53 =10'b0;

   // m121_54 = W*in
   wire signed [9:0] m121_54;
   assign m121_54 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_55 = W*in
   wire signed [9:0] m121_55;
   assign m121_55 =10'b0;

   // m121_56 = W*in
   wire signed [9:0] m121_56;
   assign m121_56 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_57 = W*in
   wire signed [9:0] m121_57;
   assign m121_57 =10'b0;

   // m121_58 = W*in
   wire signed [9:0] m121_58;
   assign m121_58 =10'b0;

   // m121_59 = W*in
   wire signed [9:0] m121_59;
   assign m121_59 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_60 = W*in
   wire signed [9:0] m121_60;
   assign m121_60 =10'b0;

   // m121_61 = W*in
   wire signed [9:0] m121_61;
   assign m121_61 =10'b0;

   // m121_62 = W*in
   wire signed [9:0] m121_62;
   assign m121_62 =10'b0;

   // m121_63 = W*in
   wire signed [9:0] m121_63;
   assign m121_63 =10'b0;

   // m121_64 = W*in
   wire signed [9:0] m121_64;
   assign m121_64 =10'b0;

   // m121_65 = W*in
   wire signed [9:0] m121_65;
   assign m121_65 =10'b0;

   // m121_66 = W*in
   wire signed [9:0] m121_66;
   assign m121_66 =10'b0;

   // m121_67 = W*in
   wire signed [9:0] m121_67;
   assign m121_67 =10'b0;

   // m121_68 = W*in
   wire signed [9:0] m121_68;
   assign m121_68 =10'b0;

   // m121_69 = W*in
   wire signed [9:0] m121_69;
   assign m121_69 =10'b0;

   // m121_70 = W*in
   wire signed [9:0] m121_70;
   assign m121_70 ={ {4{in121[5]}} , in121[5:0] };

   // m121_71 = W*in
   wire signed [9:0] m121_71;
   assign m121_71 ={ {4{in121[5]}} , in121[5:0] };

   // m121_72 = W*in
   wire signed [9:0] m121_72;
   assign m121_72 ={ {5{in121[5]}} , in121[5:1] };

   // m121_73 = W*in
   wire signed [9:0] m121_73;
   assign m121_73 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_74 = W*in
   wire signed [9:0] m121_74;
   assign m121_74 ={ {4{in121[5]}} , in121[5:0] };

   // m121_75 = W*in
   wire signed [9:0] m121_75;
   assign m121_75 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_76 = W*in
   wire signed [9:0] m121_76;
   assign m121_76 =10'b0;

   // m121_77 = W*in
   wire signed [9:0] m121_77;
   assign m121_77 =10'b0;

   // m121_78 = W*in
   wire signed [9:0] m121_78;
   assign m121_78 =10'b0;

   // m121_79 = W*in
   wire signed [9:0] m121_79;
   assign m121_79 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_80 = W*in
   wire signed [9:0] m121_80;
   assign m121_80 =10'b0;

   // m121_81 = W*in
   wire signed [9:0] m121_81;
   assign m121_81 =10'b0;

   // m121_82 = W*in
   wire signed [9:0] m121_82;
   assign m121_82 =10'b0;

   // m121_83 = W*in
   wire signed [9:0] m121_83;
   assign m121_83 ={ {5{neg121[5]}} , neg121[5:1] };

   // m121_84 = W*in
   wire signed [9:0] m121_84;
   assign m121_84 =10'b0;

   // m121_85 = W*in
   wire signed [9:0] m121_85;
   assign m121_85 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_86 = W*in
   wire signed [9:0] m121_86;
   assign m121_86 ={ {4{in121[5]}} , in121[5:0] };

   // m121_87 = W*in
   wire signed [9:0] m121_87;
   assign m121_87 ={ {4{in121[5]}} , in121[5:0] };

   // m121_88 = W*in
   wire signed [9:0] m121_88;
   assign m121_88 =10'b0;

   // m121_89 = W*in
   wire signed [9:0] m121_89;
   assign m121_89 =10'b0;

   // m121_90 = W*in
   wire signed [9:0] m121_90;
   assign m121_90 =10'b0;

   // m121_91 = W*in
   wire signed [9:0] m121_91;
   assign m121_91 =10'b0;

   // m121_92 = W*in
   wire signed [9:0] m121_92;
   assign m121_92 ={ {4{in121[5]}} , in121[5:0] };

   // m121_93 = W*in
   wire signed [9:0] m121_93;
   assign m121_93 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_94 = W*in
   wire signed [9:0] m121_94;
   assign m121_94 =10'b0;

   // m121_95 = W*in
   wire signed [9:0] m121_95;
   assign m121_95 =10'b0;

   // m121_96 = W*in
   wire signed [9:0] m121_96;
   assign m121_96 =10'b0;

   // m121_97 = W*in
   wire signed [9:0] m121_97;
   assign m121_97 ={ {4{in121[5]}} , in121[5:0] };

   // m121_98 = W*in
   wire signed [9:0] m121_98;
   assign m121_98 =10'b0;

   // m121_99 = W*in
   wire signed [9:0] m121_99;
   assign m121_99 =10'b0;

   // m121_100 = W*in
   wire signed [9:0] m121_100;
   assign m121_100 =10'b0;

   // m121_101 = W*in
   wire signed [9:0] m121_101;
   assign m121_101 =10'b0;

   // m121_102 = W*in
   wire signed [9:0] m121_102;
   assign m121_102 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_103 = W*in
   wire signed [9:0] m121_103;
   assign m121_103 =10'b0;

   // m121_104 = W*in
   wire signed [9:0] m121_104;
   assign m121_104 =10'b0;

   // m121_105 = W*in
   wire signed [9:0] m121_105;
   assign m121_105 =10'b0;

   // m121_106 = W*in
   wire signed [9:0] m121_106;
   assign m121_106 ={ {5{neg121[5]}} , neg121[5:1] };

   // m121_107 = W*in
   wire signed [9:0] m121_107;
   assign m121_107 =10'b0;

   // m121_108 = W*in
   wire signed [9:0] m121_108;
   assign m121_108 =10'b0;

   // m121_109 = W*in
   wire signed [9:0] m121_109;
   assign m121_109 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_110 = W*in
   wire signed [9:0] m121_110;
   assign m121_110 =10'b0;

   // m121_111 = W*in
   wire signed [9:0] m121_111;
   assign m121_111 ={ {4{neg121[5]}} , neg121[5:0] };

   // m121_112 = W*in
   wire signed [9:0] m121_112;
   assign m121_112 =10'b0;

   // m121_113 = W*in
   wire signed [9:0] m121_113;
   assign m121_113 ={ {5{neg121[5]}} , neg121[5:1] };

   // m121_114 = W*in
   wire signed [9:0] m121_114;
   assign m121_114 =10'b0;

   // m121_115 = W*in
   wire signed [9:0] m121_115;
   assign m121_115 =10'b0;

   // m121_116 = W*in
   wire signed [9:0] m121_116;
   assign m121_116 =10'b0;

   // m121_117 = W*in
   wire signed [9:0] m121_117;
   assign m121_117 =10'b0;

   // m122_1 = W*in
   wire signed [9:0] m122_1;
   assign m122_1 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_2 = W*in
   wire signed [9:0] m122_2;
   assign m122_2 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_3 = W*in
   wire signed [9:0] m122_3;
   assign m122_3 =10'b0;

   // m122_4 = W*in
   wire signed [9:0] m122_4;
   assign m122_4 =10'b0;

   // m122_5 = W*in
   wire signed [9:0] m122_5;
   assign m122_5 =10'b0;

   // m122_6 = W*in
   wire signed [9:0] m122_6;
   assign m122_6 =10'b0;

   // m122_7 = W*in
   wire signed [9:0] m122_7;
   assign m122_7 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_8 = W*in
   wire signed [9:0] m122_8;
   assign m122_8 =10'b0;

   // m122_9 = W*in
   wire signed [9:0] m122_9;
   assign m122_9 =10'b0;

   // m122_10 = W*in
   wire signed [9:0] m122_10;
   assign m122_10 =10'b0;

   // m122_11 = W*in
   wire signed [9:0] m122_11;
   assign m122_11 =10'b0;

   // m122_12 = W*in
   wire signed [9:0] m122_12;
   assign m122_12 ={ {4{in122[5]}} , in122[5:0] };

   // m122_13 = W*in
   wire signed [9:0] m122_13;
   assign m122_13 =10'b0;

   // m122_14 = W*in
   wire signed [9:0] m122_14;
   assign m122_14 =10'b0;

   // m122_15 = W*in
   wire signed [9:0] m122_15;
   assign m122_15 ={ {4{in122[5]}} , in122[5:0] };

   // m122_16 = W*in
   wire signed [9:0] m122_16;
   assign m122_16 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_17 = W*in
   wire signed [9:0] m122_17;
   assign m122_17 =10'b0;

   // m122_18 = W*in
   wire signed [9:0] m122_18;
   assign m122_18 ={ {4{in122[5]}} , in122[5:0] };

   // m122_19 = W*in
   wire signed [9:0] m122_19;
   assign m122_19 =10'b0;

   // m122_20 = W*in
   wire signed [9:0] m122_20;
   assign m122_20 =10'b0;

   // m122_21 = W*in
   wire signed [9:0] m122_21;
   assign m122_21 =10'b0;

   // m122_22 = W*in
   wire signed [9:0] m122_22;
   assign m122_22 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_23 = W*in
   wire signed [9:0] m122_23;
   assign m122_23 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_24 = W*in
   wire signed [9:0] m122_24;
   assign m122_24 =10'b0;

   // m122_25 = W*in
   wire signed [9:0] m122_25;
   assign m122_25 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_26 = W*in
   wire signed [9:0] m122_26;
   assign m122_26 =10'b0;

   // m122_27 = W*in
   wire signed [9:0] m122_27;
   assign m122_27 =10'b0;

   // m122_28 = W*in
   wire signed [9:0] m122_28;
   assign m122_28 =10'b0;

   // m122_29 = W*in
   wire signed [9:0] m122_29;
   assign m122_29 ={ {5{neg122[5]}} , neg122[5:1] };

   // m122_30 = W*in
   wire signed [9:0] m122_30;
   assign m122_30 =10'b0;

   // m122_31 = W*in
   wire signed [9:0] m122_31;
   assign m122_31 ={ {5{neg122[5]}} , neg122[5:1] };

   // m122_32 = W*in
   wire signed [9:0] m122_32;
   assign m122_32 =10'b0;

   // m122_33 = W*in
   wire signed [9:0] m122_33;
   assign m122_33 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_34 = W*in
   wire signed [9:0] m122_34;
   assign m122_34 =10'b0;

   // m122_35 = W*in
   wire signed [9:0] m122_35;
   assign m122_35 =10'b0;

   // m122_36 = W*in
   wire signed [9:0] m122_36;
   assign m122_36 =10'b0;

   // m122_37 = W*in
   wire signed [9:0] m122_37;
   assign m122_37 =10'b0;

   // m122_38 = W*in
   wire signed [9:0] m122_38;
   assign m122_38 =10'b0;

   // m122_39 = W*in
   wire signed [9:0] m122_39;
   assign m122_39 =10'b0;

   // m122_40 = W*in
   wire signed [9:0] m122_40;
   assign m122_40 =10'b0;

   // m122_41 = W*in
   wire signed [9:0] m122_41;
   assign m122_41 =10'b0;

   // m122_42 = W*in
   wire signed [9:0] m122_42;
   assign m122_42 =10'b0;

   // m122_43 = W*in
   wire signed [9:0] m122_43;
   assign m122_43 ={ {4{in122[5]}} , in122[5:0] };

   // m122_44 = W*in
   wire signed [9:0] m122_44;
   assign m122_44 =10'b0;

   // m122_45 = W*in
   wire signed [9:0] m122_45;
   assign m122_45 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_46 = W*in
   wire signed [9:0] m122_46;
   assign m122_46 ={ {4{in122[5]}} , in122[5:0] };

   // m122_47 = W*in
   wire signed [9:0] m122_47;
   assign m122_47 ={ {5{neg122[5]}} , neg122[5:1] };

   // m122_48 = W*in
   wire signed [9:0] m122_48;
   assign m122_48 =10'b0;

   // m122_49 = W*in
   wire signed [9:0] m122_49;
   assign m122_49 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_50 = W*in
   wire signed [9:0] m122_50;
   assign m122_50 =10'b0;

   // m122_51 = W*in
   wire signed [9:0] m122_51;
   assign m122_51 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_52 = W*in
   wire signed [9:0] m122_52;
   assign m122_52 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_53 = W*in
   wire signed [9:0] m122_53;
   assign m122_53 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_54 = W*in
   wire signed [9:0] m122_54;
   assign m122_54 =10'b0;

   // m122_55 = W*in
   wire signed [9:0] m122_55;
   assign m122_55 =10'b0;

   // m122_56 = W*in
   wire signed [9:0] m122_56;
   assign m122_56 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_57 = W*in
   wire signed [9:0] m122_57;
   assign m122_57 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_58 = W*in
   wire signed [9:0] m122_58;
   assign m122_58 =10'b0;

   // m122_59 = W*in
   wire signed [9:0] m122_59;
   assign m122_59 =10'b0;

   // m122_60 = W*in
   wire signed [9:0] m122_60;
   assign m122_60 ={ {4{in122[5]}} , in122[5:0] };

   // m122_61 = W*in
   wire signed [9:0] m122_61;
   assign m122_61 =10'b0;

   // m122_62 = W*in
   wire signed [9:0] m122_62;
   assign m122_62 =10'b0;

   // m122_63 = W*in
   wire signed [9:0] m122_63;
   assign m122_63 ={ {4{in122[5]}} , in122[5:0] };

   // m122_64 = W*in
   wire signed [9:0] m122_64;
   assign m122_64 =10'b0;

   // m122_65 = W*in
   wire signed [9:0] m122_65;
   assign m122_65 =10'b0;

   // m122_66 = W*in
   wire signed [9:0] m122_66;
   assign m122_66 ={ {4{in122[5]}} , in122[5:0] };

   // m122_67 = W*in
   wire signed [9:0] m122_67;
   assign m122_67 =10'b0;

   // m122_68 = W*in
   wire signed [9:0] m122_68;
   assign m122_68 =10'b0;

   // m122_69 = W*in
   wire signed [9:0] m122_69;
   assign m122_69 =10'b0;

   // m122_70 = W*in
   wire signed [9:0] m122_70;
   assign m122_70 ={ {5{in122[5]}} , in122[5:1] };

   // m122_71 = W*in
   wire signed [9:0] m122_71;
   assign m122_71 =10'b0;

   // m122_72 = W*in
   wire signed [9:0] m122_72;
   assign m122_72 =10'b0;

   // m122_73 = W*in
   wire signed [9:0] m122_73;
   assign m122_73 =10'b0;

   // m122_74 = W*in
   wire signed [9:0] m122_74;
   assign m122_74 ={ {4{in122[5]}} , in122[5:0] };

   // m122_75 = W*in
   wire signed [9:0] m122_75;
   assign m122_75 =10'b0;

   // m122_76 = W*in
   wire signed [9:0] m122_76;
   assign m122_76 =10'b0;

   // m122_77 = W*in
   wire signed [9:0] m122_77;
   assign m122_77 =10'b0;

   // m122_78 = W*in
   wire signed [9:0] m122_78;
   assign m122_78 =10'b0;

   // m122_79 = W*in
   wire signed [9:0] m122_79;
   assign m122_79 =10'b0;

   // m122_80 = W*in
   wire signed [9:0] m122_80;
   assign m122_80 =10'b0;

   // m122_81 = W*in
   wire signed [9:0] m122_81;
   assign m122_81 =10'b0;

   // m122_82 = W*in
   wire signed [9:0] m122_82;
   assign m122_82 =10'b0;

   // m122_83 = W*in
   wire signed [9:0] m122_83;
   assign m122_83 =10'b0;

   // m122_84 = W*in
   wire signed [9:0] m122_84;
   assign m122_84 =10'b0;

   // m122_85 = W*in
   wire signed [9:0] m122_85;
   assign m122_85 ={ {5{neg122[5]}} , neg122[5:1] };

   // m122_86 = W*in
   wire signed [9:0] m122_86;
   assign m122_86 ={ {4{in122[5]}} , in122[5:0] };

   // m122_87 = W*in
   wire signed [9:0] m122_87;
   assign m122_87 =10'b0;

   // m122_88 = W*in
   wire signed [9:0] m122_88;
   assign m122_88 ={ {4{in122[5]}} , in122[5:0] };

   // m122_89 = W*in
   wire signed [9:0] m122_89;
   assign m122_89 =10'b0;

   // m122_90 = W*in
   wire signed [9:0] m122_90;
   assign m122_90 =10'b0;

   // m122_91 = W*in
   wire signed [9:0] m122_91;
   assign m122_91 =10'b0;

   // m122_92 = W*in
   wire signed [9:0] m122_92;
   assign m122_92 ={ {4{in122[5]}} , in122[5:0] };

   // m122_93 = W*in
   wire signed [9:0] m122_93;
   assign m122_93 =10'b0;

   // m122_94 = W*in
   wire signed [9:0] m122_94;
   assign m122_94 ={ {4{in122[5]}} , in122[5:0] };

   // m122_95 = W*in
   wire signed [9:0] m122_95;
   assign m122_95 =10'b0;

   // m122_96 = W*in
   wire signed [9:0] m122_96;
   assign m122_96 =10'b0;

   // m122_97 = W*in
   wire signed [9:0] m122_97;
   assign m122_97 ={ {4{in122[5]}} , in122[5:0] };

   // m122_98 = W*in
   wire signed [9:0] m122_98;
   assign m122_98 =10'b0;

   // m122_99 = W*in
   wire signed [9:0] m122_99;
   assign m122_99 ={ {4{in122[5]}} , in122[5:0] };

   // m122_100 = W*in
   wire signed [9:0] m122_100;
   assign m122_100 ={ {4{in122[5]}} , in122[5:0] };

   // m122_101 = W*in
   wire signed [9:0] m122_101;
   assign m122_101 ={ {5{in122[5]}} , in122[5:1] };

   // m122_102 = W*in
   wire signed [9:0] m122_102;
   assign m122_102 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_103 = W*in
   wire signed [9:0] m122_103;
   assign m122_103 =10'b0;

   // m122_104 = W*in
   wire signed [9:0] m122_104;
   assign m122_104 ={ {4{in122[5]}} , in122[5:0] };

   // m122_105 = W*in
   wire signed [9:0] m122_105;
   assign m122_105 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_106 = W*in
   wire signed [9:0] m122_106;
   assign m122_106 ={ {4{neg122[5]}} , neg122[5:0] };

   // m122_107 = W*in
   wire signed [9:0] m122_107;
   assign m122_107 =10'b0;

   // m122_108 = W*in
   wire signed [9:0] m122_108;
   assign m122_108 =10'b0;

   // m122_109 = W*in
   wire signed [9:0] m122_109;
   assign m122_109 =10'b0;

   // m122_110 = W*in
   wire signed [9:0] m122_110;
   assign m122_110 =10'b0;

   // m122_111 = W*in
   wire signed [9:0] m122_111;
   assign m122_111 =10'b0;

   // m122_112 = W*in
   wire signed [9:0] m122_112;
   assign m122_112 ={ {4{in122[5]}} , in122[5:0] };

   // m122_113 = W*in
   wire signed [9:0] m122_113;
   assign m122_113 ={ {4{in122[5]}} , in122[5:0] };

   // m122_114 = W*in
   wire signed [9:0] m122_114;
   assign m122_114 ={ {5{neg122[5]}} , neg122[5:1] };

   // m122_115 = W*in
   wire signed [9:0] m122_115;
   assign m122_115 =10'b0;

   // m122_116 = W*in
   wire signed [9:0] m122_116;
   assign m122_116 =10'b0;

   // m122_117 = W*in
   wire signed [9:0] m122_117;
   assign m122_117 =10'b0;

   // m123_1 = W*in
   wire signed [9:0] m123_1;
   assign m123_1 =10'b0;

   // m123_2 = W*in
   wire signed [9:0] m123_2;
   assign m123_2 =10'b0;

   // m123_3 = W*in
   wire signed [9:0] m123_3;
   assign m123_3 =10'b0;

   // m123_4 = W*in
   wire signed [9:0] m123_4;
   assign m123_4 =10'b0;

   // m123_5 = W*in
   wire signed [9:0] m123_5;
   assign m123_5 =10'b0;

   // m123_6 = W*in
   wire signed [9:0] m123_6;
   assign m123_6 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_7 = W*in
   wire signed [9:0] m123_7;
   assign m123_7 =10'b0;

   // m123_8 = W*in
   wire signed [9:0] m123_8;
   assign m123_8 =10'b0;

   // m123_9 = W*in
   wire signed [9:0] m123_9;
   assign m123_9 =10'b0;

   // m123_10 = W*in
   wire signed [9:0] m123_10;
   assign m123_10 =10'b0;

   // m123_11 = W*in
   wire signed [9:0] m123_11;
   assign m123_11 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_12 = W*in
   wire signed [9:0] m123_12;
   assign m123_12 =10'b0;

   // m123_13 = W*in
   wire signed [9:0] m123_13;
   assign m123_13 =10'b0;

   // m123_14 = W*in
   wire signed [9:0] m123_14;
   assign m123_14 =10'b0;

   // m123_15 = W*in
   wire signed [9:0] m123_15;
   assign m123_15 =10'b0;

   // m123_16 = W*in
   wire signed [9:0] m123_16;
   assign m123_16 =10'b0;

   // m123_17 = W*in
   wire signed [9:0] m123_17;
   assign m123_17 =10'b0;

   // m123_18 = W*in
   wire signed [9:0] m123_18;
   assign m123_18 =10'b0;

   // m123_19 = W*in
   wire signed [9:0] m123_19;
   assign m123_19 =10'b0;

   // m123_20 = W*in
   wire signed [9:0] m123_20;
   assign m123_20 ={ {5{neg123[5]}} , neg123[5:1] };

   // m123_21 = W*in
   wire signed [9:0] m123_21;
   assign m123_21 =10'b0;

   // m123_22 = W*in
   wire signed [9:0] m123_22;
   assign m123_22 ={ {5{in123[5]}} , in123[5:1] };

   // m123_23 = W*in
   wire signed [9:0] m123_23;
   assign m123_23 ={ {5{in123[5]}} , in123[5:1] };

   // m123_24 = W*in
   wire signed [9:0] m123_24;
   assign m123_24 =10'b0;

   // m123_25 = W*in
   wire signed [9:0] m123_25;
   assign m123_25 =10'b0;

   // m123_26 = W*in
   wire signed [9:0] m123_26;
   assign m123_26 ={ {5{in123[5]}} , in123[5:1] };

   // m123_27 = W*in
   wire signed [9:0] m123_27;
   assign m123_27 =10'b0;

   // m123_28 = W*in
   wire signed [9:0] m123_28;
   assign m123_28 =10'b0;

   // m123_29 = W*in
   wire signed [9:0] m123_29;
   assign m123_29 ={ {4{in123[5]}} , in123[5:0] };

   // m123_30 = W*in
   wire signed [9:0] m123_30;
   assign m123_30 =10'b0;

   // m123_31 = W*in
   wire signed [9:0] m123_31;
   assign m123_31 =10'b0;

   // m123_32 = W*in
   wire signed [9:0] m123_32;
   assign m123_32 =10'b0;

   // m123_33 = W*in
   wire signed [9:0] m123_33;
   assign m123_33 =10'b0;

   // m123_34 = W*in
   wire signed [9:0] m123_34;
   assign m123_34 =10'b0;

   // m123_35 = W*in
   wire signed [9:0] m123_35;
   assign m123_35 =10'b0;

   // m123_36 = W*in
   wire signed [9:0] m123_36;
   assign m123_36 =10'b0;

   // m123_37 = W*in
   wire signed [9:0] m123_37;
   assign m123_37 =10'b0;

   // m123_38 = W*in
   wire signed [9:0] m123_38;
   assign m123_38 =10'b0;

   // m123_39 = W*in
   wire signed [9:0] m123_39;
   assign m123_39 =10'b0;

   // m123_40 = W*in
   wire signed [9:0] m123_40;
   assign m123_40 =10'b0;

   // m123_41 = W*in
   wire signed [9:0] m123_41;
   assign m123_41 =10'b0;

   // m123_42 = W*in
   wire signed [9:0] m123_42;
   assign m123_42 =10'b0;

   // m123_43 = W*in
   wire signed [9:0] m123_43;
   assign m123_43 =10'b0;

   // m123_44 = W*in
   wire signed [9:0] m123_44;
   assign m123_44 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_45 = W*in
   wire signed [9:0] m123_45;
   assign m123_45 =10'b0;

   // m123_46 = W*in
   wire signed [9:0] m123_46;
   assign m123_46 =10'b0;

   // m123_47 = W*in
   wire signed [9:0] m123_47;
   assign m123_47 =10'b0;

   // m123_48 = W*in
   wire signed [9:0] m123_48;
   assign m123_48 =10'b0;

   // m123_49 = W*in
   wire signed [9:0] m123_49;
   assign m123_49 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_50 = W*in
   wire signed [9:0] m123_50;
   assign m123_50 =10'b0;

   // m123_51 = W*in
   wire signed [9:0] m123_51;
   assign m123_51 =10'b0;

   // m123_52 = W*in
   wire signed [9:0] m123_52;
   assign m123_52 =10'b0;

   // m123_53 = W*in
   wire signed [9:0] m123_53;
   assign m123_53 =10'b0;

   // m123_54 = W*in
   wire signed [9:0] m123_54;
   assign m123_54 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_55 = W*in
   wire signed [9:0] m123_55;
   assign m123_55 =10'b0;

   // m123_56 = W*in
   wire signed [9:0] m123_56;
   assign m123_56 =10'b0;

   // m123_57 = W*in
   wire signed [9:0] m123_57;
   assign m123_57 =10'b0;

   // m123_58 = W*in
   wire signed [9:0] m123_58;
   assign m123_58 ={ {5{neg123[5]}} , neg123[5:1] };

   // m123_59 = W*in
   wire signed [9:0] m123_59;
   assign m123_59 =10'b0;

   // m123_60 = W*in
   wire signed [9:0] m123_60;
   assign m123_60 =10'b0;

   // m123_61 = W*in
   wire signed [9:0] m123_61;
   assign m123_61 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_62 = W*in
   wire signed [9:0] m123_62;
   assign m123_62 =10'b0;

   // m123_63 = W*in
   wire signed [9:0] m123_63;
   assign m123_63 =10'b0;

   // m123_64 = W*in
   wire signed [9:0] m123_64;
   assign m123_64 =10'b0;

   // m123_65 = W*in
   wire signed [9:0] m123_65;
   assign m123_65 =10'b0;

   // m123_66 = W*in
   wire signed [9:0] m123_66;
   assign m123_66 =10'b0;

   // m123_67 = W*in
   wire signed [9:0] m123_67;
   assign m123_67 =10'b0;

   // m123_68 = W*in
   wire signed [9:0] m123_68;
   assign m123_68 =10'b0;

   // m123_69 = W*in
   wire signed [9:0] m123_69;
   assign m123_69 =10'b0;

   // m123_70 = W*in
   wire signed [9:0] m123_70;
   assign m123_70 =10'b0;

   // m123_71 = W*in
   wire signed [9:0] m123_71;
   assign m123_71 =10'b0;

   // m123_72 = W*in
   wire signed [9:0] m123_72;
   assign m123_72 =10'b0;

   // m123_73 = W*in
   wire signed [9:0] m123_73;
   assign m123_73 ={ {5{in123[5]}} , in123[5:1] };

   // m123_74 = W*in
   wire signed [9:0] m123_74;
   assign m123_74 =10'b0;

   // m123_75 = W*in
   wire signed [9:0] m123_75;
   assign m123_75 =10'b0;

   // m123_76 = W*in
   wire signed [9:0] m123_76;
   assign m123_76 =10'b0;

   // m123_77 = W*in
   wire signed [9:0] m123_77;
   assign m123_77 =10'b0;

   // m123_78 = W*in
   wire signed [9:0] m123_78;
   assign m123_78 =10'b0;

   // m123_79 = W*in
   wire signed [9:0] m123_79;
   assign m123_79 =10'b0;

   // m123_80 = W*in
   wire signed [9:0] m123_80;
   assign m123_80 =10'b0;

   // m123_81 = W*in
   wire signed [9:0] m123_81;
   assign m123_81 =10'b0;

   // m123_82 = W*in
   wire signed [9:0] m123_82;
   assign m123_82 =10'b0;

   // m123_83 = W*in
   wire signed [9:0] m123_83;
   assign m123_83 =10'b0;

   // m123_84 = W*in
   wire signed [9:0] m123_84;
   assign m123_84 =10'b0;

   // m123_85 = W*in
   wire signed [9:0] m123_85;
   assign m123_85 =10'b0;

   // m123_86 = W*in
   wire signed [9:0] m123_86;
   assign m123_86 =10'b0;

   // m123_87 = W*in
   wire signed [9:0] m123_87;
   assign m123_87 =10'b0;

   // m123_88 = W*in
   wire signed [9:0] m123_88;
   assign m123_88 =10'b0;

   // m123_89 = W*in
   wire signed [9:0] m123_89;
   assign m123_89 =10'b0;

   // m123_90 = W*in
   wire signed [9:0] m123_90;
   assign m123_90 =10'b0;

   // m123_91 = W*in
   wire signed [9:0] m123_91;
   assign m123_91 =10'b0;

   // m123_92 = W*in
   wire signed [9:0] m123_92;
   assign m123_92 =10'b0;

   // m123_93 = W*in
   wire signed [9:0] m123_93;
   assign m123_93 =10'b0;

   // m123_94 = W*in
   wire signed [9:0] m123_94;
   assign m123_94 =10'b0;

   // m123_95 = W*in
   wire signed [9:0] m123_95;
   assign m123_95 =10'b0;

   // m123_96 = W*in
   wire signed [9:0] m123_96;
   assign m123_96 ={ {4{in123[5]}} , in123[5:0] };

   // m123_97 = W*in
   wire signed [9:0] m123_97;
   assign m123_97 =10'b0;

   // m123_98 = W*in
   wire signed [9:0] m123_98;
   assign m123_98 =10'b0;

   // m123_99 = W*in
   wire signed [9:0] m123_99;
   assign m123_99 =10'b0;

   // m123_100 = W*in
   wire signed [9:0] m123_100;
   assign m123_100 =10'b0;

   // m123_101 = W*in
   wire signed [9:0] m123_101;
   assign m123_101 =10'b0;

   // m123_102 = W*in
   wire signed [9:0] m123_102;
   assign m123_102 =10'b0;

   // m123_103 = W*in
   wire signed [9:0] m123_103;
   assign m123_103 ={ {4{in123[5]}} , in123[5:0] };

   // m123_104 = W*in
   wire signed [9:0] m123_104;
   assign m123_104 =10'b0;

   // m123_105 = W*in
   wire signed [9:0] m123_105;
   assign m123_105 =10'b0;

   // m123_106 = W*in
   wire signed [9:0] m123_106;
   assign m123_106 =10'b0;

   // m123_107 = W*in
   wire signed [9:0] m123_107;
   assign m123_107 =10'b0;

   // m123_108 = W*in
   wire signed [9:0] m123_108;
   assign m123_108 =10'b0;

   // m123_109 = W*in
   wire signed [9:0] m123_109;
   assign m123_109 =10'b0;

   // m123_110 = W*in
   wire signed [9:0] m123_110;
   assign m123_110 ={ {4{neg123[5]}} , neg123[5:0] };

   // m123_111 = W*in
   wire signed [9:0] m123_111;
   assign m123_111 =10'b0;

   // m123_112 = W*in
   wire signed [9:0] m123_112;
   assign m123_112 =10'b0;

   // m123_113 = W*in
   wire signed [9:0] m123_113;
   assign m123_113 =10'b0;

   // m123_114 = W*in
   wire signed [9:0] m123_114;
   assign m123_114 =10'b0;

   // m123_115 = W*in
   wire signed [9:0] m123_115;
   assign m123_115 =10'b0;

   // m123_116 = W*in
   wire signed [9:0] m123_116;
   assign m123_116 =10'b0;

   // m123_117 = W*in
   wire signed [9:0] m123_117;
   assign m123_117 =10'b0;

   // m124_1 = W*in
   wire signed [9:0] m124_1;
   assign m124_1 =10'b0;

   // m124_2 = W*in
   wire signed [9:0] m124_2;
   assign m124_2 =10'b0;

   // m124_3 = W*in
   wire signed [9:0] m124_3;
   assign m124_3 =10'b0;

   // m124_4 = W*in
   wire signed [9:0] m124_4;
   assign m124_4 =10'b0;

   // m124_5 = W*in
   wire signed [9:0] m124_5;
   assign m124_5 =10'b0;

   // m124_6 = W*in
   wire signed [9:0] m124_6;
   assign m124_6 =10'b0;

   // m124_7 = W*in
   wire signed [9:0] m124_7;
   assign m124_7 ={ {4{in124[5]}} , in124[5:0] };

   // m124_8 = W*in
   wire signed [9:0] m124_8;
   assign m124_8 =10'b0;

   // m124_9 = W*in
   wire signed [9:0] m124_9;
   assign m124_9 =10'b0;

   // m124_10 = W*in
   wire signed [9:0] m124_10;
   assign m124_10 =10'b0;

   // m124_11 = W*in
   wire signed [9:0] m124_11;
   assign m124_11 =10'b0;

   // m124_12 = W*in
   wire signed [9:0] m124_12;
   assign m124_12 =10'b0;

   // m124_13 = W*in
   wire signed [9:0] m124_13;
   assign m124_13 ={ {4{in124[5]}} , in124[5:0] };

   // m124_14 = W*in
   wire signed [9:0] m124_14;
   assign m124_14 =10'b0;

   // m124_15 = W*in
   wire signed [9:0] m124_15;
   assign m124_15 =10'b0;

   // m124_16 = W*in
   wire signed [9:0] m124_16;
   assign m124_16 =10'b0;

   // m124_17 = W*in
   wire signed [9:0] m124_17;
   assign m124_17 =10'b0;

   // m124_18 = W*in
   wire signed [9:0] m124_18;
   assign m124_18 ={ {5{neg124[5]}} , neg124[5:1] };

   // m124_19 = W*in
   wire signed [9:0] m124_19;
   assign m124_19 ={ {5{neg124[5]}} , neg124[5:1] };

   // m124_20 = W*in
   wire signed [9:0] m124_20;
   assign m124_20 =10'b0;

   // m124_21 = W*in
   wire signed [9:0] m124_21;
   assign m124_21 ={ {5{in124[5]}} , in124[5:1] };

   // m124_22 = W*in
   wire signed [9:0] m124_22;
   assign m124_22 ={ {5{in124[5]}} , in124[5:1] };

   // m124_23 = W*in
   wire signed [9:0] m124_23;
   assign m124_23 ={ {5{in124[5]}} , in124[5:1] };

   // m124_24 = W*in
   wire signed [9:0] m124_24;
   assign m124_24 =10'b0;

   // m124_25 = W*in
   wire signed [9:0] m124_25;
   assign m124_25 =10'b0;

   // m124_26 = W*in
   wire signed [9:0] m124_26;
   assign m124_26 =10'b0;

   // m124_27 = W*in
   wire signed [9:0] m124_27;
   assign m124_27 =10'b0;

   // m124_28 = W*in
   wire signed [9:0] m124_28;
   assign m124_28 =10'b0;

   // m124_29 = W*in
   wire signed [9:0] m124_29;
   assign m124_29 =10'b0;

   // m124_30 = W*in
   wire signed [9:0] m124_30;
   assign m124_30 =10'b0;

   // m124_31 = W*in
   wire signed [9:0] m124_31;
   assign m124_31 ={ {5{neg124[5]}} , neg124[5:1] };

   // m124_32 = W*in
   wire signed [9:0] m124_32;
   assign m124_32 =10'b0;

   // m124_33 = W*in
   wire signed [9:0] m124_33;
   assign m124_33 ={ {4{in124[5]}} , in124[5:0] };

   // m124_34 = W*in
   wire signed [9:0] m124_34;
   assign m124_34 =10'b0;

   // m124_35 = W*in
   wire signed [9:0] m124_35;
   assign m124_35 =10'b0;

   // m124_36 = W*in
   wire signed [9:0] m124_36;
   assign m124_36 =10'b0;

   // m124_37 = W*in
   wire signed [9:0] m124_37;
   assign m124_37 =10'b0;

   // m124_38 = W*in
   wire signed [9:0] m124_38;
   assign m124_38 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_39 = W*in
   wire signed [9:0] m124_39;
   assign m124_39 =10'b0;

   // m124_40 = W*in
   wire signed [9:0] m124_40;
   assign m124_40 =10'b0;

   // m124_41 = W*in
   wire signed [9:0] m124_41;
   assign m124_41 ={ {4{in124[5]}} , in124[5:0] };

   // m124_42 = W*in
   wire signed [9:0] m124_42;
   assign m124_42 =10'b0;

   // m124_43 = W*in
   wire signed [9:0] m124_43;
   assign m124_43 =10'b0;

   // m124_44 = W*in
   wire signed [9:0] m124_44;
   assign m124_44 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_45 = W*in
   wire signed [9:0] m124_45;
   assign m124_45 ={ {4{in124[5]}} , in124[5:0] };

   // m124_46 = W*in
   wire signed [9:0] m124_46;
   assign m124_46 =10'b0;

   // m124_47 = W*in
   wire signed [9:0] m124_47;
   assign m124_47 =10'b0;

   // m124_48 = W*in
   wire signed [9:0] m124_48;
   assign m124_48 =10'b0;

   // m124_49 = W*in
   wire signed [9:0] m124_49;
   assign m124_49 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_50 = W*in
   wire signed [9:0] m124_50;
   assign m124_50 =10'b0;

   // m124_51 = W*in
   wire signed [9:0] m124_51;
   assign m124_51 =10'b0;

   // m124_52 = W*in
   wire signed [9:0] m124_52;
   assign m124_52 =10'b0;

   // m124_53 = W*in
   wire signed [9:0] m124_53;
   assign m124_53 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_54 = W*in
   wire signed [9:0] m124_54;
   assign m124_54 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_55 = W*in
   wire signed [9:0] m124_55;
   assign m124_55 =10'b0;

   // m124_56 = W*in
   wire signed [9:0] m124_56;
   assign m124_56 =10'b0;

   // m124_57 = W*in
   wire signed [9:0] m124_57;
   assign m124_57 =10'b0;

   // m124_58 = W*in
   wire signed [9:0] m124_58;
   assign m124_58 =10'b0;

   // m124_59 = W*in
   wire signed [9:0] m124_59;
   assign m124_59 =10'b0;

   // m124_60 = W*in
   wire signed [9:0] m124_60;
   assign m124_60 =10'b0;

   // m124_61 = W*in
   wire signed [9:0] m124_61;
   assign m124_61 =10'b0;

   // m124_62 = W*in
   wire signed [9:0] m124_62;
   assign m124_62 =10'b0;

   // m124_63 = W*in
   wire signed [9:0] m124_63;
   assign m124_63 =10'b0;

   // m124_64 = W*in
   wire signed [9:0] m124_64;
   assign m124_64 =10'b0;

   // m124_65 = W*in
   wire signed [9:0] m124_65;
   assign m124_65 =10'b0;

   // m124_66 = W*in
   wire signed [9:0] m124_66;
   assign m124_66 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_67 = W*in
   wire signed [9:0] m124_67;
   assign m124_67 =10'b0;

   // m124_68 = W*in
   wire signed [9:0] m124_68;
   assign m124_68 =10'b0;

   // m124_69 = W*in
   wire signed [9:0] m124_69;
   assign m124_69 ={ {5{in124[5]}} , in124[5:1] };

   // m124_70 = W*in
   wire signed [9:0] m124_70;
   assign m124_70 =10'b0;

   // m124_71 = W*in
   wire signed [9:0] m124_71;
   assign m124_71 ={ {5{neg124[5]}} , neg124[5:1] };

   // m124_72 = W*in
   wire signed [9:0] m124_72;
   assign m124_72 =10'b0;

   // m124_73 = W*in
   wire signed [9:0] m124_73;
   assign m124_73 ={ {5{in124[5]}} , in124[5:1] };

   // m124_74 = W*in
   wire signed [9:0] m124_74;
   assign m124_74 ={ {5{neg124[5]}} , neg124[5:1] };

   // m124_75 = W*in
   wire signed [9:0] m124_75;
   assign m124_75 =10'b0;

   // m124_76 = W*in
   wire signed [9:0] m124_76;
   assign m124_76 =10'b0;

   // m124_77 = W*in
   wire signed [9:0] m124_77;
   assign m124_77 =10'b0;

   // m124_78 = W*in
   wire signed [9:0] m124_78;
   assign m124_78 ={ {5{in124[5]}} , in124[5:1] };

   // m124_79 = W*in
   wire signed [9:0] m124_79;
   assign m124_79 =10'b0;

   // m124_80 = W*in
   wire signed [9:0] m124_80;
   assign m124_80 =10'b0;

   // m124_81 = W*in
   wire signed [9:0] m124_81;
   assign m124_81 =10'b0;

   // m124_82 = W*in
   wire signed [9:0] m124_82;
   assign m124_82 ={ {4{in124[5]}} , in124[5:0] };

   // m124_83 = W*in
   wire signed [9:0] m124_83;
   assign m124_83 =10'b0;

   // m124_84 = W*in
   wire signed [9:0] m124_84;
   assign m124_84 =10'b0;

   // m124_85 = W*in
   wire signed [9:0] m124_85;
   assign m124_85 =10'b0;

   // m124_86 = W*in
   wire signed [9:0] m124_86;
   assign m124_86 =10'b0;

   // m124_87 = W*in
   wire signed [9:0] m124_87;
   assign m124_87 =10'b0;

   // m124_88 = W*in
   wire signed [9:0] m124_88;
   assign m124_88 =10'b0;

   // m124_89 = W*in
   wire signed [9:0] m124_89;
   assign m124_89 =10'b0;

   // m124_90 = W*in
   wire signed [9:0] m124_90;
   assign m124_90 =10'b0;

   // m124_91 = W*in
   wire signed [9:0] m124_91;
   assign m124_91 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_92 = W*in
   wire signed [9:0] m124_92;
   assign m124_92 =10'b0;

   // m124_93 = W*in
   wire signed [9:0] m124_93;
   assign m124_93 =10'b0;

   // m124_94 = W*in
   wire signed [9:0] m124_94;
   assign m124_94 =10'b0;

   // m124_95 = W*in
   wire signed [9:0] m124_95;
   assign m124_95 =10'b0;

   // m124_96 = W*in
   wire signed [9:0] m124_96;
   assign m124_96 =10'b0;

   // m124_97 = W*in
   wire signed [9:0] m124_97;
   assign m124_97 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_98 = W*in
   wire signed [9:0] m124_98;
   assign m124_98 =10'b0;

   // m124_99 = W*in
   wire signed [9:0] m124_99;
   assign m124_99 =10'b0;

   // m124_100 = W*in
   wire signed [9:0] m124_100;
   assign m124_100 =10'b0;

   // m124_101 = W*in
   wire signed [9:0] m124_101;
   assign m124_101 =10'b0;

   // m124_102 = W*in
   wire signed [9:0] m124_102;
   assign m124_102 =10'b0;

   // m124_103 = W*in
   wire signed [9:0] m124_103;
   assign m124_103 =10'b0;

   // m124_104 = W*in
   wire signed [9:0] m124_104;
   assign m124_104 =10'b0;

   // m124_105 = W*in
   wire signed [9:0] m124_105;
   assign m124_105 =10'b0;

   // m124_106 = W*in
   wire signed [9:0] m124_106;
   assign m124_106 =10'b0;

   // m124_107 = W*in
   wire signed [9:0] m124_107;
   assign m124_107 =10'b0;

   // m124_108 = W*in
   wire signed [9:0] m124_108;
   assign m124_108 ={ {4{in124[5]}} , in124[5:0] };

   // m124_109 = W*in
   wire signed [9:0] m124_109;
   assign m124_109 ={ {5{in124[5]}} , in124[5:1] };

   // m124_110 = W*in
   wire signed [9:0] m124_110;
   assign m124_110 ={ {4{neg124[5]}} , neg124[5:0] };

   // m124_111 = W*in
   wire signed [9:0] m124_111;
   assign m124_111 =10'b0;

   // m124_112 = W*in
   wire signed [9:0] m124_112;
   assign m124_112 =10'b0;

   // m124_113 = W*in
   wire signed [9:0] m124_113;
   assign m124_113 =10'b0;

   // m124_114 = W*in
   wire signed [9:0] m124_114;
   assign m124_114 ={ {5{in124[5]}} , in124[5:1] };

   // m124_115 = W*in
   wire signed [9:0] m124_115;
   assign m124_115 =10'b0;

   // m124_116 = W*in
   wire signed [9:0] m124_116;
   assign m124_116 ={ {4{in124[5]}} , in124[5:0] };

   // m124_117 = W*in
   wire signed [9:0] m124_117;
   assign m124_117 =10'b0;

   // m125_1 = W*in
   wire signed [9:0] m125_1;
   assign m125_1 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_2 = W*in
   wire signed [9:0] m125_2;
   assign m125_2 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_3 = W*in
   wire signed [9:0] m125_3;
   assign m125_3 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_4 = W*in
   wire signed [9:0] m125_4;
   assign m125_4 =10'b0;

   // m125_5 = W*in
   wire signed [9:0] m125_5;
   assign m125_5 ={ {4{in125[5]}} , in125[5:0] };

   // m125_6 = W*in
   wire signed [9:0] m125_6;
   assign m125_6 =10'b0;

   // m125_7 = W*in
   wire signed [9:0] m125_7;
   assign m125_7 ={ {4{in125[5]}} , in125[5:0] };

   // m125_8 = W*in
   wire signed [9:0] m125_8;
   assign m125_8 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_9 = W*in
   wire signed [9:0] m125_9;
   assign m125_9 =10'b0;

   // m125_10 = W*in
   wire signed [9:0] m125_10;
   assign m125_10 =10'b0;

   // m125_11 = W*in
   wire signed [9:0] m125_11;
   assign m125_11 =10'b0;

   // m125_12 = W*in
   wire signed [9:0] m125_12;
   assign m125_12 =10'b0;

   // m125_13 = W*in
   wire signed [9:0] m125_13;
   assign m125_13 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_14 = W*in
   wire signed [9:0] m125_14;
   assign m125_14 =10'b0;

   // m125_15 = W*in
   wire signed [9:0] m125_15;
   assign m125_15 =10'b0;

   // m125_16 = W*in
   wire signed [9:0] m125_16;
   assign m125_16 =10'b0;

   // m125_17 = W*in
   wire signed [9:0] m125_17;
   assign m125_17 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_18 = W*in
   wire signed [9:0] m125_18;
   assign m125_18 =10'b0;

   // m125_19 = W*in
   wire signed [9:0] m125_19;
   assign m125_19 ={ {5{neg125[5]}} , neg125[5:1] };

   // m125_20 = W*in
   wire signed [9:0] m125_20;
   assign m125_20 ={ {5{in125[5]}} , in125[5:1] };

   // m125_21 = W*in
   wire signed [9:0] m125_21;
   assign m125_21 =10'b0;

   // m125_22 = W*in
   wire signed [9:0] m125_22;
   assign m125_22 =10'b0;

   // m125_23 = W*in
   wire signed [9:0] m125_23;
   assign m125_23 ={ {5{neg125[5]}} , neg125[5:1] };

   // m125_24 = W*in
   wire signed [9:0] m125_24;
   assign m125_24 =10'b0;

   // m125_25 = W*in
   wire signed [9:0] m125_25;
   assign m125_25 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_26 = W*in
   wire signed [9:0] m125_26;
   assign m125_26 =10'b0;

   // m125_27 = W*in
   wire signed [9:0] m125_27;
   assign m125_27 =10'b0;

   // m125_28 = W*in
   wire signed [9:0] m125_28;
   assign m125_28 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_29 = W*in
   wire signed [9:0] m125_29;
   assign m125_29 =10'b0;

   // m125_30 = W*in
   wire signed [9:0] m125_30;
   assign m125_30 =10'b0;

   // m125_31 = W*in
   wire signed [9:0] m125_31;
   assign m125_31 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_32 = W*in
   wire signed [9:0] m125_32;
   assign m125_32 =10'b0;

   // m125_33 = W*in
   wire signed [9:0] m125_33;
   assign m125_33 =10'b0;

   // m125_34 = W*in
   wire signed [9:0] m125_34;
   assign m125_34 =10'b0;

   // m125_35 = W*in
   wire signed [9:0] m125_35;
   assign m125_35 ={ {4{in125[5]}} , in125[5:0] };

   // m125_36 = W*in
   wire signed [9:0] m125_36;
   assign m125_36 =10'b0;

   // m125_37 = W*in
   wire signed [9:0] m125_37;
   assign m125_37 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_38 = W*in
   wire signed [9:0] m125_38;
   assign m125_38 ={ {4{in125[5]}} , in125[5:0] };

   // m125_39 = W*in
   wire signed [9:0] m125_39;
   assign m125_39 ={ {4{in125[5]}} , in125[5:0] };

   // m125_40 = W*in
   wire signed [9:0] m125_40;
   assign m125_40 =10'b0;

   // m125_41 = W*in
   wire signed [9:0] m125_41;
   assign m125_41 =10'b0;

   // m125_42 = W*in
   wire signed [9:0] m125_42;
   assign m125_42 =10'b0;

   // m125_43 = W*in
   wire signed [9:0] m125_43;
   assign m125_43 =10'b0;

   // m125_44 = W*in
   wire signed [9:0] m125_44;
   assign m125_44 =10'b0;

   // m125_45 = W*in
   wire signed [9:0] m125_45;
   assign m125_45 =10'b0;

   // m125_46 = W*in
   wire signed [9:0] m125_46;
   assign m125_46 =10'b0;

   // m125_47 = W*in
   wire signed [9:0] m125_47;
   assign m125_47 =10'b0;

   // m125_48 = W*in
   wire signed [9:0] m125_48;
   assign m125_48 =10'b0;

   // m125_49 = W*in
   wire signed [9:0] m125_49;
   assign m125_49 =10'b0;

   // m125_50 = W*in
   wire signed [9:0] m125_50;
   assign m125_50 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_51 = W*in
   wire signed [9:0] m125_51;
   assign m125_51 =10'b0;

   // m125_52 = W*in
   wire signed [9:0] m125_52;
   assign m125_52 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_53 = W*in
   wire signed [9:0] m125_53;
   assign m125_53 =10'b0;

   // m125_54 = W*in
   wire signed [9:0] m125_54;
   assign m125_54 =10'b0;

   // m125_55 = W*in
   wire signed [9:0] m125_55;
   assign m125_55 =10'b0;

   // m125_56 = W*in
   wire signed [9:0] m125_56;
   assign m125_56 =10'b0;

   // m125_57 = W*in
   wire signed [9:0] m125_57;
   assign m125_57 =10'b0;

   // m125_58 = W*in
   wire signed [9:0] m125_58;
   assign m125_58 =10'b0;

   // m125_59 = W*in
   wire signed [9:0] m125_59;
   assign m125_59 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_60 = W*in
   wire signed [9:0] m125_60;
   assign m125_60 =10'b0;

   // m125_61 = W*in
   wire signed [9:0] m125_61;
   assign m125_61 =10'b0;

   // m125_62 = W*in
   wire signed [9:0] m125_62;
   assign m125_62 =10'b0;

   // m125_63 = W*in
   wire signed [9:0] m125_63;
   assign m125_63 =10'b0;

   // m125_64 = W*in
   wire signed [9:0] m125_64;
   assign m125_64 =10'b0;

   // m125_65 = W*in
   wire signed [9:0] m125_65;
   assign m125_65 =10'b0;

   // m125_66 = W*in
   wire signed [9:0] m125_66;
   assign m125_66 =10'b0;

   // m125_67 = W*in
   wire signed [9:0] m125_67;
   assign m125_67 =10'b0;

   // m125_68 = W*in
   wire signed [9:0] m125_68;
   assign m125_68 =10'b0;

   // m125_69 = W*in
   wire signed [9:0] m125_69;
   assign m125_69 =10'b0;

   // m125_70 = W*in
   wire signed [9:0] m125_70;
   assign m125_70 =10'b0;

   // m125_71 = W*in
   wire signed [9:0] m125_71;
   assign m125_71 =10'b0;

   // m125_72 = W*in
   wire signed [9:0] m125_72;
   assign m125_72 ={ {4{in125[5]}} , in125[5:0] };

   // m125_73 = W*in
   wire signed [9:0] m125_73;
   assign m125_73 =10'b0;

   // m125_74 = W*in
   wire signed [9:0] m125_74;
   assign m125_74 =10'b0;

   // m125_75 = W*in
   wire signed [9:0] m125_75;
   assign m125_75 =10'b0;

   // m125_76 = W*in
   wire signed [9:0] m125_76;
   assign m125_76 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_77 = W*in
   wire signed [9:0] m125_77;
   assign m125_77 =10'b0;

   // m125_78 = W*in
   wire signed [9:0] m125_78;
   assign m125_78 ={ {4{in125[5]}} , in125[5:0] };

   // m125_79 = W*in
   wire signed [9:0] m125_79;
   assign m125_79 =10'b0;

   // m125_80 = W*in
   wire signed [9:0] m125_80;
   assign m125_80 =10'b0;

   // m125_81 = W*in
   wire signed [9:0] m125_81;
   assign m125_81 ={ {5{neg125[5]}} , neg125[5:1] };

   // m125_82 = W*in
   wire signed [9:0] m125_82;
   assign m125_82 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_83 = W*in
   wire signed [9:0] m125_83;
   assign m125_83 =10'b0;

   // m125_84 = W*in
   wire signed [9:0] m125_84;
   assign m125_84 =10'b0;

   // m125_85 = W*in
   wire signed [9:0] m125_85;
   assign m125_85 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_86 = W*in
   wire signed [9:0] m125_86;
   assign m125_86 =10'b0;

   // m125_87 = W*in
   wire signed [9:0] m125_87;
   assign m125_87 =10'b0;

   // m125_88 = W*in
   wire signed [9:0] m125_88;
   assign m125_88 =10'b0;

   // m125_89 = W*in
   wire signed [9:0] m125_89;
   assign m125_89 =10'b0;

   // m125_90 = W*in
   wire signed [9:0] m125_90;
   assign m125_90 =10'b0;

   // m125_91 = W*in
   wire signed [9:0] m125_91;
   assign m125_91 =10'b0;

   // m125_92 = W*in
   wire signed [9:0] m125_92;
   assign m125_92 =10'b0;

   // m125_93 = W*in
   wire signed [9:0] m125_93;
   assign m125_93 =10'b0;

   // m125_94 = W*in
   wire signed [9:0] m125_94;
   assign m125_94 =10'b0;

   // m125_95 = W*in
   wire signed [9:0] m125_95;
   assign m125_95 =10'b0;

   // m125_96 = W*in
   wire signed [9:0] m125_96;
   assign m125_96 =10'b0;

   // m125_97 = W*in
   wire signed [9:0] m125_97;
   assign m125_97 =10'b0;

   // m125_98 = W*in
   wire signed [9:0] m125_98;
   assign m125_98 =10'b0;

   // m125_99 = W*in
   wire signed [9:0] m125_99;
   assign m125_99 =10'b0;

   // m125_100 = W*in
   wire signed [9:0] m125_100;
   assign m125_100 =10'b0;

   // m125_101 = W*in
   wire signed [9:0] m125_101;
   assign m125_101 =10'b0;

   // m125_102 = W*in
   wire signed [9:0] m125_102;
   assign m125_102 =10'b0;

   // m125_103 = W*in
   wire signed [9:0] m125_103;
   assign m125_103 =10'b0;

   // m125_104 = W*in
   wire signed [9:0] m125_104;
   assign m125_104 =10'b0;

   // m125_105 = W*in
   wire signed [9:0] m125_105;
   assign m125_105 =10'b0;

   // m125_106 = W*in
   wire signed [9:0] m125_106;
   assign m125_106 =10'b0;

   // m125_107 = W*in
   wire signed [9:0] m125_107;
   assign m125_107 =10'b0;

   // m125_108 = W*in
   wire signed [9:0] m125_108;
   assign m125_108 ={ {5{neg125[5]}} , neg125[5:1] };

   // m125_109 = W*in
   wire signed [9:0] m125_109;
   assign m125_109 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_110 = W*in
   wire signed [9:0] m125_110;
   assign m125_110 =10'b0;

   // m125_111 = W*in
   wire signed [9:0] m125_111;
   assign m125_111 =10'b0;

   // m125_112 = W*in
   wire signed [9:0] m125_112;
   assign m125_112 =10'b0;

   // m125_113 = W*in
   wire signed [9:0] m125_113;
   assign m125_113 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_114 = W*in
   wire signed [9:0] m125_114;
   assign m125_114 =10'b0;

   // m125_115 = W*in
   wire signed [9:0] m125_115;
   assign m125_115 ={ {5{in125[5]}} , in125[5:1] };

   // m125_116 = W*in
   wire signed [9:0] m125_116;
   assign m125_116 ={ {4{neg125[5]}} , neg125[5:0] };

   // m125_117 = W*in
   wire signed [9:0] m125_117;
   assign m125_117 =10'b0;

   // m126_1 = W*in
   wire signed [9:0] m126_1;
   assign m126_1 ={ {3{neg126[5]}} , neg126 , {1{1'b0}} };

   // m126_2 = W*in
   wire signed [9:0] m126_2;
   assign m126_2 =10'b0;

   // m126_3 = W*in
   wire signed [9:0] m126_3;
   assign m126_3 =10'b0;

   // m126_4 = W*in
   wire signed [9:0] m126_4;
   assign m126_4 =10'b0;

   // m126_5 = W*in
   wire signed [9:0] m126_5;
   assign m126_5 =10'b0;

   // m126_6 = W*in
   wire signed [9:0] m126_6;
   assign m126_6 ={ {4{in126[5]}} , in126[5:0] };

   // m126_7 = W*in
   wire signed [9:0] m126_7;
   assign m126_7 ={ {4{in126[5]}} , in126[5:0] };

   // m126_8 = W*in
   wire signed [9:0] m126_8;
   assign m126_8 =10'b0;

   // m126_9 = W*in
   wire signed [9:0] m126_9;
   assign m126_9 =10'b0;

   // m126_10 = W*in
   wire signed [9:0] m126_10;
   assign m126_10 =10'b0;

   // m126_11 = W*in
   wire signed [9:0] m126_11;
   assign m126_11 =10'b0;

   // m126_12 = W*in
   wire signed [9:0] m126_12;
   assign m126_12 =10'b0;

   // m126_13 = W*in
   wire signed [9:0] m126_13;
   assign m126_13 =10'b0;

   // m126_14 = W*in
   wire signed [9:0] m126_14;
   assign m126_14 =10'b0;

   // m126_15 = W*in
   wire signed [9:0] m126_15;
   assign m126_15 ={ {5{neg126[5]}} , neg126[5:1] };

   // m126_16 = W*in
   wire signed [9:0] m126_16;
   assign m126_16 =10'b0;

   // m126_17 = W*in
   wire signed [9:0] m126_17;
   assign m126_17 =10'b0;

   // m126_18 = W*in
   wire signed [9:0] m126_18;
   assign m126_18 =10'b0;

   // m126_19 = W*in
   wire signed [9:0] m126_19;
   assign m126_19 =10'b0;

   // m126_20 = W*in
   wire signed [9:0] m126_20;
   assign m126_20 =10'b0;

   // m126_21 = W*in
   wire signed [9:0] m126_21;
   assign m126_21 =10'b0;

   // m126_22 = W*in
   wire signed [9:0] m126_22;
   assign m126_22 =10'b0;

   // m126_23 = W*in
   wire signed [9:0] m126_23;
   assign m126_23 ={ {5{neg126[5]}} , neg126[5:1] };

   // m126_24 = W*in
   wire signed [9:0] m126_24;
   assign m126_24 =10'b0;

   // m126_25 = W*in
   wire signed [9:0] m126_25;
   assign m126_25 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_26 = W*in
   wire signed [9:0] m126_26;
   assign m126_26 =10'b0;

   // m126_27 = W*in
   wire signed [9:0] m126_27;
   assign m126_27 =10'b0;

   // m126_28 = W*in
   wire signed [9:0] m126_28;
   assign m126_28 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_29 = W*in
   wire signed [9:0] m126_29;
   assign m126_29 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_30 = W*in
   wire signed [9:0] m126_30;
   assign m126_30 =10'b0;

   // m126_31 = W*in
   wire signed [9:0] m126_31;
   assign m126_31 ={ {5{neg126[5]}} , neg126[5:1] };

   // m126_32 = W*in
   wire signed [9:0] m126_32;
   assign m126_32 ={ {4{in126[5]}} , in126[5:0] };

   // m126_33 = W*in
   wire signed [9:0] m126_33;
   assign m126_33 =10'b0;

   // m126_34 = W*in
   wire signed [9:0] m126_34;
   assign m126_34 ={ {4{in126[5]}} , in126[5:0] };

   // m126_35 = W*in
   wire signed [9:0] m126_35;
   assign m126_35 =10'b0;

   // m126_36 = W*in
   wire signed [9:0] m126_36;
   assign m126_36 =10'b0;

   // m126_37 = W*in
   wire signed [9:0] m126_37;
   assign m126_37 =10'b0;

   // m126_38 = W*in
   wire signed [9:0] m126_38;
   assign m126_38 =10'b0;

   // m126_39 = W*in
   wire signed [9:0] m126_39;
   assign m126_39 ={ {4{in126[5]}} , in126[5:0] };

   // m126_40 = W*in
   wire signed [9:0] m126_40;
   assign m126_40 =10'b0;

   // m126_41 = W*in
   wire signed [9:0] m126_41;
   assign m126_41 =10'b0;

   // m126_42 = W*in
   wire signed [9:0] m126_42;
   assign m126_42 =10'b0;

   // m126_43 = W*in
   wire signed [9:0] m126_43;
   assign m126_43 =10'b0;

   // m126_44 = W*in
   wire signed [9:0] m126_44;
   assign m126_44 =10'b0;

   // m126_45 = W*in
   wire signed [9:0] m126_45;
   assign m126_45 =10'b0;

   // m126_46 = W*in
   wire signed [9:0] m126_46;
   assign m126_46 =10'b0;

   // m126_47 = W*in
   wire signed [9:0] m126_47;
   assign m126_47 ={ {4{in126[5]}} , in126[5:0] };

   // m126_48 = W*in
   wire signed [9:0] m126_48;
   assign m126_48 =10'b0;

   // m126_49 = W*in
   wire signed [9:0] m126_49;
   assign m126_49 =10'b0;

   // m126_50 = W*in
   wire signed [9:0] m126_50;
   assign m126_50 =10'b0;

   // m126_51 = W*in
   wire signed [9:0] m126_51;
   assign m126_51 ={ {4{in126[5]}} , in126[5:0] };

   // m126_52 = W*in
   wire signed [9:0] m126_52;
   assign m126_52 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_53 = W*in
   wire signed [9:0] m126_53;
   assign m126_53 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_54 = W*in
   wire signed [9:0] m126_54;
   assign m126_54 ={ {4{in126[5]}} , in126[5:0] };

   // m126_55 = W*in
   wire signed [9:0] m126_55;
   assign m126_55 =10'b0;

   // m126_56 = W*in
   wire signed [9:0] m126_56;
   assign m126_56 =10'b0;

   // m126_57 = W*in
   wire signed [9:0] m126_57;
   assign m126_57 =10'b0;

   // m126_58 = W*in
   wire signed [9:0] m126_58;
   assign m126_58 ={ {5{in126[5]}} , in126[5:1] };

   // m126_59 = W*in
   wire signed [9:0] m126_59;
   assign m126_59 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_60 = W*in
   wire signed [9:0] m126_60;
   assign m126_60 =10'b0;

   // m126_61 = W*in
   wire signed [9:0] m126_61;
   assign m126_61 =10'b0;

   // m126_62 = W*in
   wire signed [9:0] m126_62;
   assign m126_62 =10'b0;

   // m126_63 = W*in
   wire signed [9:0] m126_63;
   assign m126_63 =10'b0;

   // m126_64 = W*in
   wire signed [9:0] m126_64;
   assign m126_64 =10'b0;

   // m126_65 = W*in
   wire signed [9:0] m126_65;
   assign m126_65 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_66 = W*in
   wire signed [9:0] m126_66;
   assign m126_66 =10'b0;

   // m126_67 = W*in
   wire signed [9:0] m126_67;
   assign m126_67 =10'b0;

   // m126_68 = W*in
   wire signed [9:0] m126_68;
   assign m126_68 =10'b0;

   // m126_69 = W*in
   wire signed [9:0] m126_69;
   assign m126_69 =10'b0;

   // m126_70 = W*in
   wire signed [9:0] m126_70;
   assign m126_70 =10'b0;

   // m126_71 = W*in
   wire signed [9:0] m126_71;
   assign m126_71 =10'b0;

   // m126_72 = W*in
   wire signed [9:0] m126_72;
   assign m126_72 ={ {5{in126[5]}} , in126[5:1] };

   // m126_73 = W*in
   wire signed [9:0] m126_73;
   assign m126_73 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_74 = W*in
   wire signed [9:0] m126_74;
   assign m126_74 ={ {4{in126[5]}} , in126[5:0] };

   // m126_75 = W*in
   wire signed [9:0] m126_75;
   assign m126_75 =10'b0;

   // m126_76 = W*in
   wire signed [9:0] m126_76;
   assign m126_76 =10'b0;

   // m126_77 = W*in
   wire signed [9:0] m126_77;
   assign m126_77 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_78 = W*in
   wire signed [9:0] m126_78;
   assign m126_78 ={ {4{in126[5]}} , in126[5:0] };

   // m126_79 = W*in
   wire signed [9:0] m126_79;
   assign m126_79 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_80 = W*in
   wire signed [9:0] m126_80;
   assign m126_80 ={ {5{neg126[5]}} , neg126[5:1] };

   // m126_81 = W*in
   wire signed [9:0] m126_81;
   assign m126_81 ={ {5{neg126[5]}} , neg126[5:1] };

   // m126_82 = W*in
   wire signed [9:0] m126_82;
   assign m126_82 =10'b0;

   // m126_83 = W*in
   wire signed [9:0] m126_83;
   assign m126_83 ={ {4{in126[5]}} , in126[5:0] };

   // m126_84 = W*in
   wire signed [9:0] m126_84;
   assign m126_84 =10'b0;

   // m126_85 = W*in
   wire signed [9:0] m126_85;
   assign m126_85 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_86 = W*in
   wire signed [9:0] m126_86;
   assign m126_86 =10'b0;

   // m126_87 = W*in
   wire signed [9:0] m126_87;
   assign m126_87 ={ {4{in126[5]}} , in126[5:0] };

   // m126_88 = W*in
   wire signed [9:0] m126_88;
   assign m126_88 =10'b0;

   // m126_89 = W*in
   wire signed [9:0] m126_89;
   assign m126_89 =10'b0;

   // m126_90 = W*in
   wire signed [9:0] m126_90;
   assign m126_90 =10'b0;

   // m126_91 = W*in
   wire signed [9:0] m126_91;
   assign m126_91 =10'b0;

   // m126_92 = W*in
   wire signed [9:0] m126_92;
   assign m126_92 ={ {4{in126[5]}} , in126[5:0] };

   // m126_93 = W*in
   wire signed [9:0] m126_93;
   assign m126_93 =10'b0;

   // m126_94 = W*in
   wire signed [9:0] m126_94;
   assign m126_94 =10'b0;

   // m126_95 = W*in
   wire signed [9:0] m126_95;
   assign m126_95 =10'b0;

   // m126_96 = W*in
   wire signed [9:0] m126_96;
   assign m126_96 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_97 = W*in
   wire signed [9:0] m126_97;
   assign m126_97 =10'b0;

   // m126_98 = W*in
   wire signed [9:0] m126_98;
   assign m126_98 =10'b0;

   // m126_99 = W*in
   wire signed [9:0] m126_99;
   assign m126_99 ={ {4{in126[5]}} , in126[5:0] };

   // m126_100 = W*in
   wire signed [9:0] m126_100;
   assign m126_100 =10'b0;

   // m126_101 = W*in
   wire signed [9:0] m126_101;
   assign m126_101 =10'b0;

   // m126_102 = W*in
   wire signed [9:0] m126_102;
   assign m126_102 ={ {4{in126[5]}} , in126[5:0] };

   // m126_103 = W*in
   wire signed [9:0] m126_103;
   assign m126_103 =10'b0;

   // m126_104 = W*in
   wire signed [9:0] m126_104;
   assign m126_104 =10'b0;

   // m126_105 = W*in
   wire signed [9:0] m126_105;
   assign m126_105 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_106 = W*in
   wire signed [9:0] m126_106;
   assign m126_106 =10'b0;

   // m126_107 = W*in
   wire signed [9:0] m126_107;
   assign m126_107 =10'b0;

   // m126_108 = W*in
   wire signed [9:0] m126_108;
   assign m126_108 ={ {5{neg126[5]}} , neg126[5:1] };

   // m126_109 = W*in
   wire signed [9:0] m126_109;
   assign m126_109 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_110 = W*in
   wire signed [9:0] m126_110;
   assign m126_110 =10'b0;

   // m126_111 = W*in
   wire signed [9:0] m126_111;
   assign m126_111 =10'b0;

   // m126_112 = W*in
   wire signed [9:0] m126_112;
   assign m126_112 ={ {4{in126[5]}} , in126[5:0] };

   // m126_113 = W*in
   wire signed [9:0] m126_113;
   assign m126_113 =10'b0;

   // m126_114 = W*in
   wire signed [9:0] m126_114;
   assign m126_114 =10'b0;

   // m126_115 = W*in
   wire signed [9:0] m126_115;
   assign m126_115 ={ {5{in126[5]}} , in126[5:1] };

   // m126_116 = W*in
   wire signed [9:0] m126_116;
   assign m126_116 ={ {4{neg126[5]}} , neg126[5:0] };

   // m126_117 = W*in
   wire signed [9:0] m126_117;
   assign m126_117 =10'b0;

   // m127_1 = W*in
   wire signed [9:0] m127_1;
   assign m127_1 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_2 = W*in
   wire signed [9:0] m127_2;
   assign m127_2 =10'b0;

   // m127_3 = W*in
   wire signed [9:0] m127_3;
   assign m127_3 =10'b0;

   // m127_4 = W*in
   wire signed [9:0] m127_4;
   assign m127_4 =10'b0;

   // m127_5 = W*in
   wire signed [9:0] m127_5;
   assign m127_5 =10'b0;

   // m127_6 = W*in
   wire signed [9:0] m127_6;
   assign m127_6 ={ {4{in127[5]}} , in127[5:0] };

   // m127_7 = W*in
   wire signed [9:0] m127_7;
   assign m127_7 =10'b0;

   // m127_8 = W*in
   wire signed [9:0] m127_8;
   assign m127_8 =10'b0;

   // m127_9 = W*in
   wire signed [9:0] m127_9;
   assign m127_9 =10'b0;

   // m127_10 = W*in
   wire signed [9:0] m127_10;
   assign m127_10 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_11 = W*in
   wire signed [9:0] m127_11;
   assign m127_11 =10'b0;

   // m127_12 = W*in
   wire signed [9:0] m127_12;
   assign m127_12 =10'b0;

   // m127_13 = W*in
   wire signed [9:0] m127_13;
   assign m127_13 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_14 = W*in
   wire signed [9:0] m127_14;
   assign m127_14 =10'b0;

   // m127_15 = W*in
   wire signed [9:0] m127_15;
   assign m127_15 =10'b0;

   // m127_16 = W*in
   wire signed [9:0] m127_16;
   assign m127_16 =10'b0;

   // m127_17 = W*in
   wire signed [9:0] m127_17;
   assign m127_17 =10'b0;

   // m127_18 = W*in
   wire signed [9:0] m127_18;
   assign m127_18 ={ {5{in127[5]}} , in127[5:1] };

   // m127_19 = W*in
   wire signed [9:0] m127_19;
   assign m127_19 =10'b0;

   // m127_20 = W*in
   wire signed [9:0] m127_20;
   assign m127_20 ={ {5{in127[5]}} , in127[5:1] };

   // m127_21 = W*in
   wire signed [9:0] m127_21;
   assign m127_21 =10'b0;

   // m127_22 = W*in
   wire signed [9:0] m127_22;
   assign m127_22 =10'b0;

   // m127_23 = W*in
   wire signed [9:0] m127_23;
   assign m127_23 ={ {4{in127[5]}} , in127[5:0] };

   // m127_24 = W*in
   wire signed [9:0] m127_24;
   assign m127_24 =10'b0;

   // m127_25 = W*in
   wire signed [9:0] m127_25;
   assign m127_25 =10'b0;

   // m127_26 = W*in
   wire signed [9:0] m127_26;
   assign m127_26 ={ {5{in127[5]}} , in127[5:1] };

   // m127_27 = W*in
   wire signed [9:0] m127_27;
   assign m127_27 =10'b0;

   // m127_28 = W*in
   wire signed [9:0] m127_28;
   assign m127_28 =10'b0;

   // m127_29 = W*in
   wire signed [9:0] m127_29;
   assign m127_29 =10'b0;

   // m127_30 = W*in
   wire signed [9:0] m127_30;
   assign m127_30 ={ {5{in127[5]}} , in127[5:1] };

   // m127_31 = W*in
   wire signed [9:0] m127_31;
   assign m127_31 ={ {5{neg127[5]}} , neg127[5:1] };

   // m127_32 = W*in
   wire signed [9:0] m127_32;
   assign m127_32 =10'b0;

   // m127_33 = W*in
   wire signed [9:0] m127_33;
   assign m127_33 =10'b0;

   // m127_34 = W*in
   wire signed [9:0] m127_34;
   assign m127_34 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_35 = W*in
   wire signed [9:0] m127_35;
   assign m127_35 ={ {5{in127[5]}} , in127[5:1] };

   // m127_36 = W*in
   wire signed [9:0] m127_36;
   assign m127_36 =10'b0;

   // m127_37 = W*in
   wire signed [9:0] m127_37;
   assign m127_37 ={ {5{neg127[5]}} , neg127[5:1] };

   // m127_38 = W*in
   wire signed [9:0] m127_38;
   assign m127_38 ={ {4{in127[5]}} , in127[5:0] };

   // m127_39 = W*in
   wire signed [9:0] m127_39;
   assign m127_39 =10'b0;

   // m127_40 = W*in
   wire signed [9:0] m127_40;
   assign m127_40 =10'b0;

   // m127_41 = W*in
   wire signed [9:0] m127_41;
   assign m127_41 =10'b0;

   // m127_42 = W*in
   wire signed [9:0] m127_42;
   assign m127_42 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_43 = W*in
   wire signed [9:0] m127_43;
   assign m127_43 =10'b0;

   // m127_44 = W*in
   wire signed [9:0] m127_44;
   assign m127_44 =10'b0;

   // m127_45 = W*in
   wire signed [9:0] m127_45;
   assign m127_45 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_46 = W*in
   wire signed [9:0] m127_46;
   assign m127_46 =10'b0;

   // m127_47 = W*in
   wire signed [9:0] m127_47;
   assign m127_47 =10'b0;

   // m127_48 = W*in
   wire signed [9:0] m127_48;
   assign m127_48 =10'b0;

   // m127_49 = W*in
   wire signed [9:0] m127_49;
   assign m127_49 =10'b0;

   // m127_50 = W*in
   wire signed [9:0] m127_50;
   assign m127_50 =10'b0;

   // m127_51 = W*in
   wire signed [9:0] m127_51;
   assign m127_51 =10'b0;

   // m127_52 = W*in
   wire signed [9:0] m127_52;
   assign m127_52 =10'b0;

   // m127_53 = W*in
   wire signed [9:0] m127_53;
   assign m127_53 =10'b0;

   // m127_54 = W*in
   wire signed [9:0] m127_54;
   assign m127_54 =10'b0;

   // m127_55 = W*in
   wire signed [9:0] m127_55;
   assign m127_55 =10'b0;

   // m127_56 = W*in
   wire signed [9:0] m127_56;
   assign m127_56 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_57 = W*in
   wire signed [9:0] m127_57;
   assign m127_57 =10'b0;

   // m127_58 = W*in
   wire signed [9:0] m127_58;
   assign m127_58 =10'b0;

   // m127_59 = W*in
   wire signed [9:0] m127_59;
   assign m127_59 =10'b0;

   // m127_60 = W*in
   wire signed [9:0] m127_60;
   assign m127_60 =10'b0;

   // m127_61 = W*in
   wire signed [9:0] m127_61;
   assign m127_61 ={ {5{neg127[5]}} , neg127[5:1] };

   // m127_62 = W*in
   wire signed [9:0] m127_62;
   assign m127_62 =10'b0;

   // m127_63 = W*in
   wire signed [9:0] m127_63;
   assign m127_63 ={ {4{in127[5]}} , in127[5:0] };

   // m127_64 = W*in
   wire signed [9:0] m127_64;
   assign m127_64 =10'b0;

   // m127_65 = W*in
   wire signed [9:0] m127_65;
   assign m127_65 =10'b0;

   // m127_66 = W*in
   wire signed [9:0] m127_66;
   assign m127_66 =10'b0;

   // m127_67 = W*in
   wire signed [9:0] m127_67;
   assign m127_67 =10'b0;

   // m127_68 = W*in
   wire signed [9:0] m127_68;
   assign m127_68 ={ {4{in127[5]}} , in127[5:0] };

   // m127_69 = W*in
   wire signed [9:0] m127_69;
   assign m127_69 =10'b0;

   // m127_70 = W*in
   wire signed [9:0] m127_70;
   assign m127_70 =10'b0;

   // m127_71 = W*in
   wire signed [9:0] m127_71;
   assign m127_71 =10'b0;

   // m127_72 = W*in
   wire signed [9:0] m127_72;
   assign m127_72 =10'b0;

   // m127_73 = W*in
   wire signed [9:0] m127_73;
   assign m127_73 ={ {5{neg127[5]}} , neg127[5:1] };

   // m127_74 = W*in
   wire signed [9:0] m127_74;
   assign m127_74 ={ {4{in127[5]}} , in127[5:0] };

   // m127_75 = W*in
   wire signed [9:0] m127_75;
   assign m127_75 =10'b0;

   // m127_76 = W*in
   wire signed [9:0] m127_76;
   assign m127_76 =10'b0;

   // m127_77 = W*in
   wire signed [9:0] m127_77;
   assign m127_77 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_78 = W*in
   wire signed [9:0] m127_78;
   assign m127_78 ={ {5{in127[5]}} , in127[5:1] };

   // m127_79 = W*in
   wire signed [9:0] m127_79;
   assign m127_79 =10'b0;

   // m127_80 = W*in
   wire signed [9:0] m127_80;
   assign m127_80 =10'b0;

   // m127_81 = W*in
   wire signed [9:0] m127_81;
   assign m127_81 =10'b0;

   // m127_82 = W*in
   wire signed [9:0] m127_82;
   assign m127_82 =10'b0;

   // m127_83 = W*in
   wire signed [9:0] m127_83;
   assign m127_83 =10'b0;

   // m127_84 = W*in
   wire signed [9:0] m127_84;
   assign m127_84 =10'b0;

   // m127_85 = W*in
   wire signed [9:0] m127_85;
   assign m127_85 =10'b0;

   // m127_86 = W*in
   wire signed [9:0] m127_86;
   assign m127_86 ={ {5{in127[5]}} , in127[5:1] };

   // m127_87 = W*in
   wire signed [9:0] m127_87;
   assign m127_87 =10'b0;

   // m127_88 = W*in
   wire signed [9:0] m127_88;
   assign m127_88 =10'b0;

   // m127_89 = W*in
   wire signed [9:0] m127_89;
   assign m127_89 ={ {4{neg127[5]}} , neg127[5:0] };

   // m127_90 = W*in
   wire signed [9:0] m127_90;
   assign m127_90 =10'b0;

   // m127_91 = W*in
   wire signed [9:0] m127_91;
   assign m127_91 =10'b0;

   // m127_92 = W*in
   wire signed [9:0] m127_92;
   assign m127_92 =10'b0;

   // m127_93 = W*in
   wire signed [9:0] m127_93;
   assign m127_93 =10'b0;

   // m127_94 = W*in
   wire signed [9:0] m127_94;
   assign m127_94 ={ {3{in127[5]}} , in127 , {1{1'b0}} };

   // m127_95 = W*in
   wire signed [9:0] m127_95;
   assign m127_95 =10'b0;

   // m127_96 = W*in
   wire signed [9:0] m127_96;
   assign m127_96 =10'b0;

   // m127_97 = W*in
   wire signed [9:0] m127_97;
   assign m127_97 =10'b0;

   // m127_98 = W*in
   wire signed [9:0] m127_98;
   assign m127_98 =10'b0;

   // m127_99 = W*in
   wire signed [9:0] m127_99;
   assign m127_99 =10'b0;

   // m127_100 = W*in
   wire signed [9:0] m127_100;
   assign m127_100 =10'b0;

   // m127_101 = W*in
   wire signed [9:0] m127_101;
   assign m127_101 =10'b0;

   // m127_102 = W*in
   wire signed [9:0] m127_102;
   assign m127_102 =10'b0;

   // m127_103 = W*in
   wire signed [9:0] m127_103;
   assign m127_103 =10'b0;

   // m127_104 = W*in
   wire signed [9:0] m127_104;
   assign m127_104 =10'b0;

   // m127_105 = W*in
   wire signed [9:0] m127_105;
   assign m127_105 =10'b0;

   // m127_106 = W*in
   wire signed [9:0] m127_106;
   assign m127_106 =10'b0;

   // m127_107 = W*in
   wire signed [9:0] m127_107;
   assign m127_107 =10'b0;

   // m127_108 = W*in
   wire signed [9:0] m127_108;
   assign m127_108 ={ {5{in127[5]}} , in127[5:1] };

   // m127_109 = W*in
   wire signed [9:0] m127_109;
   assign m127_109 =10'b0;

   // m127_110 = W*in
   wire signed [9:0] m127_110;
   assign m127_110 =10'b0;

   // m127_111 = W*in
   wire signed [9:0] m127_111;
   assign m127_111 =10'b0;

   // m127_112 = W*in
   wire signed [9:0] m127_112;
   assign m127_112 ={ {4{in127[5]}} , in127[5:0] };

   // m127_113 = W*in
   wire signed [9:0] m127_113;
   assign m127_113 =10'b0;

   // m127_114 = W*in
   wire signed [9:0] m127_114;
   assign m127_114 =10'b0;

   // m127_115 = W*in
   wire signed [9:0] m127_115;
   assign m127_115 =10'b0;

   // m127_116 = W*in
   wire signed [9:0] m127_116;
   assign m127_116 =10'b0;

   // m127_117 = W*in
   wire signed [9:0] m127_117;
   assign m127_117 =10'b0;

   // m128_1 = W*in
   wire signed [9:0] m128_1;
   assign m128_1 =10'b0;

   // m128_2 = W*in
   wire signed [9:0] m128_2;
   assign m128_2 =10'b0;

   // m128_3 = W*in
   wire signed [9:0] m128_3;
   assign m128_3 =10'b0;

   // m128_4 = W*in
   wire signed [9:0] m128_4;
   assign m128_4 =10'b0;

   // m128_5 = W*in
   wire signed [9:0] m128_5;
   assign m128_5 =10'b0;

   // m128_6 = W*in
   wire signed [9:0] m128_6;
   assign m128_6 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_7 = W*in
   wire signed [9:0] m128_7;
   assign m128_7 =10'b0;

   // m128_8 = W*in
   wire signed [9:0] m128_8;
   assign m128_8 =10'b0;

   // m128_9 = W*in
   wire signed [9:0] m128_9;
   assign m128_9 =10'b0;

   // m128_10 = W*in
   wire signed [9:0] m128_10;
   assign m128_10 =10'b0;

   // m128_11 = W*in
   wire signed [9:0] m128_11;
   assign m128_11 =10'b0;

   // m128_12 = W*in
   wire signed [9:0] m128_12;
   assign m128_12 =10'b0;

   // m128_13 = W*in
   wire signed [9:0] m128_13;
   assign m128_13 =10'b0;

   // m128_14 = W*in
   wire signed [9:0] m128_14;
   assign m128_14 =10'b0;

   // m128_15 = W*in
   wire signed [9:0] m128_15;
   assign m128_15 =10'b0;

   // m128_16 = W*in
   wire signed [9:0] m128_16;
   assign m128_16 ={ {4{in128[5]}} , in128[5:0] };

   // m128_17 = W*in
   wire signed [9:0] m128_17;
   assign m128_17 =10'b0;

   // m128_18 = W*in
   wire signed [9:0] m128_18;
   assign m128_18 =10'b0;

   // m128_19 = W*in
   wire signed [9:0] m128_19;
   assign m128_19 =10'b0;

   // m128_20 = W*in
   wire signed [9:0] m128_20;
   assign m128_20 =10'b0;

   // m128_21 = W*in
   wire signed [9:0] m128_21;
   assign m128_21 ={ {5{in128[5]}} , in128[5:1] };

   // m128_22 = W*in
   wire signed [9:0] m128_22;
   assign m128_22 ={ {5{in128[5]}} , in128[5:1] };

   // m128_23 = W*in
   wire signed [9:0] m128_23;
   assign m128_23 =10'b0;

   // m128_24 = W*in
   wire signed [9:0] m128_24;
   assign m128_24 =10'b0;

   // m128_25 = W*in
   wire signed [9:0] m128_25;
   assign m128_25 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_26 = W*in
   wire signed [9:0] m128_26;
   assign m128_26 =10'b0;

   // m128_27 = W*in
   wire signed [9:0] m128_27;
   assign m128_27 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_28 = W*in
   wire signed [9:0] m128_28;
   assign m128_28 =10'b0;

   // m128_29 = W*in
   wire signed [9:0] m128_29;
   assign m128_29 =10'b0;

   // m128_30 = W*in
   wire signed [9:0] m128_30;
   assign m128_30 =10'b0;

   // m128_31 = W*in
   wire signed [9:0] m128_31;
   assign m128_31 ={ {5{in128[5]}} , in128[5:1] };

   // m128_32 = W*in
   wire signed [9:0] m128_32;
   assign m128_32 =10'b0;

   // m128_33 = W*in
   wire signed [9:0] m128_33;
   assign m128_33 =10'b0;

   // m128_34 = W*in
   wire signed [9:0] m128_34;
   assign m128_34 =10'b0;

   // m128_35 = W*in
   wire signed [9:0] m128_35;
   assign m128_35 =10'b0;

   // m128_36 = W*in
   wire signed [9:0] m128_36;
   assign m128_36 ={ {5{in128[5]}} , in128[5:1] };

   // m128_37 = W*in
   wire signed [9:0] m128_37;
   assign m128_37 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_38 = W*in
   wire signed [9:0] m128_38;
   assign m128_38 =10'b0;

   // m128_39 = W*in
   wire signed [9:0] m128_39;
   assign m128_39 =10'b0;

   // m128_40 = W*in
   wire signed [9:0] m128_40;
   assign m128_40 =10'b0;

   // m128_41 = W*in
   wire signed [9:0] m128_41;
   assign m128_41 =10'b0;

   // m128_42 = W*in
   wire signed [9:0] m128_42;
   assign m128_42 =10'b0;

   // m128_43 = W*in
   wire signed [9:0] m128_43;
   assign m128_43 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_44 = W*in
   wire signed [9:0] m128_44;
   assign m128_44 =10'b0;

   // m128_45 = W*in
   wire signed [9:0] m128_45;
   assign m128_45 ={ {4{in128[5]}} , in128[5:0] };

   // m128_46 = W*in
   wire signed [9:0] m128_46;
   assign m128_46 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_47 = W*in
   wire signed [9:0] m128_47;
   assign m128_47 =10'b0;

   // m128_48 = W*in
   wire signed [9:0] m128_48;
   assign m128_48 =10'b0;

   // m128_49 = W*in
   wire signed [9:0] m128_49;
   assign m128_49 =10'b0;

   // m128_50 = W*in
   wire signed [9:0] m128_50;
   assign m128_50 =10'b0;

   // m128_51 = W*in
   wire signed [9:0] m128_51;
   assign m128_51 =10'b0;

   // m128_52 = W*in
   wire signed [9:0] m128_52;
   assign m128_52 =10'b0;

   // m128_53 = W*in
   wire signed [9:0] m128_53;
   assign m128_53 =10'b0;

   // m128_54 = W*in
   wire signed [9:0] m128_54;
   assign m128_54 =10'b0;

   // m128_55 = W*in
   wire signed [9:0] m128_55;
   assign m128_55 =10'b0;

   // m128_56 = W*in
   wire signed [9:0] m128_56;
   assign m128_56 =10'b0;

   // m128_57 = W*in
   wire signed [9:0] m128_57;
   assign m128_57 =10'b0;

   // m128_58 = W*in
   wire signed [9:0] m128_58;
   assign m128_58 ={ {5{neg128[5]}} , neg128[5:1] };

   // m128_59 = W*in
   wire signed [9:0] m128_59;
   assign m128_59 =10'b0;

   // m128_60 = W*in
   wire signed [9:0] m128_60;
   assign m128_60 =10'b0;

   // m128_61 = W*in
   wire signed [9:0] m128_61;
   assign m128_61 =10'b0;

   // m128_62 = W*in
   wire signed [9:0] m128_62;
   assign m128_62 =10'b0;

   // m128_63 = W*in
   wire signed [9:0] m128_63;
   assign m128_63 =10'b0;

   // m128_64 = W*in
   wire signed [9:0] m128_64;
   assign m128_64 ={ {5{in128[5]}} , in128[5:1] };

   // m128_65 = W*in
   wire signed [9:0] m128_65;
   assign m128_65 =10'b0;

   // m128_66 = W*in
   wire signed [9:0] m128_66;
   assign m128_66 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_67 = W*in
   wire signed [9:0] m128_67;
   assign m128_67 =10'b0;

   // m128_68 = W*in
   wire signed [9:0] m128_68;
   assign m128_68 ={ {5{in128[5]}} , in128[5:1] };

   // m128_69 = W*in
   wire signed [9:0] m128_69;
   assign m128_69 =10'b0;

   // m128_70 = W*in
   wire signed [9:0] m128_70;
   assign m128_70 =10'b0;

   // m128_71 = W*in
   wire signed [9:0] m128_71;
   assign m128_71 ={ {5{neg128[5]}} , neg128[5:1] };

   // m128_72 = W*in
   wire signed [9:0] m128_72;
   assign m128_72 =10'b0;

   // m128_73 = W*in
   wire signed [9:0] m128_73;
   assign m128_73 =10'b0;

   // m128_74 = W*in
   wire signed [9:0] m128_74;
   assign m128_74 ={ {5{neg128[5]}} , neg128[5:1] };

   // m128_75 = W*in
   wire signed [9:0] m128_75;
   assign m128_75 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_76 = W*in
   wire signed [9:0] m128_76;
   assign m128_76 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_77 = W*in
   wire signed [9:0] m128_77;
   assign m128_77 ={ {4{in128[5]}} , in128[5:0] };

   // m128_78 = W*in
   wire signed [9:0] m128_78;
   assign m128_78 ={ {5{neg128[5]}} , neg128[5:1] };

   // m128_79 = W*in
   wire signed [9:0] m128_79;
   assign m128_79 =10'b0;

   // m128_80 = W*in
   wire signed [9:0] m128_80;
   assign m128_80 ={ {4{in128[5]}} , in128[5:0] };

   // m128_81 = W*in
   wire signed [9:0] m128_81;
   assign m128_81 =10'b0;

   // m128_82 = W*in
   wire signed [9:0] m128_82;
   assign m128_82 =10'b0;

   // m128_83 = W*in
   wire signed [9:0] m128_83;
   assign m128_83 =10'b0;

   // m128_84 = W*in
   wire signed [9:0] m128_84;
   assign m128_84 =10'b0;

   // m128_85 = W*in
   wire signed [9:0] m128_85;
   assign m128_85 =10'b0;

   // m128_86 = W*in
   wire signed [9:0] m128_86;
   assign m128_86 ={ {5{in128[5]}} , in128[5:1] };

   // m128_87 = W*in
   wire signed [9:0] m128_87;
   assign m128_87 =10'b0;

   // m128_88 = W*in
   wire signed [9:0] m128_88;
   assign m128_88 =10'b0;

   // m128_89 = W*in
   wire signed [9:0] m128_89;
   assign m128_89 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_90 = W*in
   wire signed [9:0] m128_90;
   assign m128_90 ={ {4{in128[5]}} , in128[5:0] };

   // m128_91 = W*in
   wire signed [9:0] m128_91;
   assign m128_91 ={ {4{in128[5]}} , in128[5:0] };

   // m128_92 = W*in
   wire signed [9:0] m128_92;
   assign m128_92 =10'b0;

   // m128_93 = W*in
   wire signed [9:0] m128_93;
   assign m128_93 =10'b0;

   // m128_94 = W*in
   wire signed [9:0] m128_94;
   assign m128_94 =10'b0;

   // m128_95 = W*in
   wire signed [9:0] m128_95;
   assign m128_95 =10'b0;

   // m128_96 = W*in
   wire signed [9:0] m128_96;
   assign m128_96 =10'b0;

   // m128_97 = W*in
   wire signed [9:0] m128_97;
   assign m128_97 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_98 = W*in
   wire signed [9:0] m128_98;
   assign m128_98 ={ {4{in128[5]}} , in128[5:0] };

   // m128_99 = W*in
   wire signed [9:0] m128_99;
   assign m128_99 =10'b0;

   // m128_100 = W*in
   wire signed [9:0] m128_100;
   assign m128_100 ={ {4{neg128[5]}} , neg128[5:0] };

   // m128_101 = W*in
   wire signed [9:0] m128_101;
   assign m128_101 =10'b0;

   // m128_102 = W*in
   wire signed [9:0] m128_102;
   assign m128_102 =10'b0;

   // m128_103 = W*in
   wire signed [9:0] m128_103;
   assign m128_103 =10'b0;

   // m128_104 = W*in
   wire signed [9:0] m128_104;
   assign m128_104 =10'b0;

   // m128_105 = W*in
   wire signed [9:0] m128_105;
   assign m128_105 =10'b0;

   // m128_106 = W*in
   wire signed [9:0] m128_106;
   assign m128_106 =10'b0;

   // m128_107 = W*in
   wire signed [9:0] m128_107;
   assign m128_107 =10'b0;

   // m128_108 = W*in
   wire signed [9:0] m128_108;
   assign m128_108 ={ {5{neg128[5]}} , neg128[5:1] };

   // m128_109 = W*in
   wire signed [9:0] m128_109;
   assign m128_109 =10'b0;

   // m128_110 = W*in
   wire signed [9:0] m128_110;
   assign m128_110 =10'b0;

   // m128_111 = W*in
   wire signed [9:0] m128_111;
   assign m128_111 =10'b0;

   // m128_112 = W*in
   wire signed [9:0] m128_112;
   assign m128_112 =10'b0;

   // m128_113 = W*in
   wire signed [9:0] m128_113;
   assign m128_113 =10'b0;

   // m128_114 = W*in
   wire signed [9:0] m128_114;
   assign m128_114 =10'b0;

   // m128_115 = W*in
   wire signed [9:0] m128_115;
   assign m128_115 =10'b0;

   // m128_116 = W*in
   wire signed [9:0] m128_116;
   assign m128_116 =10'b0;

   // m128_117 = W*in
   wire signed [9:0] m128_117;
   assign m128_117 ={ {4{neg128[5]}} , neg128[5:0] };

   // m129_1 = W*in
   wire signed [9:0] m129_1;
   assign m129_1 =10'b0;

   // m129_2 = W*in
   wire signed [9:0] m129_2;
   assign m129_2 =10'b0;

   // m129_3 = W*in
   wire signed [9:0] m129_3;
   assign m129_3 =10'b0;

   // m129_4 = W*in
   wire signed [9:0] m129_4;
   assign m129_4 =10'b0;

   // m129_5 = W*in
   wire signed [9:0] m129_5;
   assign m129_5 =10'b0;

   // m129_6 = W*in
   wire signed [9:0] m129_6;
   assign m129_6 =10'b0;

   // m129_7 = W*in
   wire signed [9:0] m129_7;
   assign m129_7 ={ {3{in129[5]}} , in129 , {1{1'b0}} };

   // m129_8 = W*in
   wire signed [9:0] m129_8;
   assign m129_8 =10'b0;

   // m129_9 = W*in
   wire signed [9:0] m129_9;
   assign m129_9 =10'b0;

   // m129_10 = W*in
   wire signed [9:0] m129_10;
   assign m129_10 =10'b0;

   // m129_11 = W*in
   wire signed [9:0] m129_11;
   assign m129_11 =10'b0;

   // m129_12 = W*in
   wire signed [9:0] m129_12;
   assign m129_12 =10'b0;

   // m129_13 = W*in
   wire signed [9:0] m129_13;
   assign m129_13 ={ {4{in129[5]}} , in129[5:0] };

   // m129_14 = W*in
   wire signed [9:0] m129_14;
   assign m129_14 =10'b0;

   // m129_15 = W*in
   wire signed [9:0] m129_15;
   assign m129_15 =10'b0;

   // m129_16 = W*in
   wire signed [9:0] m129_16;
   assign m129_16 ={ {4{in129[5]}} , in129[5:0] };

   // m129_17 = W*in
   wire signed [9:0] m129_17;
   assign m129_17 =10'b0;

   // m129_18 = W*in
   wire signed [9:0] m129_18;
   assign m129_18 =10'b0;

   // m129_19 = W*in
   wire signed [9:0] m129_19;
   assign m129_19 =10'b0;

   // m129_20 = W*in
   wire signed [9:0] m129_20;
   assign m129_20 =10'b0;

   // m129_21 = W*in
   wire signed [9:0] m129_21;
   assign m129_21 =10'b0;

   // m129_22 = W*in
   wire signed [9:0] m129_22;
   assign m129_22 =10'b0;

   // m129_23 = W*in
   wire signed [9:0] m129_23;
   assign m129_23 =10'b0;

   // m129_24 = W*in
   wire signed [9:0] m129_24;
   assign m129_24 =10'b0;

   // m129_25 = W*in
   wire signed [9:0] m129_25;
   assign m129_25 =10'b0;

   // m129_26 = W*in
   wire signed [9:0] m129_26;
   assign m129_26 =10'b0;

   // m129_27 = W*in
   wire signed [9:0] m129_27;
   assign m129_27 =10'b0;

   // m129_28 = W*in
   wire signed [9:0] m129_28;
   assign m129_28 =10'b0;

   // m129_29 = W*in
   wire signed [9:0] m129_29;
   assign m129_29 =10'b0;

   // m129_30 = W*in
   wire signed [9:0] m129_30;
   assign m129_30 =10'b0;

   // m129_31 = W*in
   wire signed [9:0] m129_31;
   assign m129_31 =10'b0;

   // m129_32 = W*in
   wire signed [9:0] m129_32;
   assign m129_32 =10'b0;

   // m129_33 = W*in
   wire signed [9:0] m129_33;
   assign m129_33 ={ {4{in129[5]}} , in129[5:0] };

   // m129_34 = W*in
   wire signed [9:0] m129_34;
   assign m129_34 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_35 = W*in
   wire signed [9:0] m129_35;
   assign m129_35 =10'b0;

   // m129_36 = W*in
   wire signed [9:0] m129_36;
   assign m129_36 ={ {4{in129[5]}} , in129[5:0] };

   // m129_37 = W*in
   wire signed [9:0] m129_37;
   assign m129_37 =10'b0;

   // m129_38 = W*in
   wire signed [9:0] m129_38;
   assign m129_38 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_39 = W*in
   wire signed [9:0] m129_39;
   assign m129_39 =10'b0;

   // m129_40 = W*in
   wire signed [9:0] m129_40;
   assign m129_40 =10'b0;

   // m129_41 = W*in
   wire signed [9:0] m129_41;
   assign m129_41 =10'b0;

   // m129_42 = W*in
   wire signed [9:0] m129_42;
   assign m129_42 ={ {4{in129[5]}} , in129[5:0] };

   // m129_43 = W*in
   wire signed [9:0] m129_43;
   assign m129_43 =10'b0;

   // m129_44 = W*in
   wire signed [9:0] m129_44;
   assign m129_44 =10'b0;

   // m129_45 = W*in
   wire signed [9:0] m129_45;
   assign m129_45 ={ {4{in129[5]}} , in129[5:0] };

   // m129_46 = W*in
   wire signed [9:0] m129_46;
   assign m129_46 =10'b0;

   // m129_47 = W*in
   wire signed [9:0] m129_47;
   assign m129_47 =10'b0;

   // m129_48 = W*in
   wire signed [9:0] m129_48;
   assign m129_48 =10'b0;

   // m129_49 = W*in
   wire signed [9:0] m129_49;
   assign m129_49 =10'b0;

   // m129_50 = W*in
   wire signed [9:0] m129_50;
   assign m129_50 =10'b0;

   // m129_51 = W*in
   wire signed [9:0] m129_51;
   assign m129_51 ={ {4{in129[5]}} , in129[5:0] };

   // m129_52 = W*in
   wire signed [9:0] m129_52;
   assign m129_52 =10'b0;

   // m129_53 = W*in
   wire signed [9:0] m129_53;
   assign m129_53 =10'b0;

   // m129_54 = W*in
   wire signed [9:0] m129_54;
   assign m129_54 =10'b0;

   // m129_55 = W*in
   wire signed [9:0] m129_55;
   assign m129_55 =10'b0;

   // m129_56 = W*in
   wire signed [9:0] m129_56;
   assign m129_56 ={ {4{in129[5]}} , in129[5:0] };

   // m129_57 = W*in
   wire signed [9:0] m129_57;
   assign m129_57 =10'b0;

   // m129_58 = W*in
   wire signed [9:0] m129_58;
   assign m129_58 =10'b0;

   // m129_59 = W*in
   wire signed [9:0] m129_59;
   assign m129_59 =10'b0;

   // m129_60 = W*in
   wire signed [9:0] m129_60;
   assign m129_60 =10'b0;

   // m129_61 = W*in
   wire signed [9:0] m129_61;
   assign m129_61 =10'b0;

   // m129_62 = W*in
   wire signed [9:0] m129_62;
   assign m129_62 =10'b0;

   // m129_63 = W*in
   wire signed [9:0] m129_63;
   assign m129_63 =10'b0;

   // m129_64 = W*in
   wire signed [9:0] m129_64;
   assign m129_64 =10'b0;

   // m129_65 = W*in
   wire signed [9:0] m129_65;
   assign m129_65 =10'b0;

   // m129_66 = W*in
   wire signed [9:0] m129_66;
   assign m129_66 ={ {5{neg129[5]}} , neg129[5:1] };

   // m129_67 = W*in
   wire signed [9:0] m129_67;
   assign m129_67 =10'b0;

   // m129_68 = W*in
   wire signed [9:0] m129_68;
   assign m129_68 =10'b0;

   // m129_69 = W*in
   wire signed [9:0] m129_69;
   assign m129_69 ={ {5{neg129[5]}} , neg129[5:1] };

   // m129_70 = W*in
   wire signed [9:0] m129_70;
   assign m129_70 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_71 = W*in
   wire signed [9:0] m129_71;
   assign m129_71 ={ {5{neg129[5]}} , neg129[5:1] };

   // m129_72 = W*in
   wire signed [9:0] m129_72;
   assign m129_72 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_73 = W*in
   wire signed [9:0] m129_73;
   assign m129_73 ={ {4{in129[5]}} , in129[5:0] };

   // m129_74 = W*in
   wire signed [9:0] m129_74;
   assign m129_74 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_75 = W*in
   wire signed [9:0] m129_75;
   assign m129_75 =10'b0;

   // m129_76 = W*in
   wire signed [9:0] m129_76;
   assign m129_76 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_77 = W*in
   wire signed [9:0] m129_77;
   assign m129_77 =10'b0;

   // m129_78 = W*in
   wire signed [9:0] m129_78;
   assign m129_78 =10'b0;

   // m129_79 = W*in
   wire signed [9:0] m129_79;
   assign m129_79 =10'b0;

   // m129_80 = W*in
   wire signed [9:0] m129_80;
   assign m129_80 =10'b0;

   // m129_81 = W*in
   wire signed [9:0] m129_81;
   assign m129_81 =10'b0;

   // m129_82 = W*in
   wire signed [9:0] m129_82;
   assign m129_82 ={ {5{neg129[5]}} , neg129[5:1] };

   // m129_83 = W*in
   wire signed [9:0] m129_83;
   assign m129_83 =10'b0;

   // m129_84 = W*in
   wire signed [9:0] m129_84;
   assign m129_84 =10'b0;

   // m129_85 = W*in
   wire signed [9:0] m129_85;
   assign m129_85 =10'b0;

   // m129_86 = W*in
   wire signed [9:0] m129_86;
   assign m129_86 =10'b0;

   // m129_87 = W*in
   wire signed [9:0] m129_87;
   assign m129_87 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_88 = W*in
   wire signed [9:0] m129_88;
   assign m129_88 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_89 = W*in
   wire signed [9:0] m129_89;
   assign m129_89 =10'b0;

   // m129_90 = W*in
   wire signed [9:0] m129_90;
   assign m129_90 =10'b0;

   // m129_91 = W*in
   wire signed [9:0] m129_91;
   assign m129_91 =10'b0;

   // m129_92 = W*in
   wire signed [9:0] m129_92;
   assign m129_92 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_93 = W*in
   wire signed [9:0] m129_93;
   assign m129_93 =10'b0;

   // m129_94 = W*in
   wire signed [9:0] m129_94;
   assign m129_94 =10'b0;

   // m129_95 = W*in
   wire signed [9:0] m129_95;
   assign m129_95 =10'b0;

   // m129_96 = W*in
   wire signed [9:0] m129_96;
   assign m129_96 =10'b0;

   // m129_97 = W*in
   wire signed [9:0] m129_97;
   assign m129_97 =10'b0;

   // m129_98 = W*in
   wire signed [9:0] m129_98;
   assign m129_98 =10'b0;

   // m129_99 = W*in
   wire signed [9:0] m129_99;
   assign m129_99 ={ {4{neg129[5]}} , neg129[5:0] };

   // m129_100 = W*in
   wire signed [9:0] m129_100;
   assign m129_100 =10'b0;

   // m129_101 = W*in
   wire signed [9:0] m129_101;
   assign m129_101 =10'b0;

   // m129_102 = W*in
   wire signed [9:0] m129_102;
   assign m129_102 ={ {4{in129[5]}} , in129[5:0] };

   // m129_103 = W*in
   wire signed [9:0] m129_103;
   assign m129_103 =10'b0;

   // m129_104 = W*in
   wire signed [9:0] m129_104;
   assign m129_104 =10'b0;

   // m129_105 = W*in
   wire signed [9:0] m129_105;
   assign m129_105 =10'b0;

   // m129_106 = W*in
   wire signed [9:0] m129_106;
   assign m129_106 =10'b0;

   // m129_107 = W*in
   wire signed [9:0] m129_107;
   assign m129_107 =10'b0;

   // m129_108 = W*in
   wire signed [9:0] m129_108;
   assign m129_108 =10'b0;

   // m129_109 = W*in
   wire signed [9:0] m129_109;
   assign m129_109 =10'b0;

   // m129_110 = W*in
   wire signed [9:0] m129_110;
   assign m129_110 =10'b0;

   // m129_111 = W*in
   wire signed [9:0] m129_111;
   assign m129_111 =10'b0;

   // m129_112 = W*in
   wire signed [9:0] m129_112;
   assign m129_112 =10'b0;

   // m129_113 = W*in
   wire signed [9:0] m129_113;
   assign m129_113 =10'b0;

   // m129_114 = W*in
   wire signed [9:0] m129_114;
   assign m129_114 =10'b0;

   // m129_115 = W*in
   wire signed [9:0] m129_115;
   assign m129_115 =10'b0;

   // m129_116 = W*in
   wire signed [9:0] m129_116;
   assign m129_116 =10'b0;

   // m129_117 = W*in
   wire signed [9:0] m129_117;
   assign m129_117 =10'b0;

   // m130_1 = W*in
   wire signed [9:0] m130_1;
   assign m130_1 =10'b0;

   // m130_2 = W*in
   wire signed [9:0] m130_2;
   assign m130_2 =10'b0;

   // m130_3 = W*in
   wire signed [9:0] m130_3;
   assign m130_3 =10'b0;

   // m130_4 = W*in
   wire signed [9:0] m130_4;
   assign m130_4 =10'b0;

   // m130_5 = W*in
   wire signed [9:0] m130_5;
   assign m130_5 =10'b0;

   // m130_6 = W*in
   wire signed [9:0] m130_6;
   assign m130_6 =10'b0;

   // m130_7 = W*in
   wire signed [9:0] m130_7;
   assign m130_7 =10'b0;

   // m130_8 = W*in
   wire signed [9:0] m130_8;
   assign m130_8 =10'b0;

   // m130_9 = W*in
   wire signed [9:0] m130_9;
   assign m130_9 =10'b0;

   // m130_10 = W*in
   wire signed [9:0] m130_10;
   assign m130_10 =10'b0;

   // m130_11 = W*in
   wire signed [9:0] m130_11;
   assign m130_11 =10'b0;

   // m130_12 = W*in
   wire signed [9:0] m130_12;
   assign m130_12 =10'b0;

   // m130_13 = W*in
   wire signed [9:0] m130_13;
   assign m130_13 =10'b0;

   // m130_14 = W*in
   wire signed [9:0] m130_14;
   assign m130_14 =10'b0;

   // m130_15 = W*in
   wire signed [9:0] m130_15;
   assign m130_15 =10'b0;

   // m130_16 = W*in
   wire signed [9:0] m130_16;
   assign m130_16 =10'b0;

   // m130_17 = W*in
   wire signed [9:0] m130_17;
   assign m130_17 =10'b0;

   // m130_18 = W*in
   wire signed [9:0] m130_18;
   assign m130_18 ={ {5{neg130[5]}} , neg130[5:1] };

   // m130_19 = W*in
   wire signed [9:0] m130_19;
   assign m130_19 =10'b0;

   // m130_20 = W*in
   wire signed [9:0] m130_20;
   assign m130_20 ={ {5{in130[5]}} , in130[5:1] };

   // m130_21 = W*in
   wire signed [9:0] m130_21;
   assign m130_21 =10'b0;

   // m130_22 = W*in
   wire signed [9:0] m130_22;
   assign m130_22 =10'b0;

   // m130_23 = W*in
   wire signed [9:0] m130_23;
   assign m130_23 =10'b0;

   // m130_24 = W*in
   wire signed [9:0] m130_24;
   assign m130_24 =10'b0;

   // m130_25 = W*in
   wire signed [9:0] m130_25;
   assign m130_25 ={ {4{in130[5]}} , in130[5:0] };

   // m130_26 = W*in
   wire signed [9:0] m130_26;
   assign m130_26 ={ {5{in130[5]}} , in130[5:1] };

   // m130_27 = W*in
   wire signed [9:0] m130_27;
   assign m130_27 ={ {5{in130[5]}} , in130[5:1] };

   // m130_28 = W*in
   wire signed [9:0] m130_28;
   assign m130_28 ={ {4{in130[5]}} , in130[5:0] };

   // m130_29 = W*in
   wire signed [9:0] m130_29;
   assign m130_29 ={ {5{neg130[5]}} , neg130[5:1] };

   // m130_30 = W*in
   wire signed [9:0] m130_30;
   assign m130_30 =10'b0;

   // m130_31 = W*in
   wire signed [9:0] m130_31;
   assign m130_31 =10'b0;

   // m130_32 = W*in
   wire signed [9:0] m130_32;
   assign m130_32 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_33 = W*in
   wire signed [9:0] m130_33;
   assign m130_33 ={ {4{in130[5]}} , in130[5:0] };

   // m130_34 = W*in
   wire signed [9:0] m130_34;
   assign m130_34 =10'b0;

   // m130_35 = W*in
   wire signed [9:0] m130_35;
   assign m130_35 =10'b0;

   // m130_36 = W*in
   wire signed [9:0] m130_36;
   assign m130_36 ={ {5{in130[5]}} , in130[5:1] };

   // m130_37 = W*in
   wire signed [9:0] m130_37;
   assign m130_37 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_38 = W*in
   wire signed [9:0] m130_38;
   assign m130_38 =10'b0;

   // m130_39 = W*in
   wire signed [9:0] m130_39;
   assign m130_39 =10'b0;

   // m130_40 = W*in
   wire signed [9:0] m130_40;
   assign m130_40 =10'b0;

   // m130_41 = W*in
   wire signed [9:0] m130_41;
   assign m130_41 =10'b0;

   // m130_42 = W*in
   wire signed [9:0] m130_42;
   assign m130_42 ={ {4{in130[5]}} , in130[5:0] };

   // m130_43 = W*in
   wire signed [9:0] m130_43;
   assign m130_43 =10'b0;

   // m130_44 = W*in
   wire signed [9:0] m130_44;
   assign m130_44 ={ {4{in130[5]}} , in130[5:0] };

   // m130_45 = W*in
   wire signed [9:0] m130_45;
   assign m130_45 =10'b0;

   // m130_46 = W*in
   wire signed [9:0] m130_46;
   assign m130_46 =10'b0;

   // m130_47 = W*in
   wire signed [9:0] m130_47;
   assign m130_47 =10'b0;

   // m130_48 = W*in
   wire signed [9:0] m130_48;
   assign m130_48 =10'b0;

   // m130_49 = W*in
   wire signed [9:0] m130_49;
   assign m130_49 =10'b0;

   // m130_50 = W*in
   wire signed [9:0] m130_50;
   assign m130_50 =10'b0;

   // m130_51 = W*in
   wire signed [9:0] m130_51;
   assign m130_51 =10'b0;

   // m130_52 = W*in
   wire signed [9:0] m130_52;
   assign m130_52 =10'b0;

   // m130_53 = W*in
   wire signed [9:0] m130_53;
   assign m130_53 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_54 = W*in
   wire signed [9:0] m130_54;
   assign m130_54 =10'b0;

   // m130_55 = W*in
   wire signed [9:0] m130_55;
   assign m130_55 =10'b0;

   // m130_56 = W*in
   wire signed [9:0] m130_56;
   assign m130_56 =10'b0;

   // m130_57 = W*in
   wire signed [9:0] m130_57;
   assign m130_57 =10'b0;

   // m130_58 = W*in
   wire signed [9:0] m130_58;
   assign m130_58 =10'b0;

   // m130_59 = W*in
   wire signed [9:0] m130_59;
   assign m130_59 ={ {3{in130[5]}} , in130 , {1{1'b0}} };

   // m130_60 = W*in
   wire signed [9:0] m130_60;
   assign m130_60 =10'b0;

   // m130_61 = W*in
   wire signed [9:0] m130_61;
   assign m130_61 =10'b0;

   // m130_62 = W*in
   wire signed [9:0] m130_62;
   assign m130_62 =10'b0;

   // m130_63 = W*in
   wire signed [9:0] m130_63;
   assign m130_63 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_64 = W*in
   wire signed [9:0] m130_64;
   assign m130_64 ={ {4{in130[5]}} , in130[5:0] };

   // m130_65 = W*in
   wire signed [9:0] m130_65;
   assign m130_65 ={ {5{in130[5]}} , in130[5:1] };

   // m130_66 = W*in
   wire signed [9:0] m130_66;
   assign m130_66 =10'b0;

   // m130_67 = W*in
   wire signed [9:0] m130_67;
   assign m130_67 =10'b0;

   // m130_68 = W*in
   wire signed [9:0] m130_68;
   assign m130_68 =10'b0;

   // m130_69 = W*in
   wire signed [9:0] m130_69;
   assign m130_69 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_70 = W*in
   wire signed [9:0] m130_70;
   assign m130_70 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_71 = W*in
   wire signed [9:0] m130_71;
   assign m130_71 =10'b0;

   // m130_72 = W*in
   wire signed [9:0] m130_72;
   assign m130_72 ={ {5{neg130[5]}} , neg130[5:1] };

   // m130_73 = W*in
   wire signed [9:0] m130_73;
   assign m130_73 ={ {5{in130[5]}} , in130[5:1] };

   // m130_74 = W*in
   wire signed [9:0] m130_74;
   assign m130_74 =10'b0;

   // m130_75 = W*in
   wire signed [9:0] m130_75;
   assign m130_75 =10'b0;

   // m130_76 = W*in
   wire signed [9:0] m130_76;
   assign m130_76 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_77 = W*in
   wire signed [9:0] m130_77;
   assign m130_77 =10'b0;

   // m130_78 = W*in
   wire signed [9:0] m130_78;
   assign m130_78 ={ {5{in130[5]}} , in130[5:1] };

   // m130_79 = W*in
   wire signed [9:0] m130_79;
   assign m130_79 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_80 = W*in
   wire signed [9:0] m130_80;
   assign m130_80 =10'b0;

   // m130_81 = W*in
   wire signed [9:0] m130_81;
   assign m130_81 ={ {4{in130[5]}} , in130[5:0] };

   // m130_82 = W*in
   wire signed [9:0] m130_82;
   assign m130_82 ={ {5{neg130[5]}} , neg130[5:1] };

   // m130_83 = W*in
   wire signed [9:0] m130_83;
   assign m130_83 =10'b0;

   // m130_84 = W*in
   wire signed [9:0] m130_84;
   assign m130_84 =10'b0;

   // m130_85 = W*in
   wire signed [9:0] m130_85;
   assign m130_85 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_86 = W*in
   wire signed [9:0] m130_86;
   assign m130_86 =10'b0;

   // m130_87 = W*in
   wire signed [9:0] m130_87;
   assign m130_87 =10'b0;

   // m130_88 = W*in
   wire signed [9:0] m130_88;
   assign m130_88 =10'b0;

   // m130_89 = W*in
   wire signed [9:0] m130_89;
   assign m130_89 =10'b0;

   // m130_90 = W*in
   wire signed [9:0] m130_90;
   assign m130_90 =10'b0;

   // m130_91 = W*in
   wire signed [9:0] m130_91;
   assign m130_91 =10'b0;

   // m130_92 = W*in
   wire signed [9:0] m130_92;
   assign m130_92 =10'b0;

   // m130_93 = W*in
   wire signed [9:0] m130_93;
   assign m130_93 =10'b0;

   // m130_94 = W*in
   wire signed [9:0] m130_94;
   assign m130_94 =10'b0;

   // m130_95 = W*in
   wire signed [9:0] m130_95;
   assign m130_95 =10'b0;

   // m130_96 = W*in
   wire signed [9:0] m130_96;
   assign m130_96 =10'b0;

   // m130_97 = W*in
   wire signed [9:0] m130_97;
   assign m130_97 ={ {4{in130[5]}} , in130[5:0] };

   // m130_98 = W*in
   wire signed [9:0] m130_98;
   assign m130_98 =10'b0;

   // m130_99 = W*in
   wire signed [9:0] m130_99;
   assign m130_99 =10'b0;

   // m130_100 = W*in
   wire signed [9:0] m130_100;
   assign m130_100 =10'b0;

   // m130_101 = W*in
   wire signed [9:0] m130_101;
   assign m130_101 =10'b0;

   // m130_102 = W*in
   wire signed [9:0] m130_102;
   assign m130_102 ={ {4{in130[5]}} , in130[5:0] };

   // m130_103 = W*in
   wire signed [9:0] m130_103;
   assign m130_103 =10'b0;

   // m130_104 = W*in
   wire signed [9:0] m130_104;
   assign m130_104 =10'b0;

   // m130_105 = W*in
   wire signed [9:0] m130_105;
   assign m130_105 =10'b0;

   // m130_106 = W*in
   wire signed [9:0] m130_106;
   assign m130_106 =10'b0;

   // m130_107 = W*in
   wire signed [9:0] m130_107;
   assign m130_107 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_108 = W*in
   wire signed [9:0] m130_108;
   assign m130_108 =10'b0;

   // m130_109 = W*in
   wire signed [9:0] m130_109;
   assign m130_109 =10'b0;

   // m130_110 = W*in
   wire signed [9:0] m130_110;
   assign m130_110 ={ {4{in130[5]}} , in130[5:0] };

   // m130_111 = W*in
   wire signed [9:0] m130_111;
   assign m130_111 =10'b0;

   // m130_112 = W*in
   wire signed [9:0] m130_112;
   assign m130_112 =10'b0;

   // m130_113 = W*in
   wire signed [9:0] m130_113;
   assign m130_113 =10'b0;

   // m130_114 = W*in
   wire signed [9:0] m130_114;
   assign m130_114 ={ {5{in130[5]}} , in130[5:1] };

   // m130_115 = W*in
   wire signed [9:0] m130_115;
   assign m130_115 =10'b0;

   // m130_116 = W*in
   wire signed [9:0] m130_116;
   assign m130_116 ={ {4{neg130[5]}} , neg130[5:0] };

   // m130_117 = W*in
   wire signed [9:0] m130_117;
   assign m130_117 =10'b0;

   // m131_1 = W*in
   wire signed [9:0] m131_1;
   assign m131_1 ={ {4{in131[5]}} , in131[5:0] };

   // m131_2 = W*in
   wire signed [9:0] m131_2;
   assign m131_2 =10'b0;

   // m131_3 = W*in
   wire signed [9:0] m131_3;
   assign m131_3 =10'b0;

   // m131_4 = W*in
   wire signed [9:0] m131_4;
   assign m131_4 =10'b0;

   // m131_5 = W*in
   wire signed [9:0] m131_5;
   assign m131_5 =10'b0;

   // m131_6 = W*in
   wire signed [9:0] m131_6;
   assign m131_6 =10'b0;

   // m131_7 = W*in
   wire signed [9:0] m131_7;
   assign m131_7 ={ {4{in131[5]}} , in131[5:0] };

   // m131_8 = W*in
   wire signed [9:0] m131_8;
   assign m131_8 =10'b0;

   // m131_9 = W*in
   wire signed [9:0] m131_9;
   assign m131_9 =10'b0;

   // m131_10 = W*in
   wire signed [9:0] m131_10;
   assign m131_10 =10'b0;

   // m131_11 = W*in
   wire signed [9:0] m131_11;
   assign m131_11 ={ {5{neg131[5]}} , neg131[5:1] };

   // m131_12 = W*in
   wire signed [9:0] m131_12;
   assign m131_12 =10'b0;

   // m131_13 = W*in
   wire signed [9:0] m131_13;
   assign m131_13 =10'b0;

   // m131_14 = W*in
   wire signed [9:0] m131_14;
   assign m131_14 =10'b0;

   // m131_15 = W*in
   wire signed [9:0] m131_15;
   assign m131_15 =10'b0;

   // m131_16 = W*in
   wire signed [9:0] m131_16;
   assign m131_16 =10'b0;

   // m131_17 = W*in
   wire signed [9:0] m131_17;
   assign m131_17 ={ {4{in131[5]}} , in131[5:0] };

   // m131_18 = W*in
   wire signed [9:0] m131_18;
   assign m131_18 ={ {4{in131[5]}} , in131[5:0] };

   // m131_19 = W*in
   wire signed [9:0] m131_19;
   assign m131_19 =10'b0;

   // m131_20 = W*in
   wire signed [9:0] m131_20;
   assign m131_20 =10'b0;

   // m131_21 = W*in
   wire signed [9:0] m131_21;
   assign m131_21 ={ {5{neg131[5]}} , neg131[5:1] };

   // m131_22 = W*in
   wire signed [9:0] m131_22;
   assign m131_22 ={ {5{in131[5]}} , in131[5:1] };

   // m131_23 = W*in
   wire signed [9:0] m131_23;
   assign m131_23 =10'b0;

   // m131_24 = W*in
   wire signed [9:0] m131_24;
   assign m131_24 =10'b0;

   // m131_25 = W*in
   wire signed [9:0] m131_25;
   assign m131_25 ={ {4{in131[5]}} , in131[5:0] };

   // m131_26 = W*in
   wire signed [9:0] m131_26;
   assign m131_26 =10'b0;

   // m131_27 = W*in
   wire signed [9:0] m131_27;
   assign m131_27 ={ {3{in131[5]}} , in131 , {1{1'b0}} };

   // m131_28 = W*in
   wire signed [9:0] m131_28;
   assign m131_28 ={ {4{in131[5]}} , in131[5:0] };

   // m131_29 = W*in
   wire signed [9:0] m131_29;
   assign m131_29 ={ {5{in131[5]}} , in131[5:1] };

   // m131_30 = W*in
   wire signed [9:0] m131_30;
   assign m131_30 =10'b0;

   // m131_31 = W*in
   wire signed [9:0] m131_31;
   assign m131_31 =10'b0;

   // m131_32 = W*in
   wire signed [9:0] m131_32;
   assign m131_32 =10'b0;

   // m131_33 = W*in
   wire signed [9:0] m131_33;
   assign m131_33 ={ {4{in131[5]}} , in131[5:0] };

   // m131_34 = W*in
   wire signed [9:0] m131_34;
   assign m131_34 =10'b0;

   // m131_35 = W*in
   wire signed [9:0] m131_35;
   assign m131_35 =10'b0;

   // m131_36 = W*in
   wire signed [9:0] m131_36;
   assign m131_36 ={ {4{in131[5]}} , in131[5:0] };

   // m131_37 = W*in
   wire signed [9:0] m131_37;
   assign m131_37 =10'b0;

   // m131_38 = W*in
   wire signed [9:0] m131_38;
   assign m131_38 =10'b0;

   // m131_39 = W*in
   wire signed [9:0] m131_39;
   assign m131_39 =10'b0;

   // m131_40 = W*in
   wire signed [9:0] m131_40;
   assign m131_40 =10'b0;

   // m131_41 = W*in
   wire signed [9:0] m131_41;
   assign m131_41 =10'b0;

   // m131_42 = W*in
   wire signed [9:0] m131_42;
   assign m131_42 =10'b0;

   // m131_43 = W*in
   wire signed [9:0] m131_43;
   assign m131_43 =10'b0;

   // m131_44 = W*in
   wire signed [9:0] m131_44;
   assign m131_44 =10'b0;

   // m131_45 = W*in
   wire signed [9:0] m131_45;
   assign m131_45 =10'b0;

   // m131_46 = W*in
   wire signed [9:0] m131_46;
   assign m131_46 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_47 = W*in
   wire signed [9:0] m131_47;
   assign m131_47 =10'b0;

   // m131_48 = W*in
   wire signed [9:0] m131_48;
   assign m131_48 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_49 = W*in
   wire signed [9:0] m131_49;
   assign m131_49 =10'b0;

   // m131_50 = W*in
   wire signed [9:0] m131_50;
   assign m131_50 =10'b0;

   // m131_51 = W*in
   wire signed [9:0] m131_51;
   assign m131_51 =10'b0;

   // m131_52 = W*in
   wire signed [9:0] m131_52;
   assign m131_52 =10'b0;

   // m131_53 = W*in
   wire signed [9:0] m131_53;
   assign m131_53 =10'b0;

   // m131_54 = W*in
   wire signed [9:0] m131_54;
   assign m131_54 =10'b0;

   // m131_55 = W*in
   wire signed [9:0] m131_55;
   assign m131_55 =10'b0;

   // m131_56 = W*in
   wire signed [9:0] m131_56;
   assign m131_56 =10'b0;

   // m131_57 = W*in
   wire signed [9:0] m131_57;
   assign m131_57 =10'b0;

   // m131_58 = W*in
   wire signed [9:0] m131_58;
   assign m131_58 =10'b0;

   // m131_59 = W*in
   wire signed [9:0] m131_59;
   assign m131_59 ={ {4{in131[5]}} , in131[5:0] };

   // m131_60 = W*in
   wire signed [9:0] m131_60;
   assign m131_60 ={ {4{in131[5]}} , in131[5:0] };

   // m131_61 = W*in
   wire signed [9:0] m131_61;
   assign m131_61 =10'b0;

   // m131_62 = W*in
   wire signed [9:0] m131_62;
   assign m131_62 =10'b0;

   // m131_63 = W*in
   wire signed [9:0] m131_63;
   assign m131_63 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_64 = W*in
   wire signed [9:0] m131_64;
   assign m131_64 ={ {5{in131[5]}} , in131[5:1] };

   // m131_65 = W*in
   wire signed [9:0] m131_65;
   assign m131_65 =10'b0;

   // m131_66 = W*in
   wire signed [9:0] m131_66;
   assign m131_66 ={ {5{in131[5]}} , in131[5:1] };

   // m131_67 = W*in
   wire signed [9:0] m131_67;
   assign m131_67 =10'b0;

   // m131_68 = W*in
   wire signed [9:0] m131_68;
   assign m131_68 =10'b0;

   // m131_69 = W*in
   wire signed [9:0] m131_69;
   assign m131_69 ={ {5{neg131[5]}} , neg131[5:1] };

   // m131_70 = W*in
   wire signed [9:0] m131_70;
   assign m131_70 =10'b0;

   // m131_71 = W*in
   wire signed [9:0] m131_71;
   assign m131_71 =10'b0;

   // m131_72 = W*in
   wire signed [9:0] m131_72;
   assign m131_72 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_73 = W*in
   wire signed [9:0] m131_73;
   assign m131_73 =10'b0;

   // m131_74 = W*in
   wire signed [9:0] m131_74;
   assign m131_74 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_75 = W*in
   wire signed [9:0] m131_75;
   assign m131_75 =10'b0;

   // m131_76 = W*in
   wire signed [9:0] m131_76;
   assign m131_76 =10'b0;

   // m131_77 = W*in
   wire signed [9:0] m131_77;
   assign m131_77 ={ {4{in131[5]}} , in131[5:0] };

   // m131_78 = W*in
   wire signed [9:0] m131_78;
   assign m131_78 =10'b0;

   // m131_79 = W*in
   wire signed [9:0] m131_79;
   assign m131_79 =10'b0;

   // m131_80 = W*in
   wire signed [9:0] m131_80;
   assign m131_80 =10'b0;

   // m131_81 = W*in
   wire signed [9:0] m131_81;
   assign m131_81 ={ {4{in131[5]}} , in131[5:0] };

   // m131_82 = W*in
   wire signed [9:0] m131_82;
   assign m131_82 =10'b0;

   // m131_83 = W*in
   wire signed [9:0] m131_83;
   assign m131_83 =10'b0;

   // m131_84 = W*in
   wire signed [9:0] m131_84;
   assign m131_84 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_85 = W*in
   wire signed [9:0] m131_85;
   assign m131_85 =10'b0;

   // m131_86 = W*in
   wire signed [9:0] m131_86;
   assign m131_86 =10'b0;

   // m131_87 = W*in
   wire signed [9:0] m131_87;
   assign m131_87 =10'b0;

   // m131_88 = W*in
   wire signed [9:0] m131_88;
   assign m131_88 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_89 = W*in
   wire signed [9:0] m131_89;
   assign m131_89 ={ {3{neg131[5]}} , neg131 , {1{1'b0}} };

   // m131_90 = W*in
   wire signed [9:0] m131_90;
   assign m131_90 =10'b0;

   // m131_91 = W*in
   wire signed [9:0] m131_91;
   assign m131_91 ={ {4{in131[5]}} , in131[5:0] };

   // m131_92 = W*in
   wire signed [9:0] m131_92;
   assign m131_92 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_93 = W*in
   wire signed [9:0] m131_93;
   assign m131_93 =10'b0;

   // m131_94 = W*in
   wire signed [9:0] m131_94;
   assign m131_94 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_95 = W*in
   wire signed [9:0] m131_95;
   assign m131_95 =10'b0;

   // m131_96 = W*in
   wire signed [9:0] m131_96;
   assign m131_96 =10'b0;

   // m131_97 = W*in
   wire signed [9:0] m131_97;
   assign m131_97 ={ {4{in131[5]}} , in131[5:0] };

   // m131_98 = W*in
   wire signed [9:0] m131_98;
   assign m131_98 =10'b0;

   // m131_99 = W*in
   wire signed [9:0] m131_99;
   assign m131_99 =10'b0;

   // m131_100 = W*in
   wire signed [9:0] m131_100;
   assign m131_100 =10'b0;

   // m131_101 = W*in
   wire signed [9:0] m131_101;
   assign m131_101 =10'b0;

   // m131_102 = W*in
   wire signed [9:0] m131_102;
   assign m131_102 =10'b0;

   // m131_103 = W*in
   wire signed [9:0] m131_103;
   assign m131_103 =10'b0;

   // m131_104 = W*in
   wire signed [9:0] m131_104;
   assign m131_104 =10'b0;

   // m131_105 = W*in
   wire signed [9:0] m131_105;
   assign m131_105 =10'b0;

   // m131_106 = W*in
   wire signed [9:0] m131_106;
   assign m131_106 =10'b0;

   // m131_107 = W*in
   wire signed [9:0] m131_107;
   assign m131_107 =10'b0;

   // m131_108 = W*in
   wire signed [9:0] m131_108;
   assign m131_108 ={ {4{neg131[5]}} , neg131[5:0] };

   // m131_109 = W*in
   wire signed [9:0] m131_109;
   assign m131_109 =10'b0;

   // m131_110 = W*in
   wire signed [9:0] m131_110;
   assign m131_110 ={ {4{in131[5]}} , in131[5:0] };

   // m131_111 = W*in
   wire signed [9:0] m131_111;
   assign m131_111 =10'b0;

   // m131_112 = W*in
   wire signed [9:0] m131_112;
   assign m131_112 =10'b0;

   // m131_113 = W*in
   wire signed [9:0] m131_113;
   assign m131_113 =10'b0;

   // m131_114 = W*in
   wire signed [9:0] m131_114;
   assign m131_114 ={ {4{in131[5]}} , in131[5:0] };

   // m131_115 = W*in
   wire signed [9:0] m131_115;
   assign m131_115 =10'b0;

   // m131_116 = W*in
   wire signed [9:0] m131_116;
   assign m131_116 =10'b0;

   // m131_117 = W*in
   wire signed [9:0] m131_117;
   assign m131_117 =10'b0;

   // m132_1 = W*in
   wire signed [9:0] m132_1;
   assign m132_1 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_2 = W*in
   wire signed [9:0] m132_2;
   assign m132_2 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_3 = W*in
   wire signed [9:0] m132_3;
   assign m132_3 =10'b0;

   // m132_4 = W*in
   wire signed [9:0] m132_4;
   assign m132_4 =10'b0;

   // m132_5 = W*in
   wire signed [9:0] m132_5;
   assign m132_5 =10'b0;

   // m132_6 = W*in
   wire signed [9:0] m132_6;
   assign m132_6 =10'b0;

   // m132_7 = W*in
   wire signed [9:0] m132_7;
   assign m132_7 =10'b0;

   // m132_8 = W*in
   wire signed [9:0] m132_8;
   assign m132_8 =10'b0;

   // m132_9 = W*in
   wire signed [9:0] m132_9;
   assign m132_9 =10'b0;

   // m132_10 = W*in
   wire signed [9:0] m132_10;
   assign m132_10 =10'b0;

   // m132_11 = W*in
   wire signed [9:0] m132_11;
   assign m132_11 =10'b0;

   // m132_12 = W*in
   wire signed [9:0] m132_12;
   assign m132_12 =10'b0;

   // m132_13 = W*in
   wire signed [9:0] m132_13;
   assign m132_13 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_14 = W*in
   wire signed [9:0] m132_14;
   assign m132_14 =10'b0;

   // m132_15 = W*in
   wire signed [9:0] m132_15;
   assign m132_15 =10'b0;

   // m132_16 = W*in
   wire signed [9:0] m132_16;
   assign m132_16 =10'b0;

   // m132_17 = W*in
   wire signed [9:0] m132_17;
   assign m132_17 =10'b0;

   // m132_18 = W*in
   wire signed [9:0] m132_18;
   assign m132_18 =10'b0;

   // m132_19 = W*in
   wire signed [9:0] m132_19;
   assign m132_19 ={ {5{in132[5]}} , in132[5:1] };

   // m132_20 = W*in
   wire signed [9:0] m132_20;
   assign m132_20 ={ {4{in132[5]}} , in132[5:0] };

   // m132_21 = W*in
   wire signed [9:0] m132_21;
   assign m132_21 =10'b0;

   // m132_22 = W*in
   wire signed [9:0] m132_22;
   assign m132_22 ={ {5{neg132[5]}} , neg132[5:1] };

   // m132_23 = W*in
   wire signed [9:0] m132_23;
   assign m132_23 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_24 = W*in
   wire signed [9:0] m132_24;
   assign m132_24 ={ {3{neg132[5]}} , neg132 , {1{1'b0}} };

   // m132_25 = W*in
   wire signed [9:0] m132_25;
   assign m132_25 =10'b0;

   // m132_26 = W*in
   wire signed [9:0] m132_26;
   assign m132_26 =10'b0;

   // m132_27 = W*in
   wire signed [9:0] m132_27;
   assign m132_27 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_28 = W*in
   wire signed [9:0] m132_28;
   assign m132_28 =10'b0;

   // m132_29 = W*in
   wire signed [9:0] m132_29;
   assign m132_29 =10'b0;

   // m132_30 = W*in
   wire signed [9:0] m132_30;
   assign m132_30 ={ {4{in132[5]}} , in132[5:0] };

   // m132_31 = W*in
   wire signed [9:0] m132_31;
   assign m132_31 =10'b0;

   // m132_32 = W*in
   wire signed [9:0] m132_32;
   assign m132_32 =10'b0;

   // m132_33 = W*in
   wire signed [9:0] m132_33;
   assign m132_33 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_34 = W*in
   wire signed [9:0] m132_34;
   assign m132_34 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_35 = W*in
   wire signed [9:0] m132_35;
   assign m132_35 ={ {4{in132[5]}} , in132[5:0] };

   // m132_36 = W*in
   wire signed [9:0] m132_36;
   assign m132_36 =10'b0;

   // m132_37 = W*in
   wire signed [9:0] m132_37;
   assign m132_37 =10'b0;

   // m132_38 = W*in
   wire signed [9:0] m132_38;
   assign m132_38 =10'b0;

   // m132_39 = W*in
   wire signed [9:0] m132_39;
   assign m132_39 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_40 = W*in
   wire signed [9:0] m132_40;
   assign m132_40 =10'b0;

   // m132_41 = W*in
   wire signed [9:0] m132_41;
   assign m132_41 =10'b0;

   // m132_42 = W*in
   wire signed [9:0] m132_42;
   assign m132_42 ={ {4{in132[5]}} , in132[5:0] };

   // m132_43 = W*in
   wire signed [9:0] m132_43;
   assign m132_43 =10'b0;

   // m132_44 = W*in
   wire signed [9:0] m132_44;
   assign m132_44 ={ {4{in132[5]}} , in132[5:0] };

   // m132_45 = W*in
   wire signed [9:0] m132_45;
   assign m132_45 =10'b0;

   // m132_46 = W*in
   wire signed [9:0] m132_46;
   assign m132_46 =10'b0;

   // m132_47 = W*in
   wire signed [9:0] m132_47;
   assign m132_47 =10'b0;

   // m132_48 = W*in
   wire signed [9:0] m132_48;
   assign m132_48 =10'b0;

   // m132_49 = W*in
   wire signed [9:0] m132_49;
   assign m132_49 ={ {4{in132[5]}} , in132[5:0] };

   // m132_50 = W*in
   wire signed [9:0] m132_50;
   assign m132_50 =10'b0;

   // m132_51 = W*in
   wire signed [9:0] m132_51;
   assign m132_51 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_52 = W*in
   wire signed [9:0] m132_52;
   assign m132_52 ={ {4{in132[5]}} , in132[5:0] };

   // m132_53 = W*in
   wire signed [9:0] m132_53;
   assign m132_53 ={ {4{in132[5]}} , in132[5:0] };

   // m132_54 = W*in
   wire signed [9:0] m132_54;
   assign m132_54 =10'b0;

   // m132_55 = W*in
   wire signed [9:0] m132_55;
   assign m132_55 =10'b0;

   // m132_56 = W*in
   wire signed [9:0] m132_56;
   assign m132_56 =10'b0;

   // m132_57 = W*in
   wire signed [9:0] m132_57;
   assign m132_57 =10'b0;

   // m132_58 = W*in
   wire signed [9:0] m132_58;
   assign m132_58 =10'b0;

   // m132_59 = W*in
   wire signed [9:0] m132_59;
   assign m132_59 =10'b0;

   // m132_60 = W*in
   wire signed [9:0] m132_60;
   assign m132_60 =10'b0;

   // m132_61 = W*in
   wire signed [9:0] m132_61;
   assign m132_61 ={ {3{in132[5]}} , in132 , {1{1'b0}} };

   // m132_62 = W*in
   wire signed [9:0] m132_62;
   assign m132_62 =10'b0;

   // m132_63 = W*in
   wire signed [9:0] m132_63;
   assign m132_63 ={ {4{in132[5]}} , in132[5:0] };

   // m132_64 = W*in
   wire signed [9:0] m132_64;
   assign m132_64 =10'b0;

   // m132_65 = W*in
   wire signed [9:0] m132_65;
   assign m132_65 =10'b0;

   // m132_66 = W*in
   wire signed [9:0] m132_66;
   assign m132_66 =10'b0;

   // m132_67 = W*in
   wire signed [9:0] m132_67;
   assign m132_67 ={ {4{in132[5]}} , in132[5:0] };

   // m132_68 = W*in
   wire signed [9:0] m132_68;
   assign m132_68 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_69 = W*in
   wire signed [9:0] m132_69;
   assign m132_69 =10'b0;

   // m132_70 = W*in
   wire signed [9:0] m132_70;
   assign m132_70 =10'b0;

   // m132_71 = W*in
   wire signed [9:0] m132_71;
   assign m132_71 =10'b0;

   // m132_72 = W*in
   wire signed [9:0] m132_72;
   assign m132_72 =10'b0;

   // m132_73 = W*in
   wire signed [9:0] m132_73;
   assign m132_73 ={ {5{neg132[5]}} , neg132[5:1] };

   // m132_74 = W*in
   wire signed [9:0] m132_74;
   assign m132_74 =10'b0;

   // m132_75 = W*in
   wire signed [9:0] m132_75;
   assign m132_75 ={ {5{in132[5]}} , in132[5:1] };

   // m132_76 = W*in
   wire signed [9:0] m132_76;
   assign m132_76 ={ {4{in132[5]}} , in132[5:0] };

   // m132_77 = W*in
   wire signed [9:0] m132_77;
   assign m132_77 =10'b0;

   // m132_78 = W*in
   wire signed [9:0] m132_78;
   assign m132_78 =10'b0;

   // m132_79 = W*in
   wire signed [9:0] m132_79;
   assign m132_79 =10'b0;

   // m132_80 = W*in
   wire signed [9:0] m132_80;
   assign m132_80 =10'b0;

   // m132_81 = W*in
   wire signed [9:0] m132_81;
   assign m132_81 ={ {4{in132[5]}} , in132[5:0] };

   // m132_82 = W*in
   wire signed [9:0] m132_82;
   assign m132_82 ={ {3{in132[5]}} , in132 , {1{1'b0}} };

   // m132_83 = W*in
   wire signed [9:0] m132_83;
   assign m132_83 =10'b0;

   // m132_84 = W*in
   wire signed [9:0] m132_84;
   assign m132_84 =10'b0;

   // m132_85 = W*in
   wire signed [9:0] m132_85;
   assign m132_85 =10'b0;

   // m132_86 = W*in
   wire signed [9:0] m132_86;
   assign m132_86 =10'b0;

   // m132_87 = W*in
   wire signed [9:0] m132_87;
   assign m132_87 =10'b0;

   // m132_88 = W*in
   wire signed [9:0] m132_88;
   assign m132_88 =10'b0;

   // m132_89 = W*in
   wire signed [9:0] m132_89;
   assign m132_89 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_90 = W*in
   wire signed [9:0] m132_90;
   assign m132_90 =10'b0;

   // m132_91 = W*in
   wire signed [9:0] m132_91;
   assign m132_91 ={ {4{in132[5]}} , in132[5:0] };

   // m132_92 = W*in
   wire signed [9:0] m132_92;
   assign m132_92 =10'b0;

   // m132_93 = W*in
   wire signed [9:0] m132_93;
   assign m132_93 =10'b0;

   // m132_94 = W*in
   wire signed [9:0] m132_94;
   assign m132_94 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_95 = W*in
   wire signed [9:0] m132_95;
   assign m132_95 =10'b0;

   // m132_96 = W*in
   wire signed [9:0] m132_96;
   assign m132_96 =10'b0;

   // m132_97 = W*in
   wire signed [9:0] m132_97;
   assign m132_97 ={ {4{in132[5]}} , in132[5:0] };

   // m132_98 = W*in
   wire signed [9:0] m132_98;
   assign m132_98 =10'b0;

   // m132_99 = W*in
   wire signed [9:0] m132_99;
   assign m132_99 =10'b0;

   // m132_100 = W*in
   wire signed [9:0] m132_100;
   assign m132_100 =10'b0;

   // m132_101 = W*in
   wire signed [9:0] m132_101;
   assign m132_101 =10'b0;

   // m132_102 = W*in
   wire signed [9:0] m132_102;
   assign m132_102 =10'b0;

   // m132_103 = W*in
   wire signed [9:0] m132_103;
   assign m132_103 =10'b0;

   // m132_104 = W*in
   wire signed [9:0] m132_104;
   assign m132_104 =10'b0;

   // m132_105 = W*in
   wire signed [9:0] m132_105;
   assign m132_105 =10'b0;

   // m132_106 = W*in
   wire signed [9:0] m132_106;
   assign m132_106 ={ {4{in132[5]}} , in132[5:0] };

   // m132_107 = W*in
   wire signed [9:0] m132_107;
   assign m132_107 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_108 = W*in
   wire signed [9:0] m132_108;
   assign m132_108 =10'b0;

   // m132_109 = W*in
   wire signed [9:0] m132_109;
   assign m132_109 =10'b0;

   // m132_110 = W*in
   wire signed [9:0] m132_110;
   assign m132_110 =10'b0;

   // m132_111 = W*in
   wire signed [9:0] m132_111;
   assign m132_111 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_112 = W*in
   wire signed [9:0] m132_112;
   assign m132_112 =10'b0;

   // m132_113 = W*in
   wire signed [9:0] m132_113;
   assign m132_113 =10'b0;

   // m132_114 = W*in
   wire signed [9:0] m132_114;
   assign m132_114 ={ {4{neg132[5]}} , neg132[5:0] };

   // m132_115 = W*in
   wire signed [9:0] m132_115;
   assign m132_115 ={ {4{in132[5]}} , in132[5:0] };

   // m132_116 = W*in
   wire signed [9:0] m132_116;
   assign m132_116 =10'b0;

   // m132_117 = W*in
   wire signed [9:0] m132_117;
   assign m132_117 ={ {4{in132[5]}} , in132[5:0] };

   // m133_1 = W*in
   wire signed [9:0] m133_1;
   assign m133_1 =10'b0;

   // m133_2 = W*in
   wire signed [9:0] m133_2;
   assign m133_2 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_3 = W*in
   wire signed [9:0] m133_3;
   assign m133_3 =10'b0;

   // m133_4 = W*in
   wire signed [9:0] m133_4;
   assign m133_4 =10'b0;

   // m133_5 = W*in
   wire signed [9:0] m133_5;
   assign m133_5 =10'b0;

   // m133_6 = W*in
   wire signed [9:0] m133_6;
   assign m133_6 =10'b0;

   // m133_7 = W*in
   wire signed [9:0] m133_7;
   assign m133_7 =10'b0;

   // m133_8 = W*in
   wire signed [9:0] m133_8;
   assign m133_8 =10'b0;

   // m133_9 = W*in
   wire signed [9:0] m133_9;
   assign m133_9 =10'b0;

   // m133_10 = W*in
   wire signed [9:0] m133_10;
   assign m133_10 =10'b0;

   // m133_11 = W*in
   wire signed [9:0] m133_11;
   assign m133_11 =10'b0;

   // m133_12 = W*in
   wire signed [9:0] m133_12;
   assign m133_12 =10'b0;

   // m133_13 = W*in
   wire signed [9:0] m133_13;
   assign m133_13 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_14 = W*in
   wire signed [9:0] m133_14;
   assign m133_14 ={ {4{in133[5]}} , in133[5:0] };

   // m133_15 = W*in
   wire signed [9:0] m133_15;
   assign m133_15 =10'b0;

   // m133_16 = W*in
   wire signed [9:0] m133_16;
   assign m133_16 ={ {4{in133[5]}} , in133[5:0] };

   // m133_17 = W*in
   wire signed [9:0] m133_17;
   assign m133_17 ={ {5{neg133[5]}} , neg133[5:1] };

   // m133_18 = W*in
   wire signed [9:0] m133_18;
   assign m133_18 ={ {4{in133[5]}} , in133[5:0] };

   // m133_19 = W*in
   wire signed [9:0] m133_19;
   assign m133_19 =10'b0;

   // m133_20 = W*in
   wire signed [9:0] m133_20;
   assign m133_20 =10'b0;

   // m133_21 = W*in
   wire signed [9:0] m133_21;
   assign m133_21 =10'b0;

   // m133_22 = W*in
   wire signed [9:0] m133_22;
   assign m133_22 ={ {5{neg133[5]}} , neg133[5:1] };

   // m133_23 = W*in
   wire signed [9:0] m133_23;
   assign m133_23 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_24 = W*in
   wire signed [9:0] m133_24;
   assign m133_24 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_25 = W*in
   wire signed [9:0] m133_25;
   assign m133_25 =10'b0;

   // m133_26 = W*in
   wire signed [9:0] m133_26;
   assign m133_26 ={ {4{in133[5]}} , in133[5:0] };

   // m133_27 = W*in
   wire signed [9:0] m133_27;
   assign m133_27 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_28 = W*in
   wire signed [9:0] m133_28;
   assign m133_28 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_29 = W*in
   wire signed [9:0] m133_29;
   assign m133_29 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_30 = W*in
   wire signed [9:0] m133_30;
   assign m133_30 ={ {5{in133[5]}} , in133[5:1] };

   // m133_31 = W*in
   wire signed [9:0] m133_31;
   assign m133_31 =10'b0;

   // m133_32 = W*in
   wire signed [9:0] m133_32;
   assign m133_32 =10'b0;

   // m133_33 = W*in
   wire signed [9:0] m133_33;
   assign m133_33 =10'b0;

   // m133_34 = W*in
   wire signed [9:0] m133_34;
   assign m133_34 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_35 = W*in
   wire signed [9:0] m133_35;
   assign m133_35 =10'b0;

   // m133_36 = W*in
   wire signed [9:0] m133_36;
   assign m133_36 =10'b0;

   // m133_37 = W*in
   wire signed [9:0] m133_37;
   assign m133_37 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_38 = W*in
   wire signed [9:0] m133_38;
   assign m133_38 ={ {4{in133[5]}} , in133[5:0] };

   // m133_39 = W*in
   wire signed [9:0] m133_39;
   assign m133_39 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_40 = W*in
   wire signed [9:0] m133_40;
   assign m133_40 =10'b0;

   // m133_41 = W*in
   wire signed [9:0] m133_41;
   assign m133_41 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_42 = W*in
   wire signed [9:0] m133_42;
   assign m133_42 ={ {3{in133[5]}} , in133 , {1{1'b0}} };

   // m133_43 = W*in
   wire signed [9:0] m133_43;
   assign m133_43 =10'b0;

   // m133_44 = W*in
   wire signed [9:0] m133_44;
   assign m133_44 =10'b0;

   // m133_45 = W*in
   wire signed [9:0] m133_45;
   assign m133_45 =10'b0;

   // m133_46 = W*in
   wire signed [9:0] m133_46;
   assign m133_46 =10'b0;

   // m133_47 = W*in
   wire signed [9:0] m133_47;
   assign m133_47 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_48 = W*in
   wire signed [9:0] m133_48;
   assign m133_48 =10'b0;

   // m133_49 = W*in
   wire signed [9:0] m133_49;
   assign m133_49 =10'b0;

   // m133_50 = W*in
   wire signed [9:0] m133_50;
   assign m133_50 =10'b0;

   // m133_51 = W*in
   wire signed [9:0] m133_51;
   assign m133_51 =10'b0;

   // m133_52 = W*in
   wire signed [9:0] m133_52;
   assign m133_52 =10'b0;

   // m133_53 = W*in
   wire signed [9:0] m133_53;
   assign m133_53 =10'b0;

   // m133_54 = W*in
   wire signed [9:0] m133_54;
   assign m133_54 =10'b0;

   // m133_55 = W*in
   wire signed [9:0] m133_55;
   assign m133_55 =10'b0;

   // m133_56 = W*in
   wire signed [9:0] m133_56;
   assign m133_56 =10'b0;

   // m133_57 = W*in
   wire signed [9:0] m133_57;
   assign m133_57 =10'b0;

   // m133_58 = W*in
   wire signed [9:0] m133_58;
   assign m133_58 =10'b0;

   // m133_59 = W*in
   wire signed [9:0] m133_59;
   assign m133_59 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_60 = W*in
   wire signed [9:0] m133_60;
   assign m133_60 =10'b0;

   // m133_61 = W*in
   wire signed [9:0] m133_61;
   assign m133_61 ={ {4{in133[5]}} , in133[5:0] };

   // m133_62 = W*in
   wire signed [9:0] m133_62;
   assign m133_62 =10'b0;

   // m133_63 = W*in
   wire signed [9:0] m133_63;
   assign m133_63 =10'b0;

   // m133_64 = W*in
   wire signed [9:0] m133_64;
   assign m133_64 ={ {5{in133[5]}} , in133[5:1] };

   // m133_65 = W*in
   wire signed [9:0] m133_65;
   assign m133_65 ={ {5{in133[5]}} , in133[5:1] };

   // m133_66 = W*in
   wire signed [9:0] m133_66;
   assign m133_66 =10'b0;

   // m133_67 = W*in
   wire signed [9:0] m133_67;
   assign m133_67 ={ {4{in133[5]}} , in133[5:0] };

   // m133_68 = W*in
   wire signed [9:0] m133_68;
   assign m133_68 =10'b0;

   // m133_69 = W*in
   wire signed [9:0] m133_69;
   assign m133_69 =10'b0;

   // m133_70 = W*in
   wire signed [9:0] m133_70;
   assign m133_70 =10'b0;

   // m133_71 = W*in
   wire signed [9:0] m133_71;
   assign m133_71 =10'b0;

   // m133_72 = W*in
   wire signed [9:0] m133_72;
   assign m133_72 ={ {4{in133[5]}} , in133[5:0] };

   // m133_73 = W*in
   wire signed [9:0] m133_73;
   assign m133_73 =10'b0;

   // m133_74 = W*in
   wire signed [9:0] m133_74;
   assign m133_74 ={ {4{in133[5]}} , in133[5:0] };

   // m133_75 = W*in
   wire signed [9:0] m133_75;
   assign m133_75 =10'b0;

   // m133_76 = W*in
   wire signed [9:0] m133_76;
   assign m133_76 =10'b0;

   // m133_77 = W*in
   wire signed [9:0] m133_77;
   assign m133_77 =10'b0;

   // m133_78 = W*in
   wire signed [9:0] m133_78;
   assign m133_78 =10'b0;

   // m133_79 = W*in
   wire signed [9:0] m133_79;
   assign m133_79 =10'b0;

   // m133_80 = W*in
   wire signed [9:0] m133_80;
   assign m133_80 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_81 = W*in
   wire signed [9:0] m133_81;
   assign m133_81 ={ {5{in133[5]}} , in133[5:1] };

   // m133_82 = W*in
   wire signed [9:0] m133_82;
   assign m133_82 =10'b0;

   // m133_83 = W*in
   wire signed [9:0] m133_83;
   assign m133_83 =10'b0;

   // m133_84 = W*in
   wire signed [9:0] m133_84;
   assign m133_84 =10'b0;

   // m133_85 = W*in
   wire signed [9:0] m133_85;
   assign m133_85 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_86 = W*in
   wire signed [9:0] m133_86;
   assign m133_86 =10'b0;

   // m133_87 = W*in
   wire signed [9:0] m133_87;
   assign m133_87 =10'b0;

   // m133_88 = W*in
   wire signed [9:0] m133_88;
   assign m133_88 =10'b0;

   // m133_89 = W*in
   wire signed [9:0] m133_89;
   assign m133_89 ={ {3{neg133[5]}} , neg133 , {1{1'b0}} };

   // m133_90 = W*in
   wire signed [9:0] m133_90;
   assign m133_90 =10'b0;

   // m133_91 = W*in
   wire signed [9:0] m133_91;
   assign m133_91 ={ {4{in133[5]}} , in133[5:0] };

   // m133_92 = W*in
   wire signed [9:0] m133_92;
   assign m133_92 =10'b0;

   // m133_93 = W*in
   wire signed [9:0] m133_93;
   assign m133_93 =10'b0;

   // m133_94 = W*in
   wire signed [9:0] m133_94;
   assign m133_94 ={ {4{in133[5]}} , in133[5:0] };

   // m133_95 = W*in
   wire signed [9:0] m133_95;
   assign m133_95 =10'b0;

   // m133_96 = W*in
   wire signed [9:0] m133_96;
   assign m133_96 =10'b0;

   // m133_97 = W*in
   wire signed [9:0] m133_97;
   assign m133_97 ={ {4{in133[5]}} , in133[5:0] };

   // m133_98 = W*in
   wire signed [9:0] m133_98;
   assign m133_98 =10'b0;

   // m133_99 = W*in
   wire signed [9:0] m133_99;
   assign m133_99 =10'b0;

   // m133_100 = W*in
   wire signed [9:0] m133_100;
   assign m133_100 ={ {4{in133[5]}} , in133[5:0] };

   // m133_101 = W*in
   wire signed [9:0] m133_101;
   assign m133_101 =10'b0;

   // m133_102 = W*in
   wire signed [9:0] m133_102;
   assign m133_102 =10'b0;

   // m133_103 = W*in
   wire signed [9:0] m133_103;
   assign m133_103 =10'b0;

   // m133_104 = W*in
   wire signed [9:0] m133_104;
   assign m133_104 =10'b0;

   // m133_105 = W*in
   wire signed [9:0] m133_105;
   assign m133_105 =10'b0;

   // m133_106 = W*in
   wire signed [9:0] m133_106;
   assign m133_106 =10'b0;

   // m133_107 = W*in
   wire signed [9:0] m133_107;
   assign m133_107 =10'b0;

   // m133_108 = W*in
   wire signed [9:0] m133_108;
   assign m133_108 ={ {4{neg133[5]}} , neg133[5:0] };

   // m133_109 = W*in
   wire signed [9:0] m133_109;
   assign m133_109 ={ {3{neg133[5]}} , neg133 , {1{1'b0}} };

   // m133_110 = W*in
   wire signed [9:0] m133_110;
   assign m133_110 ={ {4{in133[5]}} , in133[5:0] };

   // m133_111 = W*in
   wire signed [9:0] m133_111;
   assign m133_111 =10'b0;

   // m133_112 = W*in
   wire signed [9:0] m133_112;
   assign m133_112 ={ {4{in133[5]}} , in133[5:0] };

   // m133_113 = W*in
   wire signed [9:0] m133_113;
   assign m133_113 =10'b0;

   // m133_114 = W*in
   wire signed [9:0] m133_114;
   assign m133_114 ={ {5{neg133[5]}} , neg133[5:1] };

   // m133_115 = W*in
   wire signed [9:0] m133_115;
   assign m133_115 =10'b0;

   // m133_116 = W*in
   wire signed [9:0] m133_116;
   assign m133_116 =10'b0;

   // m133_117 = W*in
   wire signed [9:0] m133_117;
   assign m133_117 =10'b0;

   // m134_1 = W*in
   wire signed [9:0] m134_1;
   assign m134_1 =10'b0;

   // m134_2 = W*in
   wire signed [9:0] m134_2;
   assign m134_2 =10'b0;

   // m134_3 = W*in
   wire signed [9:0] m134_3;
   assign m134_3 =10'b0;

   // m134_4 = W*in
   wire signed [9:0] m134_4;
   assign m134_4 =10'b0;

   // m134_5 = W*in
   wire signed [9:0] m134_5;
   assign m134_5 =10'b0;

   // m134_6 = W*in
   wire signed [9:0] m134_6;
   assign m134_6 =10'b0;

   // m134_7 = W*in
   wire signed [9:0] m134_7;
   assign m134_7 =10'b0;

   // m134_8 = W*in
   wire signed [9:0] m134_8;
   assign m134_8 =10'b0;

   // m134_9 = W*in
   wire signed [9:0] m134_9;
   assign m134_9 =10'b0;

   // m134_10 = W*in
   wire signed [9:0] m134_10;
   assign m134_10 =10'b0;

   // m134_11 = W*in
   wire signed [9:0] m134_11;
   assign m134_11 =10'b0;

   // m134_12 = W*in
   wire signed [9:0] m134_12;
   assign m134_12 =10'b0;

   // m134_13 = W*in
   wire signed [9:0] m134_13;
   assign m134_13 =10'b0;

   // m134_14 = W*in
   wire signed [9:0] m134_14;
   assign m134_14 =10'b0;

   // m134_15 = W*in
   wire signed [9:0] m134_15;
   assign m134_15 =10'b0;

   // m134_16 = W*in
   wire signed [9:0] m134_16;
   assign m134_16 =10'b0;

   // m134_17 = W*in
   wire signed [9:0] m134_17;
   assign m134_17 ={ {5{in134[5]}} , in134[5:1] };

   // m134_18 = W*in
   wire signed [9:0] m134_18;
   assign m134_18 ={ {5{in134[5]}} , in134[5:1] };

   // m134_19 = W*in
   wire signed [9:0] m134_19;
   assign m134_19 =10'b0;

   // m134_20 = W*in
   wire signed [9:0] m134_20;
   assign m134_20 =10'b0;

   // m134_21 = W*in
   wire signed [9:0] m134_21;
   assign m134_21 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_22 = W*in
   wire signed [9:0] m134_22;
   assign m134_22 =10'b0;

   // m134_23 = W*in
   wire signed [9:0] m134_23;
   assign m134_23 =10'b0;

   // m134_24 = W*in
   wire signed [9:0] m134_24;
   assign m134_24 =10'b0;

   // m134_25 = W*in
   wire signed [9:0] m134_25;
   assign m134_25 =10'b0;

   // m134_26 = W*in
   wire signed [9:0] m134_26;
   assign m134_26 ={ {5{in134[5]}} , in134[5:1] };

   // m134_27 = W*in
   wire signed [9:0] m134_27;
   assign m134_27 =10'b0;

   // m134_28 = W*in
   wire signed [9:0] m134_28;
   assign m134_28 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_29 = W*in
   wire signed [9:0] m134_29;
   assign m134_29 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_30 = W*in
   wire signed [9:0] m134_30;
   assign m134_30 =10'b0;

   // m134_31 = W*in
   wire signed [9:0] m134_31;
   assign m134_31 =10'b0;

   // m134_32 = W*in
   wire signed [9:0] m134_32;
   assign m134_32 =10'b0;

   // m134_33 = W*in
   wire signed [9:0] m134_33;
   assign m134_33 =10'b0;

   // m134_34 = W*in
   wire signed [9:0] m134_34;
   assign m134_34 =10'b0;

   // m134_35 = W*in
   wire signed [9:0] m134_35;
   assign m134_35 =10'b0;

   // m134_36 = W*in
   wire signed [9:0] m134_36;
   assign m134_36 =10'b0;

   // m134_37 = W*in
   wire signed [9:0] m134_37;
   assign m134_37 =10'b0;

   // m134_38 = W*in
   wire signed [9:0] m134_38;
   assign m134_38 ={ {4{in134[5]}} , in134[5:0] };

   // m134_39 = W*in
   wire signed [9:0] m134_39;
   assign m134_39 =10'b0;

   // m134_40 = W*in
   wire signed [9:0] m134_40;
   assign m134_40 =10'b0;

   // m134_41 = W*in
   wire signed [9:0] m134_41;
   assign m134_41 =10'b0;

   // m134_42 = W*in
   wire signed [9:0] m134_42;
   assign m134_42 =10'b0;

   // m134_43 = W*in
   wire signed [9:0] m134_43;
   assign m134_43 =10'b0;

   // m134_44 = W*in
   wire signed [9:0] m134_44;
   assign m134_44 =10'b0;

   // m134_45 = W*in
   wire signed [9:0] m134_45;
   assign m134_45 =10'b0;

   // m134_46 = W*in
   wire signed [9:0] m134_46;
   assign m134_46 =10'b0;

   // m134_47 = W*in
   wire signed [9:0] m134_47;
   assign m134_47 =10'b0;

   // m134_48 = W*in
   wire signed [9:0] m134_48;
   assign m134_48 =10'b0;

   // m134_49 = W*in
   wire signed [9:0] m134_49;
   assign m134_49 =10'b0;

   // m134_50 = W*in
   wire signed [9:0] m134_50;
   assign m134_50 ={ {4{neg134[5]}} , neg134[5:0] };

   // m134_51 = W*in
   wire signed [9:0] m134_51;
   assign m134_51 =10'b0;

   // m134_52 = W*in
   wire signed [9:0] m134_52;
   assign m134_52 =10'b0;

   // m134_53 = W*in
   wire signed [9:0] m134_53;
   assign m134_53 =10'b0;

   // m134_54 = W*in
   wire signed [9:0] m134_54;
   assign m134_54 =10'b0;

   // m134_55 = W*in
   wire signed [9:0] m134_55;
   assign m134_55 =10'b0;

   // m134_56 = W*in
   wire signed [9:0] m134_56;
   assign m134_56 =10'b0;

   // m134_57 = W*in
   wire signed [9:0] m134_57;
   assign m134_57 =10'b0;

   // m134_58 = W*in
   wire signed [9:0] m134_58;
   assign m134_58 =10'b0;

   // m134_59 = W*in
   wire signed [9:0] m134_59;
   assign m134_59 =10'b0;

   // m134_60 = W*in
   wire signed [9:0] m134_60;
   assign m134_60 =10'b0;

   // m134_61 = W*in
   wire signed [9:0] m134_61;
   assign m134_61 =10'b0;

   // m134_62 = W*in
   wire signed [9:0] m134_62;
   assign m134_62 =10'b0;

   // m134_63 = W*in
   wire signed [9:0] m134_63;
   assign m134_63 =10'b0;

   // m134_64 = W*in
   wire signed [9:0] m134_64;
   assign m134_64 ={ {4{in134[5]}} , in134[5:0] };

   // m134_65 = W*in
   wire signed [9:0] m134_65;
   assign m134_65 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_66 = W*in
   wire signed [9:0] m134_66;
   assign m134_66 =10'b0;

   // m134_67 = W*in
   wire signed [9:0] m134_67;
   assign m134_67 =10'b0;

   // m134_68 = W*in
   wire signed [9:0] m134_68;
   assign m134_68 =10'b0;

   // m134_69 = W*in
   wire signed [9:0] m134_69;
   assign m134_69 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_70 = W*in
   wire signed [9:0] m134_70;
   assign m134_70 =10'b0;

   // m134_71 = W*in
   wire signed [9:0] m134_71;
   assign m134_71 ={ {4{in134[5]}} , in134[5:0] };

   // m134_72 = W*in
   wire signed [9:0] m134_72;
   assign m134_72 ={ {5{in134[5]}} , in134[5:1] };

   // m134_73 = W*in
   wire signed [9:0] m134_73;
   assign m134_73 =10'b0;

   // m134_74 = W*in
   wire signed [9:0] m134_74;
   assign m134_74 =10'b0;

   // m134_75 = W*in
   wire signed [9:0] m134_75;
   assign m134_75 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_76 = W*in
   wire signed [9:0] m134_76;
   assign m134_76 =10'b0;

   // m134_77 = W*in
   wire signed [9:0] m134_77;
   assign m134_77 =10'b0;

   // m134_78 = W*in
   wire signed [9:0] m134_78;
   assign m134_78 =10'b0;

   // m134_79 = W*in
   wire signed [9:0] m134_79;
   assign m134_79 =10'b0;

   // m134_80 = W*in
   wire signed [9:0] m134_80;
   assign m134_80 =10'b0;

   // m134_81 = W*in
   wire signed [9:0] m134_81;
   assign m134_81 ={ {5{in134[5]}} , in134[5:1] };

   // m134_82 = W*in
   wire signed [9:0] m134_82;
   assign m134_82 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_83 = W*in
   wire signed [9:0] m134_83;
   assign m134_83 =10'b0;

   // m134_84 = W*in
   wire signed [9:0] m134_84;
   assign m134_84 =10'b0;

   // m134_85 = W*in
   wire signed [9:0] m134_85;
   assign m134_85 ={ {4{neg134[5]}} , neg134[5:0] };

   // m134_86 = W*in
   wire signed [9:0] m134_86;
   assign m134_86 =10'b0;

   // m134_87 = W*in
   wire signed [9:0] m134_87;
   assign m134_87 =10'b0;

   // m134_88 = W*in
   wire signed [9:0] m134_88;
   assign m134_88 =10'b0;

   // m134_89 = W*in
   wire signed [9:0] m134_89;
   assign m134_89 =10'b0;

   // m134_90 = W*in
   wire signed [9:0] m134_90;
   assign m134_90 =10'b0;

   // m134_91 = W*in
   wire signed [9:0] m134_91;
   assign m134_91 =10'b0;

   // m134_92 = W*in
   wire signed [9:0] m134_92;
   assign m134_92 =10'b0;

   // m134_93 = W*in
   wire signed [9:0] m134_93;
   assign m134_93 =10'b0;

   // m134_94 = W*in
   wire signed [9:0] m134_94;
   assign m134_94 =10'b0;

   // m134_95 = W*in
   wire signed [9:0] m134_95;
   assign m134_95 =10'b0;

   // m134_96 = W*in
   wire signed [9:0] m134_96;
   assign m134_96 =10'b0;

   // m134_97 = W*in
   wire signed [9:0] m134_97;
   assign m134_97 =10'b0;

   // m134_98 = W*in
   wire signed [9:0] m134_98;
   assign m134_98 =10'b0;

   // m134_99 = W*in
   wire signed [9:0] m134_99;
   assign m134_99 =10'b0;

   // m134_100 = W*in
   wire signed [9:0] m134_100;
   assign m134_100 =10'b0;

   // m134_101 = W*in
   wire signed [9:0] m134_101;
   assign m134_101 =10'b0;

   // m134_102 = W*in
   wire signed [9:0] m134_102;
   assign m134_102 =10'b0;

   // m134_103 = W*in
   wire signed [9:0] m134_103;
   assign m134_103 =10'b0;

   // m134_104 = W*in
   wire signed [9:0] m134_104;
   assign m134_104 =10'b0;

   // m134_105 = W*in
   wire signed [9:0] m134_105;
   assign m134_105 =10'b0;

   // m134_106 = W*in
   wire signed [9:0] m134_106;
   assign m134_106 =10'b0;

   // m134_107 = W*in
   wire signed [9:0] m134_107;
   assign m134_107 =10'b0;

   // m134_108 = W*in
   wire signed [9:0] m134_108;
   assign m134_108 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_109 = W*in
   wire signed [9:0] m134_109;
   assign m134_109 ={ {5{neg134[5]}} , neg134[5:1] };

   // m134_110 = W*in
   wire signed [9:0] m134_110;
   assign m134_110 ={ {4{in134[5]}} , in134[5:0] };

   // m134_111 = W*in
   wire signed [9:0] m134_111;
   assign m134_111 =10'b0;

   // m134_112 = W*in
   wire signed [9:0] m134_112;
   assign m134_112 =10'b0;

   // m134_113 = W*in
   wire signed [9:0] m134_113;
   assign m134_113 =10'b0;

   // m134_114 = W*in
   wire signed [9:0] m134_114;
   assign m134_114 =10'b0;

   // m134_115 = W*in
   wire signed [9:0] m134_115;
   assign m134_115 =10'b0;

   // m134_116 = W*in
   wire signed [9:0] m134_116;
   assign m134_116 =10'b0;

   // m134_117 = W*in
   wire signed [9:0] m134_117;
   assign m134_117 =10'b0;

   // m135_1 = W*in
   wire signed [9:0] m135_1;
   assign m135_1 =10'b0;

   // m135_2 = W*in
   wire signed [9:0] m135_2;
   assign m135_2 =10'b0;

   // m135_3 = W*in
   wire signed [9:0] m135_3;
   assign m135_3 ={ {4{in135[5]}} , in135[5:0] };

   // m135_4 = W*in
   wire signed [9:0] m135_4;
   assign m135_4 =10'b0;

   // m135_5 = W*in
   wire signed [9:0] m135_5;
   assign m135_5 =10'b0;

   // m135_6 = W*in
   wire signed [9:0] m135_6;
   assign m135_6 ={ {4{neg135[5]}} , neg135[5:0] };

   // m135_7 = W*in
   wire signed [9:0] m135_7;
   assign m135_7 =10'b0;

   // m135_8 = W*in
   wire signed [9:0] m135_8;
   assign m135_8 =10'b0;

   // m135_9 = W*in
   wire signed [9:0] m135_9;
   assign m135_9 =10'b0;

   // m135_10 = W*in
   wire signed [9:0] m135_10;
   assign m135_10 =10'b0;

   // m135_11 = W*in
   wire signed [9:0] m135_11;
   assign m135_11 =10'b0;

   // m135_12 = W*in
   wire signed [9:0] m135_12;
   assign m135_12 ={ {4{in135[5]}} , in135[5:0] };

   // m135_13 = W*in
   wire signed [9:0] m135_13;
   assign m135_13 =10'b0;

   // m135_14 = W*in
   wire signed [9:0] m135_14;
   assign m135_14 =10'b0;

   // m135_15 = W*in
   wire signed [9:0] m135_15;
   assign m135_15 =10'b0;

   // m135_16 = W*in
   wire signed [9:0] m135_16;
   assign m135_16 =10'b0;

   // m135_17 = W*in
   wire signed [9:0] m135_17;
   assign m135_17 ={ {5{in135[5]}} , in135[5:1] };

   // m135_18 = W*in
   wire signed [9:0] m135_18;
   assign m135_18 ={ {5{in135[5]}} , in135[5:1] };

   // m135_19 = W*in
   wire signed [9:0] m135_19;
   assign m135_19 =10'b0;

   // m135_20 = W*in
   wire signed [9:0] m135_20;
   assign m135_20 =10'b0;

   // m135_21 = W*in
   wire signed [9:0] m135_21;
   assign m135_21 ={ {5{neg135[5]}} , neg135[5:1] };

   // m135_22 = W*in
   wire signed [9:0] m135_22;
   assign m135_22 =10'b0;

   // m135_23 = W*in
   wire signed [9:0] m135_23;
   assign m135_23 ={ {5{in135[5]}} , in135[5:1] };

   // m135_24 = W*in
   wire signed [9:0] m135_24;
   assign m135_24 =10'b0;

   // m135_25 = W*in
   wire signed [9:0] m135_25;
   assign m135_25 =10'b0;

   // m135_26 = W*in
   wire signed [9:0] m135_26;
   assign m135_26 =10'b0;

   // m135_27 = W*in
   wire signed [9:0] m135_27;
   assign m135_27 ={ {5{in135[5]}} , in135[5:1] };

   // m135_28 = W*in
   wire signed [9:0] m135_28;
   assign m135_28 =10'b0;

   // m135_29 = W*in
   wire signed [9:0] m135_29;
   assign m135_29 =10'b0;

   // m135_30 = W*in
   wire signed [9:0] m135_30;
   assign m135_30 =10'b0;

   // m135_31 = W*in
   wire signed [9:0] m135_31;
   assign m135_31 =10'b0;

   // m135_32 = W*in
   wire signed [9:0] m135_32;
   assign m135_32 =10'b0;

   // m135_33 = W*in
   wire signed [9:0] m135_33;
   assign m135_33 =10'b0;

   // m135_34 = W*in
   wire signed [9:0] m135_34;
   assign m135_34 =10'b0;

   // m135_35 = W*in
   wire signed [9:0] m135_35;
   assign m135_35 =10'b0;

   // m135_36 = W*in
   wire signed [9:0] m135_36;
   assign m135_36 ={ {5{in135[5]}} , in135[5:1] };

   // m135_37 = W*in
   wire signed [9:0] m135_37;
   assign m135_37 =10'b0;

   // m135_38 = W*in
   wire signed [9:0] m135_38;
   assign m135_38 =10'b0;

   // m135_39 = W*in
   wire signed [9:0] m135_39;
   assign m135_39 =10'b0;

   // m135_40 = W*in
   wire signed [9:0] m135_40;
   assign m135_40 =10'b0;

   // m135_41 = W*in
   wire signed [9:0] m135_41;
   assign m135_41 =10'b0;

   // m135_42 = W*in
   wire signed [9:0] m135_42;
   assign m135_42 =10'b0;

   // m135_43 = W*in
   wire signed [9:0] m135_43;
   assign m135_43 =10'b0;

   // m135_44 = W*in
   wire signed [9:0] m135_44;
   assign m135_44 =10'b0;

   // m135_45 = W*in
   wire signed [9:0] m135_45;
   assign m135_45 =10'b0;

   // m135_46 = W*in
   wire signed [9:0] m135_46;
   assign m135_46 ={ {4{in135[5]}} , in135[5:0] };

   // m135_47 = W*in
   wire signed [9:0] m135_47;
   assign m135_47 =10'b0;

   // m135_48 = W*in
   wire signed [9:0] m135_48;
   assign m135_48 =10'b0;

   // m135_49 = W*in
   wire signed [9:0] m135_49;
   assign m135_49 =10'b0;

   // m135_50 = W*in
   wire signed [9:0] m135_50;
   assign m135_50 =10'b0;

   // m135_51 = W*in
   wire signed [9:0] m135_51;
   assign m135_51 =10'b0;

   // m135_52 = W*in
   wire signed [9:0] m135_52;
   assign m135_52 =10'b0;

   // m135_53 = W*in
   wire signed [9:0] m135_53;
   assign m135_53 =10'b0;

   // m135_54 = W*in
   wire signed [9:0] m135_54;
   assign m135_54 =10'b0;

   // m135_55 = W*in
   wire signed [9:0] m135_55;
   assign m135_55 =10'b0;

   // m135_56 = W*in
   wire signed [9:0] m135_56;
   assign m135_56 =10'b0;

   // m135_57 = W*in
   wire signed [9:0] m135_57;
   assign m135_57 =10'b0;

   // m135_58 = W*in
   wire signed [9:0] m135_58;
   assign m135_58 =10'b0;

   // m135_59 = W*in
   wire signed [9:0] m135_59;
   assign m135_59 =10'b0;

   // m135_60 = W*in
   wire signed [9:0] m135_60;
   assign m135_60 =10'b0;

   // m135_61 = W*in
   wire signed [9:0] m135_61;
   assign m135_61 =10'b0;

   // m135_62 = W*in
   wire signed [9:0] m135_62;
   assign m135_62 =10'b0;

   // m135_63 = W*in
   wire signed [9:0] m135_63;
   assign m135_63 ={ {4{neg135[5]}} , neg135[5:0] };

   // m135_64 = W*in
   wire signed [9:0] m135_64;
   assign m135_64 ={ {4{in135[5]}} , in135[5:0] };

   // m135_65 = W*in
   wire signed [9:0] m135_65;
   assign m135_65 =10'b0;

   // m135_66 = W*in
   wire signed [9:0] m135_66;
   assign m135_66 ={ {5{in135[5]}} , in135[5:1] };

   // m135_67 = W*in
   wire signed [9:0] m135_67;
   assign m135_67 ={ {4{neg135[5]}} , neg135[5:0] };

   // m135_68 = W*in
   wire signed [9:0] m135_68;
   assign m135_68 =10'b0;

   // m135_69 = W*in
   wire signed [9:0] m135_69;
   assign m135_69 ={ {4{neg135[5]}} , neg135[5:0] };

   // m135_70 = W*in
   wire signed [9:0] m135_70;
   assign m135_70 =10'b0;

   // m135_71 = W*in
   wire signed [9:0] m135_71;
   assign m135_71 =10'b0;

   // m135_72 = W*in
   wire signed [9:0] m135_72;
   assign m135_72 ={ {5{neg135[5]}} , neg135[5:1] };

   // m135_73 = W*in
   wire signed [9:0] m135_73;
   assign m135_73 ={ {5{in135[5]}} , in135[5:1] };

   // m135_74 = W*in
   wire signed [9:0] m135_74;
   assign m135_74 ={ {5{neg135[5]}} , neg135[5:1] };

   // m135_75 = W*in
   wire signed [9:0] m135_75;
   assign m135_75 =10'b0;

   // m135_76 = W*in
   wire signed [9:0] m135_76;
   assign m135_76 =10'b0;

   // m135_77 = W*in
   wire signed [9:0] m135_77;
   assign m135_77 =10'b0;

   // m135_78 = W*in
   wire signed [9:0] m135_78;
   assign m135_78 =10'b0;

   // m135_79 = W*in
   wire signed [9:0] m135_79;
   assign m135_79 =10'b0;

   // m135_80 = W*in
   wire signed [9:0] m135_80;
   assign m135_80 =10'b0;

   // m135_81 = W*in
   wire signed [9:0] m135_81;
   assign m135_81 ={ {5{in135[5]}} , in135[5:1] };

   // m135_82 = W*in
   wire signed [9:0] m135_82;
   assign m135_82 ={ {5{neg135[5]}} , neg135[5:1] };

   // m135_83 = W*in
   wire signed [9:0] m135_83;
   assign m135_83 =10'b0;

   // m135_84 = W*in
   wire signed [9:0] m135_84;
   assign m135_84 =10'b0;

   // m135_85 = W*in
   wire signed [9:0] m135_85;
   assign m135_85 =10'b0;

   // m135_86 = W*in
   wire signed [9:0] m135_86;
   assign m135_86 =10'b0;

   // m135_87 = W*in
   wire signed [9:0] m135_87;
   assign m135_87 =10'b0;

   // m135_88 = W*in
   wire signed [9:0] m135_88;
   assign m135_88 =10'b0;

   // m135_89 = W*in
   wire signed [9:0] m135_89;
   assign m135_89 =10'b0;

   // m135_90 = W*in
   wire signed [9:0] m135_90;
   assign m135_90 =10'b0;

   // m135_91 = W*in
   wire signed [9:0] m135_91;
   assign m135_91 =10'b0;

   // m135_92 = W*in
   wire signed [9:0] m135_92;
   assign m135_92 =10'b0;

   // m135_93 = W*in
   wire signed [9:0] m135_93;
   assign m135_93 ={ {4{neg135[5]}} , neg135[5:0] };

   // m135_94 = W*in
   wire signed [9:0] m135_94;
   assign m135_94 =10'b0;

   // m135_95 = W*in
   wire signed [9:0] m135_95;
   assign m135_95 =10'b0;

   // m135_96 = W*in
   wire signed [9:0] m135_96;
   assign m135_96 =10'b0;

   // m135_97 = W*in
   wire signed [9:0] m135_97;
   assign m135_97 =10'b0;

   // m135_98 = W*in
   wire signed [9:0] m135_98;
   assign m135_98 =10'b0;

   // m135_99 = W*in
   wire signed [9:0] m135_99;
   assign m135_99 =10'b0;

   // m135_100 = W*in
   wire signed [9:0] m135_100;
   assign m135_100 =10'b0;

   // m135_101 = W*in
   wire signed [9:0] m135_101;
   assign m135_101 =10'b0;

   // m135_102 = W*in
   wire signed [9:0] m135_102;
   assign m135_102 =10'b0;

   // m135_103 = W*in
   wire signed [9:0] m135_103;
   assign m135_103 ={ {4{in135[5]}} , in135[5:0] };

   // m135_104 = W*in
   wire signed [9:0] m135_104;
   assign m135_104 =10'b0;

   // m135_105 = W*in
   wire signed [9:0] m135_105;
   assign m135_105 =10'b0;

   // m135_106 = W*in
   wire signed [9:0] m135_106;
   assign m135_106 =10'b0;

   // m135_107 = W*in
   wire signed [9:0] m135_107;
   assign m135_107 ={ {5{in135[5]}} , in135[5:1] };

   // m135_108 = W*in
   wire signed [9:0] m135_108;
   assign m135_108 =10'b0;

   // m135_109 = W*in
   wire signed [9:0] m135_109;
   assign m135_109 ={ {5{in135[5]}} , in135[5:1] };

   // m135_110 = W*in
   wire signed [9:0] m135_110;
   assign m135_110 =10'b0;

   // m135_111 = W*in
   wire signed [9:0] m135_111;
   assign m135_111 =10'b0;

   // m135_112 = W*in
   wire signed [9:0] m135_112;
   assign m135_112 =10'b0;

   // m135_113 = W*in
   wire signed [9:0] m135_113;
   assign m135_113 =10'b0;

   // m135_114 = W*in
   wire signed [9:0] m135_114;
   assign m135_114 =10'b0;

   // m135_115 = W*in
   wire signed [9:0] m135_115;
   assign m135_115 =10'b0;

   // m135_116 = W*in
   wire signed [9:0] m135_116;
   assign m135_116 =10'b0;

   // m135_117 = W*in
   wire signed [9:0] m135_117;
   assign m135_117 =10'b0;

   // m136_1 = W*in
   wire signed [9:0] m136_1;
   assign m136_1 =10'b0;

   // m136_2 = W*in
   wire signed [9:0] m136_2;
   assign m136_2 =10'b0;

   // m136_3 = W*in
   wire signed [9:0] m136_3;
   assign m136_3 ={ {4{in136[5]}} , in136[5:0] };

   // m136_4 = W*in
   wire signed [9:0] m136_4;
   assign m136_4 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_5 = W*in
   wire signed [9:0] m136_5;
   assign m136_5 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_6 = W*in
   wire signed [9:0] m136_6;
   assign m136_6 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_7 = W*in
   wire signed [9:0] m136_7;
   assign m136_7 =10'b0;

   // m136_8 = W*in
   wire signed [9:0] m136_8;
   assign m136_8 =10'b0;

   // m136_9 = W*in
   wire signed [9:0] m136_9;
   assign m136_9 =10'b0;

   // m136_10 = W*in
   wire signed [9:0] m136_10;
   assign m136_10 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_11 = W*in
   wire signed [9:0] m136_11;
   assign m136_11 =10'b0;

   // m136_12 = W*in
   wire signed [9:0] m136_12;
   assign m136_12 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_13 = W*in
   wire signed [9:0] m136_13;
   assign m136_13 =10'b0;

   // m136_14 = W*in
   wire signed [9:0] m136_14;
   assign m136_14 =10'b0;

   // m136_15 = W*in
   wire signed [9:0] m136_15;
   assign m136_15 =10'b0;

   // m136_16 = W*in
   wire signed [9:0] m136_16;
   assign m136_16 =10'b0;

   // m136_17 = W*in
   wire signed [9:0] m136_17;
   assign m136_17 =10'b0;

   // m136_18 = W*in
   wire signed [9:0] m136_18;
   assign m136_18 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_19 = W*in
   wire signed [9:0] m136_19;
   assign m136_19 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_20 = W*in
   wire signed [9:0] m136_20;
   assign m136_20 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_21 = W*in
   wire signed [9:0] m136_21;
   assign m136_21 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_22 = W*in
   wire signed [9:0] m136_22;
   assign m136_22 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_23 = W*in
   wire signed [9:0] m136_23;
   assign m136_23 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_24 = W*in
   wire signed [9:0] m136_24;
   assign m136_24 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_25 = W*in
   wire signed [9:0] m136_25;
   assign m136_25 =10'b0;

   // m136_26 = W*in
   wire signed [9:0] m136_26;
   assign m136_26 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_27 = W*in
   wire signed [9:0] m136_27;
   assign m136_27 ={ {4{in136[5]}} , in136[5:0] };

   // m136_28 = W*in
   wire signed [9:0] m136_28;
   assign m136_28 ={ {5{in136[5]}} , in136[5:1] };

   // m136_29 = W*in
   wire signed [9:0] m136_29;
   assign m136_29 =10'b0;

   // m136_30 = W*in
   wire signed [9:0] m136_30;
   assign m136_30 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_31 = W*in
   wire signed [9:0] m136_31;
   assign m136_31 =10'b0;

   // m136_32 = W*in
   wire signed [9:0] m136_32;
   assign m136_32 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_33 = W*in
   wire signed [9:0] m136_33;
   assign m136_33 =10'b0;

   // m136_34 = W*in
   wire signed [9:0] m136_34;
   assign m136_34 =10'b0;

   // m136_35 = W*in
   wire signed [9:0] m136_35;
   assign m136_35 =10'b0;

   // m136_36 = W*in
   wire signed [9:0] m136_36;
   assign m136_36 ={ {5{in136[5]}} , in136[5:1] };

   // m136_37 = W*in
   wire signed [9:0] m136_37;
   assign m136_37 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_38 = W*in
   wire signed [9:0] m136_38;
   assign m136_38 =10'b0;

   // m136_39 = W*in
   wire signed [9:0] m136_39;
   assign m136_39 =10'b0;

   // m136_40 = W*in
   wire signed [9:0] m136_40;
   assign m136_40 =10'b0;

   // m136_41 = W*in
   wire signed [9:0] m136_41;
   assign m136_41 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_42 = W*in
   wire signed [9:0] m136_42;
   assign m136_42 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_43 = W*in
   wire signed [9:0] m136_43;
   assign m136_43 ={ {4{in136[5]}} , in136[5:0] };

   // m136_44 = W*in
   wire signed [9:0] m136_44;
   assign m136_44 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_45 = W*in
   wire signed [9:0] m136_45;
   assign m136_45 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_46 = W*in
   wire signed [9:0] m136_46;
   assign m136_46 ={ {4{in136[5]}} , in136[5:0] };

   // m136_47 = W*in
   wire signed [9:0] m136_47;
   assign m136_47 =10'b0;

   // m136_48 = W*in
   wire signed [9:0] m136_48;
   assign m136_48 =10'b0;

   // m136_49 = W*in
   wire signed [9:0] m136_49;
   assign m136_49 =10'b0;

   // m136_50 = W*in
   wire signed [9:0] m136_50;
   assign m136_50 =10'b0;

   // m136_51 = W*in
   wire signed [9:0] m136_51;
   assign m136_51 =10'b0;

   // m136_52 = W*in
   wire signed [9:0] m136_52;
   assign m136_52 =10'b0;

   // m136_53 = W*in
   wire signed [9:0] m136_53;
   assign m136_53 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_54 = W*in
   wire signed [9:0] m136_54;
   assign m136_54 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_55 = W*in
   wire signed [9:0] m136_55;
   assign m136_55 =10'b0;

   // m136_56 = W*in
   wire signed [9:0] m136_56;
   assign m136_56 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_57 = W*in
   wire signed [9:0] m136_57;
   assign m136_57 =10'b0;

   // m136_58 = W*in
   wire signed [9:0] m136_58;
   assign m136_58 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_59 = W*in
   wire signed [9:0] m136_59;
   assign m136_59 =10'b0;

   // m136_60 = W*in
   wire signed [9:0] m136_60;
   assign m136_60 =10'b0;

   // m136_61 = W*in
   wire signed [9:0] m136_61;
   assign m136_61 =10'b0;

   // m136_62 = W*in
   wire signed [9:0] m136_62;
   assign m136_62 =10'b0;

   // m136_63 = W*in
   wire signed [9:0] m136_63;
   assign m136_63 ={ {3{neg136[5]}} , neg136 , {1{1'b0}} };

   // m136_64 = W*in
   wire signed [9:0] m136_64;
   assign m136_64 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_65 = W*in
   wire signed [9:0] m136_65;
   assign m136_65 =10'b0;

   // m136_66 = W*in
   wire signed [9:0] m136_66;
   assign m136_66 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_67 = W*in
   wire signed [9:0] m136_67;
   assign m136_67 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_68 = W*in
   wire signed [9:0] m136_68;
   assign m136_68 =10'b0;

   // m136_69 = W*in
   wire signed [9:0] m136_69;
   assign m136_69 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_70 = W*in
   wire signed [9:0] m136_70;
   assign m136_70 =10'b0;

   // m136_71 = W*in
   wire signed [9:0] m136_71;
   assign m136_71 ={ {4{in136[5]}} , in136[5:0] };

   // m136_72 = W*in
   wire signed [9:0] m136_72;
   assign m136_72 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_73 = W*in
   wire signed [9:0] m136_73;
   assign m136_73 ={ {5{in136[5]}} , in136[5:1] };

   // m136_74 = W*in
   wire signed [9:0] m136_74;
   assign m136_74 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_75 = W*in
   wire signed [9:0] m136_75;
   assign m136_75 =10'b0;

   // m136_76 = W*in
   wire signed [9:0] m136_76;
   assign m136_76 =10'b0;

   // m136_77 = W*in
   wire signed [9:0] m136_77;
   assign m136_77 ={ {4{in136[5]}} , in136[5:0] };

   // m136_78 = W*in
   wire signed [9:0] m136_78;
   assign m136_78 =10'b0;

   // m136_79 = W*in
   wire signed [9:0] m136_79;
   assign m136_79 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_80 = W*in
   wire signed [9:0] m136_80;
   assign m136_80 =10'b0;

   // m136_81 = W*in
   wire signed [9:0] m136_81;
   assign m136_81 ={ {4{in136[5]}} , in136[5:0] };

   // m136_82 = W*in
   wire signed [9:0] m136_82;
   assign m136_82 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_83 = W*in
   wire signed [9:0] m136_83;
   assign m136_83 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_84 = W*in
   wire signed [9:0] m136_84;
   assign m136_84 =10'b0;

   // m136_85 = W*in
   wire signed [9:0] m136_85;
   assign m136_85 ={ {3{neg136[5]}} , neg136 , {1{1'b0}} };

   // m136_86 = W*in
   wire signed [9:0] m136_86;
   assign m136_86 ={ {4{in136[5]}} , in136[5:0] };

   // m136_87 = W*in
   wire signed [9:0] m136_87;
   assign m136_87 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_88 = W*in
   wire signed [9:0] m136_88;
   assign m136_88 =10'b0;

   // m136_89 = W*in
   wire signed [9:0] m136_89;
   assign m136_89 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_90 = W*in
   wire signed [9:0] m136_90;
   assign m136_90 =10'b0;

   // m136_91 = W*in
   wire signed [9:0] m136_91;
   assign m136_91 ={ {4{in136[5]}} , in136[5:0] };

   // m136_92 = W*in
   wire signed [9:0] m136_92;
   assign m136_92 =10'b0;

   // m136_93 = W*in
   wire signed [9:0] m136_93;
   assign m136_93 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_94 = W*in
   wire signed [9:0] m136_94;
   assign m136_94 ={ {4{in136[5]}} , in136[5:0] };

   // m136_95 = W*in
   wire signed [9:0] m136_95;
   assign m136_95 =10'b0;

   // m136_96 = W*in
   wire signed [9:0] m136_96;
   assign m136_96 =10'b0;

   // m136_97 = W*in
   wire signed [9:0] m136_97;
   assign m136_97 ={ {4{in136[5]}} , in136[5:0] };

   // m136_98 = W*in
   wire signed [9:0] m136_98;
   assign m136_98 =10'b0;

   // m136_99 = W*in
   wire signed [9:0] m136_99;
   assign m136_99 =10'b0;

   // m136_100 = W*in
   wire signed [9:0] m136_100;
   assign m136_100 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_101 = W*in
   wire signed [9:0] m136_101;
   assign m136_101 ={ {4{in136[5]}} , in136[5:0] };

   // m136_102 = W*in
   wire signed [9:0] m136_102;
   assign m136_102 =10'b0;

   // m136_103 = W*in
   wire signed [9:0] m136_103;
   assign m136_103 ={ {4{in136[5]}} , in136[5:0] };

   // m136_104 = W*in
   wire signed [9:0] m136_104;
   assign m136_104 ={ {4{in136[5]}} , in136[5:0] };

   // m136_105 = W*in
   wire signed [9:0] m136_105;
   assign m136_105 =10'b0;

   // m136_106 = W*in
   wire signed [9:0] m136_106;
   assign m136_106 =10'b0;

   // m136_107 = W*in
   wire signed [9:0] m136_107;
   assign m136_107 ={ {4{in136[5]}} , in136[5:0] };

   // m136_108 = W*in
   wire signed [9:0] m136_108;
   assign m136_108 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_109 = W*in
   wire signed [9:0] m136_109;
   assign m136_109 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_110 = W*in
   wire signed [9:0] m136_110;
   assign m136_110 ={ {4{in136[5]}} , in136[5:0] };

   // m136_111 = W*in
   wire signed [9:0] m136_111;
   assign m136_111 =10'b0;

   // m136_112 = W*in
   wire signed [9:0] m136_112;
   assign m136_112 ={ {3{in136[5]}} , in136 , {1{1'b0}} };

   // m136_113 = W*in
   wire signed [9:0] m136_113;
   assign m136_113 =10'b0;

   // m136_114 = W*in
   wire signed [9:0] m136_114;
   assign m136_114 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_115 = W*in
   wire signed [9:0] m136_115;
   assign m136_115 ={ {5{neg136[5]}} , neg136[5:1] };

   // m136_116 = W*in
   wire signed [9:0] m136_116;
   assign m136_116 ={ {4{neg136[5]}} , neg136[5:0] };

   // m136_117 = W*in
   wire signed [9:0] m136_117;
   assign m136_117 ={ {4{in136[5]}} , in136[5:0] };

   // m137_1 = W*in
   wire signed [9:0] m137_1;
   assign m137_1 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_2 = W*in
   wire signed [9:0] m137_2;
   assign m137_2 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_3 = W*in
   wire signed [9:0] m137_3;
   assign m137_3 =10'b0;

   // m137_4 = W*in
   wire signed [9:0] m137_4;
   assign m137_4 =10'b0;

   // m137_5 = W*in
   wire signed [9:0] m137_5;
   assign m137_5 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_6 = W*in
   wire signed [9:0] m137_6;
   assign m137_6 =10'b0;

   // m137_7 = W*in
   wire signed [9:0] m137_7;
   assign m137_7 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_8 = W*in
   wire signed [9:0] m137_8;
   assign m137_8 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_9 = W*in
   wire signed [9:0] m137_9;
   assign m137_9 =10'b0;

   // m137_10 = W*in
   wire signed [9:0] m137_10;
   assign m137_10 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_11 = W*in
   wire signed [9:0] m137_11;
   assign m137_11 =10'b0;

   // m137_12 = W*in
   wire signed [9:0] m137_12;
   assign m137_12 ={ {4{in137[5]}} , in137[5:0] };

   // m137_13 = W*in
   wire signed [9:0] m137_13;
   assign m137_13 =10'b0;

   // m137_14 = W*in
   wire signed [9:0] m137_14;
   assign m137_14 =10'b0;

   // m137_15 = W*in
   wire signed [9:0] m137_15;
   assign m137_15 =10'b0;

   // m137_16 = W*in
   wire signed [9:0] m137_16;
   assign m137_16 =10'b0;

   // m137_17 = W*in
   wire signed [9:0] m137_17;
   assign m137_17 =10'b0;

   // m137_18 = W*in
   wire signed [9:0] m137_18;
   assign m137_18 ={ {4{in137[5]}} , in137[5:0] };

   // m137_19 = W*in
   wire signed [9:0] m137_19;
   assign m137_19 =10'b0;

   // m137_20 = W*in
   wire signed [9:0] m137_20;
   assign m137_20 =10'b0;

   // m137_21 = W*in
   wire signed [9:0] m137_21;
   assign m137_21 =10'b0;

   // m137_22 = W*in
   wire signed [9:0] m137_22;
   assign m137_22 ={ {5{neg137[5]}} , neg137[5:1] };

   // m137_23 = W*in
   wire signed [9:0] m137_23;
   assign m137_23 =10'b0;

   // m137_24 = W*in
   wire signed [9:0] m137_24;
   assign m137_24 =10'b0;

   // m137_25 = W*in
   wire signed [9:0] m137_25;
   assign m137_25 =10'b0;

   // m137_26 = W*in
   wire signed [9:0] m137_26;
   assign m137_26 =10'b0;

   // m137_27 = W*in
   wire signed [9:0] m137_27;
   assign m137_27 =10'b0;

   // m137_28 = W*in
   wire signed [9:0] m137_28;
   assign m137_28 ={ {5{in137[5]}} , in137[5:1] };

   // m137_29 = W*in
   wire signed [9:0] m137_29;
   assign m137_29 =10'b0;

   // m137_30 = W*in
   wire signed [9:0] m137_30;
   assign m137_30 =10'b0;

   // m137_31 = W*in
   wire signed [9:0] m137_31;
   assign m137_31 ={ {5{neg137[5]}} , neg137[5:1] };

   // m137_32 = W*in
   wire signed [9:0] m137_32;
   assign m137_32 ={ {3{neg137[5]}} , neg137 , {1{1'b0}} };

   // m137_33 = W*in
   wire signed [9:0] m137_33;
   assign m137_33 =10'b0;

   // m137_34 = W*in
   wire signed [9:0] m137_34;
   assign m137_34 =10'b0;

   // m137_35 = W*in
   wire signed [9:0] m137_35;
   assign m137_35 =10'b0;

   // m137_36 = W*in
   wire signed [9:0] m137_36;
   assign m137_36 =10'b0;

   // m137_37 = W*in
   wire signed [9:0] m137_37;
   assign m137_37 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_38 = W*in
   wire signed [9:0] m137_38;
   assign m137_38 ={ {4{in137[5]}} , in137[5:0] };

   // m137_39 = W*in
   wire signed [9:0] m137_39;
   assign m137_39 =10'b0;

   // m137_40 = W*in
   wire signed [9:0] m137_40;
   assign m137_40 =10'b0;

   // m137_41 = W*in
   wire signed [9:0] m137_41;
   assign m137_41 =10'b0;

   // m137_42 = W*in
   wire signed [9:0] m137_42;
   assign m137_42 =10'b0;

   // m137_43 = W*in
   wire signed [9:0] m137_43;
   assign m137_43 ={ {4{in137[5]}} , in137[5:0] };

   // m137_44 = W*in
   wire signed [9:0] m137_44;
   assign m137_44 =10'b0;

   // m137_45 = W*in
   wire signed [9:0] m137_45;
   assign m137_45 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_46 = W*in
   wire signed [9:0] m137_46;
   assign m137_46 =10'b0;

   // m137_47 = W*in
   wire signed [9:0] m137_47;
   assign m137_47 =10'b0;

   // m137_48 = W*in
   wire signed [9:0] m137_48;
   assign m137_48 =10'b0;

   // m137_49 = W*in
   wire signed [9:0] m137_49;
   assign m137_49 =10'b0;

   // m137_50 = W*in
   wire signed [9:0] m137_50;
   assign m137_50 =10'b0;

   // m137_51 = W*in
   wire signed [9:0] m137_51;
   assign m137_51 ={ {3{neg137[5]}} , neg137 , {1{1'b0}} };

   // m137_52 = W*in
   wire signed [9:0] m137_52;
   assign m137_52 =10'b0;

   // m137_53 = W*in
   wire signed [9:0] m137_53;
   assign m137_53 =10'b0;

   // m137_54 = W*in
   wire signed [9:0] m137_54;
   assign m137_54 =10'b0;

   // m137_55 = W*in
   wire signed [9:0] m137_55;
   assign m137_55 =10'b0;

   // m137_56 = W*in
   wire signed [9:0] m137_56;
   assign m137_56 =10'b0;

   // m137_57 = W*in
   wire signed [9:0] m137_57;
   assign m137_57 =10'b0;

   // m137_58 = W*in
   wire signed [9:0] m137_58;
   assign m137_58 =10'b0;

   // m137_59 = W*in
   wire signed [9:0] m137_59;
   assign m137_59 =10'b0;

   // m137_60 = W*in
   wire signed [9:0] m137_60;
   assign m137_60 ={ {4{in137[5]}} , in137[5:0] };

   // m137_61 = W*in
   wire signed [9:0] m137_61;
   assign m137_61 =10'b0;

   // m137_62 = W*in
   wire signed [9:0] m137_62;
   assign m137_62 =10'b0;

   // m137_63 = W*in
   wire signed [9:0] m137_63;
   assign m137_63 =10'b0;

   // m137_64 = W*in
   wire signed [9:0] m137_64;
   assign m137_64 =10'b0;

   // m137_65 = W*in
   wire signed [9:0] m137_65;
   assign m137_65 =10'b0;

   // m137_66 = W*in
   wire signed [9:0] m137_66;
   assign m137_66 ={ {4{in137[5]}} , in137[5:0] };

   // m137_67 = W*in
   wire signed [9:0] m137_67;
   assign m137_67 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_68 = W*in
   wire signed [9:0] m137_68;
   assign m137_68 =10'b0;

   // m137_69 = W*in
   wire signed [9:0] m137_69;
   assign m137_69 =10'b0;

   // m137_70 = W*in
   wire signed [9:0] m137_70;
   assign m137_70 =10'b0;

   // m137_71 = W*in
   wire signed [9:0] m137_71;
   assign m137_71 ={ {4{in137[5]}} , in137[5:0] };

   // m137_72 = W*in
   wire signed [9:0] m137_72;
   assign m137_72 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_73 = W*in
   wire signed [9:0] m137_73;
   assign m137_73 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_74 = W*in
   wire signed [9:0] m137_74;
   assign m137_74 =10'b0;

   // m137_75 = W*in
   wire signed [9:0] m137_75;
   assign m137_75 =10'b0;

   // m137_76 = W*in
   wire signed [9:0] m137_76;
   assign m137_76 =10'b0;

   // m137_77 = W*in
   wire signed [9:0] m137_77;
   assign m137_77 =10'b0;

   // m137_78 = W*in
   wire signed [9:0] m137_78;
   assign m137_78 =10'b0;

   // m137_79 = W*in
   wire signed [9:0] m137_79;
   assign m137_79 =10'b0;

   // m137_80 = W*in
   wire signed [9:0] m137_80;
   assign m137_80 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_81 = W*in
   wire signed [9:0] m137_81;
   assign m137_81 =10'b0;

   // m137_82 = W*in
   wire signed [9:0] m137_82;
   assign m137_82 =10'b0;

   // m137_83 = W*in
   wire signed [9:0] m137_83;
   assign m137_83 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_84 = W*in
   wire signed [9:0] m137_84;
   assign m137_84 =10'b0;

   // m137_85 = W*in
   wire signed [9:0] m137_85;
   assign m137_85 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_86 = W*in
   wire signed [9:0] m137_86;
   assign m137_86 =10'b0;

   // m137_87 = W*in
   wire signed [9:0] m137_87;
   assign m137_87 =10'b0;

   // m137_88 = W*in
   wire signed [9:0] m137_88;
   assign m137_88 =10'b0;

   // m137_89 = W*in
   wire signed [9:0] m137_89;
   assign m137_89 ={ {4{neg137[5]}} , neg137[5:0] };

   // m137_90 = W*in
   wire signed [9:0] m137_90;
   assign m137_90 =10'b0;

   // m137_91 = W*in
   wire signed [9:0] m137_91;
   assign m137_91 ={ {4{in137[5]}} , in137[5:0] };

   // m137_92 = W*in
   wire signed [9:0] m137_92;
   assign m137_92 =10'b0;

   // m137_93 = W*in
   wire signed [9:0] m137_93;
   assign m137_93 =10'b0;

   // m137_94 = W*in
   wire signed [9:0] m137_94;
   assign m137_94 =10'b0;

   // m137_95 = W*in
   wire signed [9:0] m137_95;
   assign m137_95 =10'b0;

   // m137_96 = W*in
   wire signed [9:0] m137_96;
   assign m137_96 =10'b0;

   // m137_97 = W*in
   wire signed [9:0] m137_97;
   assign m137_97 ={ {4{in137[5]}} , in137[5:0] };

   // m137_98 = W*in
   wire signed [9:0] m137_98;
   assign m137_98 =10'b0;

   // m137_99 = W*in
   wire signed [9:0] m137_99;
   assign m137_99 =10'b0;

   // m137_100 = W*in
   wire signed [9:0] m137_100;
   assign m137_100 =10'b0;

   // m137_101 = W*in
   wire signed [9:0] m137_101;
   assign m137_101 =10'b0;

   // m137_102 = W*in
   wire signed [9:0] m137_102;
   assign m137_102 =10'b0;

   // m137_103 = W*in
   wire signed [9:0] m137_103;
   assign m137_103 =10'b0;

   // m137_104 = W*in
   wire signed [9:0] m137_104;
   assign m137_104 ={ {4{in137[5]}} , in137[5:0] };

   // m137_105 = W*in
   wire signed [9:0] m137_105;
   assign m137_105 =10'b0;

   // m137_106 = W*in
   wire signed [9:0] m137_106;
   assign m137_106 =10'b0;

   // m137_107 = W*in
   wire signed [9:0] m137_107;
   assign m137_107 =10'b0;

   // m137_108 = W*in
   wire signed [9:0] m137_108;
   assign m137_108 =10'b0;

   // m137_109 = W*in
   wire signed [9:0] m137_109;
   assign m137_109 =10'b0;

   // m137_110 = W*in
   wire signed [9:0] m137_110;
   assign m137_110 ={ {4{in137[5]}} , in137[5:0] };

   // m137_111 = W*in
   wire signed [9:0] m137_111;
   assign m137_111 =10'b0;

   // m137_112 = W*in
   wire signed [9:0] m137_112;
   assign m137_112 ={ {4{in137[5]}} , in137[5:0] };

   // m137_113 = W*in
   wire signed [9:0] m137_113;
   assign m137_113 =10'b0;

   // m137_114 = W*in
   wire signed [9:0] m137_114;
   assign m137_114 =10'b0;

   // m137_115 = W*in
   wire signed [9:0] m137_115;
   assign m137_115 =10'b0;

   // m137_116 = W*in
   wire signed [9:0] m137_116;
   assign m137_116 =10'b0;

   // m137_117 = W*in
   wire signed [9:0] m137_117;
   assign m137_117 =10'b0;

   // m138_1 = W*in
   wire signed [9:0] m138_1;
   assign m138_1 =10'b0;

   // m138_2 = W*in
   wire signed [9:0] m138_2;
   assign m138_2 =10'b0;

   // m138_3 = W*in
   wire signed [9:0] m138_3;
   assign m138_3 =10'b0;

   // m138_4 = W*in
   wire signed [9:0] m138_4;
   assign m138_4 =10'b0;

   // m138_5 = W*in
   wire signed [9:0] m138_5;
   assign m138_5 =10'b0;

   // m138_6 = W*in
   wire signed [9:0] m138_6;
   assign m138_6 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_7 = W*in
   wire signed [9:0] m138_7;
   assign m138_7 =10'b0;

   // m138_8 = W*in
   wire signed [9:0] m138_8;
   assign m138_8 =10'b0;

   // m138_9 = W*in
   wire signed [9:0] m138_9;
   assign m138_9 =10'b0;

   // m138_10 = W*in
   wire signed [9:0] m138_10;
   assign m138_10 =10'b0;

   // m138_11 = W*in
   wire signed [9:0] m138_11;
   assign m138_11 ={ {4{in138[5]}} , in138[5:0] };

   // m138_12 = W*in
   wire signed [9:0] m138_12;
   assign m138_12 =10'b0;

   // m138_13 = W*in
   wire signed [9:0] m138_13;
   assign m138_13 =10'b0;

   // m138_14 = W*in
   wire signed [9:0] m138_14;
   assign m138_14 =10'b0;

   // m138_15 = W*in
   wire signed [9:0] m138_15;
   assign m138_15 =10'b0;

   // m138_16 = W*in
   wire signed [9:0] m138_16;
   assign m138_16 =10'b0;

   // m138_17 = W*in
   wire signed [9:0] m138_17;
   assign m138_17 ={ {4{in138[5]}} , in138[5:0] };

   // m138_18 = W*in
   wire signed [9:0] m138_18;
   assign m138_18 =10'b0;

   // m138_19 = W*in
   wire signed [9:0] m138_19;
   assign m138_19 =10'b0;

   // m138_20 = W*in
   wire signed [9:0] m138_20;
   assign m138_20 =10'b0;

   // m138_21 = W*in
   wire signed [9:0] m138_21;
   assign m138_21 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_22 = W*in
   wire signed [9:0] m138_22;
   assign m138_22 ={ {5{in138[5]}} , in138[5:1] };

   // m138_23 = W*in
   wire signed [9:0] m138_23;
   assign m138_23 =10'b0;

   // m138_24 = W*in
   wire signed [9:0] m138_24;
   assign m138_24 =10'b0;

   // m138_25 = W*in
   wire signed [9:0] m138_25;
   assign m138_25 =10'b0;

   // m138_26 = W*in
   wire signed [9:0] m138_26;
   assign m138_26 =10'b0;

   // m138_27 = W*in
   wire signed [9:0] m138_27;
   assign m138_27 ={ {4{in138[5]}} , in138[5:0] };

   // m138_28 = W*in
   wire signed [9:0] m138_28;
   assign m138_28 =10'b0;

   // m138_29 = W*in
   wire signed [9:0] m138_29;
   assign m138_29 =10'b0;

   // m138_30 = W*in
   wire signed [9:0] m138_30;
   assign m138_30 =10'b0;

   // m138_31 = W*in
   wire signed [9:0] m138_31;
   assign m138_31 ={ {5{in138[5]}} , in138[5:1] };

   // m138_32 = W*in
   wire signed [9:0] m138_32;
   assign m138_32 =10'b0;

   // m138_33 = W*in
   wire signed [9:0] m138_33;
   assign m138_33 =10'b0;

   // m138_34 = W*in
   wire signed [9:0] m138_34;
   assign m138_34 =10'b0;

   // m138_35 = W*in
   wire signed [9:0] m138_35;
   assign m138_35 =10'b0;

   // m138_36 = W*in
   wire signed [9:0] m138_36;
   assign m138_36 ={ {5{in138[5]}} , in138[5:1] };

   // m138_37 = W*in
   wire signed [9:0] m138_37;
   assign m138_37 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_38 = W*in
   wire signed [9:0] m138_38;
   assign m138_38 =10'b0;

   // m138_39 = W*in
   wire signed [9:0] m138_39;
   assign m138_39 =10'b0;

   // m138_40 = W*in
   wire signed [9:0] m138_40;
   assign m138_40 =10'b0;

   // m138_41 = W*in
   wire signed [9:0] m138_41;
   assign m138_41 =10'b0;

   // m138_42 = W*in
   wire signed [9:0] m138_42;
   assign m138_42 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_43 = W*in
   wire signed [9:0] m138_43;
   assign m138_43 =10'b0;

   // m138_44 = W*in
   wire signed [9:0] m138_44;
   assign m138_44 =10'b0;

   // m138_45 = W*in
   wire signed [9:0] m138_45;
   assign m138_45 =10'b0;

   // m138_46 = W*in
   wire signed [9:0] m138_46;
   assign m138_46 ={ {4{in138[5]}} , in138[5:0] };

   // m138_47 = W*in
   wire signed [9:0] m138_47;
   assign m138_47 =10'b0;

   // m138_48 = W*in
   wire signed [9:0] m138_48;
   assign m138_48 =10'b0;

   // m138_49 = W*in
   wire signed [9:0] m138_49;
   assign m138_49 ={ {4{in138[5]}} , in138[5:0] };

   // m138_50 = W*in
   wire signed [9:0] m138_50;
   assign m138_50 =10'b0;

   // m138_51 = W*in
   wire signed [9:0] m138_51;
   assign m138_51 =10'b0;

   // m138_52 = W*in
   wire signed [9:0] m138_52;
   assign m138_52 =10'b0;

   // m138_53 = W*in
   wire signed [9:0] m138_53;
   assign m138_53 =10'b0;

   // m138_54 = W*in
   wire signed [9:0] m138_54;
   assign m138_54 =10'b0;

   // m138_55 = W*in
   wire signed [9:0] m138_55;
   assign m138_55 =10'b0;

   // m138_56 = W*in
   wire signed [9:0] m138_56;
   assign m138_56 =10'b0;

   // m138_57 = W*in
   wire signed [9:0] m138_57;
   assign m138_57 =10'b0;

   // m138_58 = W*in
   wire signed [9:0] m138_58;
   assign m138_58 =10'b0;

   // m138_59 = W*in
   wire signed [9:0] m138_59;
   assign m138_59 =10'b0;

   // m138_60 = W*in
   wire signed [9:0] m138_60;
   assign m138_60 =10'b0;

   // m138_61 = W*in
   wire signed [9:0] m138_61;
   assign m138_61 =10'b0;

   // m138_62 = W*in
   wire signed [9:0] m138_62;
   assign m138_62 =10'b0;

   // m138_63 = W*in
   wire signed [9:0] m138_63;
   assign m138_63 =10'b0;

   // m138_64 = W*in
   wire signed [9:0] m138_64;
   assign m138_64 =10'b0;

   // m138_65 = W*in
   wire signed [9:0] m138_65;
   assign m138_65 =10'b0;

   // m138_66 = W*in
   wire signed [9:0] m138_66;
   assign m138_66 =10'b0;

   // m138_67 = W*in
   wire signed [9:0] m138_67;
   assign m138_67 =10'b0;

   // m138_68 = W*in
   wire signed [9:0] m138_68;
   assign m138_68 =10'b0;

   // m138_69 = W*in
   wire signed [9:0] m138_69;
   assign m138_69 =10'b0;

   // m138_70 = W*in
   wire signed [9:0] m138_70;
   assign m138_70 ={ {5{neg138[5]}} , neg138[5:1] };

   // m138_71 = W*in
   wire signed [9:0] m138_71;
   assign m138_71 ={ {5{in138[5]}} , in138[5:1] };

   // m138_72 = W*in
   wire signed [9:0] m138_72;
   assign m138_72 ={ {5{in138[5]}} , in138[5:1] };

   // m138_73 = W*in
   wire signed [9:0] m138_73;
   assign m138_73 =10'b0;

   // m138_74 = W*in
   wire signed [9:0] m138_74;
   assign m138_74 =10'b0;

   // m138_75 = W*in
   wire signed [9:0] m138_75;
   assign m138_75 =10'b0;

   // m138_76 = W*in
   wire signed [9:0] m138_76;
   assign m138_76 =10'b0;

   // m138_77 = W*in
   wire signed [9:0] m138_77;
   assign m138_77 =10'b0;

   // m138_78 = W*in
   wire signed [9:0] m138_78;
   assign m138_78 =10'b0;

   // m138_79 = W*in
   wire signed [9:0] m138_79;
   assign m138_79 =10'b0;

   // m138_80 = W*in
   wire signed [9:0] m138_80;
   assign m138_80 =10'b0;

   // m138_81 = W*in
   wire signed [9:0] m138_81;
   assign m138_81 =10'b0;

   // m138_82 = W*in
   wire signed [9:0] m138_82;
   assign m138_82 =10'b0;

   // m138_83 = W*in
   wire signed [9:0] m138_83;
   assign m138_83 =10'b0;

   // m138_84 = W*in
   wire signed [9:0] m138_84;
   assign m138_84 =10'b0;

   // m138_85 = W*in
   wire signed [9:0] m138_85;
   assign m138_85 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_86 = W*in
   wire signed [9:0] m138_86;
   assign m138_86 =10'b0;

   // m138_87 = W*in
   wire signed [9:0] m138_87;
   assign m138_87 =10'b0;

   // m138_88 = W*in
   wire signed [9:0] m138_88;
   assign m138_88 =10'b0;

   // m138_89 = W*in
   wire signed [9:0] m138_89;
   assign m138_89 =10'b0;

   // m138_90 = W*in
   wire signed [9:0] m138_90;
   assign m138_90 =10'b0;

   // m138_91 = W*in
   wire signed [9:0] m138_91;
   assign m138_91 =10'b0;

   // m138_92 = W*in
   wire signed [9:0] m138_92;
   assign m138_92 =10'b0;

   // m138_93 = W*in
   wire signed [9:0] m138_93;
   assign m138_93 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_94 = W*in
   wire signed [9:0] m138_94;
   assign m138_94 =10'b0;

   // m138_95 = W*in
   wire signed [9:0] m138_95;
   assign m138_95 ={ {4{in138[5]}} , in138[5:0] };

   // m138_96 = W*in
   wire signed [9:0] m138_96;
   assign m138_96 =10'b0;

   // m138_97 = W*in
   wire signed [9:0] m138_97;
   assign m138_97 =10'b0;

   // m138_98 = W*in
   wire signed [9:0] m138_98;
   assign m138_98 =10'b0;

   // m138_99 = W*in
   wire signed [9:0] m138_99;
   assign m138_99 =10'b0;

   // m138_100 = W*in
   wire signed [9:0] m138_100;
   assign m138_100 =10'b0;

   // m138_101 = W*in
   wire signed [9:0] m138_101;
   assign m138_101 =10'b0;

   // m138_102 = W*in
   wire signed [9:0] m138_102;
   assign m138_102 =10'b0;

   // m138_103 = W*in
   wire signed [9:0] m138_103;
   assign m138_103 =10'b0;

   // m138_104 = W*in
   wire signed [9:0] m138_104;
   assign m138_104 ={ {4{in138[5]}} , in138[5:0] };

   // m138_105 = W*in
   wire signed [9:0] m138_105;
   assign m138_105 =10'b0;

   // m138_106 = W*in
   wire signed [9:0] m138_106;
   assign m138_106 =10'b0;

   // m138_107 = W*in
   wire signed [9:0] m138_107;
   assign m138_107 ={ {4{in138[5]}} , in138[5:0] };

   // m138_108 = W*in
   wire signed [9:0] m138_108;
   assign m138_108 =10'b0;

   // m138_109 = W*in
   wire signed [9:0] m138_109;
   assign m138_109 =10'b0;

   // m138_110 = W*in
   wire signed [9:0] m138_110;
   assign m138_110 =10'b0;

   // m138_111 = W*in
   wire signed [9:0] m138_111;
   assign m138_111 =10'b0;

   // m138_112 = W*in
   wire signed [9:0] m138_112;
   assign m138_112 =10'b0;

   // m138_113 = W*in
   wire signed [9:0] m138_113;
   assign m138_113 =10'b0;

   // m138_114 = W*in
   wire signed [9:0] m138_114;
   assign m138_114 ={ {5{in138[5]}} , in138[5:1] };

   // m138_115 = W*in
   wire signed [9:0] m138_115;
   assign m138_115 =10'b0;

   // m138_116 = W*in
   wire signed [9:0] m138_116;
   assign m138_116 ={ {4{neg138[5]}} , neg138[5:0] };

   // m138_117 = W*in
   wire signed [9:0] m138_117;
   assign m138_117 =10'b0;

   // m139_1 = W*in
   wire signed [9:0] m139_1;
   assign m139_1 =10'b0;

   // m139_2 = W*in
   wire signed [9:0] m139_2;
   assign m139_2 =10'b0;

   // m139_3 = W*in
   wire signed [9:0] m139_3;
   assign m139_3 =10'b0;

   // m139_4 = W*in
   wire signed [9:0] m139_4;
   assign m139_4 =10'b0;

   // m139_5 = W*in
   wire signed [9:0] m139_5;
   assign m139_5 =10'b0;

   // m139_6 = W*in
   wire signed [9:0] m139_6;
   assign m139_6 =10'b0;

   // m139_7 = W*in
   wire signed [9:0] m139_7;
   assign m139_7 =10'b0;

   // m139_8 = W*in
   wire signed [9:0] m139_8;
   assign m139_8 =10'b0;

   // m139_9 = W*in
   wire signed [9:0] m139_9;
   assign m139_9 =10'b0;

   // m139_10 = W*in
   wire signed [9:0] m139_10;
   assign m139_10 =10'b0;

   // m139_11 = W*in
   wire signed [9:0] m139_11;
   assign m139_11 =10'b0;

   // m139_12 = W*in
   wire signed [9:0] m139_12;
   assign m139_12 =10'b0;

   // m139_13 = W*in
   wire signed [9:0] m139_13;
   assign m139_13 =10'b0;

   // m139_14 = W*in
   wire signed [9:0] m139_14;
   assign m139_14 =10'b0;

   // m139_15 = W*in
   wire signed [9:0] m139_15;
   assign m139_15 =10'b0;

   // m139_16 = W*in
   wire signed [9:0] m139_16;
   assign m139_16 =10'b0;

   // m139_17 = W*in
   wire signed [9:0] m139_17;
   assign m139_17 =10'b0;

   // m139_18 = W*in
   wire signed [9:0] m139_18;
   assign m139_18 =10'b0;

   // m139_19 = W*in
   wire signed [9:0] m139_19;
   assign m139_19 =10'b0;

   // m139_20 = W*in
   wire signed [9:0] m139_20;
   assign m139_20 =10'b0;

   // m139_21 = W*in
   wire signed [9:0] m139_21;
   assign m139_21 =10'b0;

   // m139_22 = W*in
   wire signed [9:0] m139_22;
   assign m139_22 =10'b0;

   // m139_23 = W*in
   wire signed [9:0] m139_23;
   assign m139_23 ={ {5{in139[5]}} , in139[5:1] };

   // m139_24 = W*in
   wire signed [9:0] m139_24;
   assign m139_24 =10'b0;

   // m139_25 = W*in
   wire signed [9:0] m139_25;
   assign m139_25 =10'b0;

   // m139_26 = W*in
   wire signed [9:0] m139_26;
   assign m139_26 ={ {5{neg139[5]}} , neg139[5:1] };

   // m139_27 = W*in
   wire signed [9:0] m139_27;
   assign m139_27 ={ {4{in139[5]}} , in139[5:0] };

   // m139_28 = W*in
   wire signed [9:0] m139_28;
   assign m139_28 =10'b0;

   // m139_29 = W*in
   wire signed [9:0] m139_29;
   assign m139_29 =10'b0;

   // m139_30 = W*in
   wire signed [9:0] m139_30;
   assign m139_30 =10'b0;

   // m139_31 = W*in
   wire signed [9:0] m139_31;
   assign m139_31 =10'b0;

   // m139_32 = W*in
   wire signed [9:0] m139_32;
   assign m139_32 =10'b0;

   // m139_33 = W*in
   wire signed [9:0] m139_33;
   assign m139_33 =10'b0;

   // m139_34 = W*in
   wire signed [9:0] m139_34;
   assign m139_34 =10'b0;

   // m139_35 = W*in
   wire signed [9:0] m139_35;
   assign m139_35 ={ {5{in139[5]}} , in139[5:1] };

   // m139_36 = W*in
   wire signed [9:0] m139_36;
   assign m139_36 =10'b0;

   // m139_37 = W*in
   wire signed [9:0] m139_37;
   assign m139_37 =10'b0;

   // m139_38 = W*in
   wire signed [9:0] m139_38;
   assign m139_38 =10'b0;

   // m139_39 = W*in
   wire signed [9:0] m139_39;
   assign m139_39 =10'b0;

   // m139_40 = W*in
   wire signed [9:0] m139_40;
   assign m139_40 =10'b0;

   // m139_41 = W*in
   wire signed [9:0] m139_41;
   assign m139_41 =10'b0;

   // m139_42 = W*in
   wire signed [9:0] m139_42;
   assign m139_42 ={ {4{neg139[5]}} , neg139[5:0] };

   // m139_43 = W*in
   wire signed [9:0] m139_43;
   assign m139_43 =10'b0;

   // m139_44 = W*in
   wire signed [9:0] m139_44;
   assign m139_44 =10'b0;

   // m139_45 = W*in
   wire signed [9:0] m139_45;
   assign m139_45 =10'b0;

   // m139_46 = W*in
   wire signed [9:0] m139_46;
   assign m139_46 ={ {4{in139[5]}} , in139[5:0] };

   // m139_47 = W*in
   wire signed [9:0] m139_47;
   assign m139_47 =10'b0;

   // m139_48 = W*in
   wire signed [9:0] m139_48;
   assign m139_48 =10'b0;

   // m139_49 = W*in
   wire signed [9:0] m139_49;
   assign m139_49 =10'b0;

   // m139_50 = W*in
   wire signed [9:0] m139_50;
   assign m139_50 =10'b0;

   // m139_51 = W*in
   wire signed [9:0] m139_51;
   assign m139_51 =10'b0;

   // m139_52 = W*in
   wire signed [9:0] m139_52;
   assign m139_52 =10'b0;

   // m139_53 = W*in
   wire signed [9:0] m139_53;
   assign m139_53 =10'b0;

   // m139_54 = W*in
   wire signed [9:0] m139_54;
   assign m139_54 =10'b0;

   // m139_55 = W*in
   wire signed [9:0] m139_55;
   assign m139_55 =10'b0;

   // m139_56 = W*in
   wire signed [9:0] m139_56;
   assign m139_56 =10'b0;

   // m139_57 = W*in
   wire signed [9:0] m139_57;
   assign m139_57 =10'b0;

   // m139_58 = W*in
   wire signed [9:0] m139_58;
   assign m139_58 =10'b0;

   // m139_59 = W*in
   wire signed [9:0] m139_59;
   assign m139_59 =10'b0;

   // m139_60 = W*in
   wire signed [9:0] m139_60;
   assign m139_60 =10'b0;

   // m139_61 = W*in
   wire signed [9:0] m139_61;
   assign m139_61 =10'b0;

   // m139_62 = W*in
   wire signed [9:0] m139_62;
   assign m139_62 =10'b0;

   // m139_63 = W*in
   wire signed [9:0] m139_63;
   assign m139_63 =10'b0;

   // m139_64 = W*in
   wire signed [9:0] m139_64;
   assign m139_64 =10'b0;

   // m139_65 = W*in
   wire signed [9:0] m139_65;
   assign m139_65 ={ {5{neg139[5]}} , neg139[5:1] };

   // m139_66 = W*in
   wire signed [9:0] m139_66;
   assign m139_66 =10'b0;

   // m139_67 = W*in
   wire signed [9:0] m139_67;
   assign m139_67 =10'b0;

   // m139_68 = W*in
   wire signed [9:0] m139_68;
   assign m139_68 =10'b0;

   // m139_69 = W*in
   wire signed [9:0] m139_69;
   assign m139_69 =10'b0;

   // m139_70 = W*in
   wire signed [9:0] m139_70;
   assign m139_70 =10'b0;

   // m139_71 = W*in
   wire signed [9:0] m139_71;
   assign m139_71 =10'b0;

   // m139_72 = W*in
   wire signed [9:0] m139_72;
   assign m139_72 ={ {5{neg139[5]}} , neg139[5:1] };

   // m139_73 = W*in
   wire signed [9:0] m139_73;
   assign m139_73 =10'b0;

   // m139_74 = W*in
   wire signed [9:0] m139_74;
   assign m139_74 =10'b0;

   // m139_75 = W*in
   wire signed [9:0] m139_75;
   assign m139_75 =10'b0;

   // m139_76 = W*in
   wire signed [9:0] m139_76;
   assign m139_76 =10'b0;

   // m139_77 = W*in
   wire signed [9:0] m139_77;
   assign m139_77 =10'b0;

   // m139_78 = W*in
   wire signed [9:0] m139_78;
   assign m139_78 =10'b0;

   // m139_79 = W*in
   wire signed [9:0] m139_79;
   assign m139_79 =10'b0;

   // m139_80 = W*in
   wire signed [9:0] m139_80;
   assign m139_80 =10'b0;

   // m139_81 = W*in
   wire signed [9:0] m139_81;
   assign m139_81 =10'b0;

   // m139_82 = W*in
   wire signed [9:0] m139_82;
   assign m139_82 =10'b0;

   // m139_83 = W*in
   wire signed [9:0] m139_83;
   assign m139_83 =10'b0;

   // m139_84 = W*in
   wire signed [9:0] m139_84;
   assign m139_84 =10'b0;

   // m139_85 = W*in
   wire signed [9:0] m139_85;
   assign m139_85 =10'b0;

   // m139_86 = W*in
   wire signed [9:0] m139_86;
   assign m139_86 =10'b0;

   // m139_87 = W*in
   wire signed [9:0] m139_87;
   assign m139_87 =10'b0;

   // m139_88 = W*in
   wire signed [9:0] m139_88;
   assign m139_88 =10'b0;

   // m139_89 = W*in
   wire signed [9:0] m139_89;
   assign m139_89 =10'b0;

   // m139_90 = W*in
   wire signed [9:0] m139_90;
   assign m139_90 =10'b0;

   // m139_91 = W*in
   wire signed [9:0] m139_91;
   assign m139_91 =10'b0;

   // m139_92 = W*in
   wire signed [9:0] m139_92;
   assign m139_92 =10'b0;

   // m139_93 = W*in
   wire signed [9:0] m139_93;
   assign m139_93 =10'b0;

   // m139_94 = W*in
   wire signed [9:0] m139_94;
   assign m139_94 =10'b0;

   // m139_95 = W*in
   wire signed [9:0] m139_95;
   assign m139_95 =10'b0;

   // m139_96 = W*in
   wire signed [9:0] m139_96;
   assign m139_96 =10'b0;

   // m139_97 = W*in
   wire signed [9:0] m139_97;
   assign m139_97 =10'b0;

   // m139_98 = W*in
   wire signed [9:0] m139_98;
   assign m139_98 =10'b0;

   // m139_99 = W*in
   wire signed [9:0] m139_99;
   assign m139_99 =10'b0;

   // m139_100 = W*in
   wire signed [9:0] m139_100;
   assign m139_100 =10'b0;

   // m139_101 = W*in
   wire signed [9:0] m139_101;
   assign m139_101 =10'b0;

   // m139_102 = W*in
   wire signed [9:0] m139_102;
   assign m139_102 =10'b0;

   // m139_103 = W*in
   wire signed [9:0] m139_103;
   assign m139_103 =10'b0;

   // m139_104 = W*in
   wire signed [9:0] m139_104;
   assign m139_104 =10'b0;

   // m139_105 = W*in
   wire signed [9:0] m139_105;
   assign m139_105 =10'b0;

   // m139_106 = W*in
   wire signed [9:0] m139_106;
   assign m139_106 =10'b0;

   // m139_107 = W*in
   wire signed [9:0] m139_107;
   assign m139_107 ={ {5{in139[5]}} , in139[5:1] };

   // m139_108 = W*in
   wire signed [9:0] m139_108;
   assign m139_108 =10'b0;

   // m139_109 = W*in
   wire signed [9:0] m139_109;
   assign m139_109 ={ {5{in139[5]}} , in139[5:1] };

   // m139_110 = W*in
   wire signed [9:0] m139_110;
   assign m139_110 =10'b0;

   // m139_111 = W*in
   wire signed [9:0] m139_111;
   assign m139_111 =10'b0;

   // m139_112 = W*in
   wire signed [9:0] m139_112;
   assign m139_112 =10'b0;

   // m139_113 = W*in
   wire signed [9:0] m139_113;
   assign m139_113 =10'b0;

   // m139_114 = W*in
   wire signed [9:0] m139_114;
   assign m139_114 ={ {5{in139[5]}} , in139[5:1] };

   // m139_115 = W*in
   wire signed [9:0] m139_115;
   assign m139_115 =10'b0;

   // m139_116 = W*in
   wire signed [9:0] m139_116;
   assign m139_116 =10'b0;

   // m139_117 = W*in
   wire signed [9:0] m139_117;
   assign m139_117 =10'b0;

   // m140_1 = W*in
   wire signed [9:0] m140_1;
   assign m140_1 =10'b0;

   // m140_2 = W*in
   wire signed [9:0] m140_2;
   assign m140_2 =10'b0;

   // m140_3 = W*in
   wire signed [9:0] m140_3;
   assign m140_3 =10'b0;

   // m140_4 = W*in
   wire signed [9:0] m140_4;
   assign m140_4 =10'b0;

   // m140_5 = W*in
   wire signed [9:0] m140_5;
   assign m140_5 =10'b0;

   // m140_6 = W*in
   wire signed [9:0] m140_6;
   assign m140_6 =10'b0;

   // m140_7 = W*in
   wire signed [9:0] m140_7;
   assign m140_7 =10'b0;

   // m140_8 = W*in
   wire signed [9:0] m140_8;
   assign m140_8 =10'b0;

   // m140_9 = W*in
   wire signed [9:0] m140_9;
   assign m140_9 =10'b0;

   // m140_10 = W*in
   wire signed [9:0] m140_10;
   assign m140_10 =10'b0;

   // m140_11 = W*in
   wire signed [9:0] m140_11;
   assign m140_11 =10'b0;

   // m140_12 = W*in
   wire signed [9:0] m140_12;
   assign m140_12 =10'b0;

   // m140_13 = W*in
   wire signed [9:0] m140_13;
   assign m140_13 =10'b0;

   // m140_14 = W*in
   wire signed [9:0] m140_14;
   assign m140_14 ={ {4{in140[5]}} , in140[5:0] };

   // m140_15 = W*in
   wire signed [9:0] m140_15;
   assign m140_15 =10'b0;

   // m140_16 = W*in
   wire signed [9:0] m140_16;
   assign m140_16 =10'b0;

   // m140_17 = W*in
   wire signed [9:0] m140_17;
   assign m140_17 =10'b0;

   // m140_18 = W*in
   wire signed [9:0] m140_18;
   assign m140_18 ={ {5{in140[5]}} , in140[5:1] };

   // m140_19 = W*in
   wire signed [9:0] m140_19;
   assign m140_19 =10'b0;

   // m140_20 = W*in
   wire signed [9:0] m140_20;
   assign m140_20 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_21 = W*in
   wire signed [9:0] m140_21;
   assign m140_21 =10'b0;

   // m140_22 = W*in
   wire signed [9:0] m140_22;
   assign m140_22 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_23 = W*in
   wire signed [9:0] m140_23;
   assign m140_23 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_24 = W*in
   wire signed [9:0] m140_24;
   assign m140_24 =10'b0;

   // m140_25 = W*in
   wire signed [9:0] m140_25;
   assign m140_25 =10'b0;

   // m140_26 = W*in
   wire signed [9:0] m140_26;
   assign m140_26 =10'b0;

   // m140_27 = W*in
   wire signed [9:0] m140_27;
   assign m140_27 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_28 = W*in
   wire signed [9:0] m140_28;
   assign m140_28 ={ {4{neg140[5]}} , neg140[5:0] };

   // m140_29 = W*in
   wire signed [9:0] m140_29;
   assign m140_29 =10'b0;

   // m140_30 = W*in
   wire signed [9:0] m140_30;
   assign m140_30 =10'b0;

   // m140_31 = W*in
   wire signed [9:0] m140_31;
   assign m140_31 ={ {5{in140[5]}} , in140[5:1] };

   // m140_32 = W*in
   wire signed [9:0] m140_32;
   assign m140_32 =10'b0;

   // m140_33 = W*in
   wire signed [9:0] m140_33;
   assign m140_33 =10'b0;

   // m140_34 = W*in
   wire signed [9:0] m140_34;
   assign m140_34 =10'b0;

   // m140_35 = W*in
   wire signed [9:0] m140_35;
   assign m140_35 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_36 = W*in
   wire signed [9:0] m140_36;
   assign m140_36 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_37 = W*in
   wire signed [9:0] m140_37;
   assign m140_37 =10'b0;

   // m140_38 = W*in
   wire signed [9:0] m140_38;
   assign m140_38 =10'b0;

   // m140_39 = W*in
   wire signed [9:0] m140_39;
   assign m140_39 =10'b0;

   // m140_40 = W*in
   wire signed [9:0] m140_40;
   assign m140_40 =10'b0;

   // m140_41 = W*in
   wire signed [9:0] m140_41;
   assign m140_41 =10'b0;

   // m140_42 = W*in
   wire signed [9:0] m140_42;
   assign m140_42 =10'b0;

   // m140_43 = W*in
   wire signed [9:0] m140_43;
   assign m140_43 =10'b0;

   // m140_44 = W*in
   wire signed [9:0] m140_44;
   assign m140_44 =10'b0;

   // m140_45 = W*in
   wire signed [9:0] m140_45;
   assign m140_45 =10'b0;

   // m140_46 = W*in
   wire signed [9:0] m140_46;
   assign m140_46 =10'b0;

   // m140_47 = W*in
   wire signed [9:0] m140_47;
   assign m140_47 =10'b0;

   // m140_48 = W*in
   wire signed [9:0] m140_48;
   assign m140_48 =10'b0;

   // m140_49 = W*in
   wire signed [9:0] m140_49;
   assign m140_49 ={ {4{neg140[5]}} , neg140[5:0] };

   // m140_50 = W*in
   wire signed [9:0] m140_50;
   assign m140_50 =10'b0;

   // m140_51 = W*in
   wire signed [9:0] m140_51;
   assign m140_51 =10'b0;

   // m140_52 = W*in
   wire signed [9:0] m140_52;
   assign m140_52 =10'b0;

   // m140_53 = W*in
   wire signed [9:0] m140_53;
   assign m140_53 =10'b0;

   // m140_54 = W*in
   wire signed [9:0] m140_54;
   assign m140_54 =10'b0;

   // m140_55 = W*in
   wire signed [9:0] m140_55;
   assign m140_55 =10'b0;

   // m140_56 = W*in
   wire signed [9:0] m140_56;
   assign m140_56 =10'b0;

   // m140_57 = W*in
   wire signed [9:0] m140_57;
   assign m140_57 =10'b0;

   // m140_58 = W*in
   wire signed [9:0] m140_58;
   assign m140_58 =10'b0;

   // m140_59 = W*in
   wire signed [9:0] m140_59;
   assign m140_59 =10'b0;

   // m140_60 = W*in
   wire signed [9:0] m140_60;
   assign m140_60 =10'b0;

   // m140_61 = W*in
   wire signed [9:0] m140_61;
   assign m140_61 =10'b0;

   // m140_62 = W*in
   wire signed [9:0] m140_62;
   assign m140_62 =10'b0;

   // m140_63 = W*in
   wire signed [9:0] m140_63;
   assign m140_63 =10'b0;

   // m140_64 = W*in
   wire signed [9:0] m140_64;
   assign m140_64 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_65 = W*in
   wire signed [9:0] m140_65;
   assign m140_65 =10'b0;

   // m140_66 = W*in
   wire signed [9:0] m140_66;
   assign m140_66 =10'b0;

   // m140_67 = W*in
   wire signed [9:0] m140_67;
   assign m140_67 =10'b0;

   // m140_68 = W*in
   wire signed [9:0] m140_68;
   assign m140_68 =10'b0;

   // m140_69 = W*in
   wire signed [9:0] m140_69;
   assign m140_69 =10'b0;

   // m140_70 = W*in
   wire signed [9:0] m140_70;
   assign m140_70 ={ {5{in140[5]}} , in140[5:1] };

   // m140_71 = W*in
   wire signed [9:0] m140_71;
   assign m140_71 =10'b0;

   // m140_72 = W*in
   wire signed [9:0] m140_72;
   assign m140_72 =10'b0;

   // m140_73 = W*in
   wire signed [9:0] m140_73;
   assign m140_73 =10'b0;

   // m140_74 = W*in
   wire signed [9:0] m140_74;
   assign m140_74 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_75 = W*in
   wire signed [9:0] m140_75;
   assign m140_75 =10'b0;

   // m140_76 = W*in
   wire signed [9:0] m140_76;
   assign m140_76 =10'b0;

   // m140_77 = W*in
   wire signed [9:0] m140_77;
   assign m140_77 =10'b0;

   // m140_78 = W*in
   wire signed [9:0] m140_78;
   assign m140_78 =10'b0;

   // m140_79 = W*in
   wire signed [9:0] m140_79;
   assign m140_79 =10'b0;

   // m140_80 = W*in
   wire signed [9:0] m140_80;
   assign m140_80 =10'b0;

   // m140_81 = W*in
   wire signed [9:0] m140_81;
   assign m140_81 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_82 = W*in
   wire signed [9:0] m140_82;
   assign m140_82 =10'b0;

   // m140_83 = W*in
   wire signed [9:0] m140_83;
   assign m140_83 ={ {5{in140[5]}} , in140[5:1] };

   // m140_84 = W*in
   wire signed [9:0] m140_84;
   assign m140_84 =10'b0;

   // m140_85 = W*in
   wire signed [9:0] m140_85;
   assign m140_85 =10'b0;

   // m140_86 = W*in
   wire signed [9:0] m140_86;
   assign m140_86 =10'b0;

   // m140_87 = W*in
   wire signed [9:0] m140_87;
   assign m140_87 =10'b0;

   // m140_88 = W*in
   wire signed [9:0] m140_88;
   assign m140_88 =10'b0;

   // m140_89 = W*in
   wire signed [9:0] m140_89;
   assign m140_89 =10'b0;

   // m140_90 = W*in
   wire signed [9:0] m140_90;
   assign m140_90 =10'b0;

   // m140_91 = W*in
   wire signed [9:0] m140_91;
   assign m140_91 ={ {4{neg140[5]}} , neg140[5:0] };

   // m140_92 = W*in
   wire signed [9:0] m140_92;
   assign m140_92 =10'b0;

   // m140_93 = W*in
   wire signed [9:0] m140_93;
   assign m140_93 =10'b0;

   // m140_94 = W*in
   wire signed [9:0] m140_94;
   assign m140_94 =10'b0;

   // m140_95 = W*in
   wire signed [9:0] m140_95;
   assign m140_95 =10'b0;

   // m140_96 = W*in
   wire signed [9:0] m140_96;
   assign m140_96 =10'b0;

   // m140_97 = W*in
   wire signed [9:0] m140_97;
   assign m140_97 ={ {4{neg140[5]}} , neg140[5:0] };

   // m140_98 = W*in
   wire signed [9:0] m140_98;
   assign m140_98 =10'b0;

   // m140_99 = W*in
   wire signed [9:0] m140_99;
   assign m140_99 =10'b0;

   // m140_100 = W*in
   wire signed [9:0] m140_100;
   assign m140_100 =10'b0;

   // m140_101 = W*in
   wire signed [9:0] m140_101;
   assign m140_101 =10'b0;

   // m140_102 = W*in
   wire signed [9:0] m140_102;
   assign m140_102 =10'b0;

   // m140_103 = W*in
   wire signed [9:0] m140_103;
   assign m140_103 =10'b0;

   // m140_104 = W*in
   wire signed [9:0] m140_104;
   assign m140_104 =10'b0;

   // m140_105 = W*in
   wire signed [9:0] m140_105;
   assign m140_105 =10'b0;

   // m140_106 = W*in
   wire signed [9:0] m140_106;
   assign m140_106 =10'b0;

   // m140_107 = W*in
   wire signed [9:0] m140_107;
   assign m140_107 =10'b0;

   // m140_108 = W*in
   wire signed [9:0] m140_108;
   assign m140_108 ={ {4{neg140[5]}} , neg140[5:0] };

   // m140_109 = W*in
   wire signed [9:0] m140_109;
   assign m140_109 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_110 = W*in
   wire signed [9:0] m140_110;
   assign m140_110 ={ {4{neg140[5]}} , neg140[5:0] };

   // m140_111 = W*in
   wire signed [9:0] m140_111;
   assign m140_111 =10'b0;

   // m140_112 = W*in
   wire signed [9:0] m140_112;
   assign m140_112 =10'b0;

   // m140_113 = W*in
   wire signed [9:0] m140_113;
   assign m140_113 =10'b0;

   // m140_114 = W*in
   wire signed [9:0] m140_114;
   assign m140_114 ={ {5{neg140[5]}} , neg140[5:1] };

   // m140_115 = W*in
   wire signed [9:0] m140_115;
   assign m140_115 =10'b0;

   // m140_116 = W*in
   wire signed [9:0] m140_116;
   assign m140_116 =10'b0;

   // m140_117 = W*in
   wire signed [9:0] m140_117;
   assign m140_117 ={ {4{neg140[5]}} , neg140[5:0] };

   // m141_1 = W*in
   wire signed [9:0] m141_1;
   assign m141_1 =10'b0;

   // m141_2 = W*in
   wire signed [9:0] m141_2;
   assign m141_2 =10'b0;

   // m141_3 = W*in
   wire signed [9:0] m141_3;
   assign m141_3 =10'b0;

   // m141_4 = W*in
   wire signed [9:0] m141_4;
   assign m141_4 =10'b0;

   // m141_5 = W*in
   wire signed [9:0] m141_5;
   assign m141_5 =10'b0;

   // m141_6 = W*in
   wire signed [9:0] m141_6;
   assign m141_6 =10'b0;

   // m141_7 = W*in
   wire signed [9:0] m141_7;
   assign m141_7 =10'b0;

   // m141_8 = W*in
   wire signed [9:0] m141_8;
   assign m141_8 =10'b0;

   // m141_9 = W*in
   wire signed [9:0] m141_9;
   assign m141_9 =10'b0;

   // m141_10 = W*in
   wire signed [9:0] m141_10;
   assign m141_10 =10'b0;

   // m141_11 = W*in
   wire signed [9:0] m141_11;
   assign m141_11 =10'b0;

   // m141_12 = W*in
   wire signed [9:0] m141_12;
   assign m141_12 =10'b0;

   // m141_13 = W*in
   wire signed [9:0] m141_13;
   assign m141_13 =10'b0;

   // m141_14 = W*in
   wire signed [9:0] m141_14;
   assign m141_14 =10'b0;

   // m141_15 = W*in
   wire signed [9:0] m141_15;
   assign m141_15 =10'b0;

   // m141_16 = W*in
   wire signed [9:0] m141_16;
   assign m141_16 =10'b0;

   // m141_17 = W*in
   wire signed [9:0] m141_17;
   assign m141_17 =10'b0;

   // m141_18 = W*in
   wire signed [9:0] m141_18;
   assign m141_18 =10'b0;

   // m141_19 = W*in
   wire signed [9:0] m141_19;
   assign m141_19 ={ {4{in141[5]}} , in141[5:0] };

   // m141_20 = W*in
   wire signed [9:0] m141_20;
   assign m141_20 ={ {5{neg141[5]}} , neg141[5:1] };

   // m141_21 = W*in
   wire signed [9:0] m141_21;
   assign m141_21 ={ {4{in141[5]}} , in141[5:0] };

   // m141_22 = W*in
   wire signed [9:0] m141_22;
   assign m141_22 ={ {5{neg141[5]}} , neg141[5:1] };

   // m141_23 = W*in
   wire signed [9:0] m141_23;
   assign m141_23 ={ {5{neg141[5]}} , neg141[5:1] };

   // m141_24 = W*in
   wire signed [9:0] m141_24;
   assign m141_24 =10'b0;

   // m141_25 = W*in
   wire signed [9:0] m141_25;
   assign m141_25 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_26 = W*in
   wire signed [9:0] m141_26;
   assign m141_26 =10'b0;

   // m141_27 = W*in
   wire signed [9:0] m141_27;
   assign m141_27 =10'b0;

   // m141_28 = W*in
   wire signed [9:0] m141_28;
   assign m141_28 =10'b0;

   // m141_29 = W*in
   wire signed [9:0] m141_29;
   assign m141_29 ={ {4{in141[5]}} , in141[5:0] };

   // m141_30 = W*in
   wire signed [9:0] m141_30;
   assign m141_30 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_31 = W*in
   wire signed [9:0] m141_31;
   assign m141_31 ={ {5{in141[5]}} , in141[5:1] };

   // m141_32 = W*in
   wire signed [9:0] m141_32;
   assign m141_32 =10'b0;

   // m141_33 = W*in
   wire signed [9:0] m141_33;
   assign m141_33 =10'b0;

   // m141_34 = W*in
   wire signed [9:0] m141_34;
   assign m141_34 =10'b0;

   // m141_35 = W*in
   wire signed [9:0] m141_35;
   assign m141_35 =10'b0;

   // m141_36 = W*in
   wire signed [9:0] m141_36;
   assign m141_36 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_37 = W*in
   wire signed [9:0] m141_37;
   assign m141_37 ={ {4{in141[5]}} , in141[5:0] };

   // m141_38 = W*in
   wire signed [9:0] m141_38;
   assign m141_38 =10'b0;

   // m141_39 = W*in
   wire signed [9:0] m141_39;
   assign m141_39 =10'b0;

   // m141_40 = W*in
   wire signed [9:0] m141_40;
   assign m141_40 =10'b0;

   // m141_41 = W*in
   wire signed [9:0] m141_41;
   assign m141_41 =10'b0;

   // m141_42 = W*in
   wire signed [9:0] m141_42;
   assign m141_42 =10'b0;

   // m141_43 = W*in
   wire signed [9:0] m141_43;
   assign m141_43 =10'b0;

   // m141_44 = W*in
   wire signed [9:0] m141_44;
   assign m141_44 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_45 = W*in
   wire signed [9:0] m141_45;
   assign m141_45 =10'b0;

   // m141_46 = W*in
   wire signed [9:0] m141_46;
   assign m141_46 =10'b0;

   // m141_47 = W*in
   wire signed [9:0] m141_47;
   assign m141_47 =10'b0;

   // m141_48 = W*in
   wire signed [9:0] m141_48;
   assign m141_48 =10'b0;

   // m141_49 = W*in
   wire signed [9:0] m141_49;
   assign m141_49 =10'b0;

   // m141_50 = W*in
   wire signed [9:0] m141_50;
   assign m141_50 =10'b0;

   // m141_51 = W*in
   wire signed [9:0] m141_51;
   assign m141_51 =10'b0;

   // m141_52 = W*in
   wire signed [9:0] m141_52;
   assign m141_52 =10'b0;

   // m141_53 = W*in
   wire signed [9:0] m141_53;
   assign m141_53 =10'b0;

   // m141_54 = W*in
   wire signed [9:0] m141_54;
   assign m141_54 =10'b0;

   // m141_55 = W*in
   wire signed [9:0] m141_55;
   assign m141_55 =10'b0;

   // m141_56 = W*in
   wire signed [9:0] m141_56;
   assign m141_56 =10'b0;

   // m141_57 = W*in
   wire signed [9:0] m141_57;
   assign m141_57 =10'b0;

   // m141_58 = W*in
   wire signed [9:0] m141_58;
   assign m141_58 =10'b0;

   // m141_59 = W*in
   wire signed [9:0] m141_59;
   assign m141_59 =10'b0;

   // m141_60 = W*in
   wire signed [9:0] m141_60;
   assign m141_60 =10'b0;

   // m141_61 = W*in
   wire signed [9:0] m141_61;
   assign m141_61 =10'b0;

   // m141_62 = W*in
   wire signed [9:0] m141_62;
   assign m141_62 =10'b0;

   // m141_63 = W*in
   wire signed [9:0] m141_63;
   assign m141_63 =10'b0;

   // m141_64 = W*in
   wire signed [9:0] m141_64;
   assign m141_64 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_65 = W*in
   wire signed [9:0] m141_65;
   assign m141_65 =10'b0;

   // m141_66 = W*in
   wire signed [9:0] m141_66;
   assign m141_66 =10'b0;

   // m141_67 = W*in
   wire signed [9:0] m141_67;
   assign m141_67 ={ {4{in141[5]}} , in141[5:0] };

   // m141_68 = W*in
   wire signed [9:0] m141_68;
   assign m141_68 =10'b0;

   // m141_69 = W*in
   wire signed [9:0] m141_69;
   assign m141_69 ={ {4{in141[5]}} , in141[5:0] };

   // m141_70 = W*in
   wire signed [9:0] m141_70;
   assign m141_70 ={ {4{in141[5]}} , in141[5:0] };

   // m141_71 = W*in
   wire signed [9:0] m141_71;
   assign m141_71 =10'b0;

   // m141_72 = W*in
   wire signed [9:0] m141_72;
   assign m141_72 =10'b0;

   // m141_73 = W*in
   wire signed [9:0] m141_73;
   assign m141_73 =10'b0;

   // m141_74 = W*in
   wire signed [9:0] m141_74;
   assign m141_74 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_75 = W*in
   wire signed [9:0] m141_75;
   assign m141_75 ={ {5{neg141[5]}} , neg141[5:1] };

   // m141_76 = W*in
   wire signed [9:0] m141_76;
   assign m141_76 =10'b0;

   // m141_77 = W*in
   wire signed [9:0] m141_77;
   assign m141_77 =10'b0;

   // m141_78 = W*in
   wire signed [9:0] m141_78;
   assign m141_78 ={ {5{in141[5]}} , in141[5:1] };

   // m141_79 = W*in
   wire signed [9:0] m141_79;
   assign m141_79 =10'b0;

   // m141_80 = W*in
   wire signed [9:0] m141_80;
   assign m141_80 =10'b0;

   // m141_81 = W*in
   wire signed [9:0] m141_81;
   assign m141_81 ={ {5{neg141[5]}} , neg141[5:1] };

   // m141_82 = W*in
   wire signed [9:0] m141_82;
   assign m141_82 ={ {4{in141[5]}} , in141[5:0] };

   // m141_83 = W*in
   wire signed [9:0] m141_83;
   assign m141_83 =10'b0;

   // m141_84 = W*in
   wire signed [9:0] m141_84;
   assign m141_84 =10'b0;

   // m141_85 = W*in
   wire signed [9:0] m141_85;
   assign m141_85 ={ {4{in141[5]}} , in141[5:0] };

   // m141_86 = W*in
   wire signed [9:0] m141_86;
   assign m141_86 =10'b0;

   // m141_87 = W*in
   wire signed [9:0] m141_87;
   assign m141_87 =10'b0;

   // m141_88 = W*in
   wire signed [9:0] m141_88;
   assign m141_88 ={ {4{in141[5]}} , in141[5:0] };

   // m141_89 = W*in
   wire signed [9:0] m141_89;
   assign m141_89 =10'b0;

   // m141_90 = W*in
   wire signed [9:0] m141_90;
   assign m141_90 =10'b0;

   // m141_91 = W*in
   wire signed [9:0] m141_91;
   assign m141_91 =10'b0;

   // m141_92 = W*in
   wire signed [9:0] m141_92;
   assign m141_92 ={ {4{in141[5]}} , in141[5:0] };

   // m141_93 = W*in
   wire signed [9:0] m141_93;
   assign m141_93 =10'b0;

   // m141_94 = W*in
   wire signed [9:0] m141_94;
   assign m141_94 =10'b0;

   // m141_95 = W*in
   wire signed [9:0] m141_95;
   assign m141_95 =10'b0;

   // m141_96 = W*in
   wire signed [9:0] m141_96;
   assign m141_96 =10'b0;

   // m141_97 = W*in
   wire signed [9:0] m141_97;
   assign m141_97 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_98 = W*in
   wire signed [9:0] m141_98;
   assign m141_98 =10'b0;

   // m141_99 = W*in
   wire signed [9:0] m141_99;
   assign m141_99 =10'b0;

   // m141_100 = W*in
   wire signed [9:0] m141_100;
   assign m141_100 =10'b0;

   // m141_101 = W*in
   wire signed [9:0] m141_101;
   assign m141_101 =10'b0;

   // m141_102 = W*in
   wire signed [9:0] m141_102;
   assign m141_102 =10'b0;

   // m141_103 = W*in
   wire signed [9:0] m141_103;
   assign m141_103 =10'b0;

   // m141_104 = W*in
   wire signed [9:0] m141_104;
   assign m141_104 =10'b0;

   // m141_105 = W*in
   wire signed [9:0] m141_105;
   assign m141_105 =10'b0;

   // m141_106 = W*in
   wire signed [9:0] m141_106;
   assign m141_106 =10'b0;

   // m141_107 = W*in
   wire signed [9:0] m141_107;
   assign m141_107 =10'b0;

   // m141_108 = W*in
   wire signed [9:0] m141_108;
   assign m141_108 =10'b0;

   // m141_109 = W*in
   wire signed [9:0] m141_109;
   assign m141_109 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_110 = W*in
   wire signed [9:0] m141_110;
   assign m141_110 ={ {4{neg141[5]}} , neg141[5:0] };

   // m141_111 = W*in
   wire signed [9:0] m141_111;
   assign m141_111 =10'b0;

   // m141_112 = W*in
   wire signed [9:0] m141_112;
   assign m141_112 =10'b0;

   // m141_113 = W*in
   wire signed [9:0] m141_113;
   assign m141_113 =10'b0;

   // m141_114 = W*in
   wire signed [9:0] m141_114;
   assign m141_114 ={ {5{neg141[5]}} , neg141[5:1] };

   // m141_115 = W*in
   wire signed [9:0] m141_115;
   assign m141_115 =10'b0;

   // m141_116 = W*in
   wire signed [9:0] m141_116;
   assign m141_116 =10'b0;

   // m141_117 = W*in
   wire signed [9:0] m141_117;
   assign m141_117 =10'b0;

   // m142_1 = W*in
   wire signed [9:0] m142_1;
   assign m142_1 =10'b0;

   // m142_2 = W*in
   wire signed [9:0] m142_2;
   assign m142_2 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_3 = W*in
   wire signed [9:0] m142_3;
   assign m142_3 =10'b0;

   // m142_4 = W*in
   wire signed [9:0] m142_4;
   assign m142_4 =10'b0;

   // m142_5 = W*in
   wire signed [9:0] m142_5;
   assign m142_5 =10'b0;

   // m142_6 = W*in
   wire signed [9:0] m142_6;
   assign m142_6 =10'b0;

   // m142_7 = W*in
   wire signed [9:0] m142_7;
   assign m142_7 =10'b0;

   // m142_8 = W*in
   wire signed [9:0] m142_8;
   assign m142_8 =10'b0;

   // m142_9 = W*in
   wire signed [9:0] m142_9;
   assign m142_9 =10'b0;

   // m142_10 = W*in
   wire signed [9:0] m142_10;
   assign m142_10 =10'b0;

   // m142_11 = W*in
   wire signed [9:0] m142_11;
   assign m142_11 ={ {4{in142[5]}} , in142[5:0] };

   // m142_12 = W*in
   wire signed [9:0] m142_12;
   assign m142_12 =10'b0;

   // m142_13 = W*in
   wire signed [9:0] m142_13;
   assign m142_13 =10'b0;

   // m142_14 = W*in
   wire signed [9:0] m142_14;
   assign m142_14 =10'b0;

   // m142_15 = W*in
   wire signed [9:0] m142_15;
   assign m142_15 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_16 = W*in
   wire signed [9:0] m142_16;
   assign m142_16 =10'b0;

   // m142_17 = W*in
   wire signed [9:0] m142_17;
   assign m142_17 =10'b0;

   // m142_18 = W*in
   wire signed [9:0] m142_18;
   assign m142_18 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_19 = W*in
   wire signed [9:0] m142_19;
   assign m142_19 =10'b0;

   // m142_20 = W*in
   wire signed [9:0] m142_20;
   assign m142_20 =10'b0;

   // m142_21 = W*in
   wire signed [9:0] m142_21;
   assign m142_21 ={ {5{in142[5]}} , in142[5:1] };

   // m142_22 = W*in
   wire signed [9:0] m142_22;
   assign m142_22 =10'b0;

   // m142_23 = W*in
   wire signed [9:0] m142_23;
   assign m142_23 =10'b0;

   // m142_24 = W*in
   wire signed [9:0] m142_24;
   assign m142_24 =10'b0;

   // m142_25 = W*in
   wire signed [9:0] m142_25;
   assign m142_25 =10'b0;

   // m142_26 = W*in
   wire signed [9:0] m142_26;
   assign m142_26 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_27 = W*in
   wire signed [9:0] m142_27;
   assign m142_27 =10'b0;

   // m142_28 = W*in
   wire signed [9:0] m142_28;
   assign m142_28 =10'b0;

   // m142_29 = W*in
   wire signed [9:0] m142_29;
   assign m142_29 ={ {4{in142[5]}} , in142[5:0] };

   // m142_30 = W*in
   wire signed [9:0] m142_30;
   assign m142_30 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_31 = W*in
   wire signed [9:0] m142_31;
   assign m142_31 ={ {5{neg142[5]}} , neg142[5:1] };

   // m142_32 = W*in
   wire signed [9:0] m142_32;
   assign m142_32 =10'b0;

   // m142_33 = W*in
   wire signed [9:0] m142_33;
   assign m142_33 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_34 = W*in
   wire signed [9:0] m142_34;
   assign m142_34 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_35 = W*in
   wire signed [9:0] m142_35;
   assign m142_35 =10'b0;

   // m142_36 = W*in
   wire signed [9:0] m142_36;
   assign m142_36 =10'b0;

   // m142_37 = W*in
   wire signed [9:0] m142_37;
   assign m142_37 ={ {4{in142[5]}} , in142[5:0] };

   // m142_38 = W*in
   wire signed [9:0] m142_38;
   assign m142_38 ={ {4{in142[5]}} , in142[5:0] };

   // m142_39 = W*in
   wire signed [9:0] m142_39;
   assign m142_39 =10'b0;

   // m142_40 = W*in
   wire signed [9:0] m142_40;
   assign m142_40 =10'b0;

   // m142_41 = W*in
   wire signed [9:0] m142_41;
   assign m142_41 =10'b0;

   // m142_42 = W*in
   wire signed [9:0] m142_42;
   assign m142_42 =10'b0;

   // m142_43 = W*in
   wire signed [9:0] m142_43;
   assign m142_43 =10'b0;

   // m142_44 = W*in
   wire signed [9:0] m142_44;
   assign m142_44 =10'b0;

   // m142_45 = W*in
   wire signed [9:0] m142_45;
   assign m142_45 =10'b0;

   // m142_46 = W*in
   wire signed [9:0] m142_46;
   assign m142_46 =10'b0;

   // m142_47 = W*in
   wire signed [9:0] m142_47;
   assign m142_47 =10'b0;

   // m142_48 = W*in
   wire signed [9:0] m142_48;
   assign m142_48 =10'b0;

   // m142_49 = W*in
   wire signed [9:0] m142_49;
   assign m142_49 ={ {4{in142[5]}} , in142[5:0] };

   // m142_50 = W*in
   wire signed [9:0] m142_50;
   assign m142_50 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_51 = W*in
   wire signed [9:0] m142_51;
   assign m142_51 =10'b0;

   // m142_52 = W*in
   wire signed [9:0] m142_52;
   assign m142_52 =10'b0;

   // m142_53 = W*in
   wire signed [9:0] m142_53;
   assign m142_53 =10'b0;

   // m142_54 = W*in
   wire signed [9:0] m142_54;
   assign m142_54 ={ {4{in142[5]}} , in142[5:0] };

   // m142_55 = W*in
   wire signed [9:0] m142_55;
   assign m142_55 =10'b0;

   // m142_56 = W*in
   wire signed [9:0] m142_56;
   assign m142_56 =10'b0;

   // m142_57 = W*in
   wire signed [9:0] m142_57;
   assign m142_57 =10'b0;

   // m142_58 = W*in
   wire signed [9:0] m142_58;
   assign m142_58 ={ {5{in142[5]}} , in142[5:1] };

   // m142_59 = W*in
   wire signed [9:0] m142_59;
   assign m142_59 =10'b0;

   // m142_60 = W*in
   wire signed [9:0] m142_60;
   assign m142_60 =10'b0;

   // m142_61 = W*in
   wire signed [9:0] m142_61;
   assign m142_61 =10'b0;

   // m142_62 = W*in
   wire signed [9:0] m142_62;
   assign m142_62 =10'b0;

   // m142_63 = W*in
   wire signed [9:0] m142_63;
   assign m142_63 ={ {4{in142[5]}} , in142[5:0] };

   // m142_64 = W*in
   wire signed [9:0] m142_64;
   assign m142_64 =10'b0;

   // m142_65 = W*in
   wire signed [9:0] m142_65;
   assign m142_65 ={ {5{neg142[5]}} , neg142[5:1] };

   // m142_66 = W*in
   wire signed [9:0] m142_66;
   assign m142_66 =10'b0;

   // m142_67 = W*in
   wire signed [9:0] m142_67;
   assign m142_67 ={ {4{in142[5]}} , in142[5:0] };

   // m142_68 = W*in
   wire signed [9:0] m142_68;
   assign m142_68 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_69 = W*in
   wire signed [9:0] m142_69;
   assign m142_69 ={ {4{in142[5]}} , in142[5:0] };

   // m142_70 = W*in
   wire signed [9:0] m142_70;
   assign m142_70 ={ {5{in142[5]}} , in142[5:1] };

   // m142_71 = W*in
   wire signed [9:0] m142_71;
   assign m142_71 =10'b0;

   // m142_72 = W*in
   wire signed [9:0] m142_72;
   assign m142_72 =10'b0;

   // m142_73 = W*in
   wire signed [9:0] m142_73;
   assign m142_73 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_74 = W*in
   wire signed [9:0] m142_74;
   assign m142_74 =10'b0;

   // m142_75 = W*in
   wire signed [9:0] m142_75;
   assign m142_75 ={ {5{neg142[5]}} , neg142[5:1] };

   // m142_76 = W*in
   wire signed [9:0] m142_76;
   assign m142_76 =10'b0;

   // m142_77 = W*in
   wire signed [9:0] m142_77;
   assign m142_77 =10'b0;

   // m142_78 = W*in
   wire signed [9:0] m142_78;
   assign m142_78 =10'b0;

   // m142_79 = W*in
   wire signed [9:0] m142_79;
   assign m142_79 =10'b0;

   // m142_80 = W*in
   wire signed [9:0] m142_80;
   assign m142_80 =10'b0;

   // m142_81 = W*in
   wire signed [9:0] m142_81;
   assign m142_81 =10'b0;

   // m142_82 = W*in
   wire signed [9:0] m142_82;
   assign m142_82 ={ {4{in142[5]}} , in142[5:0] };

   // m142_83 = W*in
   wire signed [9:0] m142_83;
   assign m142_83 =10'b0;

   // m142_84 = W*in
   wire signed [9:0] m142_84;
   assign m142_84 =10'b0;

   // m142_85 = W*in
   wire signed [9:0] m142_85;
   assign m142_85 ={ {4{in142[5]}} , in142[5:0] };

   // m142_86 = W*in
   wire signed [9:0] m142_86;
   assign m142_86 =10'b0;

   // m142_87 = W*in
   wire signed [9:0] m142_87;
   assign m142_87 =10'b0;

   // m142_88 = W*in
   wire signed [9:0] m142_88;
   assign m142_88 =10'b0;

   // m142_89 = W*in
   wire signed [9:0] m142_89;
   assign m142_89 =10'b0;

   // m142_90 = W*in
   wire signed [9:0] m142_90;
   assign m142_90 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_91 = W*in
   wire signed [9:0] m142_91;
   assign m142_91 ={ {4{in142[5]}} , in142[5:0] };

   // m142_92 = W*in
   wire signed [9:0] m142_92;
   assign m142_92 =10'b0;

   // m142_93 = W*in
   wire signed [9:0] m142_93;
   assign m142_93 =10'b0;

   // m142_94 = W*in
   wire signed [9:0] m142_94;
   assign m142_94 =10'b0;

   // m142_95 = W*in
   wire signed [9:0] m142_95;
   assign m142_95 ={ {4{in142[5]}} , in142[5:0] };

   // m142_96 = W*in
   wire signed [9:0] m142_96;
   assign m142_96 =10'b0;

   // m142_97 = W*in
   wire signed [9:0] m142_97;
   assign m142_97 =10'b0;

   // m142_98 = W*in
   wire signed [9:0] m142_98;
   assign m142_98 =10'b0;

   // m142_99 = W*in
   wire signed [9:0] m142_99;
   assign m142_99 =10'b0;

   // m142_100 = W*in
   wire signed [9:0] m142_100;
   assign m142_100 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_101 = W*in
   wire signed [9:0] m142_101;
   assign m142_101 =10'b0;

   // m142_102 = W*in
   wire signed [9:0] m142_102;
   assign m142_102 =10'b0;

   // m142_103 = W*in
   wire signed [9:0] m142_103;
   assign m142_103 =10'b0;

   // m142_104 = W*in
   wire signed [9:0] m142_104;
   assign m142_104 =10'b0;

   // m142_105 = W*in
   wire signed [9:0] m142_105;
   assign m142_105 =10'b0;

   // m142_106 = W*in
   wire signed [9:0] m142_106;
   assign m142_106 =10'b0;

   // m142_107 = W*in
   wire signed [9:0] m142_107;
   assign m142_107 =10'b0;

   // m142_108 = W*in
   wire signed [9:0] m142_108;
   assign m142_108 =10'b0;

   // m142_109 = W*in
   wire signed [9:0] m142_109;
   assign m142_109 =10'b0;

   // m142_110 = W*in
   wire signed [9:0] m142_110;
   assign m142_110 =10'b0;

   // m142_111 = W*in
   wire signed [9:0] m142_111;
   assign m142_111 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_112 = W*in
   wire signed [9:0] m142_112;
   assign m142_112 =10'b0;

   // m142_113 = W*in
   wire signed [9:0] m142_113;
   assign m142_113 ={ {4{neg142[5]}} , neg142[5:0] };

   // m142_114 = W*in
   wire signed [9:0] m142_114;
   assign m142_114 =10'b0;

   // m142_115 = W*in
   wire signed [9:0] m142_115;
   assign m142_115 =10'b0;

   // m142_116 = W*in
   wire signed [9:0] m142_116;
   assign m142_116 =10'b0;

   // m142_117 = W*in
   wire signed [9:0] m142_117;
   assign m142_117 =10'b0;

   // m143_1 = W*in
   wire signed [9:0] m143_1;
   assign m143_1 =10'b0;

   // m143_2 = W*in
   wire signed [9:0] m143_2;
   assign m143_2 =10'b0;

   // m143_3 = W*in
   wire signed [9:0] m143_3;
   assign m143_3 =10'b0;

   // m143_4 = W*in
   wire signed [9:0] m143_4;
   assign m143_4 =10'b0;

   // m143_5 = W*in
   wire signed [9:0] m143_5;
   assign m143_5 =10'b0;

   // m143_6 = W*in
   wire signed [9:0] m143_6;
   assign m143_6 ={ {5{in143[5]}} , in143[5:1] };

   // m143_7 = W*in
   wire signed [9:0] m143_7;
   assign m143_7 =10'b0;

   // m143_8 = W*in
   wire signed [9:0] m143_8;
   assign m143_8 =10'b0;

   // m143_9 = W*in
   wire signed [9:0] m143_9;
   assign m143_9 =10'b0;

   // m143_10 = W*in
   wire signed [9:0] m143_10;
   assign m143_10 =10'b0;

   // m143_11 = W*in
   wire signed [9:0] m143_11;
   assign m143_11 =10'b0;

   // m143_12 = W*in
   wire signed [9:0] m143_12;
   assign m143_12 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_13 = W*in
   wire signed [9:0] m143_13;
   assign m143_13 =10'b0;

   // m143_14 = W*in
   wire signed [9:0] m143_14;
   assign m143_14 =10'b0;

   // m143_15 = W*in
   wire signed [9:0] m143_15;
   assign m143_15 =10'b0;

   // m143_16 = W*in
   wire signed [9:0] m143_16;
   assign m143_16 =10'b0;

   // m143_17 = W*in
   wire signed [9:0] m143_17;
   assign m143_17 =10'b0;

   // m143_18 = W*in
   wire signed [9:0] m143_18;
   assign m143_18 =10'b0;

   // m143_19 = W*in
   wire signed [9:0] m143_19;
   assign m143_19 =10'b0;

   // m143_20 = W*in
   wire signed [9:0] m143_20;
   assign m143_20 =10'b0;

   // m143_21 = W*in
   wire signed [9:0] m143_21;
   assign m143_21 ={ {4{in143[5]}} , in143[5:0] };

   // m143_22 = W*in
   wire signed [9:0] m143_22;
   assign m143_22 ={ {5{in143[5]}} , in143[5:1] };

   // m143_23 = W*in
   wire signed [9:0] m143_23;
   assign m143_23 ={ {4{in143[5]}} , in143[5:0] };

   // m143_24 = W*in
   wire signed [9:0] m143_24;
   assign m143_24 ={ {4{in143[5]}} , in143[5:0] };

   // m143_25 = W*in
   wire signed [9:0] m143_25;
   assign m143_25 =10'b0;

   // m143_26 = W*in
   wire signed [9:0] m143_26;
   assign m143_26 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_27 = W*in
   wire signed [9:0] m143_27;
   assign m143_27 =10'b0;

   // m143_28 = W*in
   wire signed [9:0] m143_28;
   assign m143_28 ={ {5{neg143[5]}} , neg143[5:1] };

   // m143_29 = W*in
   wire signed [9:0] m143_29;
   assign m143_29 =10'b0;

   // m143_30 = W*in
   wire signed [9:0] m143_30;
   assign m143_30 =10'b0;

   // m143_31 = W*in
   wire signed [9:0] m143_31;
   assign m143_31 ={ {5{neg143[5]}} , neg143[5:1] };

   // m143_32 = W*in
   wire signed [9:0] m143_32;
   assign m143_32 =10'b0;

   // m143_33 = W*in
   wire signed [9:0] m143_33;
   assign m143_33 =10'b0;

   // m143_34 = W*in
   wire signed [9:0] m143_34;
   assign m143_34 =10'b0;

   // m143_35 = W*in
   wire signed [9:0] m143_35;
   assign m143_35 =10'b0;

   // m143_36 = W*in
   wire signed [9:0] m143_36;
   assign m143_36 =10'b0;

   // m143_37 = W*in
   wire signed [9:0] m143_37;
   assign m143_37 ={ {4{in143[5]}} , in143[5:0] };

   // m143_38 = W*in
   wire signed [9:0] m143_38;
   assign m143_38 =10'b0;

   // m143_39 = W*in
   wire signed [9:0] m143_39;
   assign m143_39 =10'b0;

   // m143_40 = W*in
   wire signed [9:0] m143_40;
   assign m143_40 =10'b0;

   // m143_41 = W*in
   wire signed [9:0] m143_41;
   assign m143_41 =10'b0;

   // m143_42 = W*in
   wire signed [9:0] m143_42;
   assign m143_42 =10'b0;

   // m143_43 = W*in
   wire signed [9:0] m143_43;
   assign m143_43 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_44 = W*in
   wire signed [9:0] m143_44;
   assign m143_44 ={ {4{in143[5]}} , in143[5:0] };

   // m143_45 = W*in
   wire signed [9:0] m143_45;
   assign m143_45 =10'b0;

   // m143_46 = W*in
   wire signed [9:0] m143_46;
   assign m143_46 ={ {4{in143[5]}} , in143[5:0] };

   // m143_47 = W*in
   wire signed [9:0] m143_47;
   assign m143_47 =10'b0;

   // m143_48 = W*in
   wire signed [9:0] m143_48;
   assign m143_48 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_49 = W*in
   wire signed [9:0] m143_49;
   assign m143_49 ={ {4{in143[5]}} , in143[5:0] };

   // m143_50 = W*in
   wire signed [9:0] m143_50;
   assign m143_50 =10'b0;

   // m143_51 = W*in
   wire signed [9:0] m143_51;
   assign m143_51 =10'b0;

   // m143_52 = W*in
   wire signed [9:0] m143_52;
   assign m143_52 =10'b0;

   // m143_53 = W*in
   wire signed [9:0] m143_53;
   assign m143_53 =10'b0;

   // m143_54 = W*in
   wire signed [9:0] m143_54;
   assign m143_54 =10'b0;

   // m143_55 = W*in
   wire signed [9:0] m143_55;
   assign m143_55 =10'b0;

   // m143_56 = W*in
   wire signed [9:0] m143_56;
   assign m143_56 =10'b0;

   // m143_57 = W*in
   wire signed [9:0] m143_57;
   assign m143_57 =10'b0;

   // m143_58 = W*in
   wire signed [9:0] m143_58;
   assign m143_58 =10'b0;

   // m143_59 = W*in
   wire signed [9:0] m143_59;
   assign m143_59 =10'b0;

   // m143_60 = W*in
   wire signed [9:0] m143_60;
   assign m143_60 =10'b0;

   // m143_61 = W*in
   wire signed [9:0] m143_61;
   assign m143_61 =10'b0;

   // m143_62 = W*in
   wire signed [9:0] m143_62;
   assign m143_62 =10'b0;

   // m143_63 = W*in
   wire signed [9:0] m143_63;
   assign m143_63 ={ {4{in143[5]}} , in143[5:0] };

   // m143_64 = W*in
   wire signed [9:0] m143_64;
   assign m143_64 =10'b0;

   // m143_65 = W*in
   wire signed [9:0] m143_65;
   assign m143_65 ={ {4{in143[5]}} , in143[5:0] };

   // m143_66 = W*in
   wire signed [9:0] m143_66;
   assign m143_66 =10'b0;

   // m143_67 = W*in
   wire signed [9:0] m143_67;
   assign m143_67 ={ {4{in143[5]}} , in143[5:0] };

   // m143_68 = W*in
   wire signed [9:0] m143_68;
   assign m143_68 =10'b0;

   // m143_69 = W*in
   wire signed [9:0] m143_69;
   assign m143_69 ={ {4{in143[5]}} , in143[5:0] };

   // m143_70 = W*in
   wire signed [9:0] m143_70;
   assign m143_70 ={ {4{in143[5]}} , in143[5:0] };

   // m143_71 = W*in
   wire signed [9:0] m143_71;
   assign m143_71 =10'b0;

   // m143_72 = W*in
   wire signed [9:0] m143_72;
   assign m143_72 =10'b0;

   // m143_73 = W*in
   wire signed [9:0] m143_73;
   assign m143_73 =10'b0;

   // m143_74 = W*in
   wire signed [9:0] m143_74;
   assign m143_74 ={ {5{neg143[5]}} , neg143[5:1] };

   // m143_75 = W*in
   wire signed [9:0] m143_75;
   assign m143_75 =10'b0;

   // m143_76 = W*in
   wire signed [9:0] m143_76;
   assign m143_76 =10'b0;

   // m143_77 = W*in
   wire signed [9:0] m143_77;
   assign m143_77 =10'b0;

   // m143_78 = W*in
   wire signed [9:0] m143_78;
   assign m143_78 ={ {5{neg143[5]}} , neg143[5:1] };

   // m143_79 = W*in
   wire signed [9:0] m143_79;
   assign m143_79 =10'b0;

   // m143_80 = W*in
   wire signed [9:0] m143_80;
   assign m143_80 =10'b0;

   // m143_81 = W*in
   wire signed [9:0] m143_81;
   assign m143_81 =10'b0;

   // m143_82 = W*in
   wire signed [9:0] m143_82;
   assign m143_82 ={ {4{in143[5]}} , in143[5:0] };

   // m143_83 = W*in
   wire signed [9:0] m143_83;
   assign m143_83 =10'b0;

   // m143_84 = W*in
   wire signed [9:0] m143_84;
   assign m143_84 =10'b0;

   // m143_85 = W*in
   wire signed [9:0] m143_85;
   assign m143_85 ={ {4{in143[5]}} , in143[5:0] };

   // m143_86 = W*in
   wire signed [9:0] m143_86;
   assign m143_86 =10'b0;

   // m143_87 = W*in
   wire signed [9:0] m143_87;
   assign m143_87 =10'b0;

   // m143_88 = W*in
   wire signed [9:0] m143_88;
   assign m143_88 =10'b0;

   // m143_89 = W*in
   wire signed [9:0] m143_89;
   assign m143_89 ={ {4{in143[5]}} , in143[5:0] };

   // m143_90 = W*in
   wire signed [9:0] m143_90;
   assign m143_90 =10'b0;

   // m143_91 = W*in
   wire signed [9:0] m143_91;
   assign m143_91 =10'b0;

   // m143_92 = W*in
   wire signed [9:0] m143_92;
   assign m143_92 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_93 = W*in
   wire signed [9:0] m143_93;
   assign m143_93 ={ {4{in143[5]}} , in143[5:0] };

   // m143_94 = W*in
   wire signed [9:0] m143_94;
   assign m143_94 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_95 = W*in
   wire signed [9:0] m143_95;
   assign m143_95 =10'b0;

   // m143_96 = W*in
   wire signed [9:0] m143_96;
   assign m143_96 =10'b0;

   // m143_97 = W*in
   wire signed [9:0] m143_97;
   assign m143_97 =10'b0;

   // m143_98 = W*in
   wire signed [9:0] m143_98;
   assign m143_98 =10'b0;

   // m143_99 = W*in
   wire signed [9:0] m143_99;
   assign m143_99 =10'b0;

   // m143_100 = W*in
   wire signed [9:0] m143_100;
   assign m143_100 =10'b0;

   // m143_101 = W*in
   wire signed [9:0] m143_101;
   assign m143_101 =10'b0;

   // m143_102 = W*in
   wire signed [9:0] m143_102;
   assign m143_102 =10'b0;

   // m143_103 = W*in
   wire signed [9:0] m143_103;
   assign m143_103 =10'b0;

   // m143_104 = W*in
   wire signed [9:0] m143_104;
   assign m143_104 =10'b0;

   // m143_105 = W*in
   wire signed [9:0] m143_105;
   assign m143_105 =10'b0;

   // m143_106 = W*in
   wire signed [9:0] m143_106;
   assign m143_106 =10'b0;

   // m143_107 = W*in
   wire signed [9:0] m143_107;
   assign m143_107 ={ {5{neg143[5]}} , neg143[5:1] };

   // m143_108 = W*in
   wire signed [9:0] m143_108;
   assign m143_108 =10'b0;

   // m143_109 = W*in
   wire signed [9:0] m143_109;
   assign m143_109 ={ {4{in143[5]}} , in143[5:0] };

   // m143_110 = W*in
   wire signed [9:0] m143_110;
   assign m143_110 ={ {4{in143[5]}} , in143[5:0] };

   // m143_111 = W*in
   wire signed [9:0] m143_111;
   assign m143_111 =10'b0;

   // m143_112 = W*in
   wire signed [9:0] m143_112;
   assign m143_112 =10'b0;

   // m143_113 = W*in
   wire signed [9:0] m143_113;
   assign m143_113 ={ {4{neg143[5]}} , neg143[5:0] };

   // m143_114 = W*in
   wire signed [9:0] m143_114;
   assign m143_114 =10'b0;

   // m143_115 = W*in
   wire signed [9:0] m143_115;
   assign m143_115 =10'b0;

   // m143_116 = W*in
   wire signed [9:0] m143_116;
   assign m143_116 =10'b0;

   // m143_117 = W*in
   wire signed [9:0] m143_117;
   assign m143_117 =10'b0;

   // m144_1 = W*in
   wire signed [9:0] m144_1;
   assign m144_1 =10'b0;

   // m144_2 = W*in
   wire signed [9:0] m144_2;
   assign m144_2 =10'b0;

   // m144_3 = W*in
   wire signed [9:0] m144_3;
   assign m144_3 =10'b0;

   // m144_4 = W*in
   wire signed [9:0] m144_4;
   assign m144_4 =10'b0;

   // m144_5 = W*in
   wire signed [9:0] m144_5;
   assign m144_5 =10'b0;

   // m144_6 = W*in
   wire signed [9:0] m144_6;
   assign m144_6 =10'b0;

   // m144_7 = W*in
   wire signed [9:0] m144_7;
   assign m144_7 =10'b0;

   // m144_8 = W*in
   wire signed [9:0] m144_8;
   assign m144_8 =10'b0;

   // m144_9 = W*in
   wire signed [9:0] m144_9;
   assign m144_9 =10'b0;

   // m144_10 = W*in
   wire signed [9:0] m144_10;
   assign m144_10 =10'b0;

   // m144_11 = W*in
   wire signed [9:0] m144_11;
   assign m144_11 =10'b0;

   // m144_12 = W*in
   wire signed [9:0] m144_12;
   assign m144_12 =10'b0;

   // m144_13 = W*in
   wire signed [9:0] m144_13;
   assign m144_13 =10'b0;

   // m144_14 = W*in
   wire signed [9:0] m144_14;
   assign m144_14 =10'b0;

   // m144_15 = W*in
   wire signed [9:0] m144_15;
   assign m144_15 =10'b0;

   // m144_16 = W*in
   wire signed [9:0] m144_16;
   assign m144_16 =10'b0;

   // m144_17 = W*in
   wire signed [9:0] m144_17;
   assign m144_17 =10'b0;

   // m144_18 = W*in
   wire signed [9:0] m144_18;
   assign m144_18 =10'b0;

   // m144_19 = W*in
   wire signed [9:0] m144_19;
   assign m144_19 ={ {5{in144[5]}} , in144[5:1] };

   // m144_20 = W*in
   wire signed [9:0] m144_20;
   assign m144_20 ={ {5{in144[5]}} , in144[5:1] };

   // m144_21 = W*in
   wire signed [9:0] m144_21;
   assign m144_21 =10'b0;

   // m144_22 = W*in
   wire signed [9:0] m144_22;
   assign m144_22 =10'b0;

   // m144_23 = W*in
   wire signed [9:0] m144_23;
   assign m144_23 =10'b0;

   // m144_24 = W*in
   wire signed [9:0] m144_24;
   assign m144_24 =10'b0;

   // m144_25 = W*in
   wire signed [9:0] m144_25;
   assign m144_25 =10'b0;

   // m144_26 = W*in
   wire signed [9:0] m144_26;
   assign m144_26 ={ {5{neg144[5]}} , neg144[5:1] };

   // m144_27 = W*in
   wire signed [9:0] m144_27;
   assign m144_27 =10'b0;

   // m144_28 = W*in
   wire signed [9:0] m144_28;
   assign m144_28 =10'b0;

   // m144_29 = W*in
   wire signed [9:0] m144_29;
   assign m144_29 =10'b0;

   // m144_30 = W*in
   wire signed [9:0] m144_30;
   assign m144_30 =10'b0;

   // m144_31 = W*in
   wire signed [9:0] m144_31;
   assign m144_31 =10'b0;

   // m144_32 = W*in
   wire signed [9:0] m144_32;
   assign m144_32 =10'b0;

   // m144_33 = W*in
   wire signed [9:0] m144_33;
   assign m144_33 =10'b0;

   // m144_34 = W*in
   wire signed [9:0] m144_34;
   assign m144_34 =10'b0;

   // m144_35 = W*in
   wire signed [9:0] m144_35;
   assign m144_35 =10'b0;

   // m144_36 = W*in
   wire signed [9:0] m144_36;
   assign m144_36 =10'b0;

   // m144_37 = W*in
   wire signed [9:0] m144_37;
   assign m144_37 =10'b0;

   // m144_38 = W*in
   wire signed [9:0] m144_38;
   assign m144_38 =10'b0;

   // m144_39 = W*in
   wire signed [9:0] m144_39;
   assign m144_39 =10'b0;

   // m144_40 = W*in
   wire signed [9:0] m144_40;
   assign m144_40 =10'b0;

   // m144_41 = W*in
   wire signed [9:0] m144_41;
   assign m144_41 =10'b0;

   // m144_42 = W*in
   wire signed [9:0] m144_42;
   assign m144_42 =10'b0;

   // m144_43 = W*in
   wire signed [9:0] m144_43;
   assign m144_43 =10'b0;

   // m144_44 = W*in
   wire signed [9:0] m144_44;
   assign m144_44 =10'b0;

   // m144_45 = W*in
   wire signed [9:0] m144_45;
   assign m144_45 =10'b0;

   // m144_46 = W*in
   wire signed [9:0] m144_46;
   assign m144_46 =10'b0;

   // m144_47 = W*in
   wire signed [9:0] m144_47;
   assign m144_47 =10'b0;

   // m144_48 = W*in
   wire signed [9:0] m144_48;
   assign m144_48 =10'b0;

   // m144_49 = W*in
   wire signed [9:0] m144_49;
   assign m144_49 =10'b0;

   // m144_50 = W*in
   wire signed [9:0] m144_50;
   assign m144_50 =10'b0;

   // m144_51 = W*in
   wire signed [9:0] m144_51;
   assign m144_51 =10'b0;

   // m144_52 = W*in
   wire signed [9:0] m144_52;
   assign m144_52 =10'b0;

   // m144_53 = W*in
   wire signed [9:0] m144_53;
   assign m144_53 =10'b0;

   // m144_54 = W*in
   wire signed [9:0] m144_54;
   assign m144_54 =10'b0;

   // m144_55 = W*in
   wire signed [9:0] m144_55;
   assign m144_55 =10'b0;

   // m144_56 = W*in
   wire signed [9:0] m144_56;
   assign m144_56 =10'b0;

   // m144_57 = W*in
   wire signed [9:0] m144_57;
   assign m144_57 =10'b0;

   // m144_58 = W*in
   wire signed [9:0] m144_58;
   assign m144_58 =10'b0;

   // m144_59 = W*in
   wire signed [9:0] m144_59;
   assign m144_59 =10'b0;

   // m144_60 = W*in
   wire signed [9:0] m144_60;
   assign m144_60 =10'b0;

   // m144_61 = W*in
   wire signed [9:0] m144_61;
   assign m144_61 =10'b0;

   // m144_62 = W*in
   wire signed [9:0] m144_62;
   assign m144_62 =10'b0;

   // m144_63 = W*in
   wire signed [9:0] m144_63;
   assign m144_63 =10'b0;

   // m144_64 = W*in
   wire signed [9:0] m144_64;
   assign m144_64 =10'b0;

   // m144_65 = W*in
   wire signed [9:0] m144_65;
   assign m144_65 =10'b0;

   // m144_66 = W*in
   wire signed [9:0] m144_66;
   assign m144_66 =10'b0;

   // m144_67 = W*in
   wire signed [9:0] m144_67;
   assign m144_67 =10'b0;

   // m144_68 = W*in
   wire signed [9:0] m144_68;
   assign m144_68 =10'b0;

   // m144_69 = W*in
   wire signed [9:0] m144_69;
   assign m144_69 ={ {5{in144[5]}} , in144[5:1] };

   // m144_70 = W*in
   wire signed [9:0] m144_70;
   assign m144_70 =10'b0;

   // m144_71 = W*in
   wire signed [9:0] m144_71;
   assign m144_71 =10'b0;

   // m144_72 = W*in
   wire signed [9:0] m144_72;
   assign m144_72 ={ {5{neg144[5]}} , neg144[5:1] };

   // m144_73 = W*in
   wire signed [9:0] m144_73;
   assign m144_73 =10'b0;

   // m144_74 = W*in
   wire signed [9:0] m144_74;
   assign m144_74 =10'b0;

   // m144_75 = W*in
   wire signed [9:0] m144_75;
   assign m144_75 =10'b0;

   // m144_76 = W*in
   wire signed [9:0] m144_76;
   assign m144_76 =10'b0;

   // m144_77 = W*in
   wire signed [9:0] m144_77;
   assign m144_77 =10'b0;

   // m144_78 = W*in
   wire signed [9:0] m144_78;
   assign m144_78 =10'b0;

   // m144_79 = W*in
   wire signed [9:0] m144_79;
   assign m144_79 =10'b0;

   // m144_80 = W*in
   wire signed [9:0] m144_80;
   assign m144_80 =10'b0;

   // m144_81 = W*in
   wire signed [9:0] m144_81;
   assign m144_81 =10'b0;

   // m144_82 = W*in
   wire signed [9:0] m144_82;
   assign m144_82 =10'b0;

   // m144_83 = W*in
   wire signed [9:0] m144_83;
   assign m144_83 =10'b0;

   // m144_84 = W*in
   wire signed [9:0] m144_84;
   assign m144_84 =10'b0;

   // m144_85 = W*in
   wire signed [9:0] m144_85;
   assign m144_85 =10'b0;

   // m144_86 = W*in
   wire signed [9:0] m144_86;
   assign m144_86 =10'b0;

   // m144_87 = W*in
   wire signed [9:0] m144_87;
   assign m144_87 =10'b0;

   // m144_88 = W*in
   wire signed [9:0] m144_88;
   assign m144_88 =10'b0;

   // m144_89 = W*in
   wire signed [9:0] m144_89;
   assign m144_89 =10'b0;

   // m144_90 = W*in
   wire signed [9:0] m144_90;
   assign m144_90 =10'b0;

   // m144_91 = W*in
   wire signed [9:0] m144_91;
   assign m144_91 =10'b0;

   // m144_92 = W*in
   wire signed [9:0] m144_92;
   assign m144_92 =10'b0;

   // m144_93 = W*in
   wire signed [9:0] m144_93;
   assign m144_93 =10'b0;

   // m144_94 = W*in
   wire signed [9:0] m144_94;
   assign m144_94 =10'b0;

   // m144_95 = W*in
   wire signed [9:0] m144_95;
   assign m144_95 =10'b0;

   // m144_96 = W*in
   wire signed [9:0] m144_96;
   assign m144_96 =10'b0;

   // m144_97 = W*in
   wire signed [9:0] m144_97;
   assign m144_97 =10'b0;

   // m144_98 = W*in
   wire signed [9:0] m144_98;
   assign m144_98 =10'b0;

   // m144_99 = W*in
   wire signed [9:0] m144_99;
   assign m144_99 =10'b0;

   // m144_100 = W*in
   wire signed [9:0] m144_100;
   assign m144_100 =10'b0;

   // m144_101 = W*in
   wire signed [9:0] m144_101;
   assign m144_101 =10'b0;

   // m144_102 = W*in
   wire signed [9:0] m144_102;
   assign m144_102 =10'b0;

   // m144_103 = W*in
   wire signed [9:0] m144_103;
   assign m144_103 =10'b0;

   // m144_104 = W*in
   wire signed [9:0] m144_104;
   assign m144_104 =10'b0;

   // m144_105 = W*in
   wire signed [9:0] m144_105;
   assign m144_105 =10'b0;

   // m144_106 = W*in
   wire signed [9:0] m144_106;
   assign m144_106 =10'b0;

   // m144_107 = W*in
   wire signed [9:0] m144_107;
   assign m144_107 =10'b0;

   // m144_108 = W*in
   wire signed [9:0] m144_108;
   assign m144_108 =10'b0;

   // m144_109 = W*in
   wire signed [9:0] m144_109;
   assign m144_109 =10'b0;

   // m144_110 = W*in
   wire signed [9:0] m144_110;
   assign m144_110 =10'b0;

   // m144_111 = W*in
   wire signed [9:0] m144_111;
   assign m144_111 =10'b0;

   // m144_112 = W*in
   wire signed [9:0] m144_112;
   assign m144_112 =10'b0;

   // m144_113 = W*in
   wire signed [9:0] m144_113;
   assign m144_113 =10'b0;

   // m144_114 = W*in
   wire signed [9:0] m144_114;
   assign m144_114 =10'b0;

   // m144_115 = W*in
   wire signed [9:0] m144_115;
   assign m144_115 =10'b0;

   // m144_116 = W*in
   wire signed [9:0] m144_116;
   assign m144_116 =10'b0;

   // m144_117 = W*in
   wire signed [9:0] m144_117;
   assign m144_117 =10'b0;

   // m145_1 = W*in
   wire signed [9:0] m145_1;
   assign m145_1 =10'b0;

   // m145_2 = W*in
   wire signed [9:0] m145_2;
   assign m145_2 =10'b0;

   // m145_3 = W*in
   wire signed [9:0] m145_3;
   assign m145_3 =10'b0;

   // m145_4 = W*in
   wire signed [9:0] m145_4;
   assign m145_4 =10'b0;

   // m145_5 = W*in
   wire signed [9:0] m145_5;
   assign m145_5 =10'b0;

   // m145_6 = W*in
   wire signed [9:0] m145_6;
   assign m145_6 =10'b0;

   // m145_7 = W*in
   wire signed [9:0] m145_7;
   assign m145_7 =10'b0;

   // m145_8 = W*in
   wire signed [9:0] m145_8;
   assign m145_8 =10'b0;

   // m145_9 = W*in
   wire signed [9:0] m145_9;
   assign m145_9 =10'b0;

   // m145_10 = W*in
   wire signed [9:0] m145_10;
   assign m145_10 =10'b0;

   // m145_11 = W*in
   wire signed [9:0] m145_11;
   assign m145_11 =10'b0;

   // m145_12 = W*in
   wire signed [9:0] m145_12;
   assign m145_12 =10'b0;

   // m145_13 = W*in
   wire signed [9:0] m145_13;
   assign m145_13 =10'b0;

   // m145_14 = W*in
   wire signed [9:0] m145_14;
   assign m145_14 =10'b0;

   // m145_15 = W*in
   wire signed [9:0] m145_15;
   assign m145_15 =10'b0;

   // m145_16 = W*in
   wire signed [9:0] m145_16;
   assign m145_16 =10'b0;

   // m145_17 = W*in
   wire signed [9:0] m145_17;
   assign m145_17 =10'b0;

   // m145_18 = W*in
   wire signed [9:0] m145_18;
   assign m145_18 =10'b0;

   // m145_19 = W*in
   wire signed [9:0] m145_19;
   assign m145_19 ={ {5{in145[5]}} , in145[5:1] };

   // m145_20 = W*in
   wire signed [9:0] m145_20;
   assign m145_20 =10'b0;

   // m145_21 = W*in
   wire signed [9:0] m145_21;
   assign m145_21 =10'b0;

   // m145_22 = W*in
   wire signed [9:0] m145_22;
   assign m145_22 =10'b0;

   // m145_23 = W*in
   wire signed [9:0] m145_23;
   assign m145_23 =10'b0;

   // m145_24 = W*in
   wire signed [9:0] m145_24;
   assign m145_24 =10'b0;

   // m145_25 = W*in
   wire signed [9:0] m145_25;
   assign m145_25 =10'b0;

   // m145_26 = W*in
   wire signed [9:0] m145_26;
   assign m145_26 =10'b0;

   // m145_27 = W*in
   wire signed [9:0] m145_27;
   assign m145_27 =10'b0;

   // m145_28 = W*in
   wire signed [9:0] m145_28;
   assign m145_28 =10'b0;

   // m145_29 = W*in
   wire signed [9:0] m145_29;
   assign m145_29 =10'b0;

   // m145_30 = W*in
   wire signed [9:0] m145_30;
   assign m145_30 =10'b0;

   // m145_31 = W*in
   wire signed [9:0] m145_31;
   assign m145_31 =10'b0;

   // m145_32 = W*in
   wire signed [9:0] m145_32;
   assign m145_32 =10'b0;

   // m145_33 = W*in
   wire signed [9:0] m145_33;
   assign m145_33 =10'b0;

   // m145_34 = W*in
   wire signed [9:0] m145_34;
   assign m145_34 =10'b0;

   // m145_35 = W*in
   wire signed [9:0] m145_35;
   assign m145_35 =10'b0;

   // m145_36 = W*in
   wire signed [9:0] m145_36;
   assign m145_36 =10'b0;

   // m145_37 = W*in
   wire signed [9:0] m145_37;
   assign m145_37 =10'b0;

   // m145_38 = W*in
   wire signed [9:0] m145_38;
   assign m145_38 =10'b0;

   // m145_39 = W*in
   wire signed [9:0] m145_39;
   assign m145_39 =10'b0;

   // m145_40 = W*in
   wire signed [9:0] m145_40;
   assign m145_40 =10'b0;

   // m145_41 = W*in
   wire signed [9:0] m145_41;
   assign m145_41 =10'b0;

   // m145_42 = W*in
   wire signed [9:0] m145_42;
   assign m145_42 =10'b0;

   // m145_43 = W*in
   wire signed [9:0] m145_43;
   assign m145_43 =10'b0;

   // m145_44 = W*in
   wire signed [9:0] m145_44;
   assign m145_44 =10'b0;

   // m145_45 = W*in
   wire signed [9:0] m145_45;
   assign m145_45 =10'b0;

   // m145_46 = W*in
   wire signed [9:0] m145_46;
   assign m145_46 =10'b0;

   // m145_47 = W*in
   wire signed [9:0] m145_47;
   assign m145_47 =10'b0;

   // m145_48 = W*in
   wire signed [9:0] m145_48;
   assign m145_48 =10'b0;

   // m145_49 = W*in
   wire signed [9:0] m145_49;
   assign m145_49 =10'b0;

   // m145_50 = W*in
   wire signed [9:0] m145_50;
   assign m145_50 =10'b0;

   // m145_51 = W*in
   wire signed [9:0] m145_51;
   assign m145_51 =10'b0;

   // m145_52 = W*in
   wire signed [9:0] m145_52;
   assign m145_52 =10'b0;

   // m145_53 = W*in
   wire signed [9:0] m145_53;
   assign m145_53 =10'b0;

   // m145_54 = W*in
   wire signed [9:0] m145_54;
   assign m145_54 =10'b0;

   // m145_55 = W*in
   wire signed [9:0] m145_55;
   assign m145_55 =10'b0;

   // m145_56 = W*in
   wire signed [9:0] m145_56;
   assign m145_56 =10'b0;

   // m145_57 = W*in
   wire signed [9:0] m145_57;
   assign m145_57 =10'b0;

   // m145_58 = W*in
   wire signed [9:0] m145_58;
   assign m145_58 =10'b0;

   // m145_59 = W*in
   wire signed [9:0] m145_59;
   assign m145_59 =10'b0;

   // m145_60 = W*in
   wire signed [9:0] m145_60;
   assign m145_60 =10'b0;

   // m145_61 = W*in
   wire signed [9:0] m145_61;
   assign m145_61 =10'b0;

   // m145_62 = W*in
   wire signed [9:0] m145_62;
   assign m145_62 =10'b0;

   // m145_63 = W*in
   wire signed [9:0] m145_63;
   assign m145_63 =10'b0;

   // m145_64 = W*in
   wire signed [9:0] m145_64;
   assign m145_64 =10'b0;

   // m145_65 = W*in
   wire signed [9:0] m145_65;
   assign m145_65 =10'b0;

   // m145_66 = W*in
   wire signed [9:0] m145_66;
   assign m145_66 =10'b0;

   // m145_67 = W*in
   wire signed [9:0] m145_67;
   assign m145_67 =10'b0;

   // m145_68 = W*in
   wire signed [9:0] m145_68;
   assign m145_68 =10'b0;

   // m145_69 = W*in
   wire signed [9:0] m145_69;
   assign m145_69 =10'b0;

   // m145_70 = W*in
   wire signed [9:0] m145_70;
   assign m145_70 =10'b0;

   // m145_71 = W*in
   wire signed [9:0] m145_71;
   assign m145_71 =10'b0;

   // m145_72 = W*in
   wire signed [9:0] m145_72;
   assign m145_72 =10'b0;

   // m145_73 = W*in
   wire signed [9:0] m145_73;
   assign m145_73 =10'b0;

   // m145_74 = W*in
   wire signed [9:0] m145_74;
   assign m145_74 =10'b0;

   // m145_75 = W*in
   wire signed [9:0] m145_75;
   assign m145_75 =10'b0;

   // m145_76 = W*in
   wire signed [9:0] m145_76;
   assign m145_76 =10'b0;

   // m145_77 = W*in
   wire signed [9:0] m145_77;
   assign m145_77 =10'b0;

   // m145_78 = W*in
   wire signed [9:0] m145_78;
   assign m145_78 =10'b0;

   // m145_79 = W*in
   wire signed [9:0] m145_79;
   assign m145_79 =10'b0;

   // m145_80 = W*in
   wire signed [9:0] m145_80;
   assign m145_80 =10'b0;

   // m145_81 = W*in
   wire signed [9:0] m145_81;
   assign m145_81 =10'b0;

   // m145_82 = W*in
   wire signed [9:0] m145_82;
   assign m145_82 =10'b0;

   // m145_83 = W*in
   wire signed [9:0] m145_83;
   assign m145_83 =10'b0;

   // m145_84 = W*in
   wire signed [9:0] m145_84;
   assign m145_84 =10'b0;

   // m145_85 = W*in
   wire signed [9:0] m145_85;
   assign m145_85 =10'b0;

   // m145_86 = W*in
   wire signed [9:0] m145_86;
   assign m145_86 =10'b0;

   // m145_87 = W*in
   wire signed [9:0] m145_87;
   assign m145_87 =10'b0;

   // m145_88 = W*in
   wire signed [9:0] m145_88;
   assign m145_88 =10'b0;

   // m145_89 = W*in
   wire signed [9:0] m145_89;
   assign m145_89 =10'b0;

   // m145_90 = W*in
   wire signed [9:0] m145_90;
   assign m145_90 =10'b0;

   // m145_91 = W*in
   wire signed [9:0] m145_91;
   assign m145_91 =10'b0;

   // m145_92 = W*in
   wire signed [9:0] m145_92;
   assign m145_92 =10'b0;

   // m145_93 = W*in
   wire signed [9:0] m145_93;
   assign m145_93 =10'b0;

   // m145_94 = W*in
   wire signed [9:0] m145_94;
   assign m145_94 =10'b0;

   // m145_95 = W*in
   wire signed [9:0] m145_95;
   assign m145_95 =10'b0;

   // m145_96 = W*in
   wire signed [9:0] m145_96;
   assign m145_96 =10'b0;

   // m145_97 = W*in
   wire signed [9:0] m145_97;
   assign m145_97 =10'b0;

   // m145_98 = W*in
   wire signed [9:0] m145_98;
   assign m145_98 =10'b0;

   // m145_99 = W*in
   wire signed [9:0] m145_99;
   assign m145_99 =10'b0;

   // m145_100 = W*in
   wire signed [9:0] m145_100;
   assign m145_100 =10'b0;

   // m145_101 = W*in
   wire signed [9:0] m145_101;
   assign m145_101 =10'b0;

   // m145_102 = W*in
   wire signed [9:0] m145_102;
   assign m145_102 =10'b0;

   // m145_103 = W*in
   wire signed [9:0] m145_103;
   assign m145_103 =10'b0;

   // m145_104 = W*in
   wire signed [9:0] m145_104;
   assign m145_104 =10'b0;

   // m145_105 = W*in
   wire signed [9:0] m145_105;
   assign m145_105 =10'b0;

   // m145_106 = W*in
   wire signed [9:0] m145_106;
   assign m145_106 =10'b0;

   // m145_107 = W*in
   wire signed [9:0] m145_107;
   assign m145_107 =10'b0;

   // m145_108 = W*in
   wire signed [9:0] m145_108;
   assign m145_108 =10'b0;

   // m145_109 = W*in
   wire signed [9:0] m145_109;
   assign m145_109 =10'b0;

   // m145_110 = W*in
   wire signed [9:0] m145_110;
   assign m145_110 =10'b0;

   // m145_111 = W*in
   wire signed [9:0] m145_111;
   assign m145_111 =10'b0;

   // m145_112 = W*in
   wire signed [9:0] m145_112;
   assign m145_112 =10'b0;

   // m145_113 = W*in
   wire signed [9:0] m145_113;
   assign m145_113 =10'b0;

   // m145_114 = W*in
   wire signed [9:0] m145_114;
   assign m145_114 =10'b0;

   // m145_115 = W*in
   wire signed [9:0] m145_115;
   assign m145_115 =10'b0;

   // m145_116 = W*in
   wire signed [9:0] m145_116;
   assign m145_116 =10'b0;

   // m145_117 = W*in
   wire signed [9:0] m145_117;
   assign m145_117 =10'b0;

   // m146_1 = W*in
   wire signed [9:0] m146_1;
   assign m146_1 =10'b0;

   // m146_2 = W*in
   wire signed [9:0] m146_2;
   assign m146_2 =10'b0;

   // m146_3 = W*in
   wire signed [9:0] m146_3;
   assign m146_3 =10'b0;

   // m146_4 = W*in
   wire signed [9:0] m146_4;
   assign m146_4 =10'b0;

   // m146_5 = W*in
   wire signed [9:0] m146_5;
   assign m146_5 =10'b0;

   // m146_6 = W*in
   wire signed [9:0] m146_6;
   assign m146_6 =10'b0;

   // m146_7 = W*in
   wire signed [9:0] m146_7;
   assign m146_7 =10'b0;

   // m146_8 = W*in
   wire signed [9:0] m146_8;
   assign m146_8 =10'b0;

   // m146_9 = W*in
   wire signed [9:0] m146_9;
   assign m146_9 =10'b0;

   // m146_10 = W*in
   wire signed [9:0] m146_10;
   assign m146_10 =10'b0;

   // m146_11 = W*in
   wire signed [9:0] m146_11;
   assign m146_11 =10'b0;

   // m146_12 = W*in
   wire signed [9:0] m146_12;
   assign m146_12 =10'b0;

   // m146_13 = W*in
   wire signed [9:0] m146_13;
   assign m146_13 =10'b0;

   // m146_14 = W*in
   wire signed [9:0] m146_14;
   assign m146_14 =10'b0;

   // m146_15 = W*in
   wire signed [9:0] m146_15;
   assign m146_15 =10'b0;

   // m146_16 = W*in
   wire signed [9:0] m146_16;
   assign m146_16 =10'b0;

   // m146_17 = W*in
   wire signed [9:0] m146_17;
   assign m146_17 =10'b0;

   // m146_18 = W*in
   wire signed [9:0] m146_18;
   assign m146_18 =10'b0;

   // m146_19 = W*in
   wire signed [9:0] m146_19;
   assign m146_19 =10'b0;

   // m146_20 = W*in
   wire signed [9:0] m146_20;
   assign m146_20 =10'b0;

   // m146_21 = W*in
   wire signed [9:0] m146_21;
   assign m146_21 =10'b0;

   // m146_22 = W*in
   wire signed [9:0] m146_22;
   assign m146_22 =10'b0;

   // m146_23 = W*in
   wire signed [9:0] m146_23;
   assign m146_23 =10'b0;

   // m146_24 = W*in
   wire signed [9:0] m146_24;
   assign m146_24 =10'b0;

   // m146_25 = W*in
   wire signed [9:0] m146_25;
   assign m146_25 =10'b0;

   // m146_26 = W*in
   wire signed [9:0] m146_26;
   assign m146_26 =10'b0;

   // m146_27 = W*in
   wire signed [9:0] m146_27;
   assign m146_27 =10'b0;

   // m146_28 = W*in
   wire signed [9:0] m146_28;
   assign m146_28 =10'b0;

   // m146_29 = W*in
   wire signed [9:0] m146_29;
   assign m146_29 =10'b0;

   // m146_30 = W*in
   wire signed [9:0] m146_30;
   assign m146_30 =10'b0;

   // m146_31 = W*in
   wire signed [9:0] m146_31;
   assign m146_31 =10'b0;

   // m146_32 = W*in
   wire signed [9:0] m146_32;
   assign m146_32 =10'b0;

   // m146_33 = W*in
   wire signed [9:0] m146_33;
   assign m146_33 =10'b0;

   // m146_34 = W*in
   wire signed [9:0] m146_34;
   assign m146_34 =10'b0;

   // m146_35 = W*in
   wire signed [9:0] m146_35;
   assign m146_35 =10'b0;

   // m146_36 = W*in
   wire signed [9:0] m146_36;
   assign m146_36 =10'b0;

   // m146_37 = W*in
   wire signed [9:0] m146_37;
   assign m146_37 =10'b0;

   // m146_38 = W*in
   wire signed [9:0] m146_38;
   assign m146_38 =10'b0;

   // m146_39 = W*in
   wire signed [9:0] m146_39;
   assign m146_39 =10'b0;

   // m146_40 = W*in
   wire signed [9:0] m146_40;
   assign m146_40 =10'b0;

   // m146_41 = W*in
   wire signed [9:0] m146_41;
   assign m146_41 =10'b0;

   // m146_42 = W*in
   wire signed [9:0] m146_42;
   assign m146_42 =10'b0;

   // m146_43 = W*in
   wire signed [9:0] m146_43;
   assign m146_43 =10'b0;

   // m146_44 = W*in
   wire signed [9:0] m146_44;
   assign m146_44 =10'b0;

   // m146_45 = W*in
   wire signed [9:0] m146_45;
   assign m146_45 =10'b0;

   // m146_46 = W*in
   wire signed [9:0] m146_46;
   assign m146_46 =10'b0;

   // m146_47 = W*in
   wire signed [9:0] m146_47;
   assign m146_47 =10'b0;

   // m146_48 = W*in
   wire signed [9:0] m146_48;
   assign m146_48 =10'b0;

   // m146_49 = W*in
   wire signed [9:0] m146_49;
   assign m146_49 =10'b0;

   // m146_50 = W*in
   wire signed [9:0] m146_50;
   assign m146_50 =10'b0;

   // m146_51 = W*in
   wire signed [9:0] m146_51;
   assign m146_51 =10'b0;

   // m146_52 = W*in
   wire signed [9:0] m146_52;
   assign m146_52 =10'b0;

   // m146_53 = W*in
   wire signed [9:0] m146_53;
   assign m146_53 =10'b0;

   // m146_54 = W*in
   wire signed [9:0] m146_54;
   assign m146_54 =10'b0;

   // m146_55 = W*in
   wire signed [9:0] m146_55;
   assign m146_55 =10'b0;

   // m146_56 = W*in
   wire signed [9:0] m146_56;
   assign m146_56 =10'b0;

   // m146_57 = W*in
   wire signed [9:0] m146_57;
   assign m146_57 =10'b0;

   // m146_58 = W*in
   wire signed [9:0] m146_58;
   assign m146_58 =10'b0;

   // m146_59 = W*in
   wire signed [9:0] m146_59;
   assign m146_59 =10'b0;

   // m146_60 = W*in
   wire signed [9:0] m146_60;
   assign m146_60 =10'b0;

   // m146_61 = W*in
   wire signed [9:0] m146_61;
   assign m146_61 =10'b0;

   // m146_62 = W*in
   wire signed [9:0] m146_62;
   assign m146_62 =10'b0;

   // m146_63 = W*in
   wire signed [9:0] m146_63;
   assign m146_63 =10'b0;

   // m146_64 = W*in
   wire signed [9:0] m146_64;
   assign m146_64 =10'b0;

   // m146_65 = W*in
   wire signed [9:0] m146_65;
   assign m146_65 =10'b0;

   // m146_66 = W*in
   wire signed [9:0] m146_66;
   assign m146_66 =10'b0;

   // m146_67 = W*in
   wire signed [9:0] m146_67;
   assign m146_67 =10'b0;

   // m146_68 = W*in
   wire signed [9:0] m146_68;
   assign m146_68 =10'b0;

   // m146_69 = W*in
   wire signed [9:0] m146_69;
   assign m146_69 =10'b0;

   // m146_70 = W*in
   wire signed [9:0] m146_70;
   assign m146_70 =10'b0;

   // m146_71 = W*in
   wire signed [9:0] m146_71;
   assign m146_71 =10'b0;

   // m146_72 = W*in
   wire signed [9:0] m146_72;
   assign m146_72 =10'b0;

   // m146_73 = W*in
   wire signed [9:0] m146_73;
   assign m146_73 =10'b0;

   // m146_74 = W*in
   wire signed [9:0] m146_74;
   assign m146_74 =10'b0;

   // m146_75 = W*in
   wire signed [9:0] m146_75;
   assign m146_75 =10'b0;

   // m146_76 = W*in
   wire signed [9:0] m146_76;
   assign m146_76 =10'b0;

   // m146_77 = W*in
   wire signed [9:0] m146_77;
   assign m146_77 =10'b0;

   // m146_78 = W*in
   wire signed [9:0] m146_78;
   assign m146_78 =10'b0;

   // m146_79 = W*in
   wire signed [9:0] m146_79;
   assign m146_79 =10'b0;

   // m146_80 = W*in
   wire signed [9:0] m146_80;
   assign m146_80 =10'b0;

   // m146_81 = W*in
   wire signed [9:0] m146_81;
   assign m146_81 =10'b0;

   // m146_82 = W*in
   wire signed [9:0] m146_82;
   assign m146_82 =10'b0;

   // m146_83 = W*in
   wire signed [9:0] m146_83;
   assign m146_83 =10'b0;

   // m146_84 = W*in
   wire signed [9:0] m146_84;
   assign m146_84 =10'b0;

   // m146_85 = W*in
   wire signed [9:0] m146_85;
   assign m146_85 =10'b0;

   // m146_86 = W*in
   wire signed [9:0] m146_86;
   assign m146_86 =10'b0;

   // m146_87 = W*in
   wire signed [9:0] m146_87;
   assign m146_87 =10'b0;

   // m146_88 = W*in
   wire signed [9:0] m146_88;
   assign m146_88 =10'b0;

   // m146_89 = W*in
   wire signed [9:0] m146_89;
   assign m146_89 =10'b0;

   // m146_90 = W*in
   wire signed [9:0] m146_90;
   assign m146_90 =10'b0;

   // m146_91 = W*in
   wire signed [9:0] m146_91;
   assign m146_91 =10'b0;

   // m146_92 = W*in
   wire signed [9:0] m146_92;
   assign m146_92 =10'b0;

   // m146_93 = W*in
   wire signed [9:0] m146_93;
   assign m146_93 =10'b0;

   // m146_94 = W*in
   wire signed [9:0] m146_94;
   assign m146_94 =10'b0;

   // m146_95 = W*in
   wire signed [9:0] m146_95;
   assign m146_95 =10'b0;

   // m146_96 = W*in
   wire signed [9:0] m146_96;
   assign m146_96 =10'b0;

   // m146_97 = W*in
   wire signed [9:0] m146_97;
   assign m146_97 =10'b0;

   // m146_98 = W*in
   wire signed [9:0] m146_98;
   assign m146_98 =10'b0;

   // m146_99 = W*in
   wire signed [9:0] m146_99;
   assign m146_99 =10'b0;

   // m146_100 = W*in
   wire signed [9:0] m146_100;
   assign m146_100 =10'b0;

   // m146_101 = W*in
   wire signed [9:0] m146_101;
   assign m146_101 =10'b0;

   // m146_102 = W*in
   wire signed [9:0] m146_102;
   assign m146_102 =10'b0;

   // m146_103 = W*in
   wire signed [9:0] m146_103;
   assign m146_103 =10'b0;

   // m146_104 = W*in
   wire signed [9:0] m146_104;
   assign m146_104 =10'b0;

   // m146_105 = W*in
   wire signed [9:0] m146_105;
   assign m146_105 =10'b0;

   // m146_106 = W*in
   wire signed [9:0] m146_106;
   assign m146_106 =10'b0;

   // m146_107 = W*in
   wire signed [9:0] m146_107;
   assign m146_107 =10'b0;

   // m146_108 = W*in
   wire signed [9:0] m146_108;
   assign m146_108 =10'b0;

   // m146_109 = W*in
   wire signed [9:0] m146_109;
   assign m146_109 ={ {5{neg146[5]}} , neg146[5:1] };

   // m146_110 = W*in
   wire signed [9:0] m146_110;
   assign m146_110 =10'b0;

   // m146_111 = W*in
   wire signed [9:0] m146_111;
   assign m146_111 =10'b0;

   // m146_112 = W*in
   wire signed [9:0] m146_112;
   assign m146_112 =10'b0;

   // m146_113 = W*in
   wire signed [9:0] m146_113;
   assign m146_113 =10'b0;

   // m146_114 = W*in
   wire signed [9:0] m146_114;
   assign m146_114 =10'b0;

   // m146_115 = W*in
   wire signed [9:0] m146_115;
   assign m146_115 =10'b0;

   // m146_116 = W*in
   wire signed [9:0] m146_116;
   assign m146_116 =10'b0;

   // m146_117 = W*in
   wire signed [9:0] m146_117;
   assign m146_117 =10'b0;

   // m147_1 = W*in
   wire signed [9:0] m147_1;
   assign m147_1 =10'b0;

   // m147_2 = W*in
   wire signed [9:0] m147_2;
   assign m147_2 =10'b0;

   // m147_3 = W*in
   wire signed [9:0] m147_3;
   assign m147_3 =10'b0;

   // m147_4 = W*in
   wire signed [9:0] m147_4;
   assign m147_4 =10'b0;

   // m147_5 = W*in
   wire signed [9:0] m147_5;
   assign m147_5 =10'b0;

   // m147_6 = W*in
   wire signed [9:0] m147_6;
   assign m147_6 =10'b0;

   // m147_7 = W*in
   wire signed [9:0] m147_7;
   assign m147_7 =10'b0;

   // m147_8 = W*in
   wire signed [9:0] m147_8;
   assign m147_8 =10'b0;

   // m147_9 = W*in
   wire signed [9:0] m147_9;
   assign m147_9 =10'b0;

   // m147_10 = W*in
   wire signed [9:0] m147_10;
   assign m147_10 =10'b0;

   // m147_11 = W*in
   wire signed [9:0] m147_11;
   assign m147_11 =10'b0;

   // m147_12 = W*in
   wire signed [9:0] m147_12;
   assign m147_12 =10'b0;

   // m147_13 = W*in
   wire signed [9:0] m147_13;
   assign m147_13 =10'b0;

   // m147_14 = W*in
   wire signed [9:0] m147_14;
   assign m147_14 =10'b0;

   // m147_15 = W*in
   wire signed [9:0] m147_15;
   assign m147_15 =10'b0;

   // m147_16 = W*in
   wire signed [9:0] m147_16;
   assign m147_16 =10'b0;

   // m147_17 = W*in
   wire signed [9:0] m147_17;
   assign m147_17 =10'b0;

   // m147_18 = W*in
   wire signed [9:0] m147_18;
   assign m147_18 =10'b0;

   // m147_19 = W*in
   wire signed [9:0] m147_19;
   assign m147_19 =10'b0;

   // m147_20 = W*in
   wire signed [9:0] m147_20;
   assign m147_20 ={ {5{neg147[5]}} , neg147[5:1] };

   // m147_21 = W*in
   wire signed [9:0] m147_21;
   assign m147_21 =10'b0;

   // m147_22 = W*in
   wire signed [9:0] m147_22;
   assign m147_22 =10'b0;

   // m147_23 = W*in
   wire signed [9:0] m147_23;
   assign m147_23 =10'b0;

   // m147_24 = W*in
   wire signed [9:0] m147_24;
   assign m147_24 =10'b0;

   // m147_25 = W*in
   wire signed [9:0] m147_25;
   assign m147_25 =10'b0;

   // m147_26 = W*in
   wire signed [9:0] m147_26;
   assign m147_26 =10'b0;

   // m147_27 = W*in
   wire signed [9:0] m147_27;
   assign m147_27 ={ {5{neg147[5]}} , neg147[5:1] };

   // m147_28 = W*in
   wire signed [9:0] m147_28;
   assign m147_28 =10'b0;

   // m147_29 = W*in
   wire signed [9:0] m147_29;
   assign m147_29 =10'b0;

   // m147_30 = W*in
   wire signed [9:0] m147_30;
   assign m147_30 ={ {5{neg147[5]}} , neg147[5:1] };

   // m147_31 = W*in
   wire signed [9:0] m147_31;
   assign m147_31 =10'b0;

   // m147_32 = W*in
   wire signed [9:0] m147_32;
   assign m147_32 =10'b0;

   // m147_33 = W*in
   wire signed [9:0] m147_33;
   assign m147_33 =10'b0;

   // m147_34 = W*in
   wire signed [9:0] m147_34;
   assign m147_34 =10'b0;

   // m147_35 = W*in
   wire signed [9:0] m147_35;
   assign m147_35 =10'b0;

   // m147_36 = W*in
   wire signed [9:0] m147_36;
   assign m147_36 =10'b0;

   // m147_37 = W*in
   wire signed [9:0] m147_37;
   assign m147_37 =10'b0;

   // m147_38 = W*in
   wire signed [9:0] m147_38;
   assign m147_38 =10'b0;

   // m147_39 = W*in
   wire signed [9:0] m147_39;
   assign m147_39 =10'b0;

   // m147_40 = W*in
   wire signed [9:0] m147_40;
   assign m147_40 =10'b0;

   // m147_41 = W*in
   wire signed [9:0] m147_41;
   assign m147_41 =10'b0;

   // m147_42 = W*in
   wire signed [9:0] m147_42;
   assign m147_42 =10'b0;

   // m147_43 = W*in
   wire signed [9:0] m147_43;
   assign m147_43 =10'b0;

   // m147_44 = W*in
   wire signed [9:0] m147_44;
   assign m147_44 =10'b0;

   // m147_45 = W*in
   wire signed [9:0] m147_45;
   assign m147_45 =10'b0;

   // m147_46 = W*in
   wire signed [9:0] m147_46;
   assign m147_46 =10'b0;

   // m147_47 = W*in
   wire signed [9:0] m147_47;
   assign m147_47 =10'b0;

   // m147_48 = W*in
   wire signed [9:0] m147_48;
   assign m147_48 =10'b0;

   // m147_49 = W*in
   wire signed [9:0] m147_49;
   assign m147_49 =10'b0;

   // m147_50 = W*in
   wire signed [9:0] m147_50;
   assign m147_50 =10'b0;

   // m147_51 = W*in
   wire signed [9:0] m147_51;
   assign m147_51 =10'b0;

   // m147_52 = W*in
   wire signed [9:0] m147_52;
   assign m147_52 =10'b0;

   // m147_53 = W*in
   wire signed [9:0] m147_53;
   assign m147_53 =10'b0;

   // m147_54 = W*in
   wire signed [9:0] m147_54;
   assign m147_54 =10'b0;

   // m147_55 = W*in
   wire signed [9:0] m147_55;
   assign m147_55 =10'b0;

   // m147_56 = W*in
   wire signed [9:0] m147_56;
   assign m147_56 =10'b0;

   // m147_57 = W*in
   wire signed [9:0] m147_57;
   assign m147_57 =10'b0;

   // m147_58 = W*in
   wire signed [9:0] m147_58;
   assign m147_58 =10'b0;

   // m147_59 = W*in
   wire signed [9:0] m147_59;
   assign m147_59 =10'b0;

   // m147_60 = W*in
   wire signed [9:0] m147_60;
   assign m147_60 =10'b0;

   // m147_61 = W*in
   wire signed [9:0] m147_61;
   assign m147_61 =10'b0;

   // m147_62 = W*in
   wire signed [9:0] m147_62;
   assign m147_62 =10'b0;

   // m147_63 = W*in
   wire signed [9:0] m147_63;
   assign m147_63 =10'b0;

   // m147_64 = W*in
   wire signed [9:0] m147_64;
   assign m147_64 =10'b0;

   // m147_65 = W*in
   wire signed [9:0] m147_65;
   assign m147_65 =10'b0;

   // m147_66 = W*in
   wire signed [9:0] m147_66;
   assign m147_66 =10'b0;

   // m147_67 = W*in
   wire signed [9:0] m147_67;
   assign m147_67 =10'b0;

   // m147_68 = W*in
   wire signed [9:0] m147_68;
   assign m147_68 =10'b0;

   // m147_69 = W*in
   wire signed [9:0] m147_69;
   assign m147_69 =10'b0;

   // m147_70 = W*in
   wire signed [9:0] m147_70;
   assign m147_70 =10'b0;

   // m147_71 = W*in
   wire signed [9:0] m147_71;
   assign m147_71 =10'b0;

   // m147_72 = W*in
   wire signed [9:0] m147_72;
   assign m147_72 =10'b0;

   // m147_73 = W*in
   wire signed [9:0] m147_73;
   assign m147_73 =10'b0;

   // m147_74 = W*in
   wire signed [9:0] m147_74;
   assign m147_74 =10'b0;

   // m147_75 = W*in
   wire signed [9:0] m147_75;
   assign m147_75 =10'b0;

   // m147_76 = W*in
   wire signed [9:0] m147_76;
   assign m147_76 =10'b0;

   // m147_77 = W*in
   wire signed [9:0] m147_77;
   assign m147_77 =10'b0;

   // m147_78 = W*in
   wire signed [9:0] m147_78;
   assign m147_78 =10'b0;

   // m147_79 = W*in
   wire signed [9:0] m147_79;
   assign m147_79 =10'b0;

   // m147_80 = W*in
   wire signed [9:0] m147_80;
   assign m147_80 =10'b0;

   // m147_81 = W*in
   wire signed [9:0] m147_81;
   assign m147_81 =10'b0;

   // m147_82 = W*in
   wire signed [9:0] m147_82;
   assign m147_82 =10'b0;

   // m147_83 = W*in
   wire signed [9:0] m147_83;
   assign m147_83 =10'b0;

   // m147_84 = W*in
   wire signed [9:0] m147_84;
   assign m147_84 =10'b0;

   // m147_85 = W*in
   wire signed [9:0] m147_85;
   assign m147_85 =10'b0;

   // m147_86 = W*in
   wire signed [9:0] m147_86;
   assign m147_86 =10'b0;

   // m147_87 = W*in
   wire signed [9:0] m147_87;
   assign m147_87 =10'b0;

   // m147_88 = W*in
   wire signed [9:0] m147_88;
   assign m147_88 =10'b0;

   // m147_89 = W*in
   wire signed [9:0] m147_89;
   assign m147_89 =10'b0;

   // m147_90 = W*in
   wire signed [9:0] m147_90;
   assign m147_90 =10'b0;

   // m147_91 = W*in
   wire signed [9:0] m147_91;
   assign m147_91 =10'b0;

   // m147_92 = W*in
   wire signed [9:0] m147_92;
   assign m147_92 =10'b0;

   // m147_93 = W*in
   wire signed [9:0] m147_93;
   assign m147_93 =10'b0;

   // m147_94 = W*in
   wire signed [9:0] m147_94;
   assign m147_94 =10'b0;

   // m147_95 = W*in
   wire signed [9:0] m147_95;
   assign m147_95 =10'b0;

   // m147_96 = W*in
   wire signed [9:0] m147_96;
   assign m147_96 =10'b0;

   // m147_97 = W*in
   wire signed [9:0] m147_97;
   assign m147_97 =10'b0;

   // m147_98 = W*in
   wire signed [9:0] m147_98;
   assign m147_98 =10'b0;

   // m147_99 = W*in
   wire signed [9:0] m147_99;
   assign m147_99 =10'b0;

   // m147_100 = W*in
   wire signed [9:0] m147_100;
   assign m147_100 =10'b0;

   // m147_101 = W*in
   wire signed [9:0] m147_101;
   assign m147_101 =10'b0;

   // m147_102 = W*in
   wire signed [9:0] m147_102;
   assign m147_102 =10'b0;

   // m147_103 = W*in
   wire signed [9:0] m147_103;
   assign m147_103 =10'b0;

   // m147_104 = W*in
   wire signed [9:0] m147_104;
   assign m147_104 =10'b0;

   // m147_105 = W*in
   wire signed [9:0] m147_105;
   assign m147_105 =10'b0;

   // m147_106 = W*in
   wire signed [9:0] m147_106;
   assign m147_106 =10'b0;

   // m147_107 = W*in
   wire signed [9:0] m147_107;
   assign m147_107 =10'b0;

   // m147_108 = W*in
   wire signed [9:0] m147_108;
   assign m147_108 =10'b0;

   // m147_109 = W*in
   wire signed [9:0] m147_109;
   assign m147_109 ={ {5{neg147[5]}} , neg147[5:1] };

   // m147_110 = W*in
   wire signed [9:0] m147_110;
   assign m147_110 =10'b0;

   // m147_111 = W*in
   wire signed [9:0] m147_111;
   assign m147_111 =10'b0;

   // m147_112 = W*in
   wire signed [9:0] m147_112;
   assign m147_112 =10'b0;

   // m147_113 = W*in
   wire signed [9:0] m147_113;
   assign m147_113 =10'b0;

   // m147_114 = W*in
   wire signed [9:0] m147_114;
   assign m147_114 =10'b0;

   // m147_115 = W*in
   wire signed [9:0] m147_115;
   assign m147_115 =10'b0;

   // m147_116 = W*in
   wire signed [9:0] m147_116;
   assign m147_116 =10'b0;

   // m147_117 = W*in
   wire signed [9:0] m147_117;
   assign m147_117 =10'b0;

   // m148_1 = W*in
   wire signed [9:0] m148_1;
   assign m148_1 =10'b0;

   // m148_2 = W*in
   wire signed [9:0] m148_2;
   assign m148_2 =10'b0;

   // m148_3 = W*in
   wire signed [9:0] m148_3;
   assign m148_3 =10'b0;

   // m148_4 = W*in
   wire signed [9:0] m148_4;
   assign m148_4 =10'b0;

   // m148_5 = W*in
   wire signed [9:0] m148_5;
   assign m148_5 =10'b0;

   // m148_6 = W*in
   wire signed [9:0] m148_6;
   assign m148_6 =10'b0;

   // m148_7 = W*in
   wire signed [9:0] m148_7;
   assign m148_7 =10'b0;

   // m148_8 = W*in
   wire signed [9:0] m148_8;
   assign m148_8 =10'b0;

   // m148_9 = W*in
   wire signed [9:0] m148_9;
   assign m148_9 =10'b0;

   // m148_10 = W*in
   wire signed [9:0] m148_10;
   assign m148_10 =10'b0;

   // m148_11 = W*in
   wire signed [9:0] m148_11;
   assign m148_11 =10'b0;

   // m148_12 = W*in
   wire signed [9:0] m148_12;
   assign m148_12 =10'b0;

   // m148_13 = W*in
   wire signed [9:0] m148_13;
   assign m148_13 =10'b0;

   // m148_14 = W*in
   wire signed [9:0] m148_14;
   assign m148_14 =10'b0;

   // m148_15 = W*in
   wire signed [9:0] m148_15;
   assign m148_15 =10'b0;

   // m148_16 = W*in
   wire signed [9:0] m148_16;
   assign m148_16 =10'b0;

   // m148_17 = W*in
   wire signed [9:0] m148_17;
   assign m148_17 ={ {5{in148[5]}} , in148[5:1] };

   // m148_18 = W*in
   wire signed [9:0] m148_18;
   assign m148_18 =10'b0;

   // m148_19 = W*in
   wire signed [9:0] m148_19;
   assign m148_19 =10'b0;

   // m148_20 = W*in
   wire signed [9:0] m148_20;
   assign m148_20 ={ {4{neg148[5]}} , neg148[5:0] };

   // m148_21 = W*in
   wire signed [9:0] m148_21;
   assign m148_21 ={ {5{in148[5]}} , in148[5:1] };

   // m148_22 = W*in
   wire signed [9:0] m148_22;
   assign m148_22 =10'b0;

   // m148_23 = W*in
   wire signed [9:0] m148_23;
   assign m148_23 =10'b0;

   // m148_24 = W*in
   wire signed [9:0] m148_24;
   assign m148_24 =10'b0;

   // m148_25 = W*in
   wire signed [9:0] m148_25;
   assign m148_25 =10'b0;

   // m148_26 = W*in
   wire signed [9:0] m148_26;
   assign m148_26 =10'b0;

   // m148_27 = W*in
   wire signed [9:0] m148_27;
   assign m148_27 =10'b0;

   // m148_28 = W*in
   wire signed [9:0] m148_28;
   assign m148_28 =10'b0;

   // m148_29 = W*in
   wire signed [9:0] m148_29;
   assign m148_29 =10'b0;

   // m148_30 = W*in
   wire signed [9:0] m148_30;
   assign m148_30 ={ {5{neg148[5]}} , neg148[5:1] };

   // m148_31 = W*in
   wire signed [9:0] m148_31;
   assign m148_31 =10'b0;

   // m148_32 = W*in
   wire signed [9:0] m148_32;
   assign m148_32 =10'b0;

   // m148_33 = W*in
   wire signed [9:0] m148_33;
   assign m148_33 =10'b0;

   // m148_34 = W*in
   wire signed [9:0] m148_34;
   assign m148_34 =10'b0;

   // m148_35 = W*in
   wire signed [9:0] m148_35;
   assign m148_35 ={ {5{neg148[5]}} , neg148[5:1] };

   // m148_36 = W*in
   wire signed [9:0] m148_36;
   assign m148_36 =10'b0;

   // m148_37 = W*in
   wire signed [9:0] m148_37;
   assign m148_37 =10'b0;

   // m148_38 = W*in
   wire signed [9:0] m148_38;
   assign m148_38 =10'b0;

   // m148_39 = W*in
   wire signed [9:0] m148_39;
   assign m148_39 =10'b0;

   // m148_40 = W*in
   wire signed [9:0] m148_40;
   assign m148_40 =10'b0;

   // m148_41 = W*in
   wire signed [9:0] m148_41;
   assign m148_41 =10'b0;

   // m148_42 = W*in
   wire signed [9:0] m148_42;
   assign m148_42 =10'b0;

   // m148_43 = W*in
   wire signed [9:0] m148_43;
   assign m148_43 =10'b0;

   // m148_44 = W*in
   wire signed [9:0] m148_44;
   assign m148_44 =10'b0;

   // m148_45 = W*in
   wire signed [9:0] m148_45;
   assign m148_45 =10'b0;

   // m148_46 = W*in
   wire signed [9:0] m148_46;
   assign m148_46 =10'b0;

   // m148_47 = W*in
   wire signed [9:0] m148_47;
   assign m148_47 =10'b0;

   // m148_48 = W*in
   wire signed [9:0] m148_48;
   assign m148_48 =10'b0;

   // m148_49 = W*in
   wire signed [9:0] m148_49;
   assign m148_49 =10'b0;

   // m148_50 = W*in
   wire signed [9:0] m148_50;
   assign m148_50 =10'b0;

   // m148_51 = W*in
   wire signed [9:0] m148_51;
   assign m148_51 =10'b0;

   // m148_52 = W*in
   wire signed [9:0] m148_52;
   assign m148_52 =10'b0;

   // m148_53 = W*in
   wire signed [9:0] m148_53;
   assign m148_53 =10'b0;

   // m148_54 = W*in
   wire signed [9:0] m148_54;
   assign m148_54 =10'b0;

   // m148_55 = W*in
   wire signed [9:0] m148_55;
   assign m148_55 =10'b0;

   // m148_56 = W*in
   wire signed [9:0] m148_56;
   assign m148_56 =10'b0;

   // m148_57 = W*in
   wire signed [9:0] m148_57;
   assign m148_57 =10'b0;

   // m148_58 = W*in
   wire signed [9:0] m148_58;
   assign m148_58 =10'b0;

   // m148_59 = W*in
   wire signed [9:0] m148_59;
   assign m148_59 =10'b0;

   // m148_60 = W*in
   wire signed [9:0] m148_60;
   assign m148_60 =10'b0;

   // m148_61 = W*in
   wire signed [9:0] m148_61;
   assign m148_61 =10'b0;

   // m148_62 = W*in
   wire signed [9:0] m148_62;
   assign m148_62 =10'b0;

   // m148_63 = W*in
   wire signed [9:0] m148_63;
   assign m148_63 =10'b0;

   // m148_64 = W*in
   wire signed [9:0] m148_64;
   assign m148_64 =10'b0;

   // m148_65 = W*in
   wire signed [9:0] m148_65;
   assign m148_65 =10'b0;

   // m148_66 = W*in
   wire signed [9:0] m148_66;
   assign m148_66 ={ {5{in148[5]}} , in148[5:1] };

   // m148_67 = W*in
   wire signed [9:0] m148_67;
   assign m148_67 =10'b0;

   // m148_68 = W*in
   wire signed [9:0] m148_68;
   assign m148_68 =10'b0;

   // m148_69 = W*in
   wire signed [9:0] m148_69;
   assign m148_69 =10'b0;

   // m148_70 = W*in
   wire signed [9:0] m148_70;
   assign m148_70 ={ {5{in148[5]}} , in148[5:1] };

   // m148_71 = W*in
   wire signed [9:0] m148_71;
   assign m148_71 =10'b0;

   // m148_72 = W*in
   wire signed [9:0] m148_72;
   assign m148_72 ={ {5{in148[5]}} , in148[5:1] };

   // m148_73 = W*in
   wire signed [9:0] m148_73;
   assign m148_73 =10'b0;

   // m148_74 = W*in
   wire signed [9:0] m148_74;
   assign m148_74 =10'b0;

   // m148_75 = W*in
   wire signed [9:0] m148_75;
   assign m148_75 ={ {5{neg148[5]}} , neg148[5:1] };

   // m148_76 = W*in
   wire signed [9:0] m148_76;
   assign m148_76 =10'b0;

   // m148_77 = W*in
   wire signed [9:0] m148_77;
   assign m148_77 =10'b0;

   // m148_78 = W*in
   wire signed [9:0] m148_78;
   assign m148_78 ={ {5{neg148[5]}} , neg148[5:1] };

   // m148_79 = W*in
   wire signed [9:0] m148_79;
   assign m148_79 =10'b0;

   // m148_80 = W*in
   wire signed [9:0] m148_80;
   assign m148_80 =10'b0;

   // m148_81 = W*in
   wire signed [9:0] m148_81;
   assign m148_81 =10'b0;

   // m148_82 = W*in
   wire signed [9:0] m148_82;
   assign m148_82 =10'b0;

   // m148_83 = W*in
   wire signed [9:0] m148_83;
   assign m148_83 =10'b0;

   // m148_84 = W*in
   wire signed [9:0] m148_84;
   assign m148_84 =10'b0;

   // m148_85 = W*in
   wire signed [9:0] m148_85;
   assign m148_85 =10'b0;

   // m148_86 = W*in
   wire signed [9:0] m148_86;
   assign m148_86 =10'b0;

   // m148_87 = W*in
   wire signed [9:0] m148_87;
   assign m148_87 =10'b0;

   // m148_88 = W*in
   wire signed [9:0] m148_88;
   assign m148_88 =10'b0;

   // m148_89 = W*in
   wire signed [9:0] m148_89;
   assign m148_89 =10'b0;

   // m148_90 = W*in
   wire signed [9:0] m148_90;
   assign m148_90 =10'b0;

   // m148_91 = W*in
   wire signed [9:0] m148_91;
   assign m148_91 =10'b0;

   // m148_92 = W*in
   wire signed [9:0] m148_92;
   assign m148_92 =10'b0;

   // m148_93 = W*in
   wire signed [9:0] m148_93;
   assign m148_93 =10'b0;

   // m148_94 = W*in
   wire signed [9:0] m148_94;
   assign m148_94 =10'b0;

   // m148_95 = W*in
   wire signed [9:0] m148_95;
   assign m148_95 =10'b0;

   // m148_96 = W*in
   wire signed [9:0] m148_96;
   assign m148_96 =10'b0;

   // m148_97 = W*in
   wire signed [9:0] m148_97;
   assign m148_97 =10'b0;

   // m148_98 = W*in
   wire signed [9:0] m148_98;
   assign m148_98 =10'b0;

   // m148_99 = W*in
   wire signed [9:0] m148_99;
   assign m148_99 =10'b0;

   // m148_100 = W*in
   wire signed [9:0] m148_100;
   assign m148_100 =10'b0;

   // m148_101 = W*in
   wire signed [9:0] m148_101;
   assign m148_101 =10'b0;

   // m148_102 = W*in
   wire signed [9:0] m148_102;
   assign m148_102 =10'b0;

   // m148_103 = W*in
   wire signed [9:0] m148_103;
   assign m148_103 =10'b0;

   // m148_104 = W*in
   wire signed [9:0] m148_104;
   assign m148_104 =10'b0;

   // m148_105 = W*in
   wire signed [9:0] m148_105;
   assign m148_105 =10'b0;

   // m148_106 = W*in
   wire signed [9:0] m148_106;
   assign m148_106 =10'b0;

   // m148_107 = W*in
   wire signed [9:0] m148_107;
   assign m148_107 =10'b0;

   // m148_108 = W*in
   wire signed [9:0] m148_108;
   assign m148_108 ={ {5{neg148[5]}} , neg148[5:1] };

   // m148_109 = W*in
   wire signed [9:0] m148_109;
   assign m148_109 =10'b0;

   // m148_110 = W*in
   wire signed [9:0] m148_110;
   assign m148_110 =10'b0;

   // m148_111 = W*in
   wire signed [9:0] m148_111;
   assign m148_111 =10'b0;

   // m148_112 = W*in
   wire signed [9:0] m148_112;
   assign m148_112 =10'b0;

   // m148_113 = W*in
   wire signed [9:0] m148_113;
   assign m148_113 =10'b0;

   // m148_114 = W*in
   wire signed [9:0] m148_114;
   assign m148_114 ={ {5{neg148[5]}} , neg148[5:1] };

   // m148_115 = W*in
   wire signed [9:0] m148_115;
   assign m148_115 ={ {4{neg148[5]}} , neg148[5:0] };

   // m148_116 = W*in
   wire signed [9:0] m148_116;
   assign m148_116 =10'b0;

   // m148_117 = W*in
   wire signed [9:0] m148_117;
   assign m148_117 =10'b0;

   // m149_1 = W*in
   wire signed [9:0] m149_1;
   assign m149_1 =10'b0;

   // m149_2 = W*in
   wire signed [9:0] m149_2;
   assign m149_2 =10'b0;

   // m149_3 = W*in
   wire signed [9:0] m149_3;
   assign m149_3 =10'b0;

   // m149_4 = W*in
   wire signed [9:0] m149_4;
   assign m149_4 =10'b0;

   // m149_5 = W*in
   wire signed [9:0] m149_5;
   assign m149_5 =10'b0;

   // m149_6 = W*in
   wire signed [9:0] m149_6;
   assign m149_6 =10'b0;

   // m149_7 = W*in
   wire signed [9:0] m149_7;
   assign m149_7 =10'b0;

   // m149_8 = W*in
   wire signed [9:0] m149_8;
   assign m149_8 =10'b0;

   // m149_9 = W*in
   wire signed [9:0] m149_9;
   assign m149_9 =10'b0;

   // m149_10 = W*in
   wire signed [9:0] m149_10;
   assign m149_10 =10'b0;

   // m149_11 = W*in
   wire signed [9:0] m149_11;
   assign m149_11 =10'b0;

   // m149_12 = W*in
   wire signed [9:0] m149_12;
   assign m149_12 =10'b0;

   // m149_13 = W*in
   wire signed [9:0] m149_13;
   assign m149_13 =10'b0;

   // m149_14 = W*in
   wire signed [9:0] m149_14;
   assign m149_14 =10'b0;

   // m149_15 = W*in
   wire signed [9:0] m149_15;
   assign m149_15 =10'b0;

   // m149_16 = W*in
   wire signed [9:0] m149_16;
   assign m149_16 =10'b0;

   // m149_17 = W*in
   wire signed [9:0] m149_17;
   assign m149_17 ={ {5{neg149[5]}} , neg149[5:1] };

   // m149_18 = W*in
   wire signed [9:0] m149_18;
   assign m149_18 ={ {5{in149[5]}} , in149[5:1] };

   // m149_19 = W*in
   wire signed [9:0] m149_19;
   assign m149_19 ={ {4{neg149[5]}} , neg149[5:0] };

   // m149_20 = W*in
   wire signed [9:0] m149_20;
   assign m149_20 ={ {5{neg149[5]}} , neg149[5:1] };

   // m149_21 = W*in
   wire signed [9:0] m149_21;
   assign m149_21 ={ {5{in149[5]}} , in149[5:1] };

   // m149_22 = W*in
   wire signed [9:0] m149_22;
   assign m149_22 =10'b0;

   // m149_23 = W*in
   wire signed [9:0] m149_23;
   assign m149_23 ={ {5{in149[5]}} , in149[5:1] };

   // m149_24 = W*in
   wire signed [9:0] m149_24;
   assign m149_24 =10'b0;

   // m149_25 = W*in
   wire signed [9:0] m149_25;
   assign m149_25 =10'b0;

   // m149_26 = W*in
   wire signed [9:0] m149_26;
   assign m149_26 =10'b0;

   // m149_27 = W*in
   wire signed [9:0] m149_27;
   assign m149_27 =10'b0;

   // m149_28 = W*in
   wire signed [9:0] m149_28;
   assign m149_28 =10'b0;

   // m149_29 = W*in
   wire signed [9:0] m149_29;
   assign m149_29 ={ {4{in149[5]}} , in149[5:0] };

   // m149_30 = W*in
   wire signed [9:0] m149_30;
   assign m149_30 ={ {4{neg149[5]}} , neg149[5:0] };

   // m149_31 = W*in
   wire signed [9:0] m149_31;
   assign m149_31 =10'b0;

   // m149_32 = W*in
   wire signed [9:0] m149_32;
   assign m149_32 =10'b0;

   // m149_33 = W*in
   wire signed [9:0] m149_33;
   assign m149_33 =10'b0;

   // m149_34 = W*in
   wire signed [9:0] m149_34;
   assign m149_34 =10'b0;

   // m149_35 = W*in
   wire signed [9:0] m149_35;
   assign m149_35 ={ {5{neg149[5]}} , neg149[5:1] };

   // m149_36 = W*in
   wire signed [9:0] m149_36;
   assign m149_36 ={ {5{in149[5]}} , in149[5:1] };

   // m149_37 = W*in
   wire signed [9:0] m149_37;
   assign m149_37 =10'b0;

   // m149_38 = W*in
   wire signed [9:0] m149_38;
   assign m149_38 =10'b0;

   // m149_39 = W*in
   wire signed [9:0] m149_39;
   assign m149_39 =10'b0;

   // m149_40 = W*in
   wire signed [9:0] m149_40;
   assign m149_40 =10'b0;

   // m149_41 = W*in
   wire signed [9:0] m149_41;
   assign m149_41 =10'b0;

   // m149_42 = W*in
   wire signed [9:0] m149_42;
   assign m149_42 =10'b0;

   // m149_43 = W*in
   wire signed [9:0] m149_43;
   assign m149_43 =10'b0;

   // m149_44 = W*in
   wire signed [9:0] m149_44;
   assign m149_44 =10'b0;

   // m149_45 = W*in
   wire signed [9:0] m149_45;
   assign m149_45 =10'b0;

   // m149_46 = W*in
   wire signed [9:0] m149_46;
   assign m149_46 =10'b0;

   // m149_47 = W*in
   wire signed [9:0] m149_47;
   assign m149_47 =10'b0;

   // m149_48 = W*in
   wire signed [9:0] m149_48;
   assign m149_48 =10'b0;

   // m149_49 = W*in
   wire signed [9:0] m149_49;
   assign m149_49 =10'b0;

   // m149_50 = W*in
   wire signed [9:0] m149_50;
   assign m149_50 =10'b0;

   // m149_51 = W*in
   wire signed [9:0] m149_51;
   assign m149_51 =10'b0;

   // m149_52 = W*in
   wire signed [9:0] m149_52;
   assign m149_52 =10'b0;

   // m149_53 = W*in
   wire signed [9:0] m149_53;
   assign m149_53 =10'b0;

   // m149_54 = W*in
   wire signed [9:0] m149_54;
   assign m149_54 =10'b0;

   // m149_55 = W*in
   wire signed [9:0] m149_55;
   assign m149_55 =10'b0;

   // m149_56 = W*in
   wire signed [9:0] m149_56;
   assign m149_56 =10'b0;

   // m149_57 = W*in
   wire signed [9:0] m149_57;
   assign m149_57 =10'b0;

   // m149_58 = W*in
   wire signed [9:0] m149_58;
   assign m149_58 =10'b0;

   // m149_59 = W*in
   wire signed [9:0] m149_59;
   assign m149_59 =10'b0;

   // m149_60 = W*in
   wire signed [9:0] m149_60;
   assign m149_60 =10'b0;

   // m149_61 = W*in
   wire signed [9:0] m149_61;
   assign m149_61 =10'b0;

   // m149_62 = W*in
   wire signed [9:0] m149_62;
   assign m149_62 =10'b0;

   // m149_63 = W*in
   wire signed [9:0] m149_63;
   assign m149_63 =10'b0;

   // m149_64 = W*in
   wire signed [9:0] m149_64;
   assign m149_64 ={ {5{neg149[5]}} , neg149[5:1] };

   // m149_65 = W*in
   wire signed [9:0] m149_65;
   assign m149_65 ={ {5{neg149[5]}} , neg149[5:1] };

   // m149_66 = W*in
   wire signed [9:0] m149_66;
   assign m149_66 =10'b0;

   // m149_67 = W*in
   wire signed [9:0] m149_67;
   assign m149_67 =10'b0;

   // m149_68 = W*in
   wire signed [9:0] m149_68;
   assign m149_68 =10'b0;

   // m149_69 = W*in
   wire signed [9:0] m149_69;
   assign m149_69 =10'b0;

   // m149_70 = W*in
   wire signed [9:0] m149_70;
   assign m149_70 ={ {4{in149[5]}} , in149[5:0] };

   // m149_71 = W*in
   wire signed [9:0] m149_71;
   assign m149_71 =10'b0;

   // m149_72 = W*in
   wire signed [9:0] m149_72;
   assign m149_72 ={ {4{in149[5]}} , in149[5:0] };

   // m149_73 = W*in
   wire signed [9:0] m149_73;
   assign m149_73 =10'b0;

   // m149_74 = W*in
   wire signed [9:0] m149_74;
   assign m149_74 =10'b0;

   // m149_75 = W*in
   wire signed [9:0] m149_75;
   assign m149_75 =10'b0;

   // m149_76 = W*in
   wire signed [9:0] m149_76;
   assign m149_76 =10'b0;

   // m149_77 = W*in
   wire signed [9:0] m149_77;
   assign m149_77 =10'b0;

   // m149_78 = W*in
   wire signed [9:0] m149_78;
   assign m149_78 =10'b0;

   // m149_79 = W*in
   wire signed [9:0] m149_79;
   assign m149_79 =10'b0;

   // m149_80 = W*in
   wire signed [9:0] m149_80;
   assign m149_80 =10'b0;

   // m149_81 = W*in
   wire signed [9:0] m149_81;
   assign m149_81 =10'b0;

   // m149_82 = W*in
   wire signed [9:0] m149_82;
   assign m149_82 =10'b0;

   // m149_83 = W*in
   wire signed [9:0] m149_83;
   assign m149_83 =10'b0;

   // m149_84 = W*in
   wire signed [9:0] m149_84;
   assign m149_84 ={ {4{in149[5]}} , in149[5:0] };

   // m149_85 = W*in
   wire signed [9:0] m149_85;
   assign m149_85 =10'b0;

   // m149_86 = W*in
   wire signed [9:0] m149_86;
   assign m149_86 =10'b0;

   // m149_87 = W*in
   wire signed [9:0] m149_87;
   assign m149_87 =10'b0;

   // m149_88 = W*in
   wire signed [9:0] m149_88;
   assign m149_88 =10'b0;

   // m149_89 = W*in
   wire signed [9:0] m149_89;
   assign m149_89 ={ {4{in149[5]}} , in149[5:0] };

   // m149_90 = W*in
   wire signed [9:0] m149_90;
   assign m149_90 =10'b0;

   // m149_91 = W*in
   wire signed [9:0] m149_91;
   assign m149_91 ={ {4{neg149[5]}} , neg149[5:0] };

   // m149_92 = W*in
   wire signed [9:0] m149_92;
   assign m149_92 =10'b0;

   // m149_93 = W*in
   wire signed [9:0] m149_93;
   assign m149_93 =10'b0;

   // m149_94 = W*in
   wire signed [9:0] m149_94;
   assign m149_94 =10'b0;

   // m149_95 = W*in
   wire signed [9:0] m149_95;
   assign m149_95 =10'b0;

   // m149_96 = W*in
   wire signed [9:0] m149_96;
   assign m149_96 =10'b0;

   // m149_97 = W*in
   wire signed [9:0] m149_97;
   assign m149_97 ={ {4{neg149[5]}} , neg149[5:0] };

   // m149_98 = W*in
   wire signed [9:0] m149_98;
   assign m149_98 =10'b0;

   // m149_99 = W*in
   wire signed [9:0] m149_99;
   assign m149_99 ={ {4{in149[5]}} , in149[5:0] };

   // m149_100 = W*in
   wire signed [9:0] m149_100;
   assign m149_100 =10'b0;

   // m149_101 = W*in
   wire signed [9:0] m149_101;
   assign m149_101 =10'b0;

   // m149_102 = W*in
   wire signed [9:0] m149_102;
   assign m149_102 =10'b0;

   // m149_103 = W*in
   wire signed [9:0] m149_103;
   assign m149_103 =10'b0;

   // m149_104 = W*in
   wire signed [9:0] m149_104;
   assign m149_104 =10'b0;

   // m149_105 = W*in
   wire signed [9:0] m149_105;
   assign m149_105 =10'b0;

   // m149_106 = W*in
   wire signed [9:0] m149_106;
   assign m149_106 =10'b0;

   // m149_107 = W*in
   wire signed [9:0] m149_107;
   assign m149_107 ={ {5{neg149[5]}} , neg149[5:1] };

   // m149_108 = W*in
   wire signed [9:0] m149_108;
   assign m149_108 =10'b0;

   // m149_109 = W*in
   wire signed [9:0] m149_109;
   assign m149_109 =10'b0;

   // m149_110 = W*in
   wire signed [9:0] m149_110;
   assign m149_110 =10'b0;

   // m149_111 = W*in
   wire signed [9:0] m149_111;
   assign m149_111 =10'b0;

   // m149_112 = W*in
   wire signed [9:0] m149_112;
   assign m149_112 =10'b0;

   // m149_113 = W*in
   wire signed [9:0] m149_113;
   assign m149_113 =10'b0;

   // m149_114 = W*in
   wire signed [9:0] m149_114;
   assign m149_114 =10'b0;

   // m149_115 = W*in
   wire signed [9:0] m149_115;
   assign m149_115 =10'b0;

   // m149_116 = W*in
   wire signed [9:0] m149_116;
   assign m149_116 =10'b0;

   // m149_117 = W*in
   wire signed [9:0] m149_117;
   assign m149_117 =10'b0;

   // m150_1 = W*in
   wire signed [9:0] m150_1;
   assign m150_1 =10'b0;

   // m150_2 = W*in
   wire signed [9:0] m150_2;
   assign m150_2 =10'b0;

   // m150_3 = W*in
   wire signed [9:0] m150_3;
   assign m150_3 =10'b0;

   // m150_4 = W*in
   wire signed [9:0] m150_4;
   assign m150_4 =10'b0;

   // m150_5 = W*in
   wire signed [9:0] m150_5;
   assign m150_5 =10'b0;

   // m150_6 = W*in
   wire signed [9:0] m150_6;
   assign m150_6 =10'b0;

   // m150_7 = W*in
   wire signed [9:0] m150_7;
   assign m150_7 =10'b0;

   // m150_8 = W*in
   wire signed [9:0] m150_8;
   assign m150_8 =10'b0;

   // m150_9 = W*in
   wire signed [9:0] m150_9;
   assign m150_9 =10'b0;

   // m150_10 = W*in
   wire signed [9:0] m150_10;
   assign m150_10 =10'b0;

   // m150_11 = W*in
   wire signed [9:0] m150_11;
   assign m150_11 =10'b0;

   // m150_12 = W*in
   wire signed [9:0] m150_12;
   assign m150_12 =10'b0;

   // m150_13 = W*in
   wire signed [9:0] m150_13;
   assign m150_13 =10'b0;

   // m150_14 = W*in
   wire signed [9:0] m150_14;
   assign m150_14 =10'b0;

   // m150_15 = W*in
   wire signed [9:0] m150_15;
   assign m150_15 =10'b0;

   // m150_16 = W*in
   wire signed [9:0] m150_16;
   assign m150_16 =10'b0;

   // m150_17 = W*in
   wire signed [9:0] m150_17;
   assign m150_17 =10'b0;

   // m150_18 = W*in
   wire signed [9:0] m150_18;
   assign m150_18 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_19 = W*in
   wire signed [9:0] m150_19;
   assign m150_19 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_20 = W*in
   wire signed [9:0] m150_20;
   assign m150_20 =10'b0;

   // m150_21 = W*in
   wire signed [9:0] m150_21;
   assign m150_21 =10'b0;

   // m150_22 = W*in
   wire signed [9:0] m150_22;
   assign m150_22 =10'b0;

   // m150_23 = W*in
   wire signed [9:0] m150_23;
   assign m150_23 =10'b0;

   // m150_24 = W*in
   wire signed [9:0] m150_24;
   assign m150_24 =10'b0;

   // m150_25 = W*in
   wire signed [9:0] m150_25;
   assign m150_25 =10'b0;

   // m150_26 = W*in
   wire signed [9:0] m150_26;
   assign m150_26 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_27 = W*in
   wire signed [9:0] m150_27;
   assign m150_27 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_28 = W*in
   wire signed [9:0] m150_28;
   assign m150_28 =10'b0;

   // m150_29 = W*in
   wire signed [9:0] m150_29;
   assign m150_29 =10'b0;

   // m150_30 = W*in
   wire signed [9:0] m150_30;
   assign m150_30 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_31 = W*in
   wire signed [9:0] m150_31;
   assign m150_31 =10'b0;

   // m150_32 = W*in
   wire signed [9:0] m150_32;
   assign m150_32 =10'b0;

   // m150_33 = W*in
   wire signed [9:0] m150_33;
   assign m150_33 =10'b0;

   // m150_34 = W*in
   wire signed [9:0] m150_34;
   assign m150_34 =10'b0;

   // m150_35 = W*in
   wire signed [9:0] m150_35;
   assign m150_35 =10'b0;

   // m150_36 = W*in
   wire signed [9:0] m150_36;
   assign m150_36 =10'b0;

   // m150_37 = W*in
   wire signed [9:0] m150_37;
   assign m150_37 =10'b0;

   // m150_38 = W*in
   wire signed [9:0] m150_38;
   assign m150_38 =10'b0;

   // m150_39 = W*in
   wire signed [9:0] m150_39;
   assign m150_39 =10'b0;

   // m150_40 = W*in
   wire signed [9:0] m150_40;
   assign m150_40 =10'b0;

   // m150_41 = W*in
   wire signed [9:0] m150_41;
   assign m150_41 =10'b0;

   // m150_42 = W*in
   wire signed [9:0] m150_42;
   assign m150_42 =10'b0;

   // m150_43 = W*in
   wire signed [9:0] m150_43;
   assign m150_43 =10'b0;

   // m150_44 = W*in
   wire signed [9:0] m150_44;
   assign m150_44 =10'b0;

   // m150_45 = W*in
   wire signed [9:0] m150_45;
   assign m150_45 =10'b0;

   // m150_46 = W*in
   wire signed [9:0] m150_46;
   assign m150_46 =10'b0;

   // m150_47 = W*in
   wire signed [9:0] m150_47;
   assign m150_47 =10'b0;

   // m150_48 = W*in
   wire signed [9:0] m150_48;
   assign m150_48 =10'b0;

   // m150_49 = W*in
   wire signed [9:0] m150_49;
   assign m150_49 =10'b0;

   // m150_50 = W*in
   wire signed [9:0] m150_50;
   assign m150_50 =10'b0;

   // m150_51 = W*in
   wire signed [9:0] m150_51;
   assign m150_51 =10'b0;

   // m150_52 = W*in
   wire signed [9:0] m150_52;
   assign m150_52 =10'b0;

   // m150_53 = W*in
   wire signed [9:0] m150_53;
   assign m150_53 =10'b0;

   // m150_54 = W*in
   wire signed [9:0] m150_54;
   assign m150_54 =10'b0;

   // m150_55 = W*in
   wire signed [9:0] m150_55;
   assign m150_55 =10'b0;

   // m150_56 = W*in
   wire signed [9:0] m150_56;
   assign m150_56 =10'b0;

   // m150_57 = W*in
   wire signed [9:0] m150_57;
   assign m150_57 =10'b0;

   // m150_58 = W*in
   wire signed [9:0] m150_58;
   assign m150_58 =10'b0;

   // m150_59 = W*in
   wire signed [9:0] m150_59;
   assign m150_59 =10'b0;

   // m150_60 = W*in
   wire signed [9:0] m150_60;
   assign m150_60 =10'b0;

   // m150_61 = W*in
   wire signed [9:0] m150_61;
   assign m150_61 =10'b0;

   // m150_62 = W*in
   wire signed [9:0] m150_62;
   assign m150_62 =10'b0;

   // m150_63 = W*in
   wire signed [9:0] m150_63;
   assign m150_63 =10'b0;

   // m150_64 = W*in
   wire signed [9:0] m150_64;
   assign m150_64 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_65 = W*in
   wire signed [9:0] m150_65;
   assign m150_65 =10'b0;

   // m150_66 = W*in
   wire signed [9:0] m150_66;
   assign m150_66 =10'b0;

   // m150_67 = W*in
   wire signed [9:0] m150_67;
   assign m150_67 =10'b0;

   // m150_68 = W*in
   wire signed [9:0] m150_68;
   assign m150_68 =10'b0;

   // m150_69 = W*in
   wire signed [9:0] m150_69;
   assign m150_69 =10'b0;

   // m150_70 = W*in
   wire signed [9:0] m150_70;
   assign m150_70 ={ {5{in150[5]}} , in150[5:1] };

   // m150_71 = W*in
   wire signed [9:0] m150_71;
   assign m150_71 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_72 = W*in
   wire signed [9:0] m150_72;
   assign m150_72 =10'b0;

   // m150_73 = W*in
   wire signed [9:0] m150_73;
   assign m150_73 =10'b0;

   // m150_74 = W*in
   wire signed [9:0] m150_74;
   assign m150_74 =10'b0;

   // m150_75 = W*in
   wire signed [9:0] m150_75;
   assign m150_75 =10'b0;

   // m150_76 = W*in
   wire signed [9:0] m150_76;
   assign m150_76 =10'b0;

   // m150_77 = W*in
   wire signed [9:0] m150_77;
   assign m150_77 =10'b0;

   // m150_78 = W*in
   wire signed [9:0] m150_78;
   assign m150_78 =10'b0;

   // m150_79 = W*in
   wire signed [9:0] m150_79;
   assign m150_79 =10'b0;

   // m150_80 = W*in
   wire signed [9:0] m150_80;
   assign m150_80 =10'b0;

   // m150_81 = W*in
   wire signed [9:0] m150_81;
   assign m150_81 =10'b0;

   // m150_82 = W*in
   wire signed [9:0] m150_82;
   assign m150_82 =10'b0;

   // m150_83 = W*in
   wire signed [9:0] m150_83;
   assign m150_83 =10'b0;

   // m150_84 = W*in
   wire signed [9:0] m150_84;
   assign m150_84 =10'b0;

   // m150_85 = W*in
   wire signed [9:0] m150_85;
   assign m150_85 =10'b0;

   // m150_86 = W*in
   wire signed [9:0] m150_86;
   assign m150_86 =10'b0;

   // m150_87 = W*in
   wire signed [9:0] m150_87;
   assign m150_87 =10'b0;

   // m150_88 = W*in
   wire signed [9:0] m150_88;
   assign m150_88 =10'b0;

   // m150_89 = W*in
   wire signed [9:0] m150_89;
   assign m150_89 =10'b0;

   // m150_90 = W*in
   wire signed [9:0] m150_90;
   assign m150_90 =10'b0;

   // m150_91 = W*in
   wire signed [9:0] m150_91;
   assign m150_91 =10'b0;

   // m150_92 = W*in
   wire signed [9:0] m150_92;
   assign m150_92 =10'b0;

   // m150_93 = W*in
   wire signed [9:0] m150_93;
   assign m150_93 =10'b0;

   // m150_94 = W*in
   wire signed [9:0] m150_94;
   assign m150_94 =10'b0;

   // m150_95 = W*in
   wire signed [9:0] m150_95;
   assign m150_95 =10'b0;

   // m150_96 = W*in
   wire signed [9:0] m150_96;
   assign m150_96 =10'b0;

   // m150_97 = W*in
   wire signed [9:0] m150_97;
   assign m150_97 =10'b0;

   // m150_98 = W*in
   wire signed [9:0] m150_98;
   assign m150_98 =10'b0;

   // m150_99 = W*in
   wire signed [9:0] m150_99;
   assign m150_99 =10'b0;

   // m150_100 = W*in
   wire signed [9:0] m150_100;
   assign m150_100 =10'b0;

   // m150_101 = W*in
   wire signed [9:0] m150_101;
   assign m150_101 =10'b0;

   // m150_102 = W*in
   wire signed [9:0] m150_102;
   assign m150_102 =10'b0;

   // m150_103 = W*in
   wire signed [9:0] m150_103;
   assign m150_103 =10'b0;

   // m150_104 = W*in
   wire signed [9:0] m150_104;
   assign m150_104 =10'b0;

   // m150_105 = W*in
   wire signed [9:0] m150_105;
   assign m150_105 =10'b0;

   // m150_106 = W*in
   wire signed [9:0] m150_106;
   assign m150_106 =10'b0;

   // m150_107 = W*in
   wire signed [9:0] m150_107;
   assign m150_107 ={ {5{neg150[5]}} , neg150[5:1] };

   // m150_108 = W*in
   wire signed [9:0] m150_108;
   assign m150_108 ={ {5{in150[5]}} , in150[5:1] };

   // m150_109 = W*in
   wire signed [9:0] m150_109;
   assign m150_109 ={ {5{in150[5]}} , in150[5:1] };

   // m150_110 = W*in
   wire signed [9:0] m150_110;
   assign m150_110 =10'b0;

   // m150_111 = W*in
   wire signed [9:0] m150_111;
   assign m150_111 =10'b0;

   // m150_112 = W*in
   wire signed [9:0] m150_112;
   assign m150_112 =10'b0;

   // m150_113 = W*in
   wire signed [9:0] m150_113;
   assign m150_113 =10'b0;

   // m150_114 = W*in
   wire signed [9:0] m150_114;
   assign m150_114 =10'b0;

   // m150_115 = W*in
   wire signed [9:0] m150_115;
   assign m150_115 =10'b0;

   // m150_116 = W*in
   wire signed [9:0] m150_116;
   assign m150_116 =10'b0;

   // m150_117 = W*in
   wire signed [9:0] m150_117;
   assign m150_117 =10'b0;

   // m151_1 = W*in
   wire signed [9:0] m151_1;
   assign m151_1 =10'b0;

   // m151_2 = W*in
   wire signed [9:0] m151_2;
   assign m151_2 =10'b0;

   // m151_3 = W*in
   wire signed [9:0] m151_3;
   assign m151_3 =10'b0;

   // m151_4 = W*in
   wire signed [9:0] m151_4;
   assign m151_4 =10'b0;

   // m151_5 = W*in
   wire signed [9:0] m151_5;
   assign m151_5 =10'b0;

   // m151_6 = W*in
   wire signed [9:0] m151_6;
   assign m151_6 =10'b0;

   // m151_7 = W*in
   wire signed [9:0] m151_7;
   assign m151_7 =10'b0;

   // m151_8 = W*in
   wire signed [9:0] m151_8;
   assign m151_8 =10'b0;

   // m151_9 = W*in
   wire signed [9:0] m151_9;
   assign m151_9 =10'b0;

   // m151_10 = W*in
   wire signed [9:0] m151_10;
   assign m151_10 =10'b0;

   // m151_11 = W*in
   wire signed [9:0] m151_11;
   assign m151_11 =10'b0;

   // m151_12 = W*in
   wire signed [9:0] m151_12;
   assign m151_12 =10'b0;

   // m151_13 = W*in
   wire signed [9:0] m151_13;
   assign m151_13 =10'b0;

   // m151_14 = W*in
   wire signed [9:0] m151_14;
   assign m151_14 =10'b0;

   // m151_15 = W*in
   wire signed [9:0] m151_15;
   assign m151_15 =10'b0;

   // m151_16 = W*in
   wire signed [9:0] m151_16;
   assign m151_16 =10'b0;

   // m151_17 = W*in
   wire signed [9:0] m151_17;
   assign m151_17 =10'b0;

   // m151_18 = W*in
   wire signed [9:0] m151_18;
   assign m151_18 =10'b0;

   // m151_19 = W*in
   wire signed [9:0] m151_19;
   assign m151_19 =10'b0;

   // m151_20 = W*in
   wire signed [9:0] m151_20;
   assign m151_20 =10'b0;

   // m151_21 = W*in
   wire signed [9:0] m151_21;
   assign m151_21 =10'b0;

   // m151_22 = W*in
   wire signed [9:0] m151_22;
   assign m151_22 =10'b0;

   // m151_23 = W*in
   wire signed [9:0] m151_23;
   assign m151_23 =10'b0;

   // m151_24 = W*in
   wire signed [9:0] m151_24;
   assign m151_24 =10'b0;

   // m151_25 = W*in
   wire signed [9:0] m151_25;
   assign m151_25 =10'b0;

   // m151_26 = W*in
   wire signed [9:0] m151_26;
   assign m151_26 =10'b0;

   // m151_27 = W*in
   wire signed [9:0] m151_27;
   assign m151_27 =10'b0;

   // m151_28 = W*in
   wire signed [9:0] m151_28;
   assign m151_28 ={ {5{neg151[5]}} , neg151[5:1] };

   // m151_29 = W*in
   wire signed [9:0] m151_29;
   assign m151_29 =10'b0;

   // m151_30 = W*in
   wire signed [9:0] m151_30;
   assign m151_30 =10'b0;

   // m151_31 = W*in
   wire signed [9:0] m151_31;
   assign m151_31 =10'b0;

   // m151_32 = W*in
   wire signed [9:0] m151_32;
   assign m151_32 =10'b0;

   // m151_33 = W*in
   wire signed [9:0] m151_33;
   assign m151_33 =10'b0;

   // m151_34 = W*in
   wire signed [9:0] m151_34;
   assign m151_34 =10'b0;

   // m151_35 = W*in
   wire signed [9:0] m151_35;
   assign m151_35 =10'b0;

   // m151_36 = W*in
   wire signed [9:0] m151_36;
   assign m151_36 =10'b0;

   // m151_37 = W*in
   wire signed [9:0] m151_37;
   assign m151_37 =10'b0;

   // m151_38 = W*in
   wire signed [9:0] m151_38;
   assign m151_38 =10'b0;

   // m151_39 = W*in
   wire signed [9:0] m151_39;
   assign m151_39 =10'b0;

   // m151_40 = W*in
   wire signed [9:0] m151_40;
   assign m151_40 =10'b0;

   // m151_41 = W*in
   wire signed [9:0] m151_41;
   assign m151_41 =10'b0;

   // m151_42 = W*in
   wire signed [9:0] m151_42;
   assign m151_42 =10'b0;

   // m151_43 = W*in
   wire signed [9:0] m151_43;
   assign m151_43 =10'b0;

   // m151_44 = W*in
   wire signed [9:0] m151_44;
   assign m151_44 =10'b0;

   // m151_45 = W*in
   wire signed [9:0] m151_45;
   assign m151_45 =10'b0;

   // m151_46 = W*in
   wire signed [9:0] m151_46;
   assign m151_46 =10'b0;

   // m151_47 = W*in
   wire signed [9:0] m151_47;
   assign m151_47 =10'b0;

   // m151_48 = W*in
   wire signed [9:0] m151_48;
   assign m151_48 =10'b0;

   // m151_49 = W*in
   wire signed [9:0] m151_49;
   assign m151_49 =10'b0;

   // m151_50 = W*in
   wire signed [9:0] m151_50;
   assign m151_50 =10'b0;

   // m151_51 = W*in
   wire signed [9:0] m151_51;
   assign m151_51 =10'b0;

   // m151_52 = W*in
   wire signed [9:0] m151_52;
   assign m151_52 =10'b0;

   // m151_53 = W*in
   wire signed [9:0] m151_53;
   assign m151_53 =10'b0;

   // m151_54 = W*in
   wire signed [9:0] m151_54;
   assign m151_54 =10'b0;

   // m151_55 = W*in
   wire signed [9:0] m151_55;
   assign m151_55 =10'b0;

   // m151_56 = W*in
   wire signed [9:0] m151_56;
   assign m151_56 =10'b0;

   // m151_57 = W*in
   wire signed [9:0] m151_57;
   assign m151_57 =10'b0;

   // m151_58 = W*in
   wire signed [9:0] m151_58;
   assign m151_58 =10'b0;

   // m151_59 = W*in
   wire signed [9:0] m151_59;
   assign m151_59 =10'b0;

   // m151_60 = W*in
   wire signed [9:0] m151_60;
   assign m151_60 =10'b0;

   // m151_61 = W*in
   wire signed [9:0] m151_61;
   assign m151_61 =10'b0;

   // m151_62 = W*in
   wire signed [9:0] m151_62;
   assign m151_62 =10'b0;

   // m151_63 = W*in
   wire signed [9:0] m151_63;
   assign m151_63 =10'b0;

   // m151_64 = W*in
   wire signed [9:0] m151_64;
   assign m151_64 =10'b0;

   // m151_65 = W*in
   wire signed [9:0] m151_65;
   assign m151_65 =10'b0;

   // m151_66 = W*in
   wire signed [9:0] m151_66;
   assign m151_66 =10'b0;

   // m151_67 = W*in
   wire signed [9:0] m151_67;
   assign m151_67 =10'b0;

   // m151_68 = W*in
   wire signed [9:0] m151_68;
   assign m151_68 =10'b0;

   // m151_69 = W*in
   wire signed [9:0] m151_69;
   assign m151_69 =10'b0;

   // m151_70 = W*in
   wire signed [9:0] m151_70;
   assign m151_70 =10'b0;

   // m151_71 = W*in
   wire signed [9:0] m151_71;
   assign m151_71 =10'b0;

   // m151_72 = W*in
   wire signed [9:0] m151_72;
   assign m151_72 =10'b0;

   // m151_73 = W*in
   wire signed [9:0] m151_73;
   assign m151_73 =10'b0;

   // m151_74 = W*in
   wire signed [9:0] m151_74;
   assign m151_74 =10'b0;

   // m151_75 = W*in
   wire signed [9:0] m151_75;
   assign m151_75 =10'b0;

   // m151_76 = W*in
   wire signed [9:0] m151_76;
   assign m151_76 =10'b0;

   // m151_77 = W*in
   wire signed [9:0] m151_77;
   assign m151_77 =10'b0;

   // m151_78 = W*in
   wire signed [9:0] m151_78;
   assign m151_78 =10'b0;

   // m151_79 = W*in
   wire signed [9:0] m151_79;
   assign m151_79 =10'b0;

   // m151_80 = W*in
   wire signed [9:0] m151_80;
   assign m151_80 =10'b0;

   // m151_81 = W*in
   wire signed [9:0] m151_81;
   assign m151_81 =10'b0;

   // m151_82 = W*in
   wire signed [9:0] m151_82;
   assign m151_82 =10'b0;

   // m151_83 = W*in
   wire signed [9:0] m151_83;
   assign m151_83 =10'b0;

   // m151_84 = W*in
   wire signed [9:0] m151_84;
   assign m151_84 =10'b0;

   // m151_85 = W*in
   wire signed [9:0] m151_85;
   assign m151_85 =10'b0;

   // m151_86 = W*in
   wire signed [9:0] m151_86;
   assign m151_86 =10'b0;

   // m151_87 = W*in
   wire signed [9:0] m151_87;
   assign m151_87 =10'b0;

   // m151_88 = W*in
   wire signed [9:0] m151_88;
   assign m151_88 =10'b0;

   // m151_89 = W*in
   wire signed [9:0] m151_89;
   assign m151_89 =10'b0;

   // m151_90 = W*in
   wire signed [9:0] m151_90;
   assign m151_90 =10'b0;

   // m151_91 = W*in
   wire signed [9:0] m151_91;
   assign m151_91 =10'b0;

   // m151_92 = W*in
   wire signed [9:0] m151_92;
   assign m151_92 =10'b0;

   // m151_93 = W*in
   wire signed [9:0] m151_93;
   assign m151_93 =10'b0;

   // m151_94 = W*in
   wire signed [9:0] m151_94;
   assign m151_94 =10'b0;

   // m151_95 = W*in
   wire signed [9:0] m151_95;
   assign m151_95 =10'b0;

   // m151_96 = W*in
   wire signed [9:0] m151_96;
   assign m151_96 =10'b0;

   // m151_97 = W*in
   wire signed [9:0] m151_97;
   assign m151_97 =10'b0;

   // m151_98 = W*in
   wire signed [9:0] m151_98;
   assign m151_98 =10'b0;

   // m151_99 = W*in
   wire signed [9:0] m151_99;
   assign m151_99 =10'b0;

   // m151_100 = W*in
   wire signed [9:0] m151_100;
   assign m151_100 =10'b0;

   // m151_101 = W*in
   wire signed [9:0] m151_101;
   assign m151_101 =10'b0;

   // m151_102 = W*in
   wire signed [9:0] m151_102;
   assign m151_102 =10'b0;

   // m151_103 = W*in
   wire signed [9:0] m151_103;
   assign m151_103 =10'b0;

   // m151_104 = W*in
   wire signed [9:0] m151_104;
   assign m151_104 =10'b0;

   // m151_105 = W*in
   wire signed [9:0] m151_105;
   assign m151_105 =10'b0;

   // m151_106 = W*in
   wire signed [9:0] m151_106;
   assign m151_106 =10'b0;

   // m151_107 = W*in
   wire signed [9:0] m151_107;
   assign m151_107 =10'b0;

   // m151_108 = W*in
   wire signed [9:0] m151_108;
   assign m151_108 =10'b0;

   // m151_109 = W*in
   wire signed [9:0] m151_109;
   assign m151_109 =10'b0;

   // m151_110 = W*in
   wire signed [9:0] m151_110;
   assign m151_110 =10'b0;

   // m151_111 = W*in
   wire signed [9:0] m151_111;
   assign m151_111 =10'b0;

   // m151_112 = W*in
   wire signed [9:0] m151_112;
   assign m151_112 =10'b0;

   // m151_113 = W*in
   wire signed [9:0] m151_113;
   assign m151_113 =10'b0;

   // m151_114 = W*in
   wire signed [9:0] m151_114;
   assign m151_114 =10'b0;

   // m151_115 = W*in
   wire signed [9:0] m151_115;
   assign m151_115 =10'b0;

   // m151_116 = W*in
   wire signed [9:0] m151_116;
   assign m151_116 =10'b0;

   // m151_117 = W*in
   wire signed [9:0] m151_117;
   assign m151_117 =10'b0;

   // m152_1 = W*in
   wire signed [9:0] m152_1;
   assign m152_1 =10'b0;

   // m152_2 = W*in
   wire signed [9:0] m152_2;
   assign m152_2 =10'b0;

   // m152_3 = W*in
   wire signed [9:0] m152_3;
   assign m152_3 =10'b0;

   // m152_4 = W*in
   wire signed [9:0] m152_4;
   assign m152_4 =10'b0;

   // m152_5 = W*in
   wire signed [9:0] m152_5;
   assign m152_5 =10'b0;

   // m152_6 = W*in
   wire signed [9:0] m152_6;
   assign m152_6 =10'b0;

   // m152_7 = W*in
   wire signed [9:0] m152_7;
   assign m152_7 =10'b0;

   // m152_8 = W*in
   wire signed [9:0] m152_8;
   assign m152_8 ={ {4{neg152[5]}} , neg152[5:0] };

   // m152_9 = W*in
   wire signed [9:0] m152_9;
   assign m152_9 =10'b0;

   // m152_10 = W*in
   wire signed [9:0] m152_10;
   assign m152_10 ={ {4{in152[5]}} , in152[5:0] };

   // m152_11 = W*in
   wire signed [9:0] m152_11;
   assign m152_11 =10'b0;

   // m152_12 = W*in
   wire signed [9:0] m152_12;
   assign m152_12 =10'b0;

   // m152_13 = W*in
   wire signed [9:0] m152_13;
   assign m152_13 ={ {4{in152[5]}} , in152[5:0] };

   // m152_14 = W*in
   wire signed [9:0] m152_14;
   assign m152_14 =10'b0;

   // m152_15 = W*in
   wire signed [9:0] m152_15;
   assign m152_15 ={ {4{neg152[5]}} , neg152[5:0] };

   // m152_16 = W*in
   wire signed [9:0] m152_16;
   assign m152_16 =10'b0;

   // m152_17 = W*in
   wire signed [9:0] m152_17;
   assign m152_17 =10'b0;

   // m152_18 = W*in
   wire signed [9:0] m152_18;
   assign m152_18 =10'b0;

   // m152_19 = W*in
   wire signed [9:0] m152_19;
   assign m152_19 ={ {4{neg152[5]}} , neg152[5:0] };

   // m152_20 = W*in
   wire signed [9:0] m152_20;
   assign m152_20 ={ {5{neg152[5]}} , neg152[5:1] };

   // m152_21 = W*in
   wire signed [9:0] m152_21;
   assign m152_21 ={ {5{in152[5]}} , in152[5:1] };

   // m152_22 = W*in
   wire signed [9:0] m152_22;
   assign m152_22 =10'b0;

   // m152_23 = W*in
   wire signed [9:0] m152_23;
   assign m152_23 =10'b0;

   // m152_24 = W*in
   wire signed [9:0] m152_24;
   assign m152_24 =10'b0;

   // m152_25 = W*in
   wire signed [9:0] m152_25;
   assign m152_25 =10'b0;

   // m152_26 = W*in
   wire signed [9:0] m152_26;
   assign m152_26 ={ {4{in152[5]}} , in152[5:0] };

   // m152_27 = W*in
   wire signed [9:0] m152_27;
   assign m152_27 =10'b0;

   // m152_28 = W*in
   wire signed [9:0] m152_28;
   assign m152_28 =10'b0;

   // m152_29 = W*in
   wire signed [9:0] m152_29;
   assign m152_29 =10'b0;

   // m152_30 = W*in
   wire signed [9:0] m152_30;
   assign m152_30 =10'b0;

   // m152_31 = W*in
   wire signed [9:0] m152_31;
   assign m152_31 =10'b0;

   // m152_32 = W*in
   wire signed [9:0] m152_32;
   assign m152_32 =10'b0;

   // m152_33 = W*in
   wire signed [9:0] m152_33;
   assign m152_33 =10'b0;

   // m152_34 = W*in
   wire signed [9:0] m152_34;
   assign m152_34 =10'b0;

   // m152_35 = W*in
   wire signed [9:0] m152_35;
   assign m152_35 ={ {5{neg152[5]}} , neg152[5:1] };

   // m152_36 = W*in
   wire signed [9:0] m152_36;
   assign m152_36 =10'b0;

   // m152_37 = W*in
   wire signed [9:0] m152_37;
   assign m152_37 =10'b0;

   // m152_38 = W*in
   wire signed [9:0] m152_38;
   assign m152_38 =10'b0;

   // m152_39 = W*in
   wire signed [9:0] m152_39;
   assign m152_39 =10'b0;

   // m152_40 = W*in
   wire signed [9:0] m152_40;
   assign m152_40 =10'b0;

   // m152_41 = W*in
   wire signed [9:0] m152_41;
   assign m152_41 =10'b0;

   // m152_42 = W*in
   wire signed [9:0] m152_42;
   assign m152_42 =10'b0;

   // m152_43 = W*in
   wire signed [9:0] m152_43;
   assign m152_43 =10'b0;

   // m152_44 = W*in
   wire signed [9:0] m152_44;
   assign m152_44 =10'b0;

   // m152_45 = W*in
   wire signed [9:0] m152_45;
   assign m152_45 =10'b0;

   // m152_46 = W*in
   wire signed [9:0] m152_46;
   assign m152_46 =10'b0;

   // m152_47 = W*in
   wire signed [9:0] m152_47;
   assign m152_47 =10'b0;

   // m152_48 = W*in
   wire signed [9:0] m152_48;
   assign m152_48 =10'b0;

   // m152_49 = W*in
   wire signed [9:0] m152_49;
   assign m152_49 =10'b0;

   // m152_50 = W*in
   wire signed [9:0] m152_50;
   assign m152_50 ={ {4{neg152[5]}} , neg152[5:0] };

   // m152_51 = W*in
   wire signed [9:0] m152_51;
   assign m152_51 =10'b0;

   // m152_52 = W*in
   wire signed [9:0] m152_52;
   assign m152_52 =10'b0;

   // m152_53 = W*in
   wire signed [9:0] m152_53;
   assign m152_53 =10'b0;

   // m152_54 = W*in
   wire signed [9:0] m152_54;
   assign m152_54 =10'b0;

   // m152_55 = W*in
   wire signed [9:0] m152_55;
   assign m152_55 =10'b0;

   // m152_56 = W*in
   wire signed [9:0] m152_56;
   assign m152_56 =10'b0;

   // m152_57 = W*in
   wire signed [9:0] m152_57;
   assign m152_57 =10'b0;

   // m152_58 = W*in
   wire signed [9:0] m152_58;
   assign m152_58 =10'b0;

   // m152_59 = W*in
   wire signed [9:0] m152_59;
   assign m152_59 =10'b0;

   // m152_60 = W*in
   wire signed [9:0] m152_60;
   assign m152_60 =10'b0;

   // m152_61 = W*in
   wire signed [9:0] m152_61;
   assign m152_61 =10'b0;

   // m152_62 = W*in
   wire signed [9:0] m152_62;
   assign m152_62 =10'b0;

   // m152_63 = W*in
   wire signed [9:0] m152_63;
   assign m152_63 =10'b0;

   // m152_64 = W*in
   wire signed [9:0] m152_64;
   assign m152_64 =10'b0;

   // m152_65 = W*in
   wire signed [9:0] m152_65;
   assign m152_65 ={ {5{in152[5]}} , in152[5:1] };

   // m152_66 = W*in
   wire signed [9:0] m152_66;
   assign m152_66 ={ {5{in152[5]}} , in152[5:1] };

   // m152_67 = W*in
   wire signed [9:0] m152_67;
   assign m152_67 =10'b0;

   // m152_68 = W*in
   wire signed [9:0] m152_68;
   assign m152_68 =10'b0;

   // m152_69 = W*in
   wire signed [9:0] m152_69;
   assign m152_69 =10'b0;

   // m152_70 = W*in
   wire signed [9:0] m152_70;
   assign m152_70 =10'b0;

   // m152_71 = W*in
   wire signed [9:0] m152_71;
   assign m152_71 =10'b0;

   // m152_72 = W*in
   wire signed [9:0] m152_72;
   assign m152_72 ={ {4{in152[5]}} , in152[5:0] };

   // m152_73 = W*in
   wire signed [9:0] m152_73;
   assign m152_73 =10'b0;

   // m152_74 = W*in
   wire signed [9:0] m152_74;
   assign m152_74 =10'b0;

   // m152_75 = W*in
   wire signed [9:0] m152_75;
   assign m152_75 =10'b0;

   // m152_76 = W*in
   wire signed [9:0] m152_76;
   assign m152_76 =10'b0;

   // m152_77 = W*in
   wire signed [9:0] m152_77;
   assign m152_77 =10'b0;

   // m152_78 = W*in
   wire signed [9:0] m152_78;
   assign m152_78 ={ {4{in152[5]}} , in152[5:0] };

   // m152_79 = W*in
   wire signed [9:0] m152_79;
   assign m152_79 =10'b0;

   // m152_80 = W*in
   wire signed [9:0] m152_80;
   assign m152_80 =10'b0;

   // m152_81 = W*in
   wire signed [9:0] m152_81;
   assign m152_81 =10'b0;

   // m152_82 = W*in
   wire signed [9:0] m152_82;
   assign m152_82 =10'b0;

   // m152_83 = W*in
   wire signed [9:0] m152_83;
   assign m152_83 =10'b0;

   // m152_84 = W*in
   wire signed [9:0] m152_84;
   assign m152_84 =10'b0;

   // m152_85 = W*in
   wire signed [9:0] m152_85;
   assign m152_85 =10'b0;

   // m152_86 = W*in
   wire signed [9:0] m152_86;
   assign m152_86 ={ {4{in152[5]}} , in152[5:0] };

   // m152_87 = W*in
   wire signed [9:0] m152_87;
   assign m152_87 =10'b0;

   // m152_88 = W*in
   wire signed [9:0] m152_88;
   assign m152_88 =10'b0;

   // m152_89 = W*in
   wire signed [9:0] m152_89;
   assign m152_89 =10'b0;

   // m152_90 = W*in
   wire signed [9:0] m152_90;
   assign m152_90 =10'b0;

   // m152_91 = W*in
   wire signed [9:0] m152_91;
   assign m152_91 =10'b0;

   // m152_92 = W*in
   wire signed [9:0] m152_92;
   assign m152_92 =10'b0;

   // m152_93 = W*in
   wire signed [9:0] m152_93;
   assign m152_93 =10'b0;

   // m152_94 = W*in
   wire signed [9:0] m152_94;
   assign m152_94 =10'b0;

   // m152_95 = W*in
   wire signed [9:0] m152_95;
   assign m152_95 =10'b0;

   // m152_96 = W*in
   wire signed [9:0] m152_96;
   assign m152_96 =10'b0;

   // m152_97 = W*in
   wire signed [9:0] m152_97;
   assign m152_97 =10'b0;

   // m152_98 = W*in
   wire signed [9:0] m152_98;
   assign m152_98 =10'b0;

   // m152_99 = W*in
   wire signed [9:0] m152_99;
   assign m152_99 =10'b0;

   // m152_100 = W*in
   wire signed [9:0] m152_100;
   assign m152_100 =10'b0;

   // m152_101 = W*in
   wire signed [9:0] m152_101;
   assign m152_101 =10'b0;

   // m152_102 = W*in
   wire signed [9:0] m152_102;
   assign m152_102 ={ {4{in152[5]}} , in152[5:0] };

   // m152_103 = W*in
   wire signed [9:0] m152_103;
   assign m152_103 =10'b0;

   // m152_104 = W*in
   wire signed [9:0] m152_104;
   assign m152_104 =10'b0;

   // m152_105 = W*in
   wire signed [9:0] m152_105;
   assign m152_105 =10'b0;

   // m152_106 = W*in
   wire signed [9:0] m152_106;
   assign m152_106 =10'b0;

   // m152_107 = W*in
   wire signed [9:0] m152_107;
   assign m152_107 =10'b0;

   // m152_108 = W*in
   wire signed [9:0] m152_108;
   assign m152_108 =10'b0;

   // m152_109 = W*in
   wire signed [9:0] m152_109;
   assign m152_109 =10'b0;

   // m152_110 = W*in
   wire signed [9:0] m152_110;
   assign m152_110 =10'b0;

   // m152_111 = W*in
   wire signed [9:0] m152_111;
   assign m152_111 =10'b0;

   // m152_112 = W*in
   wire signed [9:0] m152_112;
   assign m152_112 =10'b0;

   // m152_113 = W*in
   wire signed [9:0] m152_113;
   assign m152_113 =10'b0;

   // m152_114 = W*in
   wire signed [9:0] m152_114;
   assign m152_114 ={ {5{neg152[5]}} , neg152[5:1] };

   // m152_115 = W*in
   wire signed [9:0] m152_115;
   assign m152_115 ={ {5{neg152[5]}} , neg152[5:1] };

   // m152_116 = W*in
   wire signed [9:0] m152_116;
   assign m152_116 =10'b0;

   // m152_117 = W*in
   wire signed [9:0] m152_117;
   assign m152_117 =10'b0;

   // m153_1 = W*in
   wire signed [9:0] m153_1;
   assign m153_1 =10'b0;

   // m153_2 = W*in
   wire signed [9:0] m153_2;
   assign m153_2 =10'b0;

   // m153_3 = W*in
   wire signed [9:0] m153_3;
   assign m153_3 =10'b0;

   // m153_4 = W*in
   wire signed [9:0] m153_4;
   assign m153_4 =10'b0;

   // m153_5 = W*in
   wire signed [9:0] m153_5;
   assign m153_5 =10'b0;

   // m153_6 = W*in
   wire signed [9:0] m153_6;
   assign m153_6 =10'b0;

   // m153_7 = W*in
   wire signed [9:0] m153_7;
   assign m153_7 =10'b0;

   // m153_8 = W*in
   wire signed [9:0] m153_8;
   assign m153_8 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_9 = W*in
   wire signed [9:0] m153_9;
   assign m153_9 =10'b0;

   // m153_10 = W*in
   wire signed [9:0] m153_10;
   assign m153_10 ={ {4{in153[5]}} , in153[5:0] };

   // m153_11 = W*in
   wire signed [9:0] m153_11;
   assign m153_11 =10'b0;

   // m153_12 = W*in
   wire signed [9:0] m153_12;
   assign m153_12 =10'b0;

   // m153_13 = W*in
   wire signed [9:0] m153_13;
   assign m153_13 =10'b0;

   // m153_14 = W*in
   wire signed [9:0] m153_14;
   assign m153_14 =10'b0;

   // m153_15 = W*in
   wire signed [9:0] m153_15;
   assign m153_15 =10'b0;

   // m153_16 = W*in
   wire signed [9:0] m153_16;
   assign m153_16 =10'b0;

   // m153_17 = W*in
   wire signed [9:0] m153_17;
   assign m153_17 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_18 = W*in
   wire signed [9:0] m153_18;
   assign m153_18 =10'b0;

   // m153_19 = W*in
   wire signed [9:0] m153_19;
   assign m153_19 =10'b0;

   // m153_20 = W*in
   wire signed [9:0] m153_20;
   assign m153_20 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_21 = W*in
   wire signed [9:0] m153_21;
   assign m153_21 ={ {4{in153[5]}} , in153[5:0] };

   // m153_22 = W*in
   wire signed [9:0] m153_22;
   assign m153_22 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_23 = W*in
   wire signed [9:0] m153_23;
   assign m153_23 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_24 = W*in
   wire signed [9:0] m153_24;
   assign m153_24 =10'b0;

   // m153_25 = W*in
   wire signed [9:0] m153_25;
   assign m153_25 =10'b0;

   // m153_26 = W*in
   wire signed [9:0] m153_26;
   assign m153_26 ={ {4{in153[5]}} , in153[5:0] };

   // m153_27 = W*in
   wire signed [9:0] m153_27;
   assign m153_27 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_28 = W*in
   wire signed [9:0] m153_28;
   assign m153_28 =10'b0;

   // m153_29 = W*in
   wire signed [9:0] m153_29;
   assign m153_29 =10'b0;

   // m153_30 = W*in
   wire signed [9:0] m153_30;
   assign m153_30 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_31 = W*in
   wire signed [9:0] m153_31;
   assign m153_31 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_32 = W*in
   wire signed [9:0] m153_32;
   assign m153_32 =10'b0;

   // m153_33 = W*in
   wire signed [9:0] m153_33;
   assign m153_33 =10'b0;

   // m153_34 = W*in
   wire signed [9:0] m153_34;
   assign m153_34 =10'b0;

   // m153_35 = W*in
   wire signed [9:0] m153_35;
   assign m153_35 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_36 = W*in
   wire signed [9:0] m153_36;
   assign m153_36 =10'b0;

   // m153_37 = W*in
   wire signed [9:0] m153_37;
   assign m153_37 =10'b0;

   // m153_38 = W*in
   wire signed [9:0] m153_38;
   assign m153_38 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_39 = W*in
   wire signed [9:0] m153_39;
   assign m153_39 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_40 = W*in
   wire signed [9:0] m153_40;
   assign m153_40 =10'b0;

   // m153_41 = W*in
   wire signed [9:0] m153_41;
   assign m153_41 =10'b0;

   // m153_42 = W*in
   wire signed [9:0] m153_42;
   assign m153_42 =10'b0;

   // m153_43 = W*in
   wire signed [9:0] m153_43;
   assign m153_43 =10'b0;

   // m153_44 = W*in
   wire signed [9:0] m153_44;
   assign m153_44 =10'b0;

   // m153_45 = W*in
   wire signed [9:0] m153_45;
   assign m153_45 =10'b0;

   // m153_46 = W*in
   wire signed [9:0] m153_46;
   assign m153_46 =10'b0;

   // m153_47 = W*in
   wire signed [9:0] m153_47;
   assign m153_47 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_48 = W*in
   wire signed [9:0] m153_48;
   assign m153_48 =10'b0;

   // m153_49 = W*in
   wire signed [9:0] m153_49;
   assign m153_49 =10'b0;

   // m153_50 = W*in
   wire signed [9:0] m153_50;
   assign m153_50 =10'b0;

   // m153_51 = W*in
   wire signed [9:0] m153_51;
   assign m153_51 =10'b0;

   // m153_52 = W*in
   wire signed [9:0] m153_52;
   assign m153_52 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_53 = W*in
   wire signed [9:0] m153_53;
   assign m153_53 =10'b0;

   // m153_54 = W*in
   wire signed [9:0] m153_54;
   assign m153_54 =10'b0;

   // m153_55 = W*in
   wire signed [9:0] m153_55;
   assign m153_55 =10'b0;

   // m153_56 = W*in
   wire signed [9:0] m153_56;
   assign m153_56 ={ {4{in153[5]}} , in153[5:0] };

   // m153_57 = W*in
   wire signed [9:0] m153_57;
   assign m153_57 =10'b0;

   // m153_58 = W*in
   wire signed [9:0] m153_58;
   assign m153_58 =10'b0;

   // m153_59 = W*in
   wire signed [9:0] m153_59;
   assign m153_59 =10'b0;

   // m153_60 = W*in
   wire signed [9:0] m153_60;
   assign m153_60 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_61 = W*in
   wire signed [9:0] m153_61;
   assign m153_61 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_62 = W*in
   wire signed [9:0] m153_62;
   assign m153_62 =10'b0;

   // m153_63 = W*in
   wire signed [9:0] m153_63;
   assign m153_63 ={ {4{in153[5]}} , in153[5:0] };

   // m153_64 = W*in
   wire signed [9:0] m153_64;
   assign m153_64 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_65 = W*in
   wire signed [9:0] m153_65;
   assign m153_65 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_66 = W*in
   wire signed [9:0] m153_66;
   assign m153_66 =10'b0;

   // m153_67 = W*in
   wire signed [9:0] m153_67;
   assign m153_67 =10'b0;

   // m153_68 = W*in
   wire signed [9:0] m153_68;
   assign m153_68 =10'b0;

   // m153_69 = W*in
   wire signed [9:0] m153_69;
   assign m153_69 ={ {4{in153[5]}} , in153[5:0] };

   // m153_70 = W*in
   wire signed [9:0] m153_70;
   assign m153_70 =10'b0;

   // m153_71 = W*in
   wire signed [9:0] m153_71;
   assign m153_71 =10'b0;

   // m153_72 = W*in
   wire signed [9:0] m153_72;
   assign m153_72 ={ {4{in153[5]}} , in153[5:0] };

   // m153_73 = W*in
   wire signed [9:0] m153_73;
   assign m153_73 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_74 = W*in
   wire signed [9:0] m153_74;
   assign m153_74 =10'b0;

   // m153_75 = W*in
   wire signed [9:0] m153_75;
   assign m153_75 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_76 = W*in
   wire signed [9:0] m153_76;
   assign m153_76 =10'b0;

   // m153_77 = W*in
   wire signed [9:0] m153_77;
   assign m153_77 =10'b0;

   // m153_78 = W*in
   wire signed [9:0] m153_78;
   assign m153_78 ={ {4{in153[5]}} , in153[5:0] };

   // m153_79 = W*in
   wire signed [9:0] m153_79;
   assign m153_79 =10'b0;

   // m153_80 = W*in
   wire signed [9:0] m153_80;
   assign m153_80 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_81 = W*in
   wire signed [9:0] m153_81;
   assign m153_81 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_82 = W*in
   wire signed [9:0] m153_82;
   assign m153_82 =10'b0;

   // m153_83 = W*in
   wire signed [9:0] m153_83;
   assign m153_83 =10'b0;

   // m153_84 = W*in
   wire signed [9:0] m153_84;
   assign m153_84 ={ {4{in153[5]}} , in153[5:0] };

   // m153_85 = W*in
   wire signed [9:0] m153_85;
   assign m153_85 ={ {5{in153[5]}} , in153[5:1] };

   // m153_86 = W*in
   wire signed [9:0] m153_86;
   assign m153_86 ={ {4{in153[5]}} , in153[5:0] };

   // m153_87 = W*in
   wire signed [9:0] m153_87;
   assign m153_87 =10'b0;

   // m153_88 = W*in
   wire signed [9:0] m153_88;
   assign m153_88 =10'b0;

   // m153_89 = W*in
   wire signed [9:0] m153_89;
   assign m153_89 =10'b0;

   // m153_90 = W*in
   wire signed [9:0] m153_90;
   assign m153_90 =10'b0;

   // m153_91 = W*in
   wire signed [9:0] m153_91;
   assign m153_91 =10'b0;

   // m153_92 = W*in
   wire signed [9:0] m153_92;
   assign m153_92 =10'b0;

   // m153_93 = W*in
   wire signed [9:0] m153_93;
   assign m153_93 =10'b0;

   // m153_94 = W*in
   wire signed [9:0] m153_94;
   assign m153_94 =10'b0;

   // m153_95 = W*in
   wire signed [9:0] m153_95;
   assign m153_95 =10'b0;

   // m153_96 = W*in
   wire signed [9:0] m153_96;
   assign m153_96 =10'b0;

   // m153_97 = W*in
   wire signed [9:0] m153_97;
   assign m153_97 =10'b0;

   // m153_98 = W*in
   wire signed [9:0] m153_98;
   assign m153_98 =10'b0;

   // m153_99 = W*in
   wire signed [9:0] m153_99;
   assign m153_99 =10'b0;

   // m153_100 = W*in
   wire signed [9:0] m153_100;
   assign m153_100 =10'b0;

   // m153_101 = W*in
   wire signed [9:0] m153_101;
   assign m153_101 =10'b0;

   // m153_102 = W*in
   wire signed [9:0] m153_102;
   assign m153_102 =10'b0;

   // m153_103 = W*in
   wire signed [9:0] m153_103;
   assign m153_103 =10'b0;

   // m153_104 = W*in
   wire signed [9:0] m153_104;
   assign m153_104 =10'b0;

   // m153_105 = W*in
   wire signed [9:0] m153_105;
   assign m153_105 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_106 = W*in
   wire signed [9:0] m153_106;
   assign m153_106 =10'b0;

   // m153_107 = W*in
   wire signed [9:0] m153_107;
   assign m153_107 =10'b0;

   // m153_108 = W*in
   wire signed [9:0] m153_108;
   assign m153_108 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_109 = W*in
   wire signed [9:0] m153_109;
   assign m153_109 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_110 = W*in
   wire signed [9:0] m153_110;
   assign m153_110 =10'b0;

   // m153_111 = W*in
   wire signed [9:0] m153_111;
   assign m153_111 ={ {4{in153[5]}} , in153[5:0] };

   // m153_112 = W*in
   wire signed [9:0] m153_112;
   assign m153_112 =10'b0;

   // m153_113 = W*in
   wire signed [9:0] m153_113;
   assign m153_113 =10'b0;

   // m153_114 = W*in
   wire signed [9:0] m153_114;
   assign m153_114 ={ {5{neg153[5]}} , neg153[5:1] };

   // m153_115 = W*in
   wire signed [9:0] m153_115;
   assign m153_115 ={ {4{neg153[5]}} , neg153[5:0] };

   // m153_116 = W*in
   wire signed [9:0] m153_116;
   assign m153_116 =10'b0;

   // m153_117 = W*in
   wire signed [9:0] m153_117;
   assign m153_117 ={ {4{neg153[5]}} , neg153[5:0] };

   // m154_1 = W*in
   wire signed [9:0] m154_1;
   assign m154_1 =10'b0;

   // m154_2 = W*in
   wire signed [9:0] m154_2;
   assign m154_2 =10'b0;

   // m154_3 = W*in
   wire signed [9:0] m154_3;
   assign m154_3 =10'b0;

   // m154_4 = W*in
   wire signed [9:0] m154_4;
   assign m154_4 =10'b0;

   // m154_5 = W*in
   wire signed [9:0] m154_5;
   assign m154_5 ={ {4{in154[5]}} , in154[5:0] };

   // m154_6 = W*in
   wire signed [9:0] m154_6;
   assign m154_6 ={ {4{in154[5]}} , in154[5:0] };

   // m154_7 = W*in
   wire signed [9:0] m154_7;
   assign m154_7 =10'b0;

   // m154_8 = W*in
   wire signed [9:0] m154_8;
   assign m154_8 =10'b0;

   // m154_9 = W*in
   wire signed [9:0] m154_9;
   assign m154_9 =10'b0;

   // m154_10 = W*in
   wire signed [9:0] m154_10;
   assign m154_10 ={ {4{in154[5]}} , in154[5:0] };

   // m154_11 = W*in
   wire signed [9:0] m154_11;
   assign m154_11 =10'b0;

   // m154_12 = W*in
   wire signed [9:0] m154_12;
   assign m154_12 =10'b0;

   // m154_13 = W*in
   wire signed [9:0] m154_13;
   assign m154_13 =10'b0;

   // m154_14 = W*in
   wire signed [9:0] m154_14;
   assign m154_14 =10'b0;

   // m154_15 = W*in
   wire signed [9:0] m154_15;
   assign m154_15 =10'b0;

   // m154_16 = W*in
   wire signed [9:0] m154_16;
   assign m154_16 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_17 = W*in
   wire signed [9:0] m154_17;
   assign m154_17 =10'b0;

   // m154_18 = W*in
   wire signed [9:0] m154_18;
   assign m154_18 =10'b0;

   // m154_19 = W*in
   wire signed [9:0] m154_19;
   assign m154_19 =10'b0;

   // m154_20 = W*in
   wire signed [9:0] m154_20;
   assign m154_20 ={ {5{neg154[5]}} , neg154[5:1] };

   // m154_21 = W*in
   wire signed [9:0] m154_21;
   assign m154_21 ={ {5{in154[5]}} , in154[5:1] };

   // m154_22 = W*in
   wire signed [9:0] m154_22;
   assign m154_22 =10'b0;

   // m154_23 = W*in
   wire signed [9:0] m154_23;
   assign m154_23 ={ {4{in154[5]}} , in154[5:0] };

   // m154_24 = W*in
   wire signed [9:0] m154_24;
   assign m154_24 =10'b0;

   // m154_25 = W*in
   wire signed [9:0] m154_25;
   assign m154_25 =10'b0;

   // m154_26 = W*in
   wire signed [9:0] m154_26;
   assign m154_26 =10'b0;

   // m154_27 = W*in
   wire signed [9:0] m154_27;
   assign m154_27 =10'b0;

   // m154_28 = W*in
   wire signed [9:0] m154_28;
   assign m154_28 =10'b0;

   // m154_29 = W*in
   wire signed [9:0] m154_29;
   assign m154_29 =10'b0;

   // m154_30 = W*in
   wire signed [9:0] m154_30;
   assign m154_30 ={ {5{neg154[5]}} , neg154[5:1] };

   // m154_31 = W*in
   wire signed [9:0] m154_31;
   assign m154_31 =10'b0;

   // m154_32 = W*in
   wire signed [9:0] m154_32;
   assign m154_32 ={ {4{in154[5]}} , in154[5:0] };

   // m154_33 = W*in
   wire signed [9:0] m154_33;
   assign m154_33 =10'b0;

   // m154_34 = W*in
   wire signed [9:0] m154_34;
   assign m154_34 =10'b0;

   // m154_35 = W*in
   wire signed [9:0] m154_35;
   assign m154_35 ={ {5{neg154[5]}} , neg154[5:1] };

   // m154_36 = W*in
   wire signed [9:0] m154_36;
   assign m154_36 =10'b0;

   // m154_37 = W*in
   wire signed [9:0] m154_37;
   assign m154_37 =10'b0;

   // m154_38 = W*in
   wire signed [9:0] m154_38;
   assign m154_38 =10'b0;

   // m154_39 = W*in
   wire signed [9:0] m154_39;
   assign m154_39 =10'b0;

   // m154_40 = W*in
   wire signed [9:0] m154_40;
   assign m154_40 =10'b0;

   // m154_41 = W*in
   wire signed [9:0] m154_41;
   assign m154_41 =10'b0;

   // m154_42 = W*in
   wire signed [9:0] m154_42;
   assign m154_42 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_43 = W*in
   wire signed [9:0] m154_43;
   assign m154_43 =10'b0;

   // m154_44 = W*in
   wire signed [9:0] m154_44;
   assign m154_44 =10'b0;

   // m154_45 = W*in
   wire signed [9:0] m154_45;
   assign m154_45 =10'b0;

   // m154_46 = W*in
   wire signed [9:0] m154_46;
   assign m154_46 =10'b0;

   // m154_47 = W*in
   wire signed [9:0] m154_47;
   assign m154_47 =10'b0;

   // m154_48 = W*in
   wire signed [9:0] m154_48;
   assign m154_48 ={ {4{in154[5]}} , in154[5:0] };

   // m154_49 = W*in
   wire signed [9:0] m154_49;
   assign m154_49 =10'b0;

   // m154_50 = W*in
   wire signed [9:0] m154_50;
   assign m154_50 =10'b0;

   // m154_51 = W*in
   wire signed [9:0] m154_51;
   assign m154_51 =10'b0;

   // m154_52 = W*in
   wire signed [9:0] m154_52;
   assign m154_52 =10'b0;

   // m154_53 = W*in
   wire signed [9:0] m154_53;
   assign m154_53 ={ {4{in154[5]}} , in154[5:0] };

   // m154_54 = W*in
   wire signed [9:0] m154_54;
   assign m154_54 =10'b0;

   // m154_55 = W*in
   wire signed [9:0] m154_55;
   assign m154_55 =10'b0;

   // m154_56 = W*in
   wire signed [9:0] m154_56;
   assign m154_56 =10'b0;

   // m154_57 = W*in
   wire signed [9:0] m154_57;
   assign m154_57 =10'b0;

   // m154_58 = W*in
   wire signed [9:0] m154_58;
   assign m154_58 =10'b0;

   // m154_59 = W*in
   wire signed [9:0] m154_59;
   assign m154_59 =10'b0;

   // m154_60 = W*in
   wire signed [9:0] m154_60;
   assign m154_60 =10'b0;

   // m154_61 = W*in
   wire signed [9:0] m154_61;
   assign m154_61 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_62 = W*in
   wire signed [9:0] m154_62;
   assign m154_62 =10'b0;

   // m154_63 = W*in
   wire signed [9:0] m154_63;
   assign m154_63 =10'b0;

   // m154_64 = W*in
   wire signed [9:0] m154_64;
   assign m154_64 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_65 = W*in
   wire signed [9:0] m154_65;
   assign m154_65 ={ {5{neg154[5]}} , neg154[5:1] };

   // m154_66 = W*in
   wire signed [9:0] m154_66;
   assign m154_66 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_67 = W*in
   wire signed [9:0] m154_67;
   assign m154_67 ={ {4{in154[5]}} , in154[5:0] };

   // m154_68 = W*in
   wire signed [9:0] m154_68;
   assign m154_68 =10'b0;

   // m154_69 = W*in
   wire signed [9:0] m154_69;
   assign m154_69 ={ {4{in154[5]}} , in154[5:0] };

   // m154_70 = W*in
   wire signed [9:0] m154_70;
   assign m154_70 ={ {5{in154[5]}} , in154[5:1] };

   // m154_71 = W*in
   wire signed [9:0] m154_71;
   assign m154_71 =10'b0;

   // m154_72 = W*in
   wire signed [9:0] m154_72;
   assign m154_72 ={ {4{in154[5]}} , in154[5:0] };

   // m154_73 = W*in
   wire signed [9:0] m154_73;
   assign m154_73 =10'b0;

   // m154_74 = W*in
   wire signed [9:0] m154_74;
   assign m154_74 =10'b0;

   // m154_75 = W*in
   wire signed [9:0] m154_75;
   assign m154_75 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_76 = W*in
   wire signed [9:0] m154_76;
   assign m154_76 =10'b0;

   // m154_77 = W*in
   wire signed [9:0] m154_77;
   assign m154_77 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_78 = W*in
   wire signed [9:0] m154_78;
   assign m154_78 ={ {5{in154[5]}} , in154[5:1] };

   // m154_79 = W*in
   wire signed [9:0] m154_79;
   assign m154_79 =10'b0;

   // m154_80 = W*in
   wire signed [9:0] m154_80;
   assign m154_80 =10'b0;

   // m154_81 = W*in
   wire signed [9:0] m154_81;
   assign m154_81 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_82 = W*in
   wire signed [9:0] m154_82;
   assign m154_82 =10'b0;

   // m154_83 = W*in
   wire signed [9:0] m154_83;
   assign m154_83 =10'b0;

   // m154_84 = W*in
   wire signed [9:0] m154_84;
   assign m154_84 ={ {4{in154[5]}} , in154[5:0] };

   // m154_85 = W*in
   wire signed [9:0] m154_85;
   assign m154_85 ={ {4{in154[5]}} , in154[5:0] };

   // m154_86 = W*in
   wire signed [9:0] m154_86;
   assign m154_86 =10'b0;

   // m154_87 = W*in
   wire signed [9:0] m154_87;
   assign m154_87 =10'b0;

   // m154_88 = W*in
   wire signed [9:0] m154_88;
   assign m154_88 =10'b0;

   // m154_89 = W*in
   wire signed [9:0] m154_89;
   assign m154_89 =10'b0;

   // m154_90 = W*in
   wire signed [9:0] m154_90;
   assign m154_90 =10'b0;

   // m154_91 = W*in
   wire signed [9:0] m154_91;
   assign m154_91 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_92 = W*in
   wire signed [9:0] m154_92;
   assign m154_92 =10'b0;

   // m154_93 = W*in
   wire signed [9:0] m154_93;
   assign m154_93 ={ {4{in154[5]}} , in154[5:0] };

   // m154_94 = W*in
   wire signed [9:0] m154_94;
   assign m154_94 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_95 = W*in
   wire signed [9:0] m154_95;
   assign m154_95 =10'b0;

   // m154_96 = W*in
   wire signed [9:0] m154_96;
   assign m154_96 =10'b0;

   // m154_97 = W*in
   wire signed [9:0] m154_97;
   assign m154_97 =10'b0;

   // m154_98 = W*in
   wire signed [9:0] m154_98;
   assign m154_98 =10'b0;

   // m154_99 = W*in
   wire signed [9:0] m154_99;
   assign m154_99 =10'b0;

   // m154_100 = W*in
   wire signed [9:0] m154_100;
   assign m154_100 ={ {3{neg154[5]}} , neg154 , {1{1'b0}} };

   // m154_101 = W*in
   wire signed [9:0] m154_101;
   assign m154_101 =10'b0;

   // m154_102 = W*in
   wire signed [9:0] m154_102;
   assign m154_102 =10'b0;

   // m154_103 = W*in
   wire signed [9:0] m154_103;
   assign m154_103 =10'b0;

   // m154_104 = W*in
   wire signed [9:0] m154_104;
   assign m154_104 =10'b0;

   // m154_105 = W*in
   wire signed [9:0] m154_105;
   assign m154_105 =10'b0;

   // m154_106 = W*in
   wire signed [9:0] m154_106;
   assign m154_106 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_107 = W*in
   wire signed [9:0] m154_107;
   assign m154_107 =10'b0;

   // m154_108 = W*in
   wire signed [9:0] m154_108;
   assign m154_108 ={ {5{neg154[5]}} , neg154[5:1] };

   // m154_109 = W*in
   wire signed [9:0] m154_109;
   assign m154_109 =10'b0;

   // m154_110 = W*in
   wire signed [9:0] m154_110;
   assign m154_110 =10'b0;

   // m154_111 = W*in
   wire signed [9:0] m154_111;
   assign m154_111 ={ {4{in154[5]}} , in154[5:0] };

   // m154_112 = W*in
   wire signed [9:0] m154_112;
   assign m154_112 ={ {4{neg154[5]}} , neg154[5:0] };

   // m154_113 = W*in
   wire signed [9:0] m154_113;
   assign m154_113 =10'b0;

   // m154_114 = W*in
   wire signed [9:0] m154_114;
   assign m154_114 =10'b0;

   // m154_115 = W*in
   wire signed [9:0] m154_115;
   assign m154_115 ={ {5{neg154[5]}} , neg154[5:1] };

   // m154_116 = W*in
   wire signed [9:0] m154_116;
   assign m154_116 =10'b0;

   // m154_117 = W*in
   wire signed [9:0] m154_117;
   assign m154_117 =10'b0;

   // m155_1 = W*in
   wire signed [9:0] m155_1;
   assign m155_1 =10'b0;

   // m155_2 = W*in
   wire signed [9:0] m155_2;
   assign m155_2 =10'b0;

   // m155_3 = W*in
   wire signed [9:0] m155_3;
   assign m155_3 =10'b0;

   // m155_4 = W*in
   wire signed [9:0] m155_4;
   assign m155_4 =10'b0;

   // m155_5 = W*in
   wire signed [9:0] m155_5;
   assign m155_5 =10'b0;

   // m155_6 = W*in
   wire signed [9:0] m155_6;
   assign m155_6 =10'b0;

   // m155_7 = W*in
   wire signed [9:0] m155_7;
   assign m155_7 =10'b0;

   // m155_8 = W*in
   wire signed [9:0] m155_8;
   assign m155_8 =10'b0;

   // m155_9 = W*in
   wire signed [9:0] m155_9;
   assign m155_9 =10'b0;

   // m155_10 = W*in
   wire signed [9:0] m155_10;
   assign m155_10 =10'b0;

   // m155_11 = W*in
   wire signed [9:0] m155_11;
   assign m155_11 =10'b0;

   // m155_12 = W*in
   wire signed [9:0] m155_12;
   assign m155_12 =10'b0;

   // m155_13 = W*in
   wire signed [9:0] m155_13;
   assign m155_13 =10'b0;

   // m155_14 = W*in
   wire signed [9:0] m155_14;
   assign m155_14 =10'b0;

   // m155_15 = W*in
   wire signed [9:0] m155_15;
   assign m155_15 =10'b0;

   // m155_16 = W*in
   wire signed [9:0] m155_16;
   assign m155_16 =10'b0;

   // m155_17 = W*in
   wire signed [9:0] m155_17;
   assign m155_17 =10'b0;

   // m155_18 = W*in
   wire signed [9:0] m155_18;
   assign m155_18 ={ {5{neg155[5]}} , neg155[5:1] };

   // m155_19 = W*in
   wire signed [9:0] m155_19;
   assign m155_19 =10'b0;

   // m155_20 = W*in
   wire signed [9:0] m155_20;
   assign m155_20 =10'b0;

   // m155_21 = W*in
   wire signed [9:0] m155_21;
   assign m155_21 ={ {5{in155[5]}} , in155[5:1] };

   // m155_22 = W*in
   wire signed [9:0] m155_22;
   assign m155_22 =10'b0;

   // m155_23 = W*in
   wire signed [9:0] m155_23;
   assign m155_23 ={ {5{in155[5]}} , in155[5:1] };

   // m155_24 = W*in
   wire signed [9:0] m155_24;
   assign m155_24 =10'b0;

   // m155_25 = W*in
   wire signed [9:0] m155_25;
   assign m155_25 =10'b0;

   // m155_26 = W*in
   wire signed [9:0] m155_26;
   assign m155_26 =10'b0;

   // m155_27 = W*in
   wire signed [9:0] m155_27;
   assign m155_27 =10'b0;

   // m155_28 = W*in
   wire signed [9:0] m155_28;
   assign m155_28 =10'b0;

   // m155_29 = W*in
   wire signed [9:0] m155_29;
   assign m155_29 =10'b0;

   // m155_30 = W*in
   wire signed [9:0] m155_30;
   assign m155_30 ={ {5{neg155[5]}} , neg155[5:1] };

   // m155_31 = W*in
   wire signed [9:0] m155_31;
   assign m155_31 =10'b0;

   // m155_32 = W*in
   wire signed [9:0] m155_32;
   assign m155_32 =10'b0;

   // m155_33 = W*in
   wire signed [9:0] m155_33;
   assign m155_33 =10'b0;

   // m155_34 = W*in
   wire signed [9:0] m155_34;
   assign m155_34 =10'b0;

   // m155_35 = W*in
   wire signed [9:0] m155_35;
   assign m155_35 =10'b0;

   // m155_36 = W*in
   wire signed [9:0] m155_36;
   assign m155_36 =10'b0;

   // m155_37 = W*in
   wire signed [9:0] m155_37;
   assign m155_37 =10'b0;

   // m155_38 = W*in
   wire signed [9:0] m155_38;
   assign m155_38 =10'b0;

   // m155_39 = W*in
   wire signed [9:0] m155_39;
   assign m155_39 =10'b0;

   // m155_40 = W*in
   wire signed [9:0] m155_40;
   assign m155_40 =10'b0;

   // m155_41 = W*in
   wire signed [9:0] m155_41;
   assign m155_41 =10'b0;

   // m155_42 = W*in
   wire signed [9:0] m155_42;
   assign m155_42 ={ {4{neg155[5]}} , neg155[5:0] };

   // m155_43 = W*in
   wire signed [9:0] m155_43;
   assign m155_43 =10'b0;

   // m155_44 = W*in
   wire signed [9:0] m155_44;
   assign m155_44 =10'b0;

   // m155_45 = W*in
   wire signed [9:0] m155_45;
   assign m155_45 =10'b0;

   // m155_46 = W*in
   wire signed [9:0] m155_46;
   assign m155_46 =10'b0;

   // m155_47 = W*in
   wire signed [9:0] m155_47;
   assign m155_47 =10'b0;

   // m155_48 = W*in
   wire signed [9:0] m155_48;
   assign m155_48 =10'b0;

   // m155_49 = W*in
   wire signed [9:0] m155_49;
   assign m155_49 =10'b0;

   // m155_50 = W*in
   wire signed [9:0] m155_50;
   assign m155_50 =10'b0;

   // m155_51 = W*in
   wire signed [9:0] m155_51;
   assign m155_51 =10'b0;

   // m155_52 = W*in
   wire signed [9:0] m155_52;
   assign m155_52 =10'b0;

   // m155_53 = W*in
   wire signed [9:0] m155_53;
   assign m155_53 =10'b0;

   // m155_54 = W*in
   wire signed [9:0] m155_54;
   assign m155_54 =10'b0;

   // m155_55 = W*in
   wire signed [9:0] m155_55;
   assign m155_55 =10'b0;

   // m155_56 = W*in
   wire signed [9:0] m155_56;
   assign m155_56 ={ {4{neg155[5]}} , neg155[5:0] };

   // m155_57 = W*in
   wire signed [9:0] m155_57;
   assign m155_57 =10'b0;

   // m155_58 = W*in
   wire signed [9:0] m155_58;
   assign m155_58 =10'b0;

   // m155_59 = W*in
   wire signed [9:0] m155_59;
   assign m155_59 =10'b0;

   // m155_60 = W*in
   wire signed [9:0] m155_60;
   assign m155_60 =10'b0;

   // m155_61 = W*in
   wire signed [9:0] m155_61;
   assign m155_61 ={ {4{neg155[5]}} , neg155[5:0] };

   // m155_62 = W*in
   wire signed [9:0] m155_62;
   assign m155_62 =10'b0;

   // m155_63 = W*in
   wire signed [9:0] m155_63;
   assign m155_63 =10'b0;

   // m155_64 = W*in
   wire signed [9:0] m155_64;
   assign m155_64 ={ {5{neg155[5]}} , neg155[5:1] };

   // m155_65 = W*in
   wire signed [9:0] m155_65;
   assign m155_65 =10'b0;

   // m155_66 = W*in
   wire signed [9:0] m155_66;
   assign m155_66 ={ {5{neg155[5]}} , neg155[5:1] };

   // m155_67 = W*in
   wire signed [9:0] m155_67;
   assign m155_67 ={ {4{in155[5]}} , in155[5:0] };

   // m155_68 = W*in
   wire signed [9:0] m155_68;
   assign m155_68 =10'b0;

   // m155_69 = W*in
   wire signed [9:0] m155_69;
   assign m155_69 =10'b0;

   // m155_70 = W*in
   wire signed [9:0] m155_70;
   assign m155_70 ={ {5{in155[5]}} , in155[5:1] };

   // m155_71 = W*in
   wire signed [9:0] m155_71;
   assign m155_71 =10'b0;

   // m155_72 = W*in
   wire signed [9:0] m155_72;
   assign m155_72 =10'b0;

   // m155_73 = W*in
   wire signed [9:0] m155_73;
   assign m155_73 =10'b0;

   // m155_74 = W*in
   wire signed [9:0] m155_74;
   assign m155_74 =10'b0;

   // m155_75 = W*in
   wire signed [9:0] m155_75;
   assign m155_75 ={ {5{neg155[5]}} , neg155[5:1] };

   // m155_76 = W*in
   wire signed [9:0] m155_76;
   assign m155_76 =10'b0;

   // m155_77 = W*in
   wire signed [9:0] m155_77;
   assign m155_77 =10'b0;

   // m155_78 = W*in
   wire signed [9:0] m155_78;
   assign m155_78 =10'b0;

   // m155_79 = W*in
   wire signed [9:0] m155_79;
   assign m155_79 =10'b0;

   // m155_80 = W*in
   wire signed [9:0] m155_80;
   assign m155_80 =10'b0;

   // m155_81 = W*in
   wire signed [9:0] m155_81;
   assign m155_81 ={ {5{neg155[5]}} , neg155[5:1] };

   // m155_82 = W*in
   wire signed [9:0] m155_82;
   assign m155_82 =10'b0;

   // m155_83 = W*in
   wire signed [9:0] m155_83;
   assign m155_83 =10'b0;

   // m155_84 = W*in
   wire signed [9:0] m155_84;
   assign m155_84 =10'b0;

   // m155_85 = W*in
   wire signed [9:0] m155_85;
   assign m155_85 =10'b0;

   // m155_86 = W*in
   wire signed [9:0] m155_86;
   assign m155_86 =10'b0;

   // m155_87 = W*in
   wire signed [9:0] m155_87;
   assign m155_87 =10'b0;

   // m155_88 = W*in
   wire signed [9:0] m155_88;
   assign m155_88 =10'b0;

   // m155_89 = W*in
   wire signed [9:0] m155_89;
   assign m155_89 =10'b0;

   // m155_90 = W*in
   wire signed [9:0] m155_90;
   assign m155_90 =10'b0;

   // m155_91 = W*in
   wire signed [9:0] m155_91;
   assign m155_91 =10'b0;

   // m155_92 = W*in
   wire signed [9:0] m155_92;
   assign m155_92 =10'b0;

   // m155_93 = W*in
   wire signed [9:0] m155_93;
   assign m155_93 ={ {4{in155[5]}} , in155[5:0] };

   // m155_94 = W*in
   wire signed [9:0] m155_94;
   assign m155_94 ={ {4{neg155[5]}} , neg155[5:0] };

   // m155_95 = W*in
   wire signed [9:0] m155_95;
   assign m155_95 =10'b0;

   // m155_96 = W*in
   wire signed [9:0] m155_96;
   assign m155_96 =10'b0;

   // m155_97 = W*in
   wire signed [9:0] m155_97;
   assign m155_97 =10'b0;

   // m155_98 = W*in
   wire signed [9:0] m155_98;
   assign m155_98 =10'b0;

   // m155_99 = W*in
   wire signed [9:0] m155_99;
   assign m155_99 =10'b0;

   // m155_100 = W*in
   wire signed [9:0] m155_100;
   assign m155_100 ={ {4{neg155[5]}} , neg155[5:0] };

   // m155_101 = W*in
   wire signed [9:0] m155_101;
   assign m155_101 =10'b0;

   // m155_102 = W*in
   wire signed [9:0] m155_102;
   assign m155_102 =10'b0;

   // m155_103 = W*in
   wire signed [9:0] m155_103;
   assign m155_103 =10'b0;

   // m155_104 = W*in
   wire signed [9:0] m155_104;
   assign m155_104 =10'b0;

   // m155_105 = W*in
   wire signed [9:0] m155_105;
   assign m155_105 =10'b0;

   // m155_106 = W*in
   wire signed [9:0] m155_106;
   assign m155_106 =10'b0;

   // m155_107 = W*in
   wire signed [9:0] m155_107;
   assign m155_107 =10'b0;

   // m155_108 = W*in
   wire signed [9:0] m155_108;
   assign m155_108 =10'b0;

   // m155_109 = W*in
   wire signed [9:0] m155_109;
   assign m155_109 ={ {5{in155[5]}} , in155[5:1] };

   // m155_110 = W*in
   wire signed [9:0] m155_110;
   assign m155_110 =10'b0;

   // m155_111 = W*in
   wire signed [9:0] m155_111;
   assign m155_111 =10'b0;

   // m155_112 = W*in
   wire signed [9:0] m155_112;
   assign m155_112 =10'b0;

   // m155_113 = W*in
   wire signed [9:0] m155_113;
   assign m155_113 =10'b0;

   // m155_114 = W*in
   wire signed [9:0] m155_114;
   assign m155_114 =10'b0;

   // m155_115 = W*in
   wire signed [9:0] m155_115;
   assign m155_115 =10'b0;

   // m155_116 = W*in
   wire signed [9:0] m155_116;
   assign m155_116 =10'b0;

   // m155_117 = W*in
   wire signed [9:0] m155_117;
   assign m155_117 =10'b0;

   // m156_1 = W*in
   wire signed [9:0] m156_1;
   assign m156_1 =10'b0;

   // m156_2 = W*in
   wire signed [9:0] m156_2;
   assign m156_2 =10'b0;

   // m156_3 = W*in
   wire signed [9:0] m156_3;
   assign m156_3 =10'b0;

   // m156_4 = W*in
   wire signed [9:0] m156_4;
   assign m156_4 =10'b0;

   // m156_5 = W*in
   wire signed [9:0] m156_5;
   assign m156_5 =10'b0;

   // m156_6 = W*in
   wire signed [9:0] m156_6;
   assign m156_6 =10'b0;

   // m156_7 = W*in
   wire signed [9:0] m156_7;
   assign m156_7 =10'b0;

   // m156_8 = W*in
   wire signed [9:0] m156_8;
   assign m156_8 =10'b0;

   // m156_9 = W*in
   wire signed [9:0] m156_9;
   assign m156_9 =10'b0;

   // m156_10 = W*in
   wire signed [9:0] m156_10;
   assign m156_10 =10'b0;

   // m156_11 = W*in
   wire signed [9:0] m156_11;
   assign m156_11 =10'b0;

   // m156_12 = W*in
   wire signed [9:0] m156_12;
   assign m156_12 =10'b0;

   // m156_13 = W*in
   wire signed [9:0] m156_13;
   assign m156_13 =10'b0;

   // m156_14 = W*in
   wire signed [9:0] m156_14;
   assign m156_14 =10'b0;

   // m156_15 = W*in
   wire signed [9:0] m156_15;
   assign m156_15 =10'b0;

   // m156_16 = W*in
   wire signed [9:0] m156_16;
   assign m156_16 =10'b0;

   // m156_17 = W*in
   wire signed [9:0] m156_17;
   assign m156_17 =10'b0;

   // m156_18 = W*in
   wire signed [9:0] m156_18;
   assign m156_18 =10'b0;

   // m156_19 = W*in
   wire signed [9:0] m156_19;
   assign m156_19 =10'b0;

   // m156_20 = W*in
   wire signed [9:0] m156_20;
   assign m156_20 =10'b0;

   // m156_21 = W*in
   wire signed [9:0] m156_21;
   assign m156_21 =10'b0;

   // m156_22 = W*in
   wire signed [9:0] m156_22;
   assign m156_22 =10'b0;

   // m156_23 = W*in
   wire signed [9:0] m156_23;
   assign m156_23 ={ {5{in156[5]}} , in156[5:1] };

   // m156_24 = W*in
   wire signed [9:0] m156_24;
   assign m156_24 =10'b0;

   // m156_25 = W*in
   wire signed [9:0] m156_25;
   assign m156_25 =10'b0;

   // m156_26 = W*in
   wire signed [9:0] m156_26;
   assign m156_26 =10'b0;

   // m156_27 = W*in
   wire signed [9:0] m156_27;
   assign m156_27 =10'b0;

   // m156_28 = W*in
   wire signed [9:0] m156_28;
   assign m156_28 =10'b0;

   // m156_29 = W*in
   wire signed [9:0] m156_29;
   assign m156_29 =10'b0;

   // m156_30 = W*in
   wire signed [9:0] m156_30;
   assign m156_30 =10'b0;

   // m156_31 = W*in
   wire signed [9:0] m156_31;
   assign m156_31 =10'b0;

   // m156_32 = W*in
   wire signed [9:0] m156_32;
   assign m156_32 =10'b0;

   // m156_33 = W*in
   wire signed [9:0] m156_33;
   assign m156_33 =10'b0;

   // m156_34 = W*in
   wire signed [9:0] m156_34;
   assign m156_34 =10'b0;

   // m156_35 = W*in
   wire signed [9:0] m156_35;
   assign m156_35 =10'b0;

   // m156_36 = W*in
   wire signed [9:0] m156_36;
   assign m156_36 =10'b0;

   // m156_37 = W*in
   wire signed [9:0] m156_37;
   assign m156_37 =10'b0;

   // m156_38 = W*in
   wire signed [9:0] m156_38;
   assign m156_38 =10'b0;

   // m156_39 = W*in
   wire signed [9:0] m156_39;
   assign m156_39 =10'b0;

   // m156_40 = W*in
   wire signed [9:0] m156_40;
   assign m156_40 =10'b0;

   // m156_41 = W*in
   wire signed [9:0] m156_41;
   assign m156_41 =10'b0;

   // m156_42 = W*in
   wire signed [9:0] m156_42;
   assign m156_42 =10'b0;

   // m156_43 = W*in
   wire signed [9:0] m156_43;
   assign m156_43 =10'b0;

   // m156_44 = W*in
   wire signed [9:0] m156_44;
   assign m156_44 =10'b0;

   // m156_45 = W*in
   wire signed [9:0] m156_45;
   assign m156_45 =10'b0;

   // m156_46 = W*in
   wire signed [9:0] m156_46;
   assign m156_46 =10'b0;

   // m156_47 = W*in
   wire signed [9:0] m156_47;
   assign m156_47 =10'b0;

   // m156_48 = W*in
   wire signed [9:0] m156_48;
   assign m156_48 =10'b0;

   // m156_49 = W*in
   wire signed [9:0] m156_49;
   assign m156_49 =10'b0;

   // m156_50 = W*in
   wire signed [9:0] m156_50;
   assign m156_50 =10'b0;

   // m156_51 = W*in
   wire signed [9:0] m156_51;
   assign m156_51 =10'b0;

   // m156_52 = W*in
   wire signed [9:0] m156_52;
   assign m156_52 =10'b0;

   // m156_53 = W*in
   wire signed [9:0] m156_53;
   assign m156_53 =10'b0;

   // m156_54 = W*in
   wire signed [9:0] m156_54;
   assign m156_54 =10'b0;

   // m156_55 = W*in
   wire signed [9:0] m156_55;
   assign m156_55 =10'b0;

   // m156_56 = W*in
   wire signed [9:0] m156_56;
   assign m156_56 =10'b0;

   // m156_57 = W*in
   wire signed [9:0] m156_57;
   assign m156_57 =10'b0;

   // m156_58 = W*in
   wire signed [9:0] m156_58;
   assign m156_58 =10'b0;

   // m156_59 = W*in
   wire signed [9:0] m156_59;
   assign m156_59 =10'b0;

   // m156_60 = W*in
   wire signed [9:0] m156_60;
   assign m156_60 =10'b0;

   // m156_61 = W*in
   wire signed [9:0] m156_61;
   assign m156_61 =10'b0;

   // m156_62 = W*in
   wire signed [9:0] m156_62;
   assign m156_62 =10'b0;

   // m156_63 = W*in
   wire signed [9:0] m156_63;
   assign m156_63 =10'b0;

   // m156_64 = W*in
   wire signed [9:0] m156_64;
   assign m156_64 =10'b0;

   // m156_65 = W*in
   wire signed [9:0] m156_65;
   assign m156_65 =10'b0;

   // m156_66 = W*in
   wire signed [9:0] m156_66;
   assign m156_66 =10'b0;

   // m156_67 = W*in
   wire signed [9:0] m156_67;
   assign m156_67 =10'b0;

   // m156_68 = W*in
   wire signed [9:0] m156_68;
   assign m156_68 =10'b0;

   // m156_69 = W*in
   wire signed [9:0] m156_69;
   assign m156_69 =10'b0;

   // m156_70 = W*in
   wire signed [9:0] m156_70;
   assign m156_70 =10'b0;

   // m156_71 = W*in
   wire signed [9:0] m156_71;
   assign m156_71 =10'b0;

   // m156_72 = W*in
   wire signed [9:0] m156_72;
   assign m156_72 =10'b0;

   // m156_73 = W*in
   wire signed [9:0] m156_73;
   assign m156_73 =10'b0;

   // m156_74 = W*in
   wire signed [9:0] m156_74;
   assign m156_74 =10'b0;

   // m156_75 = W*in
   wire signed [9:0] m156_75;
   assign m156_75 =10'b0;

   // m156_76 = W*in
   wire signed [9:0] m156_76;
   assign m156_76 =10'b0;

   // m156_77 = W*in
   wire signed [9:0] m156_77;
   assign m156_77 =10'b0;

   // m156_78 = W*in
   wire signed [9:0] m156_78;
   assign m156_78 =10'b0;

   // m156_79 = W*in
   wire signed [9:0] m156_79;
   assign m156_79 =10'b0;

   // m156_80 = W*in
   wire signed [9:0] m156_80;
   assign m156_80 =10'b0;

   // m156_81 = W*in
   wire signed [9:0] m156_81;
   assign m156_81 =10'b0;

   // m156_82 = W*in
   wire signed [9:0] m156_82;
   assign m156_82 =10'b0;

   // m156_83 = W*in
   wire signed [9:0] m156_83;
   assign m156_83 =10'b0;

   // m156_84 = W*in
   wire signed [9:0] m156_84;
   assign m156_84 =10'b0;

   // m156_85 = W*in
   wire signed [9:0] m156_85;
   assign m156_85 =10'b0;

   // m156_86 = W*in
   wire signed [9:0] m156_86;
   assign m156_86 =10'b0;

   // m156_87 = W*in
   wire signed [9:0] m156_87;
   assign m156_87 =10'b0;

   // m156_88 = W*in
   wire signed [9:0] m156_88;
   assign m156_88 =10'b0;

   // m156_89 = W*in
   wire signed [9:0] m156_89;
   assign m156_89 =10'b0;

   // m156_90 = W*in
   wire signed [9:0] m156_90;
   assign m156_90 =10'b0;

   // m156_91 = W*in
   wire signed [9:0] m156_91;
   assign m156_91 =10'b0;

   // m156_92 = W*in
   wire signed [9:0] m156_92;
   assign m156_92 =10'b0;

   // m156_93 = W*in
   wire signed [9:0] m156_93;
   assign m156_93 =10'b0;

   // m156_94 = W*in
   wire signed [9:0] m156_94;
   assign m156_94 =10'b0;

   // m156_95 = W*in
   wire signed [9:0] m156_95;
   assign m156_95 =10'b0;

   // m156_96 = W*in
   wire signed [9:0] m156_96;
   assign m156_96 =10'b0;

   // m156_97 = W*in
   wire signed [9:0] m156_97;
   assign m156_97 =10'b0;

   // m156_98 = W*in
   wire signed [9:0] m156_98;
   assign m156_98 =10'b0;

   // m156_99 = W*in
   wire signed [9:0] m156_99;
   assign m156_99 =10'b0;

   // m156_100 = W*in
   wire signed [9:0] m156_100;
   assign m156_100 =10'b0;

   // m156_101 = W*in
   wire signed [9:0] m156_101;
   assign m156_101 =10'b0;

   // m156_102 = W*in
   wire signed [9:0] m156_102;
   assign m156_102 =10'b0;

   // m156_103 = W*in
   wire signed [9:0] m156_103;
   assign m156_103 =10'b0;

   // m156_104 = W*in
   wire signed [9:0] m156_104;
   assign m156_104 =10'b0;

   // m156_105 = W*in
   wire signed [9:0] m156_105;
   assign m156_105 =10'b0;

   // m156_106 = W*in
   wire signed [9:0] m156_106;
   assign m156_106 =10'b0;

   // m156_107 = W*in
   wire signed [9:0] m156_107;
   assign m156_107 =10'b0;

   // m156_108 = W*in
   wire signed [9:0] m156_108;
   assign m156_108 =10'b0;

   // m156_109 = W*in
   wire signed [9:0] m156_109;
   assign m156_109 =10'b0;

   // m156_110 = W*in
   wire signed [9:0] m156_110;
   assign m156_110 =10'b0;

   // m156_111 = W*in
   wire signed [9:0] m156_111;
   assign m156_111 =10'b0;

   // m156_112 = W*in
   wire signed [9:0] m156_112;
   assign m156_112 =10'b0;

   // m156_113 = W*in
   wire signed [9:0] m156_113;
   assign m156_113 =10'b0;

   // m156_114 = W*in
   wire signed [9:0] m156_114;
   assign m156_114 =10'b0;

   // m156_115 = W*in
   wire signed [9:0] m156_115;
   assign m156_115 =10'b0;

   // m156_116 = W*in
   wire signed [9:0] m156_116;
   assign m156_116 =10'b0;

   // m156_117 = W*in
   wire signed [9:0] m156_117;
   assign m156_117 =10'b0;

   // m157_1 = W*in
   wire signed [9:0] m157_1;
   assign m157_1 =10'b0;

   // m157_2 = W*in
   wire signed [9:0] m157_2;
   assign m157_2 =10'b0;

   // m157_3 = W*in
   wire signed [9:0] m157_3;
   assign m157_3 =10'b0;

   // m157_4 = W*in
   wire signed [9:0] m157_4;
   assign m157_4 =10'b0;

   // m157_5 = W*in
   wire signed [9:0] m157_5;
   assign m157_5 =10'b0;

   // m157_6 = W*in
   wire signed [9:0] m157_6;
   assign m157_6 =10'b0;

   // m157_7 = W*in
   wire signed [9:0] m157_7;
   assign m157_7 =10'b0;

   // m157_8 = W*in
   wire signed [9:0] m157_8;
   assign m157_8 =10'b0;

   // m157_9 = W*in
   wire signed [9:0] m157_9;
   assign m157_9 =10'b0;

   // m157_10 = W*in
   wire signed [9:0] m157_10;
   assign m157_10 =10'b0;

   // m157_11 = W*in
   wire signed [9:0] m157_11;
   assign m157_11 =10'b0;

   // m157_12 = W*in
   wire signed [9:0] m157_12;
   assign m157_12 =10'b0;

   // m157_13 = W*in
   wire signed [9:0] m157_13;
   assign m157_13 =10'b0;

   // m157_14 = W*in
   wire signed [9:0] m157_14;
   assign m157_14 =10'b0;

   // m157_15 = W*in
   wire signed [9:0] m157_15;
   assign m157_15 =10'b0;

   // m157_16 = W*in
   wire signed [9:0] m157_16;
   assign m157_16 =10'b0;

   // m157_17 = W*in
   wire signed [9:0] m157_17;
   assign m157_17 ={ {5{neg157[5]}} , neg157[5:1] };

   // m157_18 = W*in
   wire signed [9:0] m157_18;
   assign m157_18 =10'b0;

   // m157_19 = W*in
   wire signed [9:0] m157_19;
   assign m157_19 =10'b0;

   // m157_20 = W*in
   wire signed [9:0] m157_20;
   assign m157_20 =10'b0;

   // m157_21 = W*in
   wire signed [9:0] m157_21;
   assign m157_21 ={ {5{neg157[5]}} , neg157[5:1] };

   // m157_22 = W*in
   wire signed [9:0] m157_22;
   assign m157_22 =10'b0;

   // m157_23 = W*in
   wire signed [9:0] m157_23;
   assign m157_23 =10'b0;

   // m157_24 = W*in
   wire signed [9:0] m157_24;
   assign m157_24 =10'b0;

   // m157_25 = W*in
   wire signed [9:0] m157_25;
   assign m157_25 =10'b0;

   // m157_26 = W*in
   wire signed [9:0] m157_26;
   assign m157_26 ={ {5{in157[5]}} , in157[5:1] };

   // m157_27 = W*in
   wire signed [9:0] m157_27;
   assign m157_27 =10'b0;

   // m157_28 = W*in
   wire signed [9:0] m157_28;
   assign m157_28 =10'b0;

   // m157_29 = W*in
   wire signed [9:0] m157_29;
   assign m157_29 =10'b0;

   // m157_30 = W*in
   wire signed [9:0] m157_30;
   assign m157_30 =10'b0;

   // m157_31 = W*in
   wire signed [9:0] m157_31;
   assign m157_31 =10'b0;

   // m157_32 = W*in
   wire signed [9:0] m157_32;
   assign m157_32 =10'b0;

   // m157_33 = W*in
   wire signed [9:0] m157_33;
   assign m157_33 =10'b0;

   // m157_34 = W*in
   wire signed [9:0] m157_34;
   assign m157_34 =10'b0;

   // m157_35 = W*in
   wire signed [9:0] m157_35;
   assign m157_35 =10'b0;

   // m157_36 = W*in
   wire signed [9:0] m157_36;
   assign m157_36 ={ {5{neg157[5]}} , neg157[5:1] };

   // m157_37 = W*in
   wire signed [9:0] m157_37;
   assign m157_37 =10'b0;

   // m157_38 = W*in
   wire signed [9:0] m157_38;
   assign m157_38 =10'b0;

   // m157_39 = W*in
   wire signed [9:0] m157_39;
   assign m157_39 =10'b0;

   // m157_40 = W*in
   wire signed [9:0] m157_40;
   assign m157_40 =10'b0;

   // m157_41 = W*in
   wire signed [9:0] m157_41;
   assign m157_41 =10'b0;

   // m157_42 = W*in
   wire signed [9:0] m157_42;
   assign m157_42 =10'b0;

   // m157_43 = W*in
   wire signed [9:0] m157_43;
   assign m157_43 =10'b0;

   // m157_44 = W*in
   wire signed [9:0] m157_44;
   assign m157_44 =10'b0;

   // m157_45 = W*in
   wire signed [9:0] m157_45;
   assign m157_45 =10'b0;

   // m157_46 = W*in
   wire signed [9:0] m157_46;
   assign m157_46 =10'b0;

   // m157_47 = W*in
   wire signed [9:0] m157_47;
   assign m157_47 =10'b0;

   // m157_48 = W*in
   wire signed [9:0] m157_48;
   assign m157_48 =10'b0;

   // m157_49 = W*in
   wire signed [9:0] m157_49;
   assign m157_49 =10'b0;

   // m157_50 = W*in
   wire signed [9:0] m157_50;
   assign m157_50 =10'b0;

   // m157_51 = W*in
   wire signed [9:0] m157_51;
   assign m157_51 =10'b0;

   // m157_52 = W*in
   wire signed [9:0] m157_52;
   assign m157_52 =10'b0;

   // m157_53 = W*in
   wire signed [9:0] m157_53;
   assign m157_53 =10'b0;

   // m157_54 = W*in
   wire signed [9:0] m157_54;
   assign m157_54 =10'b0;

   // m157_55 = W*in
   wire signed [9:0] m157_55;
   assign m157_55 =10'b0;

   // m157_56 = W*in
   wire signed [9:0] m157_56;
   assign m157_56 =10'b0;

   // m157_57 = W*in
   wire signed [9:0] m157_57;
   assign m157_57 =10'b0;

   // m157_58 = W*in
   wire signed [9:0] m157_58;
   assign m157_58 =10'b0;

   // m157_59 = W*in
   wire signed [9:0] m157_59;
   assign m157_59 =10'b0;

   // m157_60 = W*in
   wire signed [9:0] m157_60;
   assign m157_60 =10'b0;

   // m157_61 = W*in
   wire signed [9:0] m157_61;
   assign m157_61 =10'b0;

   // m157_62 = W*in
   wire signed [9:0] m157_62;
   assign m157_62 =10'b0;

   // m157_63 = W*in
   wire signed [9:0] m157_63;
   assign m157_63 =10'b0;

   // m157_64 = W*in
   wire signed [9:0] m157_64;
   assign m157_64 =10'b0;

   // m157_65 = W*in
   wire signed [9:0] m157_65;
   assign m157_65 =10'b0;

   // m157_66 = W*in
   wire signed [9:0] m157_66;
   assign m157_66 =10'b0;

   // m157_67 = W*in
   wire signed [9:0] m157_67;
   assign m157_67 =10'b0;

   // m157_68 = W*in
   wire signed [9:0] m157_68;
   assign m157_68 =10'b0;

   // m157_69 = W*in
   wire signed [9:0] m157_69;
   assign m157_69 =10'b0;

   // m157_70 = W*in
   wire signed [9:0] m157_70;
   assign m157_70 =10'b0;

   // m157_71 = W*in
   wire signed [9:0] m157_71;
   assign m157_71 =10'b0;

   // m157_72 = W*in
   wire signed [9:0] m157_72;
   assign m157_72 ={ {5{in157[5]}} , in157[5:1] };

   // m157_73 = W*in
   wire signed [9:0] m157_73;
   assign m157_73 =10'b0;

   // m157_74 = W*in
   wire signed [9:0] m157_74;
   assign m157_74 =10'b0;

   // m157_75 = W*in
   wire signed [9:0] m157_75;
   assign m157_75 =10'b0;

   // m157_76 = W*in
   wire signed [9:0] m157_76;
   assign m157_76 =10'b0;

   // m157_77 = W*in
   wire signed [9:0] m157_77;
   assign m157_77 =10'b0;

   // m157_78 = W*in
   wire signed [9:0] m157_78;
   assign m157_78 ={ {5{in157[5]}} , in157[5:1] };

   // m157_79 = W*in
   wire signed [9:0] m157_79;
   assign m157_79 =10'b0;

   // m157_80 = W*in
   wire signed [9:0] m157_80;
   assign m157_80 =10'b0;

   // m157_81 = W*in
   wire signed [9:0] m157_81;
   assign m157_81 =10'b0;

   // m157_82 = W*in
   wire signed [9:0] m157_82;
   assign m157_82 =10'b0;

   // m157_83 = W*in
   wire signed [9:0] m157_83;
   assign m157_83 =10'b0;

   // m157_84 = W*in
   wire signed [9:0] m157_84;
   assign m157_84 =10'b0;

   // m157_85 = W*in
   wire signed [9:0] m157_85;
   assign m157_85 =10'b0;

   // m157_86 = W*in
   wire signed [9:0] m157_86;
   assign m157_86 =10'b0;

   // m157_87 = W*in
   wire signed [9:0] m157_87;
   assign m157_87 =10'b0;

   // m157_88 = W*in
   wire signed [9:0] m157_88;
   assign m157_88 =10'b0;

   // m157_89 = W*in
   wire signed [9:0] m157_89;
   assign m157_89 =10'b0;

   // m157_90 = W*in
   wire signed [9:0] m157_90;
   assign m157_90 =10'b0;

   // m157_91 = W*in
   wire signed [9:0] m157_91;
   assign m157_91 =10'b0;

   // m157_92 = W*in
   wire signed [9:0] m157_92;
   assign m157_92 =10'b0;

   // m157_93 = W*in
   wire signed [9:0] m157_93;
   assign m157_93 =10'b0;

   // m157_94 = W*in
   wire signed [9:0] m157_94;
   assign m157_94 =10'b0;

   // m157_95 = W*in
   wire signed [9:0] m157_95;
   assign m157_95 =10'b0;

   // m157_96 = W*in
   wire signed [9:0] m157_96;
   assign m157_96 =10'b0;

   // m157_97 = W*in
   wire signed [9:0] m157_97;
   assign m157_97 =10'b0;

   // m157_98 = W*in
   wire signed [9:0] m157_98;
   assign m157_98 =10'b0;

   // m157_99 = W*in
   wire signed [9:0] m157_99;
   assign m157_99 =10'b0;

   // m157_100 = W*in
   wire signed [9:0] m157_100;
   assign m157_100 =10'b0;

   // m157_101 = W*in
   wire signed [9:0] m157_101;
   assign m157_101 =10'b0;

   // m157_102 = W*in
   wire signed [9:0] m157_102;
   assign m157_102 =10'b0;

   // m157_103 = W*in
   wire signed [9:0] m157_103;
   assign m157_103 =10'b0;

   // m157_104 = W*in
   wire signed [9:0] m157_104;
   assign m157_104 =10'b0;

   // m157_105 = W*in
   wire signed [9:0] m157_105;
   assign m157_105 =10'b0;

   // m157_106 = W*in
   wire signed [9:0] m157_106;
   assign m157_106 =10'b0;

   // m157_107 = W*in
   wire signed [9:0] m157_107;
   assign m157_107 =10'b0;

   // m157_108 = W*in
   wire signed [9:0] m157_108;
   assign m157_108 =10'b0;

   // m157_109 = W*in
   wire signed [9:0] m157_109;
   assign m157_109 =10'b0;

   // m157_110 = W*in
   wire signed [9:0] m157_110;
   assign m157_110 =10'b0;

   // m157_111 = W*in
   wire signed [9:0] m157_111;
   assign m157_111 =10'b0;

   // m157_112 = W*in
   wire signed [9:0] m157_112;
   assign m157_112 =10'b0;

   // m157_113 = W*in
   wire signed [9:0] m157_113;
   assign m157_113 =10'b0;

   // m157_114 = W*in
   wire signed [9:0] m157_114;
   assign m157_114 =10'b0;

   // m157_115 = W*in
   wire signed [9:0] m157_115;
   assign m157_115 =10'b0;

   // m157_116 = W*in
   wire signed [9:0] m157_116;
   assign m157_116 =10'b0;

   // m157_117 = W*in
   wire signed [9:0] m157_117;
   assign m157_117 =10'b0;

   // m158_1 = W*in
   wire signed [9:0] m158_1;
   assign m158_1 =10'b0;

   // m158_2 = W*in
   wire signed [9:0] m158_2;
   assign m158_2 =10'b0;

   // m158_3 = W*in
   wire signed [9:0] m158_3;
   assign m158_3 =10'b0;

   // m158_4 = W*in
   wire signed [9:0] m158_4;
   assign m158_4 =10'b0;

   // m158_5 = W*in
   wire signed [9:0] m158_5;
   assign m158_5 ={ {4{in158[5]}} , in158[5:0] };

   // m158_6 = W*in
   wire signed [9:0] m158_6;
   assign m158_6 ={ {4{in158[5]}} , in158[5:0] };

   // m158_7 = W*in
   wire signed [9:0] m158_7;
   assign m158_7 =10'b0;

   // m158_8 = W*in
   wire signed [9:0] m158_8;
   assign m158_8 =10'b0;

   // m158_9 = W*in
   wire signed [9:0] m158_9;
   assign m158_9 =10'b0;

   // m158_10 = W*in
   wire signed [9:0] m158_10;
   assign m158_10 =10'b0;

   // m158_11 = W*in
   wire signed [9:0] m158_11;
   assign m158_11 =10'b0;

   // m158_12 = W*in
   wire signed [9:0] m158_12;
   assign m158_12 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_13 = W*in
   wire signed [9:0] m158_13;
   assign m158_13 =10'b0;

   // m158_14 = W*in
   wire signed [9:0] m158_14;
   assign m158_14 =10'b0;

   // m158_15 = W*in
   wire signed [9:0] m158_15;
   assign m158_15 =10'b0;

   // m158_16 = W*in
   wire signed [9:0] m158_16;
   assign m158_16 =10'b0;

   // m158_17 = W*in
   wire signed [9:0] m158_17;
   assign m158_17 ={ {5{neg158[5]}} , neg158[5:1] };

   // m158_18 = W*in
   wire signed [9:0] m158_18;
   assign m158_18 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_19 = W*in
   wire signed [9:0] m158_19;
   assign m158_19 ={ {5{in158[5]}} , in158[5:1] };

   // m158_20 = W*in
   wire signed [9:0] m158_20;
   assign m158_20 =10'b0;

   // m158_21 = W*in
   wire signed [9:0] m158_21;
   assign m158_21 =10'b0;

   // m158_22 = W*in
   wire signed [9:0] m158_22;
   assign m158_22 ={ {5{neg158[5]}} , neg158[5:1] };

   // m158_23 = W*in
   wire signed [9:0] m158_23;
   assign m158_23 ={ {5{neg158[5]}} , neg158[5:1] };

   // m158_24 = W*in
   wire signed [9:0] m158_24;
   assign m158_24 =10'b0;

   // m158_25 = W*in
   wire signed [9:0] m158_25;
   assign m158_25 =10'b0;

   // m158_26 = W*in
   wire signed [9:0] m158_26;
   assign m158_26 ={ {5{in158[5]}} , in158[5:1] };

   // m158_27 = W*in
   wire signed [9:0] m158_27;
   assign m158_27 =10'b0;

   // m158_28 = W*in
   wire signed [9:0] m158_28;
   assign m158_28 ={ {4{in158[5]}} , in158[5:0] };

   // m158_29 = W*in
   wire signed [9:0] m158_29;
   assign m158_29 ={ {4{in158[5]}} , in158[5:0] };

   // m158_30 = W*in
   wire signed [9:0] m158_30;
   assign m158_30 =10'b0;

   // m158_31 = W*in
   wire signed [9:0] m158_31;
   assign m158_31 =10'b0;

   // m158_32 = W*in
   wire signed [9:0] m158_32;
   assign m158_32 =10'b0;

   // m158_33 = W*in
   wire signed [9:0] m158_33;
   assign m158_33 =10'b0;

   // m158_34 = W*in
   wire signed [9:0] m158_34;
   assign m158_34 =10'b0;

   // m158_35 = W*in
   wire signed [9:0] m158_35;
   assign m158_35 =10'b0;

   // m158_36 = W*in
   wire signed [9:0] m158_36;
   assign m158_36 ={ {5{in158[5]}} , in158[5:1] };

   // m158_37 = W*in
   wire signed [9:0] m158_37;
   assign m158_37 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_38 = W*in
   wire signed [9:0] m158_38;
   assign m158_38 =10'b0;

   // m158_39 = W*in
   wire signed [9:0] m158_39;
   assign m158_39 =10'b0;

   // m158_40 = W*in
   wire signed [9:0] m158_40;
   assign m158_40 =10'b0;

   // m158_41 = W*in
   wire signed [9:0] m158_41;
   assign m158_41 =10'b0;

   // m158_42 = W*in
   wire signed [9:0] m158_42;
   assign m158_42 =10'b0;

   // m158_43 = W*in
   wire signed [9:0] m158_43;
   assign m158_43 =10'b0;

   // m158_44 = W*in
   wire signed [9:0] m158_44;
   assign m158_44 ={ {4{in158[5]}} , in158[5:0] };

   // m158_45 = W*in
   wire signed [9:0] m158_45;
   assign m158_45 =10'b0;

   // m158_46 = W*in
   wire signed [9:0] m158_46;
   assign m158_46 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_47 = W*in
   wire signed [9:0] m158_47;
   assign m158_47 =10'b0;

   // m158_48 = W*in
   wire signed [9:0] m158_48;
   assign m158_48 ={ {4{in158[5]}} , in158[5:0] };

   // m158_49 = W*in
   wire signed [9:0] m158_49;
   assign m158_49 =10'b0;

   // m158_50 = W*in
   wire signed [9:0] m158_50;
   assign m158_50 =10'b0;

   // m158_51 = W*in
   wire signed [9:0] m158_51;
   assign m158_51 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_52 = W*in
   wire signed [9:0] m158_52;
   assign m158_52 =10'b0;

   // m158_53 = W*in
   wire signed [9:0] m158_53;
   assign m158_53 ={ {4{in158[5]}} , in158[5:0] };

   // m158_54 = W*in
   wire signed [9:0] m158_54;
   assign m158_54 =10'b0;

   // m158_55 = W*in
   wire signed [9:0] m158_55;
   assign m158_55 =10'b0;

   // m158_56 = W*in
   wire signed [9:0] m158_56;
   assign m158_56 =10'b0;

   // m158_57 = W*in
   wire signed [9:0] m158_57;
   assign m158_57 =10'b0;

   // m158_58 = W*in
   wire signed [9:0] m158_58;
   assign m158_58 ={ {5{in158[5]}} , in158[5:1] };

   // m158_59 = W*in
   wire signed [9:0] m158_59;
   assign m158_59 =10'b0;

   // m158_60 = W*in
   wire signed [9:0] m158_60;
   assign m158_60 =10'b0;

   // m158_61 = W*in
   wire signed [9:0] m158_61;
   assign m158_61 =10'b0;

   // m158_62 = W*in
   wire signed [9:0] m158_62;
   assign m158_62 =10'b0;

   // m158_63 = W*in
   wire signed [9:0] m158_63;
   assign m158_63 ={ {4{in158[5]}} , in158[5:0] };

   // m158_64 = W*in
   wire signed [9:0] m158_64;
   assign m158_64 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_65 = W*in
   wire signed [9:0] m158_65;
   assign m158_65 ={ {5{neg158[5]}} , neg158[5:1] };

   // m158_66 = W*in
   wire signed [9:0] m158_66;
   assign m158_66 =10'b0;

   // m158_67 = W*in
   wire signed [9:0] m158_67;
   assign m158_67 ={ {4{in158[5]}} , in158[5:0] };

   // m158_68 = W*in
   wire signed [9:0] m158_68;
   assign m158_68 =10'b0;

   // m158_69 = W*in
   wire signed [9:0] m158_69;
   assign m158_69 =10'b0;

   // m158_70 = W*in
   wire signed [9:0] m158_70;
   assign m158_70 =10'b0;

   // m158_71 = W*in
   wire signed [9:0] m158_71;
   assign m158_71 =10'b0;

   // m158_72 = W*in
   wire signed [9:0] m158_72;
   assign m158_72 ={ {5{in158[5]}} , in158[5:1] };

   // m158_73 = W*in
   wire signed [9:0] m158_73;
   assign m158_73 =10'b0;

   // m158_74 = W*in
   wire signed [9:0] m158_74;
   assign m158_74 =10'b0;

   // m158_75 = W*in
   wire signed [9:0] m158_75;
   assign m158_75 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_76 = W*in
   wire signed [9:0] m158_76;
   assign m158_76 =10'b0;

   // m158_77 = W*in
   wire signed [9:0] m158_77;
   assign m158_77 =10'b0;

   // m158_78 = W*in
   wire signed [9:0] m158_78;
   assign m158_78 =10'b0;

   // m158_79 = W*in
   wire signed [9:0] m158_79;
   assign m158_79 =10'b0;

   // m158_80 = W*in
   wire signed [9:0] m158_80;
   assign m158_80 =10'b0;

   // m158_81 = W*in
   wire signed [9:0] m158_81;
   assign m158_81 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_82 = W*in
   wire signed [9:0] m158_82;
   assign m158_82 =10'b0;

   // m158_83 = W*in
   wire signed [9:0] m158_83;
   assign m158_83 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_84 = W*in
   wire signed [9:0] m158_84;
   assign m158_84 =10'b0;

   // m158_85 = W*in
   wire signed [9:0] m158_85;
   assign m158_85 =10'b0;

   // m158_86 = W*in
   wire signed [9:0] m158_86;
   assign m158_86 =10'b0;

   // m158_87 = W*in
   wire signed [9:0] m158_87;
   assign m158_87 =10'b0;

   // m158_88 = W*in
   wire signed [9:0] m158_88;
   assign m158_88 =10'b0;

   // m158_89 = W*in
   wire signed [9:0] m158_89;
   assign m158_89 =10'b0;

   // m158_90 = W*in
   wire signed [9:0] m158_90;
   assign m158_90 =10'b0;

   // m158_91 = W*in
   wire signed [9:0] m158_91;
   assign m158_91 =10'b0;

   // m158_92 = W*in
   wire signed [9:0] m158_92;
   assign m158_92 =10'b0;

   // m158_93 = W*in
   wire signed [9:0] m158_93;
   assign m158_93 ={ {4{in158[5]}} , in158[5:0] };

   // m158_94 = W*in
   wire signed [9:0] m158_94;
   assign m158_94 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_95 = W*in
   wire signed [9:0] m158_95;
   assign m158_95 =10'b0;

   // m158_96 = W*in
   wire signed [9:0] m158_96;
   assign m158_96 =10'b0;

   // m158_97 = W*in
   wire signed [9:0] m158_97;
   assign m158_97 =10'b0;

   // m158_98 = W*in
   wire signed [9:0] m158_98;
   assign m158_98 =10'b0;

   // m158_99 = W*in
   wire signed [9:0] m158_99;
   assign m158_99 =10'b0;

   // m158_100 = W*in
   wire signed [9:0] m158_100;
   assign m158_100 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_101 = W*in
   wire signed [9:0] m158_101;
   assign m158_101 =10'b0;

   // m158_102 = W*in
   wire signed [9:0] m158_102;
   assign m158_102 =10'b0;

   // m158_103 = W*in
   wire signed [9:0] m158_103;
   assign m158_103 =10'b0;

   // m158_104 = W*in
   wire signed [9:0] m158_104;
   assign m158_104 =10'b0;

   // m158_105 = W*in
   wire signed [9:0] m158_105;
   assign m158_105 =10'b0;

   // m158_106 = W*in
   wire signed [9:0] m158_106;
   assign m158_106 =10'b0;

   // m158_107 = W*in
   wire signed [9:0] m158_107;
   assign m158_107 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_108 = W*in
   wire signed [9:0] m158_108;
   assign m158_108 ={ {5{neg158[5]}} , neg158[5:1] };

   // m158_109 = W*in
   wire signed [9:0] m158_109;
   assign m158_109 =10'b0;

   // m158_110 = W*in
   wire signed [9:0] m158_110;
   assign m158_110 =10'b0;

   // m158_111 = W*in
   wire signed [9:0] m158_111;
   assign m158_111 =10'b0;

   // m158_112 = W*in
   wire signed [9:0] m158_112;
   assign m158_112 ={ {4{neg158[5]}} , neg158[5:0] };

   // m158_113 = W*in
   wire signed [9:0] m158_113;
   assign m158_113 ={ {5{in158[5]}} , in158[5:1] };

   // m158_114 = W*in
   wire signed [9:0] m158_114;
   assign m158_114 ={ {5{neg158[5]}} , neg158[5:1] };

   // m158_115 = W*in
   wire signed [9:0] m158_115;
   assign m158_115 =10'b0;

   // m158_116 = W*in
   wire signed [9:0] m158_116;
   assign m158_116 =10'b0;

   // m158_117 = W*in
   wire signed [9:0] m158_117;
   assign m158_117 =10'b0;

   // m159_1 = W*in
   wire signed [9:0] m159_1;
   assign m159_1 =10'b0;

   // m159_2 = W*in
   wire signed [9:0] m159_2;
   assign m159_2 =10'b0;

   // m159_3 = W*in
   wire signed [9:0] m159_3;
   assign m159_3 =10'b0;

   // m159_4 = W*in
   wire signed [9:0] m159_4;
   assign m159_4 =10'b0;

   // m159_5 = W*in
   wire signed [9:0] m159_5;
   assign m159_5 ={ {4{in159[5]}} , in159[5:0] };

   // m159_6 = W*in
   wire signed [9:0] m159_6;
   assign m159_6 ={ {4{in159[5]}} , in159[5:0] };

   // m159_7 = W*in
   wire signed [9:0] m159_7;
   assign m159_7 =10'b0;

   // m159_8 = W*in
   wire signed [9:0] m159_8;
   assign m159_8 =10'b0;

   // m159_9 = W*in
   wire signed [9:0] m159_9;
   assign m159_9 =10'b0;

   // m159_10 = W*in
   wire signed [9:0] m159_10;
   assign m159_10 =10'b0;

   // m159_11 = W*in
   wire signed [9:0] m159_11;
   assign m159_11 ={ {5{in159[5]}} , in159[5:1] };

   // m159_12 = W*in
   wire signed [9:0] m159_12;
   assign m159_12 =10'b0;

   // m159_13 = W*in
   wire signed [9:0] m159_13;
   assign m159_13 =10'b0;

   // m159_14 = W*in
   wire signed [9:0] m159_14;
   assign m159_14 =10'b0;

   // m159_15 = W*in
   wire signed [9:0] m159_15;
   assign m159_15 =10'b0;

   // m159_16 = W*in
   wire signed [9:0] m159_16;
   assign m159_16 =10'b0;

   // m159_17 = W*in
   wire signed [9:0] m159_17;
   assign m159_17 =10'b0;

   // m159_18 = W*in
   wire signed [9:0] m159_18;
   assign m159_18 ={ {4{neg159[5]}} , neg159[5:0] };

   // m159_19 = W*in
   wire signed [9:0] m159_19;
   assign m159_19 ={ {4{in159[5]}} , in159[5:0] };

   // m159_20 = W*in
   wire signed [9:0] m159_20;
   assign m159_20 =10'b0;

   // m159_21 = W*in
   wire signed [9:0] m159_21;
   assign m159_21 =10'b0;

   // m159_22 = W*in
   wire signed [9:0] m159_22;
   assign m159_22 =10'b0;

   // m159_23 = W*in
   wire signed [9:0] m159_23;
   assign m159_23 =10'b0;

   // m159_24 = W*in
   wire signed [9:0] m159_24;
   assign m159_24 =10'b0;

   // m159_25 = W*in
   wire signed [9:0] m159_25;
   assign m159_25 =10'b0;

   // m159_26 = W*in
   wire signed [9:0] m159_26;
   assign m159_26 ={ {4{neg159[5]}} , neg159[5:0] };

   // m159_27 = W*in
   wire signed [9:0] m159_27;
   assign m159_27 =10'b0;

   // m159_28 = W*in
   wire signed [9:0] m159_28;
   assign m159_28 =10'b0;

   // m159_29 = W*in
   wire signed [9:0] m159_29;
   assign m159_29 =10'b0;

   // m159_30 = W*in
   wire signed [9:0] m159_30;
   assign m159_30 ={ {4{in159[5]}} , in159[5:0] };

   // m159_31 = W*in
   wire signed [9:0] m159_31;
   assign m159_31 =10'b0;

   // m159_32 = W*in
   wire signed [9:0] m159_32;
   assign m159_32 =10'b0;

   // m159_33 = W*in
   wire signed [9:0] m159_33;
   assign m159_33 =10'b0;

   // m159_34 = W*in
   wire signed [9:0] m159_34;
   assign m159_34 =10'b0;

   // m159_35 = W*in
   wire signed [9:0] m159_35;
   assign m159_35 =10'b0;

   // m159_36 = W*in
   wire signed [9:0] m159_36;
   assign m159_36 =10'b0;

   // m159_37 = W*in
   wire signed [9:0] m159_37;
   assign m159_37 =10'b0;

   // m159_38 = W*in
   wire signed [9:0] m159_38;
   assign m159_38 =10'b0;

   // m159_39 = W*in
   wire signed [9:0] m159_39;
   assign m159_39 =10'b0;

   // m159_40 = W*in
   wire signed [9:0] m159_40;
   assign m159_40 =10'b0;

   // m159_41 = W*in
   wire signed [9:0] m159_41;
   assign m159_41 =10'b0;

   // m159_42 = W*in
   wire signed [9:0] m159_42;
   assign m159_42 =10'b0;

   // m159_43 = W*in
   wire signed [9:0] m159_43;
   assign m159_43 =10'b0;

   // m159_44 = W*in
   wire signed [9:0] m159_44;
   assign m159_44 ={ {4{in159[5]}} , in159[5:0] };

   // m159_45 = W*in
   wire signed [9:0] m159_45;
   assign m159_45 =10'b0;

   // m159_46 = W*in
   wire signed [9:0] m159_46;
   assign m159_46 =10'b0;

   // m159_47 = W*in
   wire signed [9:0] m159_47;
   assign m159_47 =10'b0;

   // m159_48 = W*in
   wire signed [9:0] m159_48;
   assign m159_48 =10'b0;

   // m159_49 = W*in
   wire signed [9:0] m159_49;
   assign m159_49 =10'b0;

   // m159_50 = W*in
   wire signed [9:0] m159_50;
   assign m159_50 =10'b0;

   // m159_51 = W*in
   wire signed [9:0] m159_51;
   assign m159_51 =10'b0;

   // m159_52 = W*in
   wire signed [9:0] m159_52;
   assign m159_52 =10'b0;

   // m159_53 = W*in
   wire signed [9:0] m159_53;
   assign m159_53 ={ {4{in159[5]}} , in159[5:0] };

   // m159_54 = W*in
   wire signed [9:0] m159_54;
   assign m159_54 ={ {4{in159[5]}} , in159[5:0] };

   // m159_55 = W*in
   wire signed [9:0] m159_55;
   assign m159_55 =10'b0;

   // m159_56 = W*in
   wire signed [9:0] m159_56;
   assign m159_56 =10'b0;

   // m159_57 = W*in
   wire signed [9:0] m159_57;
   assign m159_57 =10'b0;

   // m159_58 = W*in
   wire signed [9:0] m159_58;
   assign m159_58 =10'b0;

   // m159_59 = W*in
   wire signed [9:0] m159_59;
   assign m159_59 =10'b0;

   // m159_60 = W*in
   wire signed [9:0] m159_60;
   assign m159_60 =10'b0;

   // m159_61 = W*in
   wire signed [9:0] m159_61;
   assign m159_61 =10'b0;

   // m159_62 = W*in
   wire signed [9:0] m159_62;
   assign m159_62 =10'b0;

   // m159_63 = W*in
   wire signed [9:0] m159_63;
   assign m159_63 ={ {4{in159[5]}} , in159[5:0] };

   // m159_64 = W*in
   wire signed [9:0] m159_64;
   assign m159_64 ={ {4{neg159[5]}} , neg159[5:0] };

   // m159_65 = W*in
   wire signed [9:0] m159_65;
   assign m159_65 =10'b0;

   // m159_66 = W*in
   wire signed [9:0] m159_66;
   assign m159_66 =10'b0;

   // m159_67 = W*in
   wire signed [9:0] m159_67;
   assign m159_67 ={ {4{in159[5]}} , in159[5:0] };

   // m159_68 = W*in
   wire signed [9:0] m159_68;
   assign m159_68 =10'b0;

   // m159_69 = W*in
   wire signed [9:0] m159_69;
   assign m159_69 ={ {5{in159[5]}} , in159[5:1] };

   // m159_70 = W*in
   wire signed [9:0] m159_70;
   assign m159_70 =10'b0;

   // m159_71 = W*in
   wire signed [9:0] m159_71;
   assign m159_71 ={ {5{neg159[5]}} , neg159[5:1] };

   // m159_72 = W*in
   wire signed [9:0] m159_72;
   assign m159_72 ={ {5{neg159[5]}} , neg159[5:1] };

   // m159_73 = W*in
   wire signed [9:0] m159_73;
   assign m159_73 ={ {5{neg159[5]}} , neg159[5:1] };

   // m159_74 = W*in
   wire signed [9:0] m159_74;
   assign m159_74 =10'b0;

   // m159_75 = W*in
   wire signed [9:0] m159_75;
   assign m159_75 ={ {5{neg159[5]}} , neg159[5:1] };

   // m159_76 = W*in
   wire signed [9:0] m159_76;
   assign m159_76 =10'b0;

   // m159_77 = W*in
   wire signed [9:0] m159_77;
   assign m159_77 =10'b0;

   // m159_78 = W*in
   wire signed [9:0] m159_78;
   assign m159_78 ={ {5{neg159[5]}} , neg159[5:1] };

   // m159_79 = W*in
   wire signed [9:0] m159_79;
   assign m159_79 =10'b0;

   // m159_80 = W*in
   wire signed [9:0] m159_80;
   assign m159_80 =10'b0;

   // m159_81 = W*in
   wire signed [9:0] m159_81;
   assign m159_81 ={ {5{neg159[5]}} , neg159[5:1] };

   // m159_82 = W*in
   wire signed [9:0] m159_82;
   assign m159_82 ={ {5{in159[5]}} , in159[5:1] };

   // m159_83 = W*in
   wire signed [9:0] m159_83;
   assign m159_83 =10'b0;

   // m159_84 = W*in
   wire signed [9:0] m159_84;
   assign m159_84 =10'b0;

   // m159_85 = W*in
   wire signed [9:0] m159_85;
   assign m159_85 =10'b0;

   // m159_86 = W*in
   wire signed [9:0] m159_86;
   assign m159_86 =10'b0;

   // m159_87 = W*in
   wire signed [9:0] m159_87;
   assign m159_87 =10'b0;

   // m159_88 = W*in
   wire signed [9:0] m159_88;
   assign m159_88 =10'b0;

   // m159_89 = W*in
   wire signed [9:0] m159_89;
   assign m159_89 =10'b0;

   // m159_90 = W*in
   wire signed [9:0] m159_90;
   assign m159_90 =10'b0;

   // m159_91 = W*in
   wire signed [9:0] m159_91;
   assign m159_91 =10'b0;

   // m159_92 = W*in
   wire signed [9:0] m159_92;
   assign m159_92 =10'b0;

   // m159_93 = W*in
   wire signed [9:0] m159_93;
   assign m159_93 ={ {4{in159[5]}} , in159[5:0] };

   // m159_94 = W*in
   wire signed [9:0] m159_94;
   assign m159_94 ={ {4{neg159[5]}} , neg159[5:0] };

   // m159_95 = W*in
   wire signed [9:0] m159_95;
   assign m159_95 =10'b0;

   // m159_96 = W*in
   wire signed [9:0] m159_96;
   assign m159_96 =10'b0;

   // m159_97 = W*in
   wire signed [9:0] m159_97;
   assign m159_97 =10'b0;

   // m159_98 = W*in
   wire signed [9:0] m159_98;
   assign m159_98 =10'b0;

   // m159_99 = W*in
   wire signed [9:0] m159_99;
   assign m159_99 =10'b0;

   // m159_100 = W*in
   wire signed [9:0] m159_100;
   assign m159_100 =10'b0;

   // m159_101 = W*in
   wire signed [9:0] m159_101;
   assign m159_101 =10'b0;

   // m159_102 = W*in
   wire signed [9:0] m159_102;
   assign m159_102 =10'b0;

   // m159_103 = W*in
   wire signed [9:0] m159_103;
   assign m159_103 =10'b0;

   // m159_104 = W*in
   wire signed [9:0] m159_104;
   assign m159_104 =10'b0;

   // m159_105 = W*in
   wire signed [9:0] m159_105;
   assign m159_105 =10'b0;

   // m159_106 = W*in
   wire signed [9:0] m159_106;
   assign m159_106 =10'b0;

   // m159_107 = W*in
   wire signed [9:0] m159_107;
   assign m159_107 =10'b0;

   // m159_108 = W*in
   wire signed [9:0] m159_108;
   assign m159_108 =10'b0;

   // m159_109 = W*in
   wire signed [9:0] m159_109;
   assign m159_109 =10'b0;

   // m159_110 = W*in
   wire signed [9:0] m159_110;
   assign m159_110 =10'b0;

   // m159_111 = W*in
   wire signed [9:0] m159_111;
   assign m159_111 =10'b0;

   // m159_112 = W*in
   wire signed [9:0] m159_112;
   assign m159_112 ={ {4{neg159[5]}} , neg159[5:0] };

   // m159_113 = W*in
   wire signed [9:0] m159_113;
   assign m159_113 =10'b0;

   // m159_114 = W*in
   wire signed [9:0] m159_114;
   assign m159_114 =10'b0;

   // m159_115 = W*in
   wire signed [9:0] m159_115;
   assign m159_115 =10'b0;

   // m159_116 = W*in
   wire signed [9:0] m159_116;
   assign m159_116 =10'b0;

   // m159_117 = W*in
   wire signed [9:0] m159_117;
   assign m159_117 =10'b0;

   // m160_1 = W*in
   wire signed [9:0] m160_1;
   assign m160_1 =10'b0;

   // m160_2 = W*in
   wire signed [9:0] m160_2;
   assign m160_2 =10'b0;

   // m160_3 = W*in
   wire signed [9:0] m160_3;
   assign m160_3 =10'b0;

   // m160_4 = W*in
   wire signed [9:0] m160_4;
   assign m160_4 =10'b0;

   // m160_5 = W*in
   wire signed [9:0] m160_5;
   assign m160_5 =10'b0;

   // m160_6 = W*in
   wire signed [9:0] m160_6;
   assign m160_6 =10'b0;

   // m160_7 = W*in
   wire signed [9:0] m160_7;
   assign m160_7 =10'b0;

   // m160_8 = W*in
   wire signed [9:0] m160_8;
   assign m160_8 =10'b0;

   // m160_9 = W*in
   wire signed [9:0] m160_9;
   assign m160_9 =10'b0;

   // m160_10 = W*in
   wire signed [9:0] m160_10;
   assign m160_10 =10'b0;

   // m160_11 = W*in
   wire signed [9:0] m160_11;
   assign m160_11 =10'b0;

   // m160_12 = W*in
   wire signed [9:0] m160_12;
   assign m160_12 =10'b0;

   // m160_13 = W*in
   wire signed [9:0] m160_13;
   assign m160_13 =10'b0;

   // m160_14 = W*in
   wire signed [9:0] m160_14;
   assign m160_14 =10'b0;

   // m160_15 = W*in
   wire signed [9:0] m160_15;
   assign m160_15 =10'b0;

   // m160_16 = W*in
   wire signed [9:0] m160_16;
   assign m160_16 =10'b0;

   // m160_17 = W*in
   wire signed [9:0] m160_17;
   assign m160_17 =10'b0;

   // m160_18 = W*in
   wire signed [9:0] m160_18;
   assign m160_18 =10'b0;

   // m160_19 = W*in
   wire signed [9:0] m160_19;
   assign m160_19 =10'b0;

   // m160_20 = W*in
   wire signed [9:0] m160_20;
   assign m160_20 =10'b0;

   // m160_21 = W*in
   wire signed [9:0] m160_21;
   assign m160_21 ={ {5{neg160[5]}} , neg160[5:1] };

   // m160_22 = W*in
   wire signed [9:0] m160_22;
   assign m160_22 ={ {5{in160[5]}} , in160[5:1] };

   // m160_23 = W*in
   wire signed [9:0] m160_23;
   assign m160_23 ={ {5{in160[5]}} , in160[5:1] };

   // m160_24 = W*in
   wire signed [9:0] m160_24;
   assign m160_24 =10'b0;

   // m160_25 = W*in
   wire signed [9:0] m160_25;
   assign m160_25 =10'b0;

   // m160_26 = W*in
   wire signed [9:0] m160_26;
   assign m160_26 =10'b0;

   // m160_27 = W*in
   wire signed [9:0] m160_27;
   assign m160_27 =10'b0;

   // m160_28 = W*in
   wire signed [9:0] m160_28;
   assign m160_28 =10'b0;

   // m160_29 = W*in
   wire signed [9:0] m160_29;
   assign m160_29 =10'b0;

   // m160_30 = W*in
   wire signed [9:0] m160_30;
   assign m160_30 =10'b0;

   // m160_31 = W*in
   wire signed [9:0] m160_31;
   assign m160_31 =10'b0;

   // m160_32 = W*in
   wire signed [9:0] m160_32;
   assign m160_32 =10'b0;

   // m160_33 = W*in
   wire signed [9:0] m160_33;
   assign m160_33 =10'b0;

   // m160_34 = W*in
   wire signed [9:0] m160_34;
   assign m160_34 =10'b0;

   // m160_35 = W*in
   wire signed [9:0] m160_35;
   assign m160_35 =10'b0;

   // m160_36 = W*in
   wire signed [9:0] m160_36;
   assign m160_36 =10'b0;

   // m160_37 = W*in
   wire signed [9:0] m160_37;
   assign m160_37 =10'b0;

   // m160_38 = W*in
   wire signed [9:0] m160_38;
   assign m160_38 =10'b0;

   // m160_39 = W*in
   wire signed [9:0] m160_39;
   assign m160_39 =10'b0;

   // m160_40 = W*in
   wire signed [9:0] m160_40;
   assign m160_40 =10'b0;

   // m160_41 = W*in
   wire signed [9:0] m160_41;
   assign m160_41 =10'b0;

   // m160_42 = W*in
   wire signed [9:0] m160_42;
   assign m160_42 =10'b0;

   // m160_43 = W*in
   wire signed [9:0] m160_43;
   assign m160_43 =10'b0;

   // m160_44 = W*in
   wire signed [9:0] m160_44;
   assign m160_44 =10'b0;

   // m160_45 = W*in
   wire signed [9:0] m160_45;
   assign m160_45 =10'b0;

   // m160_46 = W*in
   wire signed [9:0] m160_46;
   assign m160_46 =10'b0;

   // m160_47 = W*in
   wire signed [9:0] m160_47;
   assign m160_47 =10'b0;

   // m160_48 = W*in
   wire signed [9:0] m160_48;
   assign m160_48 =10'b0;

   // m160_49 = W*in
   wire signed [9:0] m160_49;
   assign m160_49 =10'b0;

   // m160_50 = W*in
   wire signed [9:0] m160_50;
   assign m160_50 =10'b0;

   // m160_51 = W*in
   wire signed [9:0] m160_51;
   assign m160_51 =10'b0;

   // m160_52 = W*in
   wire signed [9:0] m160_52;
   assign m160_52 =10'b0;

   // m160_53 = W*in
   wire signed [9:0] m160_53;
   assign m160_53 =10'b0;

   // m160_54 = W*in
   wire signed [9:0] m160_54;
   assign m160_54 =10'b0;

   // m160_55 = W*in
   wire signed [9:0] m160_55;
   assign m160_55 =10'b0;

   // m160_56 = W*in
   wire signed [9:0] m160_56;
   assign m160_56 =10'b0;

   // m160_57 = W*in
   wire signed [9:0] m160_57;
   assign m160_57 =10'b0;

   // m160_58 = W*in
   wire signed [9:0] m160_58;
   assign m160_58 =10'b0;

   // m160_59 = W*in
   wire signed [9:0] m160_59;
   assign m160_59 =10'b0;

   // m160_60 = W*in
   wire signed [9:0] m160_60;
   assign m160_60 =10'b0;

   // m160_61 = W*in
   wire signed [9:0] m160_61;
   assign m160_61 =10'b0;

   // m160_62 = W*in
   wire signed [9:0] m160_62;
   assign m160_62 =10'b0;

   // m160_63 = W*in
   wire signed [9:0] m160_63;
   assign m160_63 =10'b0;

   // m160_64 = W*in
   wire signed [9:0] m160_64;
   assign m160_64 =10'b0;

   // m160_65 = W*in
   wire signed [9:0] m160_65;
   assign m160_65 =10'b0;

   // m160_66 = W*in
   wire signed [9:0] m160_66;
   assign m160_66 ={ {5{in160[5]}} , in160[5:1] };

   // m160_67 = W*in
   wire signed [9:0] m160_67;
   assign m160_67 =10'b0;

   // m160_68 = W*in
   wire signed [9:0] m160_68;
   assign m160_68 =10'b0;

   // m160_69 = W*in
   wire signed [9:0] m160_69;
   assign m160_69 ={ {4{neg160[5]}} , neg160[5:0] };

   // m160_70 = W*in
   wire signed [9:0] m160_70;
   assign m160_70 ={ {5{neg160[5]}} , neg160[5:1] };

   // m160_71 = W*in
   wire signed [9:0] m160_71;
   assign m160_71 =10'b0;

   // m160_72 = W*in
   wire signed [9:0] m160_72;
   assign m160_72 ={ {4{neg160[5]}} , neg160[5:0] };

   // m160_73 = W*in
   wire signed [9:0] m160_73;
   assign m160_73 =10'b0;

   // m160_74 = W*in
   wire signed [9:0] m160_74;
   assign m160_74 ={ {5{neg160[5]}} , neg160[5:1] };

   // m160_75 = W*in
   wire signed [9:0] m160_75;
   assign m160_75 =10'b0;

   // m160_76 = W*in
   wire signed [9:0] m160_76;
   assign m160_76 =10'b0;

   // m160_77 = W*in
   wire signed [9:0] m160_77;
   assign m160_77 =10'b0;

   // m160_78 = W*in
   wire signed [9:0] m160_78;
   assign m160_78 =10'b0;

   // m160_79 = W*in
   wire signed [9:0] m160_79;
   assign m160_79 =10'b0;

   // m160_80 = W*in
   wire signed [9:0] m160_80;
   assign m160_80 =10'b0;

   // m160_81 = W*in
   wire signed [9:0] m160_81;
   assign m160_81 =10'b0;

   // m160_82 = W*in
   wire signed [9:0] m160_82;
   assign m160_82 ={ {4{neg160[5]}} , neg160[5:0] };

   // m160_83 = W*in
   wire signed [9:0] m160_83;
   assign m160_83 =10'b0;

   // m160_84 = W*in
   wire signed [9:0] m160_84;
   assign m160_84 =10'b0;

   // m160_85 = W*in
   wire signed [9:0] m160_85;
   assign m160_85 =10'b0;

   // m160_86 = W*in
   wire signed [9:0] m160_86;
   assign m160_86 =10'b0;

   // m160_87 = W*in
   wire signed [9:0] m160_87;
   assign m160_87 =10'b0;

   // m160_88 = W*in
   wire signed [9:0] m160_88;
   assign m160_88 =10'b0;

   // m160_89 = W*in
   wire signed [9:0] m160_89;
   assign m160_89 =10'b0;

   // m160_90 = W*in
   wire signed [9:0] m160_90;
   assign m160_90 =10'b0;

   // m160_91 = W*in
   wire signed [9:0] m160_91;
   assign m160_91 =10'b0;

   // m160_92 = W*in
   wire signed [9:0] m160_92;
   assign m160_92 =10'b0;

   // m160_93 = W*in
   wire signed [9:0] m160_93;
   assign m160_93 =10'b0;

   // m160_94 = W*in
   wire signed [9:0] m160_94;
   assign m160_94 =10'b0;

   // m160_95 = W*in
   wire signed [9:0] m160_95;
   assign m160_95 =10'b0;

   // m160_96 = W*in
   wire signed [9:0] m160_96;
   assign m160_96 =10'b0;

   // m160_97 = W*in
   wire signed [9:0] m160_97;
   assign m160_97 =10'b0;

   // m160_98 = W*in
   wire signed [9:0] m160_98;
   assign m160_98 =10'b0;

   // m160_99 = W*in
   wire signed [9:0] m160_99;
   assign m160_99 =10'b0;

   // m160_100 = W*in
   wire signed [9:0] m160_100;
   assign m160_100 =10'b0;

   // m160_101 = W*in
   wire signed [9:0] m160_101;
   assign m160_101 =10'b0;

   // m160_102 = W*in
   wire signed [9:0] m160_102;
   assign m160_102 =10'b0;

   // m160_103 = W*in
   wire signed [9:0] m160_103;
   assign m160_103 =10'b0;

   // m160_104 = W*in
   wire signed [9:0] m160_104;
   assign m160_104 =10'b0;

   // m160_105 = W*in
   wire signed [9:0] m160_105;
   assign m160_105 =10'b0;

   // m160_106 = W*in
   wire signed [9:0] m160_106;
   assign m160_106 =10'b0;

   // m160_107 = W*in
   wire signed [9:0] m160_107;
   assign m160_107 =10'b0;

   // m160_108 = W*in
   wire signed [9:0] m160_108;
   assign m160_108 ={ {5{in160[5]}} , in160[5:1] };

   // m160_109 = W*in
   wire signed [9:0] m160_109;
   assign m160_109 =10'b0;

   // m160_110 = W*in
   wire signed [9:0] m160_110;
   assign m160_110 =10'b0;

   // m160_111 = W*in
   wire signed [9:0] m160_111;
   assign m160_111 =10'b0;

   // m160_112 = W*in
   wire signed [9:0] m160_112;
   assign m160_112 =10'b0;

   // m160_113 = W*in
   wire signed [9:0] m160_113;
   assign m160_113 =10'b0;

   // m160_114 = W*in
   wire signed [9:0] m160_114;
   assign m160_114 =10'b0;

   // m160_115 = W*in
   wire signed [9:0] m160_115;
   assign m160_115 =10'b0;

   // m160_116 = W*in
   wire signed [9:0] m160_116;
   assign m160_116 =10'b0;

   // m160_117 = W*in
   wire signed [9:0] m160_117;
   assign m160_117 =10'b0;

   // m161_1 = W*in
   wire signed [9:0] m161_1;
   assign m161_1 =10'b0;

   // m161_2 = W*in
   wire signed [9:0] m161_2;
   assign m161_2 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_3 = W*in
   wire signed [9:0] m161_3;
   assign m161_3 =10'b0;

   // m161_4 = W*in
   wire signed [9:0] m161_4;
   assign m161_4 =10'b0;

   // m161_5 = W*in
   wire signed [9:0] m161_5;
   assign m161_5 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_6 = W*in
   wire signed [9:0] m161_6;
   assign m161_6 =10'b0;

   // m161_7 = W*in
   wire signed [9:0] m161_7;
   assign m161_7 =10'b0;

   // m161_8 = W*in
   wire signed [9:0] m161_8;
   assign m161_8 =10'b0;

   // m161_9 = W*in
   wire signed [9:0] m161_9;
   assign m161_9 =10'b0;

   // m161_10 = W*in
   wire signed [9:0] m161_10;
   assign m161_10 =10'b0;

   // m161_11 = W*in
   wire signed [9:0] m161_11;
   assign m161_11 =10'b0;

   // m161_12 = W*in
   wire signed [9:0] m161_12;
   assign m161_12 ={ {4{in161[5]}} , in161[5:0] };

   // m161_13 = W*in
   wire signed [9:0] m161_13;
   assign m161_13 =10'b0;

   // m161_14 = W*in
   wire signed [9:0] m161_14;
   assign m161_14 =10'b0;

   // m161_15 = W*in
   wire signed [9:0] m161_15;
   assign m161_15 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_16 = W*in
   wire signed [9:0] m161_16;
   assign m161_16 =10'b0;

   // m161_17 = W*in
   wire signed [9:0] m161_17;
   assign m161_17 =10'b0;

   // m161_18 = W*in
   wire signed [9:0] m161_18;
   assign m161_18 =10'b0;

   // m161_19 = W*in
   wire signed [9:0] m161_19;
   assign m161_19 =10'b0;

   // m161_20 = W*in
   wire signed [9:0] m161_20;
   assign m161_20 ={ {5{in161[5]}} , in161[5:1] };

   // m161_21 = W*in
   wire signed [9:0] m161_21;
   assign m161_21 =10'b0;

   // m161_22 = W*in
   wire signed [9:0] m161_22;
   assign m161_22 ={ {4{in161[5]}} , in161[5:0] };

   // m161_23 = W*in
   wire signed [9:0] m161_23;
   assign m161_23 ={ {4{in161[5]}} , in161[5:0] };

   // m161_24 = W*in
   wire signed [9:0] m161_24;
   assign m161_24 =10'b0;

   // m161_25 = W*in
   wire signed [9:0] m161_25;
   assign m161_25 =10'b0;

   // m161_26 = W*in
   wire signed [9:0] m161_26;
   assign m161_26 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_27 = W*in
   wire signed [9:0] m161_27;
   assign m161_27 =10'b0;

   // m161_28 = W*in
   wire signed [9:0] m161_28;
   assign m161_28 =10'b0;

   // m161_29 = W*in
   wire signed [9:0] m161_29;
   assign m161_29 ={ {4{in161[5]}} , in161[5:0] };

   // m161_30 = W*in
   wire signed [9:0] m161_30;
   assign m161_30 =10'b0;

   // m161_31 = W*in
   wire signed [9:0] m161_31;
   assign m161_31 ={ {5{neg161[5]}} , neg161[5:1] };

   // m161_32 = W*in
   wire signed [9:0] m161_32;
   assign m161_32 =10'b0;

   // m161_33 = W*in
   wire signed [9:0] m161_33;
   assign m161_33 =10'b0;

   // m161_34 = W*in
   wire signed [9:0] m161_34;
   assign m161_34 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_35 = W*in
   wire signed [9:0] m161_35;
   assign m161_35 ={ {5{in161[5]}} , in161[5:1] };

   // m161_36 = W*in
   wire signed [9:0] m161_36;
   assign m161_36 ={ {5{neg161[5]}} , neg161[5:1] };

   // m161_37 = W*in
   wire signed [9:0] m161_37;
   assign m161_37 =10'b0;

   // m161_38 = W*in
   wire signed [9:0] m161_38;
   assign m161_38 =10'b0;

   // m161_39 = W*in
   wire signed [9:0] m161_39;
   assign m161_39 ={ {4{in161[5]}} , in161[5:0] };

   // m161_40 = W*in
   wire signed [9:0] m161_40;
   assign m161_40 =10'b0;

   // m161_41 = W*in
   wire signed [9:0] m161_41;
   assign m161_41 =10'b0;

   // m161_42 = W*in
   wire signed [9:0] m161_42;
   assign m161_42 =10'b0;

   // m161_43 = W*in
   wire signed [9:0] m161_43;
   assign m161_43 =10'b0;

   // m161_44 = W*in
   wire signed [9:0] m161_44;
   assign m161_44 =10'b0;

   // m161_45 = W*in
   wire signed [9:0] m161_45;
   assign m161_45 =10'b0;

   // m161_46 = W*in
   wire signed [9:0] m161_46;
   assign m161_46 ={ {4{in161[5]}} , in161[5:0] };

   // m161_47 = W*in
   wire signed [9:0] m161_47;
   assign m161_47 =10'b0;

   // m161_48 = W*in
   wire signed [9:0] m161_48;
   assign m161_48 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_49 = W*in
   wire signed [9:0] m161_49;
   assign m161_49 =10'b0;

   // m161_50 = W*in
   wire signed [9:0] m161_50;
   assign m161_50 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_51 = W*in
   wire signed [9:0] m161_51;
   assign m161_51 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_52 = W*in
   wire signed [9:0] m161_52;
   assign m161_52 =10'b0;

   // m161_53 = W*in
   wire signed [9:0] m161_53;
   assign m161_53 =10'b0;

   // m161_54 = W*in
   wire signed [9:0] m161_54;
   assign m161_54 =10'b0;

   // m161_55 = W*in
   wire signed [9:0] m161_55;
   assign m161_55 =10'b0;

   // m161_56 = W*in
   wire signed [9:0] m161_56;
   assign m161_56 =10'b0;

   // m161_57 = W*in
   wire signed [9:0] m161_57;
   assign m161_57 =10'b0;

   // m161_58 = W*in
   wire signed [9:0] m161_58;
   assign m161_58 =10'b0;

   // m161_59 = W*in
   wire signed [9:0] m161_59;
   assign m161_59 =10'b0;

   // m161_60 = W*in
   wire signed [9:0] m161_60;
   assign m161_60 =10'b0;

   // m161_61 = W*in
   wire signed [9:0] m161_61;
   assign m161_61 =10'b0;

   // m161_62 = W*in
   wire signed [9:0] m161_62;
   assign m161_62 =10'b0;

   // m161_63 = W*in
   wire signed [9:0] m161_63;
   assign m161_63 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_64 = W*in
   wire signed [9:0] m161_64;
   assign m161_64 =10'b0;

   // m161_65 = W*in
   wire signed [9:0] m161_65;
   assign m161_65 =10'b0;

   // m161_66 = W*in
   wire signed [9:0] m161_66;
   assign m161_66 ={ {4{in161[5]}} , in161[5:0] };

   // m161_67 = W*in
   wire signed [9:0] m161_67;
   assign m161_67 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_68 = W*in
   wire signed [9:0] m161_68;
   assign m161_68 =10'b0;

   // m161_69 = W*in
   wire signed [9:0] m161_69;
   assign m161_69 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_70 = W*in
   wire signed [9:0] m161_70;
   assign m161_70 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_71 = W*in
   wire signed [9:0] m161_71;
   assign m161_71 =10'b0;

   // m161_72 = W*in
   wire signed [9:0] m161_72;
   assign m161_72 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_73 = W*in
   wire signed [9:0] m161_73;
   assign m161_73 ={ {5{neg161[5]}} , neg161[5:1] };

   // m161_74 = W*in
   wire signed [9:0] m161_74;
   assign m161_74 =10'b0;

   // m161_75 = W*in
   wire signed [9:0] m161_75;
   assign m161_75 =10'b0;

   // m161_76 = W*in
   wire signed [9:0] m161_76;
   assign m161_76 =10'b0;

   // m161_77 = W*in
   wire signed [9:0] m161_77;
   assign m161_77 =10'b0;

   // m161_78 = W*in
   wire signed [9:0] m161_78;
   assign m161_78 =10'b0;

   // m161_79 = W*in
   wire signed [9:0] m161_79;
   assign m161_79 ={ {4{in161[5]}} , in161[5:0] };

   // m161_80 = W*in
   wire signed [9:0] m161_80;
   assign m161_80 =10'b0;

   // m161_81 = W*in
   wire signed [9:0] m161_81;
   assign m161_81 ={ {4{in161[5]}} , in161[5:0] };

   // m161_82 = W*in
   wire signed [9:0] m161_82;
   assign m161_82 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_83 = W*in
   wire signed [9:0] m161_83;
   assign m161_83 =10'b0;

   // m161_84 = W*in
   wire signed [9:0] m161_84;
   assign m161_84 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_85 = W*in
   wire signed [9:0] m161_85;
   assign m161_85 =10'b0;

   // m161_86 = W*in
   wire signed [9:0] m161_86;
   assign m161_86 =10'b0;

   // m161_87 = W*in
   wire signed [9:0] m161_87;
   assign m161_87 =10'b0;

   // m161_88 = W*in
   wire signed [9:0] m161_88;
   assign m161_88 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_89 = W*in
   wire signed [9:0] m161_89;
   assign m161_89 =10'b0;

   // m161_90 = W*in
   wire signed [9:0] m161_90;
   assign m161_90 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_91 = W*in
   wire signed [9:0] m161_91;
   assign m161_91 =10'b0;

   // m161_92 = W*in
   wire signed [9:0] m161_92;
   assign m161_92 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_93 = W*in
   wire signed [9:0] m161_93;
   assign m161_93 =10'b0;

   // m161_94 = W*in
   wire signed [9:0] m161_94;
   assign m161_94 ={ {4{in161[5]}} , in161[5:0] };

   // m161_95 = W*in
   wire signed [9:0] m161_95;
   assign m161_95 ={ {4{in161[5]}} , in161[5:0] };

   // m161_96 = W*in
   wire signed [9:0] m161_96;
   assign m161_96 =10'b0;

   // m161_97 = W*in
   wire signed [9:0] m161_97;
   assign m161_97 ={ {4{in161[5]}} , in161[5:0] };

   // m161_98 = W*in
   wire signed [9:0] m161_98;
   assign m161_98 =10'b0;

   // m161_99 = W*in
   wire signed [9:0] m161_99;
   assign m161_99 =10'b0;

   // m161_100 = W*in
   wire signed [9:0] m161_100;
   assign m161_100 ={ {4{in161[5]}} , in161[5:0] };

   // m161_101 = W*in
   wire signed [9:0] m161_101;
   assign m161_101 =10'b0;

   // m161_102 = W*in
   wire signed [9:0] m161_102;
   assign m161_102 =10'b0;

   // m161_103 = W*in
   wire signed [9:0] m161_103;
   assign m161_103 =10'b0;

   // m161_104 = W*in
   wire signed [9:0] m161_104;
   assign m161_104 =10'b0;

   // m161_105 = W*in
   wire signed [9:0] m161_105;
   assign m161_105 =10'b0;

   // m161_106 = W*in
   wire signed [9:0] m161_106;
   assign m161_106 =10'b0;

   // m161_107 = W*in
   wire signed [9:0] m161_107;
   assign m161_107 =10'b0;

   // m161_108 = W*in
   wire signed [9:0] m161_108;
   assign m161_108 =10'b0;

   // m161_109 = W*in
   wire signed [9:0] m161_109;
   assign m161_109 ={ {4{in161[5]}} , in161[5:0] };

   // m161_110 = W*in
   wire signed [9:0] m161_110;
   assign m161_110 ={ {4{in161[5]}} , in161[5:0] };

   // m161_111 = W*in
   wire signed [9:0] m161_111;
   assign m161_111 ={ {4{neg161[5]}} , neg161[5:0] };

   // m161_112 = W*in
   wire signed [9:0] m161_112;
   assign m161_112 ={ {4{in161[5]}} , in161[5:0] };

   // m161_113 = W*in
   wire signed [9:0] m161_113;
   assign m161_113 =10'b0;

   // m161_114 = W*in
   wire signed [9:0] m161_114;
   assign m161_114 ={ {5{in161[5]}} , in161[5:1] };

   // m161_115 = W*in
   wire signed [9:0] m161_115;
   assign m161_115 =10'b0;

   // m161_116 = W*in
   wire signed [9:0] m161_116;
   assign m161_116 =10'b0;

   // m161_117 = W*in
   wire signed [9:0] m161_117;
   assign m161_117 ={ {4{in161[5]}} , in161[5:0] };

   // m162_1 = W*in
   wire signed [9:0] m162_1;
   assign m162_1 =10'b0;

   // m162_2 = W*in
   wire signed [9:0] m162_2;
   assign m162_2 =10'b0;

   // m162_3 = W*in
   wire signed [9:0] m162_3;
   assign m162_3 =10'b0;

   // m162_4 = W*in
   wire signed [9:0] m162_4;
   assign m162_4 =10'b0;

   // m162_5 = W*in
   wire signed [9:0] m162_5;
   assign m162_5 =10'b0;

   // m162_6 = W*in
   wire signed [9:0] m162_6;
   assign m162_6 ={ {4{in162[5]}} , in162[5:0] };

   // m162_7 = W*in
   wire signed [9:0] m162_7;
   assign m162_7 =10'b0;

   // m162_8 = W*in
   wire signed [9:0] m162_8;
   assign m162_8 =10'b0;

   // m162_9 = W*in
   wire signed [9:0] m162_9;
   assign m162_9 =10'b0;

   // m162_10 = W*in
   wire signed [9:0] m162_10;
   assign m162_10 =10'b0;

   // m162_11 = W*in
   wire signed [9:0] m162_11;
   assign m162_11 =10'b0;

   // m162_12 = W*in
   wire signed [9:0] m162_12;
   assign m162_12 ={ {4{in162[5]}} , in162[5:0] };

   // m162_13 = W*in
   wire signed [9:0] m162_13;
   assign m162_13 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_14 = W*in
   wire signed [9:0] m162_14;
   assign m162_14 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_15 = W*in
   wire signed [9:0] m162_15;
   assign m162_15 =10'b0;

   // m162_16 = W*in
   wire signed [9:0] m162_16;
   assign m162_16 =10'b0;

   // m162_17 = W*in
   wire signed [9:0] m162_17;
   assign m162_17 ={ {5{in162[5]}} , in162[5:1] };

   // m162_18 = W*in
   wire signed [9:0] m162_18;
   assign m162_18 =10'b0;

   // m162_19 = W*in
   wire signed [9:0] m162_19;
   assign m162_19 =10'b0;

   // m162_20 = W*in
   wire signed [9:0] m162_20;
   assign m162_20 ={ {4{in162[5]}} , in162[5:0] };

   // m162_21 = W*in
   wire signed [9:0] m162_21;
   assign m162_21 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_22 = W*in
   wire signed [9:0] m162_22;
   assign m162_22 ={ {5{in162[5]}} , in162[5:1] };

   // m162_23 = W*in
   wire signed [9:0] m162_23;
   assign m162_23 ={ {4{in162[5]}} , in162[5:0] };

   // m162_24 = W*in
   wire signed [9:0] m162_24;
   assign m162_24 ={ {4{in162[5]}} , in162[5:0] };

   // m162_25 = W*in
   wire signed [9:0] m162_25;
   assign m162_25 =10'b0;

   // m162_26 = W*in
   wire signed [9:0] m162_26;
   assign m162_26 =10'b0;

   // m162_27 = W*in
   wire signed [9:0] m162_27;
   assign m162_27 ={ {5{in162[5]}} , in162[5:1] };

   // m162_28 = W*in
   wire signed [9:0] m162_28;
   assign m162_28 =10'b0;

   // m162_29 = W*in
   wire signed [9:0] m162_29;
   assign m162_29 =10'b0;

   // m162_30 = W*in
   wire signed [9:0] m162_30;
   assign m162_30 ={ {4{in162[5]}} , in162[5:0] };

   // m162_31 = W*in
   wire signed [9:0] m162_31;
   assign m162_31 =10'b0;

   // m162_32 = W*in
   wire signed [9:0] m162_32;
   assign m162_32 =10'b0;

   // m162_33 = W*in
   wire signed [9:0] m162_33;
   assign m162_33 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_34 = W*in
   wire signed [9:0] m162_34;
   assign m162_34 =10'b0;

   // m162_35 = W*in
   wire signed [9:0] m162_35;
   assign m162_35 ={ {4{in162[5]}} , in162[5:0] };

   // m162_36 = W*in
   wire signed [9:0] m162_36;
   assign m162_36 =10'b0;

   // m162_37 = W*in
   wire signed [9:0] m162_37;
   assign m162_37 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_38 = W*in
   wire signed [9:0] m162_38;
   assign m162_38 =10'b0;

   // m162_39 = W*in
   wire signed [9:0] m162_39;
   assign m162_39 ={ {4{in162[5]}} , in162[5:0] };

   // m162_40 = W*in
   wire signed [9:0] m162_40;
   assign m162_40 =10'b0;

   // m162_41 = W*in
   wire signed [9:0] m162_41;
   assign m162_41 =10'b0;

   // m162_42 = W*in
   wire signed [9:0] m162_42;
   assign m162_42 =10'b0;

   // m162_43 = W*in
   wire signed [9:0] m162_43;
   assign m162_43 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_44 = W*in
   wire signed [9:0] m162_44;
   assign m162_44 =10'b0;

   // m162_45 = W*in
   wire signed [9:0] m162_45;
   assign m162_45 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_46 = W*in
   wire signed [9:0] m162_46;
   assign m162_46 =10'b0;

   // m162_47 = W*in
   wire signed [9:0] m162_47;
   assign m162_47 =10'b0;

   // m162_48 = W*in
   wire signed [9:0] m162_48;
   assign m162_48 ={ {3{neg162[5]}} , neg162 , {1{1'b0}} };

   // m162_49 = W*in
   wire signed [9:0] m162_49;
   assign m162_49 =10'b0;

   // m162_50 = W*in
   wire signed [9:0] m162_50;
   assign m162_50 =10'b0;

   // m162_51 = W*in
   wire signed [9:0] m162_51;
   assign m162_51 =10'b0;

   // m162_52 = W*in
   wire signed [9:0] m162_52;
   assign m162_52 =10'b0;

   // m162_53 = W*in
   wire signed [9:0] m162_53;
   assign m162_53 =10'b0;

   // m162_54 = W*in
   wire signed [9:0] m162_54;
   assign m162_54 =10'b0;

   // m162_55 = W*in
   wire signed [9:0] m162_55;
   assign m162_55 =10'b0;

   // m162_56 = W*in
   wire signed [9:0] m162_56;
   assign m162_56 =10'b0;

   // m162_57 = W*in
   wire signed [9:0] m162_57;
   assign m162_57 =10'b0;

   // m162_58 = W*in
   wire signed [9:0] m162_58;
   assign m162_58 =10'b0;

   // m162_59 = W*in
   wire signed [9:0] m162_59;
   assign m162_59 =10'b0;

   // m162_60 = W*in
   wire signed [9:0] m162_60;
   assign m162_60 =10'b0;

   // m162_61 = W*in
   wire signed [9:0] m162_61;
   assign m162_61 ={ {4{in162[5]}} , in162[5:0] };

   // m162_62 = W*in
   wire signed [9:0] m162_62;
   assign m162_62 =10'b0;

   // m162_63 = W*in
   wire signed [9:0] m162_63;
   assign m162_63 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_64 = W*in
   wire signed [9:0] m162_64;
   assign m162_64 ={ {4{in162[5]}} , in162[5:0] };

   // m162_65 = W*in
   wire signed [9:0] m162_65;
   assign m162_65 =10'b0;

   // m162_66 = W*in
   wire signed [9:0] m162_66;
   assign m162_66 ={ {4{in162[5]}} , in162[5:0] };

   // m162_67 = W*in
   wire signed [9:0] m162_67;
   assign m162_67 =10'b0;

   // m162_68 = W*in
   wire signed [9:0] m162_68;
   assign m162_68 =10'b0;

   // m162_69 = W*in
   wire signed [9:0] m162_69;
   assign m162_69 ={ {3{neg162[5]}} , neg162 , {1{1'b0}} };

   // m162_70 = W*in
   wire signed [9:0] m162_70;
   assign m162_70 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_71 = W*in
   wire signed [9:0] m162_71;
   assign m162_71 =10'b0;

   // m162_72 = W*in
   wire signed [9:0] m162_72;
   assign m162_72 ={ {3{neg162[5]}} , neg162 , {1{1'b0}} };

   // m162_73 = W*in
   wire signed [9:0] m162_73;
   assign m162_73 =10'b0;

   // m162_74 = W*in
   wire signed [9:0] m162_74;
   assign m162_74 ={ {4{in162[5]}} , in162[5:0] };

   // m162_75 = W*in
   wire signed [9:0] m162_75;
   assign m162_75 =10'b0;

   // m162_76 = W*in
   wire signed [9:0] m162_76;
   assign m162_76 =10'b0;

   // m162_77 = W*in
   wire signed [9:0] m162_77;
   assign m162_77 =10'b0;

   // m162_78 = W*in
   wire signed [9:0] m162_78;
   assign m162_78 =10'b0;

   // m162_79 = W*in
   wire signed [9:0] m162_79;
   assign m162_79 =10'b0;

   // m162_80 = W*in
   wire signed [9:0] m162_80;
   assign m162_80 =10'b0;

   // m162_81 = W*in
   wire signed [9:0] m162_81;
   assign m162_81 ={ {5{in162[5]}} , in162[5:1] };

   // m162_82 = W*in
   wire signed [9:0] m162_82;
   assign m162_82 ={ {3{neg162[5]}} , neg162 , {1{1'b0}} };

   // m162_83 = W*in
   wire signed [9:0] m162_83;
   assign m162_83 =10'b0;

   // m162_84 = W*in
   wire signed [9:0] m162_84;
   assign m162_84 ={ {3{neg162[5]}} , neg162 , {1{1'b0}} };

   // m162_85 = W*in
   wire signed [9:0] m162_85;
   assign m162_85 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_86 = W*in
   wire signed [9:0] m162_86;
   assign m162_86 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_87 = W*in
   wire signed [9:0] m162_87;
   assign m162_87 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_88 = W*in
   wire signed [9:0] m162_88;
   assign m162_88 =10'b0;

   // m162_89 = W*in
   wire signed [9:0] m162_89;
   assign m162_89 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_90 = W*in
   wire signed [9:0] m162_90;
   assign m162_90 =10'b0;

   // m162_91 = W*in
   wire signed [9:0] m162_91;
   assign m162_91 ={ {4{in162[5]}} , in162[5:0] };

   // m162_92 = W*in
   wire signed [9:0] m162_92;
   assign m162_92 =10'b0;

   // m162_93 = W*in
   wire signed [9:0] m162_93;
   assign m162_93 =10'b0;

   // m162_94 = W*in
   wire signed [9:0] m162_94;
   assign m162_94 ={ {4{in162[5]}} , in162[5:0] };

   // m162_95 = W*in
   wire signed [9:0] m162_95;
   assign m162_95 =10'b0;

   // m162_96 = W*in
   wire signed [9:0] m162_96;
   assign m162_96 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_97 = W*in
   wire signed [9:0] m162_97;
   assign m162_97 ={ {4{in162[5]}} , in162[5:0] };

   // m162_98 = W*in
   wire signed [9:0] m162_98;
   assign m162_98 ={ {4{in162[5]}} , in162[5:0] };

   // m162_99 = W*in
   wire signed [9:0] m162_99;
   assign m162_99 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_100 = W*in
   wire signed [9:0] m162_100;
   assign m162_100 =10'b0;

   // m162_101 = W*in
   wire signed [9:0] m162_101;
   assign m162_101 =10'b0;

   // m162_102 = W*in
   wire signed [9:0] m162_102;
   assign m162_102 =10'b0;

   // m162_103 = W*in
   wire signed [9:0] m162_103;
   assign m162_103 =10'b0;

   // m162_104 = W*in
   wire signed [9:0] m162_104;
   assign m162_104 ={ {4{in162[5]}} , in162[5:0] };

   // m162_105 = W*in
   wire signed [9:0] m162_105;
   assign m162_105 =10'b0;

   // m162_106 = W*in
   wire signed [9:0] m162_106;
   assign m162_106 =10'b0;

   // m162_107 = W*in
   wire signed [9:0] m162_107;
   assign m162_107 =10'b0;

   // m162_108 = W*in
   wire signed [9:0] m162_108;
   assign m162_108 =10'b0;

   // m162_109 = W*in
   wire signed [9:0] m162_109;
   assign m162_109 =10'b0;

   // m162_110 = W*in
   wire signed [9:0] m162_110;
   assign m162_110 ={ {5{neg162[5]}} , neg162[5:1] };

   // m162_111 = W*in
   wire signed [9:0] m162_111;
   assign m162_111 ={ {4{neg162[5]}} , neg162[5:0] };

   // m162_112 = W*in
   wire signed [9:0] m162_112;
   assign m162_112 ={ {4{in162[5]}} , in162[5:0] };

   // m162_113 = W*in
   wire signed [9:0] m162_113;
   assign m162_113 =10'b0;

   // m162_114 = W*in
   wire signed [9:0] m162_114;
   assign m162_114 =10'b0;

   // m162_115 = W*in
   wire signed [9:0] m162_115;
   assign m162_115 ={ {4{in162[5]}} , in162[5:0] };

   // m162_116 = W*in
   wire signed [9:0] m162_116;
   assign m162_116 =10'b0;

   // m162_117 = W*in
   wire signed [9:0] m162_117;
   assign m162_117 =10'b0;

   // m163_1 = W*in
   wire signed [9:0] m163_1;
   assign m163_1 ={ {4{in163[5]}} , in163[5:0] };

   // m163_2 = W*in
   wire signed [9:0] m163_2;
   assign m163_2 =10'b0;

   // m163_3 = W*in
   wire signed [9:0] m163_3;
   assign m163_3 =10'b0;

   // m163_4 = W*in
   wire signed [9:0] m163_4;
   assign m163_4 =10'b0;

   // m163_5 = W*in
   wire signed [9:0] m163_5;
   assign m163_5 =10'b0;

   // m163_6 = W*in
   wire signed [9:0] m163_6;
   assign m163_6 =10'b0;

   // m163_7 = W*in
   wire signed [9:0] m163_7;
   assign m163_7 =10'b0;

   // m163_8 = W*in
   wire signed [9:0] m163_8;
   assign m163_8 =10'b0;

   // m163_9 = W*in
   wire signed [9:0] m163_9;
   assign m163_9 =10'b0;

   // m163_10 = W*in
   wire signed [9:0] m163_10;
   assign m163_10 =10'b0;

   // m163_11 = W*in
   wire signed [9:0] m163_11;
   assign m163_11 =10'b0;

   // m163_12 = W*in
   wire signed [9:0] m163_12;
   assign m163_12 =10'b0;

   // m163_13 = W*in
   wire signed [9:0] m163_13;
   assign m163_13 =10'b0;

   // m163_14 = W*in
   wire signed [9:0] m163_14;
   assign m163_14 =10'b0;

   // m163_15 = W*in
   wire signed [9:0] m163_15;
   assign m163_15 =10'b0;

   // m163_16 = W*in
   wire signed [9:0] m163_16;
   assign m163_16 =10'b0;

   // m163_17 = W*in
   wire signed [9:0] m163_17;
   assign m163_17 =10'b0;

   // m163_18 = W*in
   wire signed [9:0] m163_18;
   assign m163_18 =10'b0;

   // m163_19 = W*in
   wire signed [9:0] m163_19;
   assign m163_19 =10'b0;

   // m163_20 = W*in
   wire signed [9:0] m163_20;
   assign m163_20 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_21 = W*in
   wire signed [9:0] m163_21;
   assign m163_21 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_22 = W*in
   wire signed [9:0] m163_22;
   assign m163_22 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_23 = W*in
   wire signed [9:0] m163_23;
   assign m163_23 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_24 = W*in
   wire signed [9:0] m163_24;
   assign m163_24 =10'b0;

   // m163_25 = W*in
   wire signed [9:0] m163_25;
   assign m163_25 =10'b0;

   // m163_26 = W*in
   wire signed [9:0] m163_26;
   assign m163_26 =10'b0;

   // m163_27 = W*in
   wire signed [9:0] m163_27;
   assign m163_27 ={ {5{in163[5]}} , in163[5:1] };

   // m163_28 = W*in
   wire signed [9:0] m163_28;
   assign m163_28 ={ {5{in163[5]}} , in163[5:1] };

   // m163_29 = W*in
   wire signed [9:0] m163_29;
   assign m163_29 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_30 = W*in
   wire signed [9:0] m163_30;
   assign m163_30 =10'b0;

   // m163_31 = W*in
   wire signed [9:0] m163_31;
   assign m163_31 =10'b0;

   // m163_32 = W*in
   wire signed [9:0] m163_32;
   assign m163_32 =10'b0;

   // m163_33 = W*in
   wire signed [9:0] m163_33;
   assign m163_33 =10'b0;

   // m163_34 = W*in
   wire signed [9:0] m163_34;
   assign m163_34 =10'b0;

   // m163_35 = W*in
   wire signed [9:0] m163_35;
   assign m163_35 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_36 = W*in
   wire signed [9:0] m163_36;
   assign m163_36 =10'b0;

   // m163_37 = W*in
   wire signed [9:0] m163_37;
   assign m163_37 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_38 = W*in
   wire signed [9:0] m163_38;
   assign m163_38 =10'b0;

   // m163_39 = W*in
   wire signed [9:0] m163_39;
   assign m163_39 =10'b0;

   // m163_40 = W*in
   wire signed [9:0] m163_40;
   assign m163_40 =10'b0;

   // m163_41 = W*in
   wire signed [9:0] m163_41;
   assign m163_41 =10'b0;

   // m163_42 = W*in
   wire signed [9:0] m163_42;
   assign m163_42 =10'b0;

   // m163_43 = W*in
   wire signed [9:0] m163_43;
   assign m163_43 ={ {4{in163[5]}} , in163[5:0] };

   // m163_44 = W*in
   wire signed [9:0] m163_44;
   assign m163_44 =10'b0;

   // m163_45 = W*in
   wire signed [9:0] m163_45;
   assign m163_45 =10'b0;

   // m163_46 = W*in
   wire signed [9:0] m163_46;
   assign m163_46 =10'b0;

   // m163_47 = W*in
   wire signed [9:0] m163_47;
   assign m163_47 =10'b0;

   // m163_48 = W*in
   wire signed [9:0] m163_48;
   assign m163_48 =10'b0;

   // m163_49 = W*in
   wire signed [9:0] m163_49;
   assign m163_49 =10'b0;

   // m163_50 = W*in
   wire signed [9:0] m163_50;
   assign m163_50 =10'b0;

   // m163_51 = W*in
   wire signed [9:0] m163_51;
   assign m163_51 ={ {4{in163[5]}} , in163[5:0] };

   // m163_52 = W*in
   wire signed [9:0] m163_52;
   assign m163_52 =10'b0;

   // m163_53 = W*in
   wire signed [9:0] m163_53;
   assign m163_53 =10'b0;

   // m163_54 = W*in
   wire signed [9:0] m163_54;
   assign m163_54 =10'b0;

   // m163_55 = W*in
   wire signed [9:0] m163_55;
   assign m163_55 =10'b0;

   // m163_56 = W*in
   wire signed [9:0] m163_56;
   assign m163_56 =10'b0;

   // m163_57 = W*in
   wire signed [9:0] m163_57;
   assign m163_57 =10'b0;

   // m163_58 = W*in
   wire signed [9:0] m163_58;
   assign m163_58 =10'b0;

   // m163_59 = W*in
   wire signed [9:0] m163_59;
   assign m163_59 =10'b0;

   // m163_60 = W*in
   wire signed [9:0] m163_60;
   assign m163_60 =10'b0;

   // m163_61 = W*in
   wire signed [9:0] m163_61;
   assign m163_61 =10'b0;

   // m163_62 = W*in
   wire signed [9:0] m163_62;
   assign m163_62 =10'b0;

   // m163_63 = W*in
   wire signed [9:0] m163_63;
   assign m163_63 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_64 = W*in
   wire signed [9:0] m163_64;
   assign m163_64 =10'b0;

   // m163_65 = W*in
   wire signed [9:0] m163_65;
   assign m163_65 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_66 = W*in
   wire signed [9:0] m163_66;
   assign m163_66 =10'b0;

   // m163_67 = W*in
   wire signed [9:0] m163_67;
   assign m163_67 =10'b0;

   // m163_68 = W*in
   wire signed [9:0] m163_68;
   assign m163_68 =10'b0;

   // m163_69 = W*in
   wire signed [9:0] m163_69;
   assign m163_69 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_70 = W*in
   wire signed [9:0] m163_70;
   assign m163_70 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_71 = W*in
   wire signed [9:0] m163_71;
   assign m163_71 ={ {5{in163[5]}} , in163[5:1] };

   // m163_72 = W*in
   wire signed [9:0] m163_72;
   assign m163_72 =10'b0;

   // m163_73 = W*in
   wire signed [9:0] m163_73;
   assign m163_73 =10'b0;

   // m163_74 = W*in
   wire signed [9:0] m163_74;
   assign m163_74 ={ {4{in163[5]}} , in163[5:0] };

   // m163_75 = W*in
   wire signed [9:0] m163_75;
   assign m163_75 =10'b0;

   // m163_76 = W*in
   wire signed [9:0] m163_76;
   assign m163_76 =10'b0;

   // m163_77 = W*in
   wire signed [9:0] m163_77;
   assign m163_77 =10'b0;

   // m163_78 = W*in
   wire signed [9:0] m163_78;
   assign m163_78 =10'b0;

   // m163_79 = W*in
   wire signed [9:0] m163_79;
   assign m163_79 =10'b0;

   // m163_80 = W*in
   wire signed [9:0] m163_80;
   assign m163_80 =10'b0;

   // m163_81 = W*in
   wire signed [9:0] m163_81;
   assign m163_81 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_82 = W*in
   wire signed [9:0] m163_82;
   assign m163_82 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_83 = W*in
   wire signed [9:0] m163_83;
   assign m163_83 ={ {5{in163[5]}} , in163[5:1] };

   // m163_84 = W*in
   wire signed [9:0] m163_84;
   assign m163_84 =10'b0;

   // m163_85 = W*in
   wire signed [9:0] m163_85;
   assign m163_85 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_86 = W*in
   wire signed [9:0] m163_86;
   assign m163_86 =10'b0;

   // m163_87 = W*in
   wire signed [9:0] m163_87;
   assign m163_87 =10'b0;

   // m163_88 = W*in
   wire signed [9:0] m163_88;
   assign m163_88 =10'b0;

   // m163_89 = W*in
   wire signed [9:0] m163_89;
   assign m163_89 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_90 = W*in
   wire signed [9:0] m163_90;
   assign m163_90 =10'b0;

   // m163_91 = W*in
   wire signed [9:0] m163_91;
   assign m163_91 =10'b0;

   // m163_92 = W*in
   wire signed [9:0] m163_92;
   assign m163_92 ={ {4{in163[5]}} , in163[5:0] };

   // m163_93 = W*in
   wire signed [9:0] m163_93;
   assign m163_93 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_94 = W*in
   wire signed [9:0] m163_94;
   assign m163_94 =10'b0;

   // m163_95 = W*in
   wire signed [9:0] m163_95;
   assign m163_95 =10'b0;

   // m163_96 = W*in
   wire signed [9:0] m163_96;
   assign m163_96 =10'b0;

   // m163_97 = W*in
   wire signed [9:0] m163_97;
   assign m163_97 =10'b0;

   // m163_98 = W*in
   wire signed [9:0] m163_98;
   assign m163_98 =10'b0;

   // m163_99 = W*in
   wire signed [9:0] m163_99;
   assign m163_99 =10'b0;

   // m163_100 = W*in
   wire signed [9:0] m163_100;
   assign m163_100 =10'b0;

   // m163_101 = W*in
   wire signed [9:0] m163_101;
   assign m163_101 =10'b0;

   // m163_102 = W*in
   wire signed [9:0] m163_102;
   assign m163_102 =10'b0;

   // m163_103 = W*in
   wire signed [9:0] m163_103;
   assign m163_103 =10'b0;

   // m163_104 = W*in
   wire signed [9:0] m163_104;
   assign m163_104 =10'b0;

   // m163_105 = W*in
   wire signed [9:0] m163_105;
   assign m163_105 =10'b0;

   // m163_106 = W*in
   wire signed [9:0] m163_106;
   assign m163_106 =10'b0;

   // m163_107 = W*in
   wire signed [9:0] m163_107;
   assign m163_107 ={ {4{in163[5]}} , in163[5:0] };

   // m163_108 = W*in
   wire signed [9:0] m163_108;
   assign m163_108 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_109 = W*in
   wire signed [9:0] m163_109;
   assign m163_109 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_110 = W*in
   wire signed [9:0] m163_110;
   assign m163_110 =10'b0;

   // m163_111 = W*in
   wire signed [9:0] m163_111;
   assign m163_111 =10'b0;

   // m163_112 = W*in
   wire signed [9:0] m163_112;
   assign m163_112 =10'b0;

   // m163_113 = W*in
   wire signed [9:0] m163_113;
   assign m163_113 ={ {4{in163[5]}} , in163[5:0] };

   // m163_114 = W*in
   wire signed [9:0] m163_114;
   assign m163_114 ={ {5{neg163[5]}} , neg163[5:1] };

   // m163_115 = W*in
   wire signed [9:0] m163_115;
   assign m163_115 =10'b0;

   // m163_116 = W*in
   wire signed [9:0] m163_116;
   assign m163_116 ={ {4{neg163[5]}} , neg163[5:0] };

   // m163_117 = W*in
   wire signed [9:0] m163_117;
   assign m163_117 =10'b0;

   // m164_1 = W*in
   wire signed [9:0] m164_1;
   assign m164_1 =10'b0;

   // m164_2 = W*in
   wire signed [9:0] m164_2;
   assign m164_2 =10'b0;

   // m164_3 = W*in
   wire signed [9:0] m164_3;
   assign m164_3 =10'b0;

   // m164_4 = W*in
   wire signed [9:0] m164_4;
   assign m164_4 =10'b0;

   // m164_5 = W*in
   wire signed [9:0] m164_5;
   assign m164_5 =10'b0;

   // m164_6 = W*in
   wire signed [9:0] m164_6;
   assign m164_6 =10'b0;

   // m164_7 = W*in
   wire signed [9:0] m164_7;
   assign m164_7 =10'b0;

   // m164_8 = W*in
   wire signed [9:0] m164_8;
   assign m164_8 =10'b0;

   // m164_9 = W*in
   wire signed [9:0] m164_9;
   assign m164_9 =10'b0;

   // m164_10 = W*in
   wire signed [9:0] m164_10;
   assign m164_10 =10'b0;

   // m164_11 = W*in
   wire signed [9:0] m164_11;
   assign m164_11 =10'b0;

   // m164_12 = W*in
   wire signed [9:0] m164_12;
   assign m164_12 =10'b0;

   // m164_13 = W*in
   wire signed [9:0] m164_13;
   assign m164_13 =10'b0;

   // m164_14 = W*in
   wire signed [9:0] m164_14;
   assign m164_14 =10'b0;

   // m164_15 = W*in
   wire signed [9:0] m164_15;
   assign m164_15 =10'b0;

   // m164_16 = W*in
   wire signed [9:0] m164_16;
   assign m164_16 =10'b0;

   // m164_17 = W*in
   wire signed [9:0] m164_17;
   assign m164_17 =10'b0;

   // m164_18 = W*in
   wire signed [9:0] m164_18;
   assign m164_18 =10'b0;

   // m164_19 = W*in
   wire signed [9:0] m164_19;
   assign m164_19 =10'b0;

   // m164_20 = W*in
   wire signed [9:0] m164_20;
   assign m164_20 =10'b0;

   // m164_21 = W*in
   wire signed [9:0] m164_21;
   assign m164_21 =10'b0;

   // m164_22 = W*in
   wire signed [9:0] m164_22;
   assign m164_22 =10'b0;

   // m164_23 = W*in
   wire signed [9:0] m164_23;
   assign m164_23 =10'b0;

   // m164_24 = W*in
   wire signed [9:0] m164_24;
   assign m164_24 =10'b0;

   // m164_25 = W*in
   wire signed [9:0] m164_25;
   assign m164_25 ={ {4{in164[5]}} , in164[5:0] };

   // m164_26 = W*in
   wire signed [9:0] m164_26;
   assign m164_26 =10'b0;

   // m164_27 = W*in
   wire signed [9:0] m164_27;
   assign m164_27 =10'b0;

   // m164_28 = W*in
   wire signed [9:0] m164_28;
   assign m164_28 ={ {5{in164[5]}} , in164[5:1] };

   // m164_29 = W*in
   wire signed [9:0] m164_29;
   assign m164_29 =10'b0;

   // m164_30 = W*in
   wire signed [9:0] m164_30;
   assign m164_30 =10'b0;

   // m164_31 = W*in
   wire signed [9:0] m164_31;
   assign m164_31 =10'b0;

   // m164_32 = W*in
   wire signed [9:0] m164_32;
   assign m164_32 =10'b0;

   // m164_33 = W*in
   wire signed [9:0] m164_33;
   assign m164_33 =10'b0;

   // m164_34 = W*in
   wire signed [9:0] m164_34;
   assign m164_34 =10'b0;

   // m164_35 = W*in
   wire signed [9:0] m164_35;
   assign m164_35 =10'b0;

   // m164_36 = W*in
   wire signed [9:0] m164_36;
   assign m164_36 =10'b0;

   // m164_37 = W*in
   wire signed [9:0] m164_37;
   assign m164_37 =10'b0;

   // m164_38 = W*in
   wire signed [9:0] m164_38;
   assign m164_38 =10'b0;

   // m164_39 = W*in
   wire signed [9:0] m164_39;
   assign m164_39 =10'b0;

   // m164_40 = W*in
   wire signed [9:0] m164_40;
   assign m164_40 =10'b0;

   // m164_41 = W*in
   wire signed [9:0] m164_41;
   assign m164_41 =10'b0;

   // m164_42 = W*in
   wire signed [9:0] m164_42;
   assign m164_42 =10'b0;

   // m164_43 = W*in
   wire signed [9:0] m164_43;
   assign m164_43 ={ {4{in164[5]}} , in164[5:0] };

   // m164_44 = W*in
   wire signed [9:0] m164_44;
   assign m164_44 =10'b0;

   // m164_45 = W*in
   wire signed [9:0] m164_45;
   assign m164_45 =10'b0;

   // m164_46 = W*in
   wire signed [9:0] m164_46;
   assign m164_46 =10'b0;

   // m164_47 = W*in
   wire signed [9:0] m164_47;
   assign m164_47 =10'b0;

   // m164_48 = W*in
   wire signed [9:0] m164_48;
   assign m164_48 ={ {4{in164[5]}} , in164[5:0] };

   // m164_49 = W*in
   wire signed [9:0] m164_49;
   assign m164_49 =10'b0;

   // m164_50 = W*in
   wire signed [9:0] m164_50;
   assign m164_50 =10'b0;

   // m164_51 = W*in
   wire signed [9:0] m164_51;
   assign m164_51 =10'b0;

   // m164_52 = W*in
   wire signed [9:0] m164_52;
   assign m164_52 =10'b0;

   // m164_53 = W*in
   wire signed [9:0] m164_53;
   assign m164_53 =10'b0;

   // m164_54 = W*in
   wire signed [9:0] m164_54;
   assign m164_54 =10'b0;

   // m164_55 = W*in
   wire signed [9:0] m164_55;
   assign m164_55 =10'b0;

   // m164_56 = W*in
   wire signed [9:0] m164_56;
   assign m164_56 =10'b0;

   // m164_57 = W*in
   wire signed [9:0] m164_57;
   assign m164_57 =10'b0;

   // m164_58 = W*in
   wire signed [9:0] m164_58;
   assign m164_58 =10'b0;

   // m164_59 = W*in
   wire signed [9:0] m164_59;
   assign m164_59 =10'b0;

   // m164_60 = W*in
   wire signed [9:0] m164_60;
   assign m164_60 =10'b0;

   // m164_61 = W*in
   wire signed [9:0] m164_61;
   assign m164_61 =10'b0;

   // m164_62 = W*in
   wire signed [9:0] m164_62;
   assign m164_62 =10'b0;

   // m164_63 = W*in
   wire signed [9:0] m164_63;
   assign m164_63 =10'b0;

   // m164_64 = W*in
   wire signed [9:0] m164_64;
   assign m164_64 =10'b0;

   // m164_65 = W*in
   wire signed [9:0] m164_65;
   assign m164_65 =10'b0;

   // m164_66 = W*in
   wire signed [9:0] m164_66;
   assign m164_66 ={ {5{neg164[5]}} , neg164[5:1] };

   // m164_67 = W*in
   wire signed [9:0] m164_67;
   assign m164_67 =10'b0;

   // m164_68 = W*in
   wire signed [9:0] m164_68;
   assign m164_68 =10'b0;

   // m164_69 = W*in
   wire signed [9:0] m164_69;
   assign m164_69 =10'b0;

   // m164_70 = W*in
   wire signed [9:0] m164_70;
   assign m164_70 =10'b0;

   // m164_71 = W*in
   wire signed [9:0] m164_71;
   assign m164_71 =10'b0;

   // m164_72 = W*in
   wire signed [9:0] m164_72;
   assign m164_72 ={ {5{in164[5]}} , in164[5:1] };

   // m164_73 = W*in
   wire signed [9:0] m164_73;
   assign m164_73 =10'b0;

   // m164_74 = W*in
   wire signed [9:0] m164_74;
   assign m164_74 =10'b0;

   // m164_75 = W*in
   wire signed [9:0] m164_75;
   assign m164_75 =10'b0;

   // m164_76 = W*in
   wire signed [9:0] m164_76;
   assign m164_76 =10'b0;

   // m164_77 = W*in
   wire signed [9:0] m164_77;
   assign m164_77 =10'b0;

   // m164_78 = W*in
   wire signed [9:0] m164_78;
   assign m164_78 ={ {5{in164[5]}} , in164[5:1] };

   // m164_79 = W*in
   wire signed [9:0] m164_79;
   assign m164_79 =10'b0;

   // m164_80 = W*in
   wire signed [9:0] m164_80;
   assign m164_80 =10'b0;

   // m164_81 = W*in
   wire signed [9:0] m164_81;
   assign m164_81 =10'b0;

   // m164_82 = W*in
   wire signed [9:0] m164_82;
   assign m164_82 =10'b0;

   // m164_83 = W*in
   wire signed [9:0] m164_83;
   assign m164_83 =10'b0;

   // m164_84 = W*in
   wire signed [9:0] m164_84;
   assign m164_84 =10'b0;

   // m164_85 = W*in
   wire signed [9:0] m164_85;
   assign m164_85 =10'b0;

   // m164_86 = W*in
   wire signed [9:0] m164_86;
   assign m164_86 =10'b0;

   // m164_87 = W*in
   wire signed [9:0] m164_87;
   assign m164_87 =10'b0;

   // m164_88 = W*in
   wire signed [9:0] m164_88;
   assign m164_88 =10'b0;

   // m164_89 = W*in
   wire signed [9:0] m164_89;
   assign m164_89 =10'b0;

   // m164_90 = W*in
   wire signed [9:0] m164_90;
   assign m164_90 =10'b0;

   // m164_91 = W*in
   wire signed [9:0] m164_91;
   assign m164_91 =10'b0;

   // m164_92 = W*in
   wire signed [9:0] m164_92;
   assign m164_92 =10'b0;

   // m164_93 = W*in
   wire signed [9:0] m164_93;
   assign m164_93 =10'b0;

   // m164_94 = W*in
   wire signed [9:0] m164_94;
   assign m164_94 =10'b0;

   // m164_95 = W*in
   wire signed [9:0] m164_95;
   assign m164_95 =10'b0;

   // m164_96 = W*in
   wire signed [9:0] m164_96;
   assign m164_96 =10'b0;

   // m164_97 = W*in
   wire signed [9:0] m164_97;
   assign m164_97 =10'b0;

   // m164_98 = W*in
   wire signed [9:0] m164_98;
   assign m164_98 =10'b0;

   // m164_99 = W*in
   wire signed [9:0] m164_99;
   assign m164_99 =10'b0;

   // m164_100 = W*in
   wire signed [9:0] m164_100;
   assign m164_100 =10'b0;

   // m164_101 = W*in
   wire signed [9:0] m164_101;
   assign m164_101 =10'b0;

   // m164_102 = W*in
   wire signed [9:0] m164_102;
   assign m164_102 =10'b0;

   // m164_103 = W*in
   wire signed [9:0] m164_103;
   assign m164_103 =10'b0;

   // m164_104 = W*in
   wire signed [9:0] m164_104;
   assign m164_104 =10'b0;

   // m164_105 = W*in
   wire signed [9:0] m164_105;
   assign m164_105 =10'b0;

   // m164_106 = W*in
   wire signed [9:0] m164_106;
   assign m164_106 =10'b0;

   // m164_107 = W*in
   wire signed [9:0] m164_107;
   assign m164_107 =10'b0;

   // m164_108 = W*in
   wire signed [9:0] m164_108;
   assign m164_108 ={ {5{neg164[5]}} , neg164[5:1] };

   // m164_109 = W*in
   wire signed [9:0] m164_109;
   assign m164_109 ={ {5{neg164[5]}} , neg164[5:1] };

   // m164_110 = W*in
   wire signed [9:0] m164_110;
   assign m164_110 =10'b0;

   // m164_111 = W*in
   wire signed [9:0] m164_111;
   assign m164_111 =10'b0;

   // m164_112 = W*in
   wire signed [9:0] m164_112;
   assign m164_112 =10'b0;

   // m164_113 = W*in
   wire signed [9:0] m164_113;
   assign m164_113 =10'b0;

   // m164_114 = W*in
   wire signed [9:0] m164_114;
   assign m164_114 =10'b0;

   // m164_115 = W*in
   wire signed [9:0] m164_115;
   assign m164_115 =10'b0;

   // m164_116 = W*in
   wire signed [9:0] m164_116;
   assign m164_116 =10'b0;

   // m164_117 = W*in
   wire signed [9:0] m164_117;
   assign m164_117 =10'b0;

   // m165_1 = W*in
   wire signed [9:0] m165_1;
   assign m165_1 =10'b0;

   // m165_2 = W*in
   wire signed [9:0] m165_2;
   assign m165_2 =10'b0;

   // m165_3 = W*in
   wire signed [9:0] m165_3;
   assign m165_3 =10'b0;

   // m165_4 = W*in
   wire signed [9:0] m165_4;
   assign m165_4 =10'b0;

   // m165_5 = W*in
   wire signed [9:0] m165_5;
   assign m165_5 =10'b0;

   // m165_6 = W*in
   wire signed [9:0] m165_6;
   assign m165_6 =10'b0;

   // m165_7 = W*in
   wire signed [9:0] m165_7;
   assign m165_7 =10'b0;

   // m165_8 = W*in
   wire signed [9:0] m165_8;
   assign m165_8 =10'b0;

   // m165_9 = W*in
   wire signed [9:0] m165_9;
   assign m165_9 =10'b0;

   // m165_10 = W*in
   wire signed [9:0] m165_10;
   assign m165_10 =10'b0;

   // m165_11 = W*in
   wire signed [9:0] m165_11;
   assign m165_11 =10'b0;

   // m165_12 = W*in
   wire signed [9:0] m165_12;
   assign m165_12 =10'b0;

   // m165_13 = W*in
   wire signed [9:0] m165_13;
   assign m165_13 =10'b0;

   // m165_14 = W*in
   wire signed [9:0] m165_14;
   assign m165_14 =10'b0;

   // m165_15 = W*in
   wire signed [9:0] m165_15;
   assign m165_15 =10'b0;

   // m165_16 = W*in
   wire signed [9:0] m165_16;
   assign m165_16 =10'b0;

   // m165_17 = W*in
   wire signed [9:0] m165_17;
   assign m165_17 =10'b0;

   // m165_18 = W*in
   wire signed [9:0] m165_18;
   assign m165_18 =10'b0;

   // m165_19 = W*in
   wire signed [9:0] m165_19;
   assign m165_19 =10'b0;

   // m165_20 = W*in
   wire signed [9:0] m165_20;
   assign m165_20 ={ {5{in165[5]}} , in165[5:1] };

   // m165_21 = W*in
   wire signed [9:0] m165_21;
   assign m165_21 =10'b0;

   // m165_22 = W*in
   wire signed [9:0] m165_22;
   assign m165_22 ={ {5{neg165[5]}} , neg165[5:1] };

   // m165_23 = W*in
   wire signed [9:0] m165_23;
   assign m165_23 =10'b0;

   // m165_24 = W*in
   wire signed [9:0] m165_24;
   assign m165_24 =10'b0;

   // m165_25 = W*in
   wire signed [9:0] m165_25;
   assign m165_25 =10'b0;

   // m165_26 = W*in
   wire signed [9:0] m165_26;
   assign m165_26 ={ {5{neg165[5]}} , neg165[5:1] };

   // m165_27 = W*in
   wire signed [9:0] m165_27;
   assign m165_27 ={ {5{neg165[5]}} , neg165[5:1] };

   // m165_28 = W*in
   wire signed [9:0] m165_28;
   assign m165_28 =10'b0;

   // m165_29 = W*in
   wire signed [9:0] m165_29;
   assign m165_29 =10'b0;

   // m165_30 = W*in
   wire signed [9:0] m165_30;
   assign m165_30 ={ {4{in165[5]}} , in165[5:0] };

   // m165_31 = W*in
   wire signed [9:0] m165_31;
   assign m165_31 =10'b0;

   // m165_32 = W*in
   wire signed [9:0] m165_32;
   assign m165_32 =10'b0;

   // m165_33 = W*in
   wire signed [9:0] m165_33;
   assign m165_33 =10'b0;

   // m165_34 = W*in
   wire signed [9:0] m165_34;
   assign m165_34 =10'b0;

   // m165_35 = W*in
   wire signed [9:0] m165_35;
   assign m165_35 ={ {5{in165[5]}} , in165[5:1] };

   // m165_36 = W*in
   wire signed [9:0] m165_36;
   assign m165_36 =10'b0;

   // m165_37 = W*in
   wire signed [9:0] m165_37;
   assign m165_37 =10'b0;

   // m165_38 = W*in
   wire signed [9:0] m165_38;
   assign m165_38 =10'b0;

   // m165_39 = W*in
   wire signed [9:0] m165_39;
   assign m165_39 =10'b0;

   // m165_40 = W*in
   wire signed [9:0] m165_40;
   assign m165_40 =10'b0;

   // m165_41 = W*in
   wire signed [9:0] m165_41;
   assign m165_41 =10'b0;

   // m165_42 = W*in
   wire signed [9:0] m165_42;
   assign m165_42 ={ {4{in165[5]}} , in165[5:0] };

   // m165_43 = W*in
   wire signed [9:0] m165_43;
   assign m165_43 =10'b0;

   // m165_44 = W*in
   wire signed [9:0] m165_44;
   assign m165_44 =10'b0;

   // m165_45 = W*in
   wire signed [9:0] m165_45;
   assign m165_45 =10'b0;

   // m165_46 = W*in
   wire signed [9:0] m165_46;
   assign m165_46 =10'b0;

   // m165_47 = W*in
   wire signed [9:0] m165_47;
   assign m165_47 =10'b0;

   // m165_48 = W*in
   wire signed [9:0] m165_48;
   assign m165_48 =10'b0;

   // m165_49 = W*in
   wire signed [9:0] m165_49;
   assign m165_49 =10'b0;

   // m165_50 = W*in
   wire signed [9:0] m165_50;
   assign m165_50 =10'b0;

   // m165_51 = W*in
   wire signed [9:0] m165_51;
   assign m165_51 =10'b0;

   // m165_52 = W*in
   wire signed [9:0] m165_52;
   assign m165_52 =10'b0;

   // m165_53 = W*in
   wire signed [9:0] m165_53;
   assign m165_53 =10'b0;

   // m165_54 = W*in
   wire signed [9:0] m165_54;
   assign m165_54 =10'b0;

   // m165_55 = W*in
   wire signed [9:0] m165_55;
   assign m165_55 =10'b0;

   // m165_56 = W*in
   wire signed [9:0] m165_56;
   assign m165_56 =10'b0;

   // m165_57 = W*in
   wire signed [9:0] m165_57;
   assign m165_57 =10'b0;

   // m165_58 = W*in
   wire signed [9:0] m165_58;
   assign m165_58 =10'b0;

   // m165_59 = W*in
   wire signed [9:0] m165_59;
   assign m165_59 =10'b0;

   // m165_60 = W*in
   wire signed [9:0] m165_60;
   assign m165_60 =10'b0;

   // m165_61 = W*in
   wire signed [9:0] m165_61;
   assign m165_61 =10'b0;

   // m165_62 = W*in
   wire signed [9:0] m165_62;
   assign m165_62 =10'b0;

   // m165_63 = W*in
   wire signed [9:0] m165_63;
   assign m165_63 =10'b0;

   // m165_64 = W*in
   wire signed [9:0] m165_64;
   assign m165_64 ={ {5{in165[5]}} , in165[5:1] };

   // m165_65 = W*in
   wire signed [9:0] m165_65;
   assign m165_65 ={ {5{in165[5]}} , in165[5:1] };

   // m165_66 = W*in
   wire signed [9:0] m165_66;
   assign m165_66 ={ {5{in165[5]}} , in165[5:1] };

   // m165_67 = W*in
   wire signed [9:0] m165_67;
   assign m165_67 =10'b0;

   // m165_68 = W*in
   wire signed [9:0] m165_68;
   assign m165_68 =10'b0;

   // m165_69 = W*in
   wire signed [9:0] m165_69;
   assign m165_69 =10'b0;

   // m165_70 = W*in
   wire signed [9:0] m165_70;
   assign m165_70 =10'b0;

   // m165_71 = W*in
   wire signed [9:0] m165_71;
   assign m165_71 ={ {5{neg165[5]}} , neg165[5:1] };

   // m165_72 = W*in
   wire signed [9:0] m165_72;
   assign m165_72 =10'b0;

   // m165_73 = W*in
   wire signed [9:0] m165_73;
   assign m165_73 =10'b0;

   // m165_74 = W*in
   wire signed [9:0] m165_74;
   assign m165_74 =10'b0;

   // m165_75 = W*in
   wire signed [9:0] m165_75;
   assign m165_75 =10'b0;

   // m165_76 = W*in
   wire signed [9:0] m165_76;
   assign m165_76 =10'b0;

   // m165_77 = W*in
   wire signed [9:0] m165_77;
   assign m165_77 =10'b0;

   // m165_78 = W*in
   wire signed [9:0] m165_78;
   assign m165_78 ={ {5{neg165[5]}} , neg165[5:1] };

   // m165_79 = W*in
   wire signed [9:0] m165_79;
   assign m165_79 =10'b0;

   // m165_80 = W*in
   wire signed [9:0] m165_80;
   assign m165_80 =10'b0;

   // m165_81 = W*in
   wire signed [9:0] m165_81;
   assign m165_81 =10'b0;

   // m165_82 = W*in
   wire signed [9:0] m165_82;
   assign m165_82 =10'b0;

   // m165_83 = W*in
   wire signed [9:0] m165_83;
   assign m165_83 ={ {5{neg165[5]}} , neg165[5:1] };

   // m165_84 = W*in
   wire signed [9:0] m165_84;
   assign m165_84 =10'b0;

   // m165_85 = W*in
   wire signed [9:0] m165_85;
   assign m165_85 =10'b0;

   // m165_86 = W*in
   wire signed [9:0] m165_86;
   assign m165_86 =10'b0;

   // m165_87 = W*in
   wire signed [9:0] m165_87;
   assign m165_87 =10'b0;

   // m165_88 = W*in
   wire signed [9:0] m165_88;
   assign m165_88 =10'b0;

   // m165_89 = W*in
   wire signed [9:0] m165_89;
   assign m165_89 =10'b0;

   // m165_90 = W*in
   wire signed [9:0] m165_90;
   assign m165_90 =10'b0;

   // m165_91 = W*in
   wire signed [9:0] m165_91;
   assign m165_91 =10'b0;

   // m165_92 = W*in
   wire signed [9:0] m165_92;
   assign m165_92 =10'b0;

   // m165_93 = W*in
   wire signed [9:0] m165_93;
   assign m165_93 =10'b0;

   // m165_94 = W*in
   wire signed [9:0] m165_94;
   assign m165_94 ={ {4{in165[5]}} , in165[5:0] };

   // m165_95 = W*in
   wire signed [9:0] m165_95;
   assign m165_95 =10'b0;

   // m165_96 = W*in
   wire signed [9:0] m165_96;
   assign m165_96 =10'b0;

   // m165_97 = W*in
   wire signed [9:0] m165_97;
   assign m165_97 =10'b0;

   // m165_98 = W*in
   wire signed [9:0] m165_98;
   assign m165_98 =10'b0;

   // m165_99 = W*in
   wire signed [9:0] m165_99;
   assign m165_99 =10'b0;

   // m165_100 = W*in
   wire signed [9:0] m165_100;
   assign m165_100 =10'b0;

   // m165_101 = W*in
   wire signed [9:0] m165_101;
   assign m165_101 =10'b0;

   // m165_102 = W*in
   wire signed [9:0] m165_102;
   assign m165_102 =10'b0;

   // m165_103 = W*in
   wire signed [9:0] m165_103;
   assign m165_103 =10'b0;

   // m165_104 = W*in
   wire signed [9:0] m165_104;
   assign m165_104 =10'b0;

   // m165_105 = W*in
   wire signed [9:0] m165_105;
   assign m165_105 =10'b0;

   // m165_106 = W*in
   wire signed [9:0] m165_106;
   assign m165_106 =10'b0;

   // m165_107 = W*in
   wire signed [9:0] m165_107;
   assign m165_107 =10'b0;

   // m165_108 = W*in
   wire signed [9:0] m165_108;
   assign m165_108 ={ {4{in165[5]}} , in165[5:0] };

   // m165_109 = W*in
   wire signed [9:0] m165_109;
   assign m165_109 =10'b0;

   // m165_110 = W*in
   wire signed [9:0] m165_110;
   assign m165_110 =10'b0;

   // m165_111 = W*in
   wire signed [9:0] m165_111;
   assign m165_111 =10'b0;

   // m165_112 = W*in
   wire signed [9:0] m165_112;
   assign m165_112 =10'b0;

   // m165_113 = W*in
   wire signed [9:0] m165_113;
   assign m165_113 =10'b0;

   // m165_114 = W*in
   wire signed [9:0] m165_114;
   assign m165_114 =10'b0;

   // m165_115 = W*in
   wire signed [9:0] m165_115;
   assign m165_115 =10'b0;

   // m165_116 = W*in
   wire signed [9:0] m165_116;
   assign m165_116 ={ {4{in165[5]}} , in165[5:0] };

   // m165_117 = W*in
   wire signed [9:0] m165_117;
   assign m165_117 =10'b0;

   // m166_1 = W*in
   wire signed [9:0] m166_1;
   assign m166_1 ={ {4{in166[5]}} , in166[5:0] };

   // m166_2 = W*in
   wire signed [9:0] m166_2;
   assign m166_2 ={ {4{in166[5]}} , in166[5:0] };

   // m166_3 = W*in
   wire signed [9:0] m166_3;
   assign m166_3 =10'b0;

   // m166_4 = W*in
   wire signed [9:0] m166_4;
   assign m166_4 =10'b0;

   // m166_5 = W*in
   wire signed [9:0] m166_5;
   assign m166_5 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_6 = W*in
   wire signed [9:0] m166_6;
   assign m166_6 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_7 = W*in
   wire signed [9:0] m166_7;
   assign m166_7 =10'b0;

   // m166_8 = W*in
   wire signed [9:0] m166_8;
   assign m166_8 =10'b0;

   // m166_9 = W*in
   wire signed [9:0] m166_9;
   assign m166_9 =10'b0;

   // m166_10 = W*in
   wire signed [9:0] m166_10;
   assign m166_10 =10'b0;

   // m166_11 = W*in
   wire signed [9:0] m166_11;
   assign m166_11 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_12 = W*in
   wire signed [9:0] m166_12;
   assign m166_12 =10'b0;

   // m166_13 = W*in
   wire signed [9:0] m166_13;
   assign m166_13 ={ {4{in166[5]}} , in166[5:0] };

   // m166_14 = W*in
   wire signed [9:0] m166_14;
   assign m166_14 =10'b0;

   // m166_15 = W*in
   wire signed [9:0] m166_15;
   assign m166_15 =10'b0;

   // m166_16 = W*in
   wire signed [9:0] m166_16;
   assign m166_16 ={ {4{in166[5]}} , in166[5:0] };

   // m166_17 = W*in
   wire signed [9:0] m166_17;
   assign m166_17 =10'b0;

   // m166_18 = W*in
   wire signed [9:0] m166_18;
   assign m166_18 =10'b0;

   // m166_19 = W*in
   wire signed [9:0] m166_19;
   assign m166_19 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_20 = W*in
   wire signed [9:0] m166_20;
   assign m166_20 =10'b0;

   // m166_21 = W*in
   wire signed [9:0] m166_21;
   assign m166_21 =10'b0;

   // m166_22 = W*in
   wire signed [9:0] m166_22;
   assign m166_22 =10'b0;

   // m166_23 = W*in
   wire signed [9:0] m166_23;
   assign m166_23 =10'b0;

   // m166_24 = W*in
   wire signed [9:0] m166_24;
   assign m166_24 =10'b0;

   // m166_25 = W*in
   wire signed [9:0] m166_25;
   assign m166_25 =10'b0;

   // m166_26 = W*in
   wire signed [9:0] m166_26;
   assign m166_26 =10'b0;

   // m166_27 = W*in
   wire signed [9:0] m166_27;
   assign m166_27 ={ {5{in166[5]}} , in166[5:1] };

   // m166_28 = W*in
   wire signed [9:0] m166_28;
   assign m166_28 ={ {5{in166[5]}} , in166[5:1] };

   // m166_29 = W*in
   wire signed [9:0] m166_29;
   assign m166_29 =10'b0;

   // m166_30 = W*in
   wire signed [9:0] m166_30;
   assign m166_30 =10'b0;

   // m166_31 = W*in
   wire signed [9:0] m166_31;
   assign m166_31 =10'b0;

   // m166_32 = W*in
   wire signed [9:0] m166_32;
   assign m166_32 =10'b0;

   // m166_33 = W*in
   wire signed [9:0] m166_33;
   assign m166_33 =10'b0;

   // m166_34 = W*in
   wire signed [9:0] m166_34;
   assign m166_34 =10'b0;

   // m166_35 = W*in
   wire signed [9:0] m166_35;
   assign m166_35 ={ {5{neg166[5]}} , neg166[5:1] };

   // m166_36 = W*in
   wire signed [9:0] m166_36;
   assign m166_36 =10'b0;

   // m166_37 = W*in
   wire signed [9:0] m166_37;
   assign m166_37 ={ {4{in166[5]}} , in166[5:0] };

   // m166_38 = W*in
   wire signed [9:0] m166_38;
   assign m166_38 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_39 = W*in
   wire signed [9:0] m166_39;
   assign m166_39 =10'b0;

   // m166_40 = W*in
   wire signed [9:0] m166_40;
   assign m166_40 =10'b0;

   // m166_41 = W*in
   wire signed [9:0] m166_41;
   assign m166_41 ={ {3{in166[5]}} , in166 , {1{1'b0}} };

   // m166_42 = W*in
   wire signed [9:0] m166_42;
   assign m166_42 =10'b0;

   // m166_43 = W*in
   wire signed [9:0] m166_43;
   assign m166_43 =10'b0;

   // m166_44 = W*in
   wire signed [9:0] m166_44;
   assign m166_44 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_45 = W*in
   wire signed [9:0] m166_45;
   assign m166_45 ={ {4{in166[5]}} , in166[5:0] };

   // m166_46 = W*in
   wire signed [9:0] m166_46;
   assign m166_46 =10'b0;

   // m166_47 = W*in
   wire signed [9:0] m166_47;
   assign m166_47 =10'b0;

   // m166_48 = W*in
   wire signed [9:0] m166_48;
   assign m166_48 =10'b0;

   // m166_49 = W*in
   wire signed [9:0] m166_49;
   assign m166_49 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_50 = W*in
   wire signed [9:0] m166_50;
   assign m166_50 =10'b0;

   // m166_51 = W*in
   wire signed [9:0] m166_51;
   assign m166_51 ={ {4{in166[5]}} , in166[5:0] };

   // m166_52 = W*in
   wire signed [9:0] m166_52;
   assign m166_52 =10'b0;

   // m166_53 = W*in
   wire signed [9:0] m166_53;
   assign m166_53 =10'b0;

   // m166_54 = W*in
   wire signed [9:0] m166_54;
   assign m166_54 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_55 = W*in
   wire signed [9:0] m166_55;
   assign m166_55 =10'b0;

   // m166_56 = W*in
   wire signed [9:0] m166_56;
   assign m166_56 ={ {4{in166[5]}} , in166[5:0] };

   // m166_57 = W*in
   wire signed [9:0] m166_57;
   assign m166_57 =10'b0;

   // m166_58 = W*in
   wire signed [9:0] m166_58;
   assign m166_58 ={ {5{neg166[5]}} , neg166[5:1] };

   // m166_59 = W*in
   wire signed [9:0] m166_59;
   assign m166_59 =10'b0;

   // m166_60 = W*in
   wire signed [9:0] m166_60;
   assign m166_60 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_61 = W*in
   wire signed [9:0] m166_61;
   assign m166_61 =10'b0;

   // m166_62 = W*in
   wire signed [9:0] m166_62;
   assign m166_62 =10'b0;

   // m166_63 = W*in
   wire signed [9:0] m166_63;
   assign m166_63 =10'b0;

   // m166_64 = W*in
   wire signed [9:0] m166_64;
   assign m166_64 =10'b0;

   // m166_65 = W*in
   wire signed [9:0] m166_65;
   assign m166_65 =10'b0;

   // m166_66 = W*in
   wire signed [9:0] m166_66;
   assign m166_66 ={ {5{in166[5]}} , in166[5:1] };

   // m166_67 = W*in
   wire signed [9:0] m166_67;
   assign m166_67 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_68 = W*in
   wire signed [9:0] m166_68;
   assign m166_68 =10'b0;

   // m166_69 = W*in
   wire signed [9:0] m166_69;
   assign m166_69 =10'b0;

   // m166_70 = W*in
   wire signed [9:0] m166_70;
   assign m166_70 =10'b0;

   // m166_71 = W*in
   wire signed [9:0] m166_71;
   assign m166_71 ={ {5{neg166[5]}} , neg166[5:1] };

   // m166_72 = W*in
   wire signed [9:0] m166_72;
   assign m166_72 =10'b0;

   // m166_73 = W*in
   wire signed [9:0] m166_73;
   assign m166_73 =10'b0;

   // m166_74 = W*in
   wire signed [9:0] m166_74;
   assign m166_74 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_75 = W*in
   wire signed [9:0] m166_75;
   assign m166_75 ={ {5{neg166[5]}} , neg166[5:1] };

   // m166_76 = W*in
   wire signed [9:0] m166_76;
   assign m166_76 =10'b0;

   // m166_77 = W*in
   wire signed [9:0] m166_77;
   assign m166_77 =10'b0;

   // m166_78 = W*in
   wire signed [9:0] m166_78;
   assign m166_78 =10'b0;

   // m166_79 = W*in
   wire signed [9:0] m166_79;
   assign m166_79 =10'b0;

   // m166_80 = W*in
   wire signed [9:0] m166_80;
   assign m166_80 =10'b0;

   // m166_81 = W*in
   wire signed [9:0] m166_81;
   assign m166_81 =10'b0;

   // m166_82 = W*in
   wire signed [9:0] m166_82;
   assign m166_82 =10'b0;

   // m166_83 = W*in
   wire signed [9:0] m166_83;
   assign m166_83 =10'b0;

   // m166_84 = W*in
   wire signed [9:0] m166_84;
   assign m166_84 =10'b0;

   // m166_85 = W*in
   wire signed [9:0] m166_85;
   assign m166_85 ={ {4{in166[5]}} , in166[5:0] };

   // m166_86 = W*in
   wire signed [9:0] m166_86;
   assign m166_86 =10'b0;

   // m166_87 = W*in
   wire signed [9:0] m166_87;
   assign m166_87 =10'b0;

   // m166_88 = W*in
   wire signed [9:0] m166_88;
   assign m166_88 =10'b0;

   // m166_89 = W*in
   wire signed [9:0] m166_89;
   assign m166_89 ={ {4{in166[5]}} , in166[5:0] };

   // m166_90 = W*in
   wire signed [9:0] m166_90;
   assign m166_90 =10'b0;

   // m166_91 = W*in
   wire signed [9:0] m166_91;
   assign m166_91 =10'b0;

   // m166_92 = W*in
   wire signed [9:0] m166_92;
   assign m166_92 =10'b0;

   // m166_93 = W*in
   wire signed [9:0] m166_93;
   assign m166_93 =10'b0;

   // m166_94 = W*in
   wire signed [9:0] m166_94;
   assign m166_94 ={ {4{in166[5]}} , in166[5:0] };

   // m166_95 = W*in
   wire signed [9:0] m166_95;
   assign m166_95 =10'b0;

   // m166_96 = W*in
   wire signed [9:0] m166_96;
   assign m166_96 ={ {4{in166[5]}} , in166[5:0] };

   // m166_97 = W*in
   wire signed [9:0] m166_97;
   assign m166_97 =10'b0;

   // m166_98 = W*in
   wire signed [9:0] m166_98;
   assign m166_98 =10'b0;

   // m166_99 = W*in
   wire signed [9:0] m166_99;
   assign m166_99 =10'b0;

   // m166_100 = W*in
   wire signed [9:0] m166_100;
   assign m166_100 =10'b0;

   // m166_101 = W*in
   wire signed [9:0] m166_101;
   assign m166_101 =10'b0;

   // m166_102 = W*in
   wire signed [9:0] m166_102;
   assign m166_102 =10'b0;

   // m166_103 = W*in
   wire signed [9:0] m166_103;
   assign m166_103 =10'b0;

   // m166_104 = W*in
   wire signed [9:0] m166_104;
   assign m166_104 =10'b0;

   // m166_105 = W*in
   wire signed [9:0] m166_105;
   assign m166_105 =10'b0;

   // m166_106 = W*in
   wire signed [9:0] m166_106;
   assign m166_106 =10'b0;

   // m166_107 = W*in
   wire signed [9:0] m166_107;
   assign m166_107 =10'b0;

   // m166_108 = W*in
   wire signed [9:0] m166_108;
   assign m166_108 ={ {4{in166[5]}} , in166[5:0] };

   // m166_109 = W*in
   wire signed [9:0] m166_109;
   assign m166_109 ={ {4{in166[5]}} , in166[5:0] };

   // m166_110 = W*in
   wire signed [9:0] m166_110;
   assign m166_110 ={ {4{neg166[5]}} , neg166[5:0] };

   // m166_111 = W*in
   wire signed [9:0] m166_111;
   assign m166_111 =10'b0;

   // m166_112 = W*in
   wire signed [9:0] m166_112;
   assign m166_112 =10'b0;

   // m166_113 = W*in
   wire signed [9:0] m166_113;
   assign m166_113 =10'b0;

   // m166_114 = W*in
   wire signed [9:0] m166_114;
   assign m166_114 ={ {5{neg166[5]}} , neg166[5:1] };

   // m166_115 = W*in
   wire signed [9:0] m166_115;
   assign m166_115 =10'b0;

   // m166_116 = W*in
   wire signed [9:0] m166_116;
   assign m166_116 ={ {4{in166[5]}} , in166[5:0] };

   // m166_117 = W*in
   wire signed [9:0] m166_117;
   assign m166_117 =10'b0;

   // m167_1 = W*in
   wire signed [9:0] m167_1;
   assign m167_1 =10'b0;

   // m167_2 = W*in
   wire signed [9:0] m167_2;
   assign m167_2 =10'b0;

   // m167_3 = W*in
   wire signed [9:0] m167_3;
   assign m167_3 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_4 = W*in
   wire signed [9:0] m167_4;
   assign m167_4 =10'b0;

   // m167_5 = W*in
   wire signed [9:0] m167_5;
   assign m167_5 =10'b0;

   // m167_6 = W*in
   wire signed [9:0] m167_6;
   assign m167_6 =10'b0;

   // m167_7 = W*in
   wire signed [9:0] m167_7;
   assign m167_7 =10'b0;

   // m167_8 = W*in
   wire signed [9:0] m167_8;
   assign m167_8 =10'b0;

   // m167_9 = W*in
   wire signed [9:0] m167_9;
   assign m167_9 =10'b0;

   // m167_10 = W*in
   wire signed [9:0] m167_10;
   assign m167_10 ={ {4{in167[5]}} , in167[5:0] };

   // m167_11 = W*in
   wire signed [9:0] m167_11;
   assign m167_11 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_12 = W*in
   wire signed [9:0] m167_12;
   assign m167_12 =10'b0;

   // m167_13 = W*in
   wire signed [9:0] m167_13;
   assign m167_13 ={ {4{in167[5]}} , in167[5:0] };

   // m167_14 = W*in
   wire signed [9:0] m167_14;
   assign m167_14 =10'b0;

   // m167_15 = W*in
   wire signed [9:0] m167_15;
   assign m167_15 =10'b0;

   // m167_16 = W*in
   wire signed [9:0] m167_16;
   assign m167_16 =10'b0;

   // m167_17 = W*in
   wire signed [9:0] m167_17;
   assign m167_17 =10'b0;

   // m167_18 = W*in
   wire signed [9:0] m167_18;
   assign m167_18 =10'b0;

   // m167_19 = W*in
   wire signed [9:0] m167_19;
   assign m167_19 ={ {5{neg167[5]}} , neg167[5:1] };

   // m167_20 = W*in
   wire signed [9:0] m167_20;
   assign m167_20 =10'b0;

   // m167_21 = W*in
   wire signed [9:0] m167_21;
   assign m167_21 =10'b0;

   // m167_22 = W*in
   wire signed [9:0] m167_22;
   assign m167_22 =10'b0;

   // m167_23 = W*in
   wire signed [9:0] m167_23;
   assign m167_23 =10'b0;

   // m167_24 = W*in
   wire signed [9:0] m167_24;
   assign m167_24 =10'b0;

   // m167_25 = W*in
   wire signed [9:0] m167_25;
   assign m167_25 =10'b0;

   // m167_26 = W*in
   wire signed [9:0] m167_26;
   assign m167_26 =10'b0;

   // m167_27 = W*in
   wire signed [9:0] m167_27;
   assign m167_27 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_28 = W*in
   wire signed [9:0] m167_28;
   assign m167_28 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_29 = W*in
   wire signed [9:0] m167_29;
   assign m167_29 =10'b0;

   // m167_30 = W*in
   wire signed [9:0] m167_30;
   assign m167_30 =10'b0;

   // m167_31 = W*in
   wire signed [9:0] m167_31;
   assign m167_31 =10'b0;

   // m167_32 = W*in
   wire signed [9:0] m167_32;
   assign m167_32 =10'b0;

   // m167_33 = W*in
   wire signed [9:0] m167_33;
   assign m167_33 =10'b0;

   // m167_34 = W*in
   wire signed [9:0] m167_34;
   assign m167_34 =10'b0;

   // m167_35 = W*in
   wire signed [9:0] m167_35;
   assign m167_35 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_36 = W*in
   wire signed [9:0] m167_36;
   assign m167_36 =10'b0;

   // m167_37 = W*in
   wire signed [9:0] m167_37;
   assign m167_37 =10'b0;

   // m167_38 = W*in
   wire signed [9:0] m167_38;
   assign m167_38 =10'b0;

   // m167_39 = W*in
   wire signed [9:0] m167_39;
   assign m167_39 =10'b0;

   // m167_40 = W*in
   wire signed [9:0] m167_40;
   assign m167_40 =10'b0;

   // m167_41 = W*in
   wire signed [9:0] m167_41;
   assign m167_41 =10'b0;

   // m167_42 = W*in
   wire signed [9:0] m167_42;
   assign m167_42 =10'b0;

   // m167_43 = W*in
   wire signed [9:0] m167_43;
   assign m167_43 =10'b0;

   // m167_44 = W*in
   wire signed [9:0] m167_44;
   assign m167_44 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_45 = W*in
   wire signed [9:0] m167_45;
   assign m167_45 ={ {4{in167[5]}} , in167[5:0] };

   // m167_46 = W*in
   wire signed [9:0] m167_46;
   assign m167_46 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_47 = W*in
   wire signed [9:0] m167_47;
   assign m167_47 =10'b0;

   // m167_48 = W*in
   wire signed [9:0] m167_48;
   assign m167_48 =10'b0;

   // m167_49 = W*in
   wire signed [9:0] m167_49;
   assign m167_49 =10'b0;

   // m167_50 = W*in
   wire signed [9:0] m167_50;
   assign m167_50 =10'b0;

   // m167_51 = W*in
   wire signed [9:0] m167_51;
   assign m167_51 ={ {4{in167[5]}} , in167[5:0] };

   // m167_52 = W*in
   wire signed [9:0] m167_52;
   assign m167_52 =10'b0;

   // m167_53 = W*in
   wire signed [9:0] m167_53;
   assign m167_53 =10'b0;

   // m167_54 = W*in
   wire signed [9:0] m167_54;
   assign m167_54 =10'b0;

   // m167_55 = W*in
   wire signed [9:0] m167_55;
   assign m167_55 =10'b0;

   // m167_56 = W*in
   wire signed [9:0] m167_56;
   assign m167_56 =10'b0;

   // m167_57 = W*in
   wire signed [9:0] m167_57;
   assign m167_57 =10'b0;

   // m167_58 = W*in
   wire signed [9:0] m167_58;
   assign m167_58 =10'b0;

   // m167_59 = W*in
   wire signed [9:0] m167_59;
   assign m167_59 =10'b0;

   // m167_60 = W*in
   wire signed [9:0] m167_60;
   assign m167_60 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_61 = W*in
   wire signed [9:0] m167_61;
   assign m167_61 =10'b0;

   // m167_62 = W*in
   wire signed [9:0] m167_62;
   assign m167_62 =10'b0;

   // m167_63 = W*in
   wire signed [9:0] m167_63;
   assign m167_63 =10'b0;

   // m167_64 = W*in
   wire signed [9:0] m167_64;
   assign m167_64 =10'b0;

   // m167_65 = W*in
   wire signed [9:0] m167_65;
   assign m167_65 =10'b0;

   // m167_66 = W*in
   wire signed [9:0] m167_66;
   assign m167_66 ={ {5{neg167[5]}} , neg167[5:1] };

   // m167_67 = W*in
   wire signed [9:0] m167_67;
   assign m167_67 =10'b0;

   // m167_68 = W*in
   wire signed [9:0] m167_68;
   assign m167_68 =10'b0;

   // m167_69 = W*in
   wire signed [9:0] m167_69;
   assign m167_69 ={ {5{neg167[5]}} , neg167[5:1] };

   // m167_70 = W*in
   wire signed [9:0] m167_70;
   assign m167_70 =10'b0;

   // m167_71 = W*in
   wire signed [9:0] m167_71;
   assign m167_71 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_72 = W*in
   wire signed [9:0] m167_72;
   assign m167_72 =10'b0;

   // m167_73 = W*in
   wire signed [9:0] m167_73;
   assign m167_73 =10'b0;

   // m167_74 = W*in
   wire signed [9:0] m167_74;
   assign m167_74 =10'b0;

   // m167_75 = W*in
   wire signed [9:0] m167_75;
   assign m167_75 =10'b0;

   // m167_76 = W*in
   wire signed [9:0] m167_76;
   assign m167_76 =10'b0;

   // m167_77 = W*in
   wire signed [9:0] m167_77;
   assign m167_77 =10'b0;

   // m167_78 = W*in
   wire signed [9:0] m167_78;
   assign m167_78 =10'b0;

   // m167_79 = W*in
   wire signed [9:0] m167_79;
   assign m167_79 =10'b0;

   // m167_80 = W*in
   wire signed [9:0] m167_80;
   assign m167_80 =10'b0;

   // m167_81 = W*in
   wire signed [9:0] m167_81;
   assign m167_81 =10'b0;

   // m167_82 = W*in
   wire signed [9:0] m167_82;
   assign m167_82 ={ {5{neg167[5]}} , neg167[5:1] };

   // m167_83 = W*in
   wire signed [9:0] m167_83;
   assign m167_83 ={ {5{in167[5]}} , in167[5:1] };

   // m167_84 = W*in
   wire signed [9:0] m167_84;
   assign m167_84 =10'b0;

   // m167_85 = W*in
   wire signed [9:0] m167_85;
   assign m167_85 ={ {4{in167[5]}} , in167[5:0] };

   // m167_86 = W*in
   wire signed [9:0] m167_86;
   assign m167_86 =10'b0;

   // m167_87 = W*in
   wire signed [9:0] m167_87;
   assign m167_87 =10'b0;

   // m167_88 = W*in
   wire signed [9:0] m167_88;
   assign m167_88 =10'b0;

   // m167_89 = W*in
   wire signed [9:0] m167_89;
   assign m167_89 =10'b0;

   // m167_90 = W*in
   wire signed [9:0] m167_90;
   assign m167_90 =10'b0;

   // m167_91 = W*in
   wire signed [9:0] m167_91;
   assign m167_91 =10'b0;

   // m167_92 = W*in
   wire signed [9:0] m167_92;
   assign m167_92 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_93 = W*in
   wire signed [9:0] m167_93;
   assign m167_93 =10'b0;

   // m167_94 = W*in
   wire signed [9:0] m167_94;
   assign m167_94 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_95 = W*in
   wire signed [9:0] m167_95;
   assign m167_95 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_96 = W*in
   wire signed [9:0] m167_96;
   assign m167_96 =10'b0;

   // m167_97 = W*in
   wire signed [9:0] m167_97;
   assign m167_97 =10'b0;

   // m167_98 = W*in
   wire signed [9:0] m167_98;
   assign m167_98 =10'b0;

   // m167_99 = W*in
   wire signed [9:0] m167_99;
   assign m167_99 =10'b0;

   // m167_100 = W*in
   wire signed [9:0] m167_100;
   assign m167_100 =10'b0;

   // m167_101 = W*in
   wire signed [9:0] m167_101;
   assign m167_101 =10'b0;

   // m167_102 = W*in
   wire signed [9:0] m167_102;
   assign m167_102 =10'b0;

   // m167_103 = W*in
   wire signed [9:0] m167_103;
   assign m167_103 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_104 = W*in
   wire signed [9:0] m167_104;
   assign m167_104 ={ {4{neg167[5]}} , neg167[5:0] };

   // m167_105 = W*in
   wire signed [9:0] m167_105;
   assign m167_105 =10'b0;

   // m167_106 = W*in
   wire signed [9:0] m167_106;
   assign m167_106 =10'b0;

   // m167_107 = W*in
   wire signed [9:0] m167_107;
   assign m167_107 =10'b0;

   // m167_108 = W*in
   wire signed [9:0] m167_108;
   assign m167_108 =10'b0;

   // m167_109 = W*in
   wire signed [9:0] m167_109;
   assign m167_109 =10'b0;

   // m167_110 = W*in
   wire signed [9:0] m167_110;
   assign m167_110 =10'b0;

   // m167_111 = W*in
   wire signed [9:0] m167_111;
   assign m167_111 =10'b0;

   // m167_112 = W*in
   wire signed [9:0] m167_112;
   assign m167_112 =10'b0;

   // m167_113 = W*in
   wire signed [9:0] m167_113;
   assign m167_113 =10'b0;

   // m167_114 = W*in
   wire signed [9:0] m167_114;
   assign m167_114 =10'b0;

   // m167_115 = W*in
   wire signed [9:0] m167_115;
   assign m167_115 =10'b0;

   // m167_116 = W*in
   wire signed [9:0] m167_116;
   assign m167_116 ={ {4{in167[5]}} , in167[5:0] };

   // m167_117 = W*in
   wire signed [9:0] m167_117;
   assign m167_117 ={ {4{neg167[5]}} , neg167[5:0] };

   // m168_1 = W*in
   wire signed [9:0] m168_1;
   assign m168_1 =10'b0;

   // m168_2 = W*in
   wire signed [9:0] m168_2;
   assign m168_2 =10'b0;

   // m168_3 = W*in
   wire signed [9:0] m168_3;
   assign m168_3 =10'b0;

   // m168_4 = W*in
   wire signed [9:0] m168_4;
   assign m168_4 =10'b0;

   // m168_5 = W*in
   wire signed [9:0] m168_5;
   assign m168_5 =10'b0;

   // m168_6 = W*in
   wire signed [9:0] m168_6;
   assign m168_6 =10'b0;

   // m168_7 = W*in
   wire signed [9:0] m168_7;
   assign m168_7 =10'b0;

   // m168_8 = W*in
   wire signed [9:0] m168_8;
   assign m168_8 =10'b0;

   // m168_9 = W*in
   wire signed [9:0] m168_9;
   assign m168_9 =10'b0;

   // m168_10 = W*in
   wire signed [9:0] m168_10;
   assign m168_10 =10'b0;

   // m168_11 = W*in
   wire signed [9:0] m168_11;
   assign m168_11 =10'b0;

   // m168_12 = W*in
   wire signed [9:0] m168_12;
   assign m168_12 =10'b0;

   // m168_13 = W*in
   wire signed [9:0] m168_13;
   assign m168_13 =10'b0;

   // m168_14 = W*in
   wire signed [9:0] m168_14;
   assign m168_14 =10'b0;

   // m168_15 = W*in
   wire signed [9:0] m168_15;
   assign m168_15 =10'b0;

   // m168_16 = W*in
   wire signed [9:0] m168_16;
   assign m168_16 =10'b0;

   // m168_17 = W*in
   wire signed [9:0] m168_17;
   assign m168_17 ={ {5{neg168[5]}} , neg168[5:1] };

   // m168_18 = W*in
   wire signed [9:0] m168_18;
   assign m168_18 =10'b0;

   // m168_19 = W*in
   wire signed [9:0] m168_19;
   assign m168_19 ={ {5{neg168[5]}} , neg168[5:1] };

   // m168_20 = W*in
   wire signed [9:0] m168_20;
   assign m168_20 =10'b0;

   // m168_21 = W*in
   wire signed [9:0] m168_21;
   assign m168_21 =10'b0;

   // m168_22 = W*in
   wire signed [9:0] m168_22;
   assign m168_22 =10'b0;

   // m168_23 = W*in
   wire signed [9:0] m168_23;
   assign m168_23 ={ {5{in168[5]}} , in168[5:1] };

   // m168_24 = W*in
   wire signed [9:0] m168_24;
   assign m168_24 =10'b0;

   // m168_25 = W*in
   wire signed [9:0] m168_25;
   assign m168_25 =10'b0;

   // m168_26 = W*in
   wire signed [9:0] m168_26;
   assign m168_26 =10'b0;

   // m168_27 = W*in
   wire signed [9:0] m168_27;
   assign m168_27 =10'b0;

   // m168_28 = W*in
   wire signed [9:0] m168_28;
   assign m168_28 ={ {5{neg168[5]}} , neg168[5:1] };

   // m168_29 = W*in
   wire signed [9:0] m168_29;
   assign m168_29 =10'b0;

   // m168_30 = W*in
   wire signed [9:0] m168_30;
   assign m168_30 =10'b0;

   // m168_31 = W*in
   wire signed [9:0] m168_31;
   assign m168_31 =10'b0;

   // m168_32 = W*in
   wire signed [9:0] m168_32;
   assign m168_32 =10'b0;

   // m168_33 = W*in
   wire signed [9:0] m168_33;
   assign m168_33 =10'b0;

   // m168_34 = W*in
   wire signed [9:0] m168_34;
   assign m168_34 =10'b0;

   // m168_35 = W*in
   wire signed [9:0] m168_35;
   assign m168_35 ={ {5{neg168[5]}} , neg168[5:1] };

   // m168_36 = W*in
   wire signed [9:0] m168_36;
   assign m168_36 =10'b0;

   // m168_37 = W*in
   wire signed [9:0] m168_37;
   assign m168_37 =10'b0;

   // m168_38 = W*in
   wire signed [9:0] m168_38;
   assign m168_38 =10'b0;

   // m168_39 = W*in
   wire signed [9:0] m168_39;
   assign m168_39 =10'b0;

   // m168_40 = W*in
   wire signed [9:0] m168_40;
   assign m168_40 =10'b0;

   // m168_41 = W*in
   wire signed [9:0] m168_41;
   assign m168_41 =10'b0;

   // m168_42 = W*in
   wire signed [9:0] m168_42;
   assign m168_42 =10'b0;

   // m168_43 = W*in
   wire signed [9:0] m168_43;
   assign m168_43 =10'b0;

   // m168_44 = W*in
   wire signed [9:0] m168_44;
   assign m168_44 =10'b0;

   // m168_45 = W*in
   wire signed [9:0] m168_45;
   assign m168_45 ={ {4{in168[5]}} , in168[5:0] };

   // m168_46 = W*in
   wire signed [9:0] m168_46;
   assign m168_46 =10'b0;

   // m168_47 = W*in
   wire signed [9:0] m168_47;
   assign m168_47 =10'b0;

   // m168_48 = W*in
   wire signed [9:0] m168_48;
   assign m168_48 =10'b0;

   // m168_49 = W*in
   wire signed [9:0] m168_49;
   assign m168_49 =10'b0;

   // m168_50 = W*in
   wire signed [9:0] m168_50;
   assign m168_50 =10'b0;

   // m168_51 = W*in
   wire signed [9:0] m168_51;
   assign m168_51 =10'b0;

   // m168_52 = W*in
   wire signed [9:0] m168_52;
   assign m168_52 =10'b0;

   // m168_53 = W*in
   wire signed [9:0] m168_53;
   assign m168_53 =10'b0;

   // m168_54 = W*in
   wire signed [9:0] m168_54;
   assign m168_54 =10'b0;

   // m168_55 = W*in
   wire signed [9:0] m168_55;
   assign m168_55 =10'b0;

   // m168_56 = W*in
   wire signed [9:0] m168_56;
   assign m168_56 =10'b0;

   // m168_57 = W*in
   wire signed [9:0] m168_57;
   assign m168_57 =10'b0;

   // m168_58 = W*in
   wire signed [9:0] m168_58;
   assign m168_58 =10'b0;

   // m168_59 = W*in
   wire signed [9:0] m168_59;
   assign m168_59 =10'b0;

   // m168_60 = W*in
   wire signed [9:0] m168_60;
   assign m168_60 ={ {4{neg168[5]}} , neg168[5:0] };

   // m168_61 = W*in
   wire signed [9:0] m168_61;
   assign m168_61 =10'b0;

   // m168_62 = W*in
   wire signed [9:0] m168_62;
   assign m168_62 =10'b0;

   // m168_63 = W*in
   wire signed [9:0] m168_63;
   assign m168_63 =10'b0;

   // m168_64 = W*in
   wire signed [9:0] m168_64;
   assign m168_64 =10'b0;

   // m168_65 = W*in
   wire signed [9:0] m168_65;
   assign m168_65 =10'b0;

   // m168_66 = W*in
   wire signed [9:0] m168_66;
   assign m168_66 =10'b0;

   // m168_67 = W*in
   wire signed [9:0] m168_67;
   assign m168_67 =10'b0;

   // m168_68 = W*in
   wire signed [9:0] m168_68;
   assign m168_68 =10'b0;

   // m168_69 = W*in
   wire signed [9:0] m168_69;
   assign m168_69 ={ {5{in168[5]}} , in168[5:1] };

   // m168_70 = W*in
   wire signed [9:0] m168_70;
   assign m168_70 =10'b0;

   // m168_71 = W*in
   wire signed [9:0] m168_71;
   assign m168_71 =10'b0;

   // m168_72 = W*in
   wire signed [9:0] m168_72;
   assign m168_72 =10'b0;

   // m168_73 = W*in
   wire signed [9:0] m168_73;
   assign m168_73 =10'b0;

   // m168_74 = W*in
   wire signed [9:0] m168_74;
   assign m168_74 =10'b0;

   // m168_75 = W*in
   wire signed [9:0] m168_75;
   assign m168_75 =10'b0;

   // m168_76 = W*in
   wire signed [9:0] m168_76;
   assign m168_76 =10'b0;

   // m168_77 = W*in
   wire signed [9:0] m168_77;
   assign m168_77 =10'b0;

   // m168_78 = W*in
   wire signed [9:0] m168_78;
   assign m168_78 ={ {5{in168[5]}} , in168[5:1] };

   // m168_79 = W*in
   wire signed [9:0] m168_79;
   assign m168_79 =10'b0;

   // m168_80 = W*in
   wire signed [9:0] m168_80;
   assign m168_80 =10'b0;

   // m168_81 = W*in
   wire signed [9:0] m168_81;
   assign m168_81 =10'b0;

   // m168_82 = W*in
   wire signed [9:0] m168_82;
   assign m168_82 =10'b0;

   // m168_83 = W*in
   wire signed [9:0] m168_83;
   assign m168_83 ={ {5{in168[5]}} , in168[5:1] };

   // m168_84 = W*in
   wire signed [9:0] m168_84;
   assign m168_84 =10'b0;

   // m168_85 = W*in
   wire signed [9:0] m168_85;
   assign m168_85 =10'b0;

   // m168_86 = W*in
   wire signed [9:0] m168_86;
   assign m168_86 =10'b0;

   // m168_87 = W*in
   wire signed [9:0] m168_87;
   assign m168_87 =10'b0;

   // m168_88 = W*in
   wire signed [9:0] m168_88;
   assign m168_88 =10'b0;

   // m168_89 = W*in
   wire signed [9:0] m168_89;
   assign m168_89 =10'b0;

   // m168_90 = W*in
   wire signed [9:0] m168_90;
   assign m168_90 =10'b0;

   // m168_91 = W*in
   wire signed [9:0] m168_91;
   assign m168_91 =10'b0;

   // m168_92 = W*in
   wire signed [9:0] m168_92;
   assign m168_92 =10'b0;

   // m168_93 = W*in
   wire signed [9:0] m168_93;
   assign m168_93 =10'b0;

   // m168_94 = W*in
   wire signed [9:0] m168_94;
   assign m168_94 =10'b0;

   // m168_95 = W*in
   wire signed [9:0] m168_95;
   assign m168_95 =10'b0;

   // m168_96 = W*in
   wire signed [9:0] m168_96;
   assign m168_96 =10'b0;

   // m168_97 = W*in
   wire signed [9:0] m168_97;
   assign m168_97 ={ {4{neg168[5]}} , neg168[5:0] };

   // m168_98 = W*in
   wire signed [9:0] m168_98;
   assign m168_98 =10'b0;

   // m168_99 = W*in
   wire signed [9:0] m168_99;
   assign m168_99 =10'b0;

   // m168_100 = W*in
   wire signed [9:0] m168_100;
   assign m168_100 =10'b0;

   // m168_101 = W*in
   wire signed [9:0] m168_101;
   assign m168_101 =10'b0;

   // m168_102 = W*in
   wire signed [9:0] m168_102;
   assign m168_102 =10'b0;

   // m168_103 = W*in
   wire signed [9:0] m168_103;
   assign m168_103 =10'b0;

   // m168_104 = W*in
   wire signed [9:0] m168_104;
   assign m168_104 =10'b0;

   // m168_105 = W*in
   wire signed [9:0] m168_105;
   assign m168_105 =10'b0;

   // m168_106 = W*in
   wire signed [9:0] m168_106;
   assign m168_106 =10'b0;

   // m168_107 = W*in
   wire signed [9:0] m168_107;
   assign m168_107 =10'b0;

   // m168_108 = W*in
   wire signed [9:0] m168_108;
   assign m168_108 =10'b0;

   // m168_109 = W*in
   wire signed [9:0] m168_109;
   assign m168_109 ={ {5{in168[5]}} , in168[5:1] };

   // m168_110 = W*in
   wire signed [9:0] m168_110;
   assign m168_110 ={ {4{neg168[5]}} , neg168[5:0] };

   // m168_111 = W*in
   wire signed [9:0] m168_111;
   assign m168_111 =10'b0;

   // m168_112 = W*in
   wire signed [9:0] m168_112;
   assign m168_112 =10'b0;

   // m168_113 = W*in
   wire signed [9:0] m168_113;
   assign m168_113 =10'b0;

   // m168_114 = W*in
   wire signed [9:0] m168_114;
   assign m168_114 =10'b0;

   // m168_115 = W*in
   wire signed [9:0] m168_115;
   assign m168_115 =10'b0;

   // m168_116 = W*in
   wire signed [9:0] m168_116;
   assign m168_116 =10'b0;

   // m168_117 = W*in
   wire signed [9:0] m168_117;
   assign m168_117 =10'b0;

   // m169_1 = W*in
   wire signed [9:0] m169_1;
   assign m169_1 =10'b0;

   // m169_2 = W*in
   wire signed [9:0] m169_2;
   assign m169_2 =10'b0;

   // m169_3 = W*in
   wire signed [9:0] m169_3;
   assign m169_3 =10'b0;

   // m169_4 = W*in
   wire signed [9:0] m169_4;
   assign m169_4 =10'b0;

   // m169_5 = W*in
   wire signed [9:0] m169_5;
   assign m169_5 =10'b0;

   // m169_6 = W*in
   wire signed [9:0] m169_6;
   assign m169_6 =10'b0;

   // m169_7 = W*in
   wire signed [9:0] m169_7;
   assign m169_7 =10'b0;

   // m169_8 = W*in
   wire signed [9:0] m169_8;
   assign m169_8 =10'b0;

   // m169_9 = W*in
   wire signed [9:0] m169_9;
   assign m169_9 =10'b0;

   // m169_10 = W*in
   wire signed [9:0] m169_10;
   assign m169_10 =10'b0;

   // m169_11 = W*in
   wire signed [9:0] m169_11;
   assign m169_11 =10'b0;

   // m169_12 = W*in
   wire signed [9:0] m169_12;
   assign m169_12 =10'b0;

   // m169_13 = W*in
   wire signed [9:0] m169_13;
   assign m169_13 =10'b0;

   // m169_14 = W*in
   wire signed [9:0] m169_14;
   assign m169_14 =10'b0;

   // m169_15 = W*in
   wire signed [9:0] m169_15;
   assign m169_15 =10'b0;

   // m169_16 = W*in
   wire signed [9:0] m169_16;
   assign m169_16 =10'b0;

   // m169_17 = W*in
   wire signed [9:0] m169_17;
   assign m169_17 =10'b0;

   // m169_18 = W*in
   wire signed [9:0] m169_18;
   assign m169_18 =10'b0;

   // m169_19 = W*in
   wire signed [9:0] m169_19;
   assign m169_19 =10'b0;

   // m169_20 = W*in
   wire signed [9:0] m169_20;
   assign m169_20 =10'b0;

   // m169_21 = W*in
   wire signed [9:0] m169_21;
   assign m169_21 =10'b0;

   // m169_22 = W*in
   wire signed [9:0] m169_22;
   assign m169_22 =10'b0;

   // m169_23 = W*in
   wire signed [9:0] m169_23;
   assign m169_23 =10'b0;

   // m169_24 = W*in
   wire signed [9:0] m169_24;
   assign m169_24 =10'b0;

   // m169_25 = W*in
   wire signed [9:0] m169_25;
   assign m169_25 =10'b0;

   // m169_26 = W*in
   wire signed [9:0] m169_26;
   assign m169_26 =10'b0;

   // m169_27 = W*in
   wire signed [9:0] m169_27;
   assign m169_27 ={ {5{in169[5]}} , in169[5:1] };

   // m169_28 = W*in
   wire signed [9:0] m169_28;
   assign m169_28 =10'b0;

   // m169_29 = W*in
   wire signed [9:0] m169_29;
   assign m169_29 =10'b0;

   // m169_30 = W*in
   wire signed [9:0] m169_30;
   assign m169_30 =10'b0;

   // m169_31 = W*in
   wire signed [9:0] m169_31;
   assign m169_31 =10'b0;

   // m169_32 = W*in
   wire signed [9:0] m169_32;
   assign m169_32 =10'b0;

   // m169_33 = W*in
   wire signed [9:0] m169_33;
   assign m169_33 =10'b0;

   // m169_34 = W*in
   wire signed [9:0] m169_34;
   assign m169_34 =10'b0;

   // m169_35 = W*in
   wire signed [9:0] m169_35;
   assign m169_35 =10'b0;

   // m169_36 = W*in
   wire signed [9:0] m169_36;
   assign m169_36 =10'b0;

   // m169_37 = W*in
   wire signed [9:0] m169_37;
   assign m169_37 =10'b0;

   // m169_38 = W*in
   wire signed [9:0] m169_38;
   assign m169_38 =10'b0;

   // m169_39 = W*in
   wire signed [9:0] m169_39;
   assign m169_39 =10'b0;

   // m169_40 = W*in
   wire signed [9:0] m169_40;
   assign m169_40 =10'b0;

   // m169_41 = W*in
   wire signed [9:0] m169_41;
   assign m169_41 =10'b0;

   // m169_42 = W*in
   wire signed [9:0] m169_42;
   assign m169_42 =10'b0;

   // m169_43 = W*in
   wire signed [9:0] m169_43;
   assign m169_43 =10'b0;

   // m169_44 = W*in
   wire signed [9:0] m169_44;
   assign m169_44 =10'b0;

   // m169_45 = W*in
   wire signed [9:0] m169_45;
   assign m169_45 =10'b0;

   // m169_46 = W*in
   wire signed [9:0] m169_46;
   assign m169_46 =10'b0;

   // m169_47 = W*in
   wire signed [9:0] m169_47;
   assign m169_47 =10'b0;

   // m169_48 = W*in
   wire signed [9:0] m169_48;
   assign m169_48 =10'b0;

   // m169_49 = W*in
   wire signed [9:0] m169_49;
   assign m169_49 =10'b0;

   // m169_50 = W*in
   wire signed [9:0] m169_50;
   assign m169_50 =10'b0;

   // m169_51 = W*in
   wire signed [9:0] m169_51;
   assign m169_51 =10'b0;

   // m169_52 = W*in
   wire signed [9:0] m169_52;
   assign m169_52 =10'b0;

   // m169_53 = W*in
   wire signed [9:0] m169_53;
   assign m169_53 =10'b0;

   // m169_54 = W*in
   wire signed [9:0] m169_54;
   assign m169_54 =10'b0;

   // m169_55 = W*in
   wire signed [9:0] m169_55;
   assign m169_55 =10'b0;

   // m169_56 = W*in
   wire signed [9:0] m169_56;
   assign m169_56 =10'b0;

   // m169_57 = W*in
   wire signed [9:0] m169_57;
   assign m169_57 =10'b0;

   // m169_58 = W*in
   wire signed [9:0] m169_58;
   assign m169_58 =10'b0;

   // m169_59 = W*in
   wire signed [9:0] m169_59;
   assign m169_59 =10'b0;

   // m169_60 = W*in
   wire signed [9:0] m169_60;
   assign m169_60 =10'b0;

   // m169_61 = W*in
   wire signed [9:0] m169_61;
   assign m169_61 =10'b0;

   // m169_62 = W*in
   wire signed [9:0] m169_62;
   assign m169_62 =10'b0;

   // m169_63 = W*in
   wire signed [9:0] m169_63;
   assign m169_63 =10'b0;

   // m169_64 = W*in
   wire signed [9:0] m169_64;
   assign m169_64 =10'b0;

   // m169_65 = W*in
   wire signed [9:0] m169_65;
   assign m169_65 =10'b0;

   // m169_66 = W*in
   wire signed [9:0] m169_66;
   assign m169_66 =10'b0;

   // m169_67 = W*in
   wire signed [9:0] m169_67;
   assign m169_67 =10'b0;

   // m169_68 = W*in
   wire signed [9:0] m169_68;
   assign m169_68 =10'b0;

   // m169_69 = W*in
   wire signed [9:0] m169_69;
   assign m169_69 =10'b0;

   // m169_70 = W*in
   wire signed [9:0] m169_70;
   assign m169_70 =10'b0;

   // m169_71 = W*in
   wire signed [9:0] m169_71;
   assign m169_71 =10'b0;

   // m169_72 = W*in
   wire signed [9:0] m169_72;
   assign m169_72 =10'b0;

   // m169_73 = W*in
   wire signed [9:0] m169_73;
   assign m169_73 =10'b0;

   // m169_74 = W*in
   wire signed [9:0] m169_74;
   assign m169_74 =10'b0;

   // m169_75 = W*in
   wire signed [9:0] m169_75;
   assign m169_75 =10'b0;

   // m169_76 = W*in
   wire signed [9:0] m169_76;
   assign m169_76 =10'b0;

   // m169_77 = W*in
   wire signed [9:0] m169_77;
   assign m169_77 =10'b0;

   // m169_78 = W*in
   wire signed [9:0] m169_78;
   assign m169_78 =10'b0;

   // m169_79 = W*in
   wire signed [9:0] m169_79;
   assign m169_79 =10'b0;

   // m169_80 = W*in
   wire signed [9:0] m169_80;
   assign m169_80 =10'b0;

   // m169_81 = W*in
   wire signed [9:0] m169_81;
   assign m169_81 =10'b0;

   // m169_82 = W*in
   wire signed [9:0] m169_82;
   assign m169_82 =10'b0;

   // m169_83 = W*in
   wire signed [9:0] m169_83;
   assign m169_83 =10'b0;

   // m169_84 = W*in
   wire signed [9:0] m169_84;
   assign m169_84 =10'b0;

   // m169_85 = W*in
   wire signed [9:0] m169_85;
   assign m169_85 =10'b0;

   // m169_86 = W*in
   wire signed [9:0] m169_86;
   assign m169_86 =10'b0;

   // m169_87 = W*in
   wire signed [9:0] m169_87;
   assign m169_87 =10'b0;

   // m169_88 = W*in
   wire signed [9:0] m169_88;
   assign m169_88 =10'b0;

   // m169_89 = W*in
   wire signed [9:0] m169_89;
   assign m169_89 =10'b0;

   // m169_90 = W*in
   wire signed [9:0] m169_90;
   assign m169_90 =10'b0;

   // m169_91 = W*in
   wire signed [9:0] m169_91;
   assign m169_91 =10'b0;

   // m169_92 = W*in
   wire signed [9:0] m169_92;
   assign m169_92 =10'b0;

   // m169_93 = W*in
   wire signed [9:0] m169_93;
   assign m169_93 =10'b0;

   // m169_94 = W*in
   wire signed [9:0] m169_94;
   assign m169_94 =10'b0;

   // m169_95 = W*in
   wire signed [9:0] m169_95;
   assign m169_95 =10'b0;

   // m169_96 = W*in
   wire signed [9:0] m169_96;
   assign m169_96 =10'b0;

   // m169_97 = W*in
   wire signed [9:0] m169_97;
   assign m169_97 =10'b0;

   // m169_98 = W*in
   wire signed [9:0] m169_98;
   assign m169_98 =10'b0;

   // m169_99 = W*in
   wire signed [9:0] m169_99;
   assign m169_99 =10'b0;

   // m169_100 = W*in
   wire signed [9:0] m169_100;
   assign m169_100 =10'b0;

   // m169_101 = W*in
   wire signed [9:0] m169_101;
   assign m169_101 =10'b0;

   // m169_102 = W*in
   wire signed [9:0] m169_102;
   assign m169_102 =10'b0;

   // m169_103 = W*in
   wire signed [9:0] m169_103;
   assign m169_103 =10'b0;

   // m169_104 = W*in
   wire signed [9:0] m169_104;
   assign m169_104 =10'b0;

   // m169_105 = W*in
   wire signed [9:0] m169_105;
   assign m169_105 =10'b0;

   // m169_106 = W*in
   wire signed [9:0] m169_106;
   assign m169_106 =10'b0;

   // m169_107 = W*in
   wire signed [9:0] m169_107;
   assign m169_107 =10'b0;

   // m169_108 = W*in
   wire signed [9:0] m169_108;
   assign m169_108 =10'b0;

   // m169_109 = W*in
   wire signed [9:0] m169_109;
   assign m169_109 =10'b0;

   // m169_110 = W*in
   wire signed [9:0] m169_110;
   assign m169_110 =10'b0;

   // m169_111 = W*in
   wire signed [9:0] m169_111;
   assign m169_111 =10'b0;

   // m169_112 = W*in
   wire signed [9:0] m169_112;
   assign m169_112 =10'b0;

   // m169_113 = W*in
   wire signed [9:0] m169_113;
   assign m169_113 =10'b0;

   // m169_114 = W*in
   wire signed [9:0] m169_114;
   assign m169_114 =10'b0;

   // m169_115 = W*in
   wire signed [9:0] m169_115;
   assign m169_115 =10'b0;

   // m169_116 = W*in
   wire signed [9:0] m169_116;
   assign m169_116 =10'b0;

   // m169_117 = W*in
   wire signed [9:0] m169_117;
   assign m169_117 =10'b0;

   // m170_1 = W*in
   wire signed [9:0] m170_1;
   assign m170_1 =10'b0;

   // m170_2 = W*in
   wire signed [9:0] m170_2;
   assign m170_2 =10'b0;

   // m170_3 = W*in
   wire signed [9:0] m170_3;
   assign m170_3 =10'b0;

   // m170_4 = W*in
   wire signed [9:0] m170_4;
   assign m170_4 =10'b0;

   // m170_5 = W*in
   wire signed [9:0] m170_5;
   assign m170_5 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_6 = W*in
   wire signed [9:0] m170_6;
   assign m170_6 =10'b0;

   // m170_7 = W*in
   wire signed [9:0] m170_7;
   assign m170_7 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_8 = W*in
   wire signed [9:0] m170_8;
   assign m170_8 =10'b0;

   // m170_9 = W*in
   wire signed [9:0] m170_9;
   assign m170_9 =10'b0;

   // m170_10 = W*in
   wire signed [9:0] m170_10;
   assign m170_10 =10'b0;

   // m170_11 = W*in
   wire signed [9:0] m170_11;
   assign m170_11 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_12 = W*in
   wire signed [9:0] m170_12;
   assign m170_12 =10'b0;

   // m170_13 = W*in
   wire signed [9:0] m170_13;
   assign m170_13 ={ {4{in170[5]}} , in170[5:0] };

   // m170_14 = W*in
   wire signed [9:0] m170_14;
   assign m170_14 ={ {4{in170[5]}} , in170[5:0] };

   // m170_15 = W*in
   wire signed [9:0] m170_15;
   assign m170_15 ={ {4{in170[5]}} , in170[5:0] };

   // m170_16 = W*in
   wire signed [9:0] m170_16;
   assign m170_16 ={ {4{in170[5]}} , in170[5:0] };

   // m170_17 = W*in
   wire signed [9:0] m170_17;
   assign m170_17 =10'b0;

   // m170_18 = W*in
   wire signed [9:0] m170_18;
   assign m170_18 ={ {4{in170[5]}} , in170[5:0] };

   // m170_19 = W*in
   wire signed [9:0] m170_19;
   assign m170_19 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_20 = W*in
   wire signed [9:0] m170_20;
   assign m170_20 ={ {5{in170[5]}} , in170[5:1] };

   // m170_21 = W*in
   wire signed [9:0] m170_21;
   assign m170_21 =10'b0;

   // m170_22 = W*in
   wire signed [9:0] m170_22;
   assign m170_22 =10'b0;

   // m170_23 = W*in
   wire signed [9:0] m170_23;
   assign m170_23 =10'b0;

   // m170_24 = W*in
   wire signed [9:0] m170_24;
   assign m170_24 =10'b0;

   // m170_25 = W*in
   wire signed [9:0] m170_25;
   assign m170_25 =10'b0;

   // m170_26 = W*in
   wire signed [9:0] m170_26;
   assign m170_26 ={ {4{in170[5]}} , in170[5:0] };

   // m170_27 = W*in
   wire signed [9:0] m170_27;
   assign m170_27 =10'b0;

   // m170_28 = W*in
   wire signed [9:0] m170_28;
   assign m170_28 =10'b0;

   // m170_29 = W*in
   wire signed [9:0] m170_29;
   assign m170_29 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_30 = W*in
   wire signed [9:0] m170_30;
   assign m170_30 ={ {4{in170[5]}} , in170[5:0] };

   // m170_31 = W*in
   wire signed [9:0] m170_31;
   assign m170_31 =10'b0;

   // m170_32 = W*in
   wire signed [9:0] m170_32;
   assign m170_32 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_33 = W*in
   wire signed [9:0] m170_33;
   assign m170_33 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_34 = W*in
   wire signed [9:0] m170_34;
   assign m170_34 =10'b0;

   // m170_35 = W*in
   wire signed [9:0] m170_35;
   assign m170_35 =10'b0;

   // m170_36 = W*in
   wire signed [9:0] m170_36;
   assign m170_36 =10'b0;

   // m170_37 = W*in
   wire signed [9:0] m170_37;
   assign m170_37 =10'b0;

   // m170_38 = W*in
   wire signed [9:0] m170_38;
   assign m170_38 =10'b0;

   // m170_39 = W*in
   wire signed [9:0] m170_39;
   assign m170_39 =10'b0;

   // m170_40 = W*in
   wire signed [9:0] m170_40;
   assign m170_40 =10'b0;

   // m170_41 = W*in
   wire signed [9:0] m170_41;
   assign m170_41 ={ {4{in170[5]}} , in170[5:0] };

   // m170_42 = W*in
   wire signed [9:0] m170_42;
   assign m170_42 ={ {3{in170[5]}} , in170 , {1{1'b0}} };

   // m170_43 = W*in
   wire signed [9:0] m170_43;
   assign m170_43 =10'b0;

   // m170_44 = W*in
   wire signed [9:0] m170_44;
   assign m170_44 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_45 = W*in
   wire signed [9:0] m170_45;
   assign m170_45 =10'b0;

   // m170_46 = W*in
   wire signed [9:0] m170_46;
   assign m170_46 =10'b0;

   // m170_47 = W*in
   wire signed [9:0] m170_47;
   assign m170_47 =10'b0;

   // m170_48 = W*in
   wire signed [9:0] m170_48;
   assign m170_48 =10'b0;

   // m170_49 = W*in
   wire signed [9:0] m170_49;
   assign m170_49 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_50 = W*in
   wire signed [9:0] m170_50;
   assign m170_50 =10'b0;

   // m170_51 = W*in
   wire signed [9:0] m170_51;
   assign m170_51 =10'b0;

   // m170_52 = W*in
   wire signed [9:0] m170_52;
   assign m170_52 =10'b0;

   // m170_53 = W*in
   wire signed [9:0] m170_53;
   assign m170_53 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_54 = W*in
   wire signed [9:0] m170_54;
   assign m170_54 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_55 = W*in
   wire signed [9:0] m170_55;
   assign m170_55 ={ {4{in170[5]}} , in170[5:0] };

   // m170_56 = W*in
   wire signed [9:0] m170_56;
   assign m170_56 =10'b0;

   // m170_57 = W*in
   wire signed [9:0] m170_57;
   assign m170_57 =10'b0;

   // m170_58 = W*in
   wire signed [9:0] m170_58;
   assign m170_58 =10'b0;

   // m170_59 = W*in
   wire signed [9:0] m170_59;
   assign m170_59 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_60 = W*in
   wire signed [9:0] m170_60;
   assign m170_60 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_61 = W*in
   wire signed [9:0] m170_61;
   assign m170_61 =10'b0;

   // m170_62 = W*in
   wire signed [9:0] m170_62;
   assign m170_62 =10'b0;

   // m170_63 = W*in
   wire signed [9:0] m170_63;
   assign m170_63 =10'b0;

   // m170_64 = W*in
   wire signed [9:0] m170_64;
   assign m170_64 ={ {4{in170[5]}} , in170[5:0] };

   // m170_65 = W*in
   wire signed [9:0] m170_65;
   assign m170_65 ={ {5{in170[5]}} , in170[5:1] };

   // m170_66 = W*in
   wire signed [9:0] m170_66;
   assign m170_66 =10'b0;

   // m170_67 = W*in
   wire signed [9:0] m170_67;
   assign m170_67 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_68 = W*in
   wire signed [9:0] m170_68;
   assign m170_68 =10'b0;

   // m170_69 = W*in
   wire signed [9:0] m170_69;
   assign m170_69 =10'b0;

   // m170_70 = W*in
   wire signed [9:0] m170_70;
   assign m170_70 =10'b0;

   // m170_71 = W*in
   wire signed [9:0] m170_71;
   assign m170_71 =10'b0;

   // m170_72 = W*in
   wire signed [9:0] m170_72;
   assign m170_72 ={ {4{in170[5]}} , in170[5:0] };

   // m170_73 = W*in
   wire signed [9:0] m170_73;
   assign m170_73 =10'b0;

   // m170_74 = W*in
   wire signed [9:0] m170_74;
   assign m170_74 ={ {4{in170[5]}} , in170[5:0] };

   // m170_75 = W*in
   wire signed [9:0] m170_75;
   assign m170_75 ={ {4{in170[5]}} , in170[5:0] };

   // m170_76 = W*in
   wire signed [9:0] m170_76;
   assign m170_76 =10'b0;

   // m170_77 = W*in
   wire signed [9:0] m170_77;
   assign m170_77 =10'b0;

   // m170_78 = W*in
   wire signed [9:0] m170_78;
   assign m170_78 =10'b0;

   // m170_79 = W*in
   wire signed [9:0] m170_79;
   assign m170_79 =10'b0;

   // m170_80 = W*in
   wire signed [9:0] m170_80;
   assign m170_80 =10'b0;

   // m170_81 = W*in
   wire signed [9:0] m170_81;
   assign m170_81 ={ {4{in170[5]}} , in170[5:0] };

   // m170_82 = W*in
   wire signed [9:0] m170_82;
   assign m170_82 =10'b0;

   // m170_83 = W*in
   wire signed [9:0] m170_83;
   assign m170_83 ={ {5{neg170[5]}} , neg170[5:1] };

   // m170_84 = W*in
   wire signed [9:0] m170_84;
   assign m170_84 =10'b0;

   // m170_85 = W*in
   wire signed [9:0] m170_85;
   assign m170_85 =10'b0;

   // m170_86 = W*in
   wire signed [9:0] m170_86;
   assign m170_86 =10'b0;

   // m170_87 = W*in
   wire signed [9:0] m170_87;
   assign m170_87 =10'b0;

   // m170_88 = W*in
   wire signed [9:0] m170_88;
   assign m170_88 =10'b0;

   // m170_89 = W*in
   wire signed [9:0] m170_89;
   assign m170_89 ={ {4{in170[5]}} , in170[5:0] };

   // m170_90 = W*in
   wire signed [9:0] m170_90;
   assign m170_90 =10'b0;

   // m170_91 = W*in
   wire signed [9:0] m170_91;
   assign m170_91 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_92 = W*in
   wire signed [9:0] m170_92;
   assign m170_92 =10'b0;

   // m170_93 = W*in
   wire signed [9:0] m170_93;
   assign m170_93 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_94 = W*in
   wire signed [9:0] m170_94;
   assign m170_94 ={ {4{in170[5]}} , in170[5:0] };

   // m170_95 = W*in
   wire signed [9:0] m170_95;
   assign m170_95 ={ {3{neg170[5]}} , neg170 , {1{1'b0}} };

   // m170_96 = W*in
   wire signed [9:0] m170_96;
   assign m170_96 ={ {4{in170[5]}} , in170[5:0] };

   // m170_97 = W*in
   wire signed [9:0] m170_97;
   assign m170_97 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_98 = W*in
   wire signed [9:0] m170_98;
   assign m170_98 =10'b0;

   // m170_99 = W*in
   wire signed [9:0] m170_99;
   assign m170_99 =10'b0;

   // m170_100 = W*in
   wire signed [9:0] m170_100;
   assign m170_100 ={ {4{in170[5]}} , in170[5:0] };

   // m170_101 = W*in
   wire signed [9:0] m170_101;
   assign m170_101 =10'b0;

   // m170_102 = W*in
   wire signed [9:0] m170_102;
   assign m170_102 ={ {4{in170[5]}} , in170[5:0] };

   // m170_103 = W*in
   wire signed [9:0] m170_103;
   assign m170_103 =10'b0;

   // m170_104 = W*in
   wire signed [9:0] m170_104;
   assign m170_104 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_105 = W*in
   wire signed [9:0] m170_105;
   assign m170_105 =10'b0;

   // m170_106 = W*in
   wire signed [9:0] m170_106;
   assign m170_106 ={ {4{in170[5]}} , in170[5:0] };

   // m170_107 = W*in
   wire signed [9:0] m170_107;
   assign m170_107 =10'b0;

   // m170_108 = W*in
   wire signed [9:0] m170_108;
   assign m170_108 ={ {4{in170[5]}} , in170[5:0] };

   // m170_109 = W*in
   wire signed [9:0] m170_109;
   assign m170_109 ={ {4{in170[5]}} , in170[5:0] };

   // m170_110 = W*in
   wire signed [9:0] m170_110;
   assign m170_110 ={ {4{neg170[5]}} , neg170[5:0] };

   // m170_111 = W*in
   wire signed [9:0] m170_111;
   assign m170_111 =10'b0;

   // m170_112 = W*in
   wire signed [9:0] m170_112;
   assign m170_112 =10'b0;

   // m170_113 = W*in
   wire signed [9:0] m170_113;
   assign m170_113 =10'b0;

   // m170_114 = W*in
   wire signed [9:0] m170_114;
   assign m170_114 =10'b0;

   // m170_115 = W*in
   wire signed [9:0] m170_115;
   assign m170_115 =10'b0;

   // m170_116 = W*in
   wire signed [9:0] m170_116;
   assign m170_116 ={ {4{in170[5]}} , in170[5:0] };

   // m170_117 = W*in
   wire signed [9:0] m170_117;
   assign m170_117 ={ {4{neg170[5]}} , neg170[5:0] };

   // m171_1 = W*in
   wire signed [9:0] m171_1;
   assign m171_1 =10'b0;

   // m171_2 = W*in
   wire signed [9:0] m171_2;
   assign m171_2 =10'b0;

   // m171_3 = W*in
   wire signed [9:0] m171_3;
   assign m171_3 =10'b0;

   // m171_4 = W*in
   wire signed [9:0] m171_4;
   assign m171_4 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_5 = W*in
   wire signed [9:0] m171_5;
   assign m171_5 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_6 = W*in
   wire signed [9:0] m171_6;
   assign m171_6 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_7 = W*in
   wire signed [9:0] m171_7;
   assign m171_7 =10'b0;

   // m171_8 = W*in
   wire signed [9:0] m171_8;
   assign m171_8 =10'b0;

   // m171_9 = W*in
   wire signed [9:0] m171_9;
   assign m171_9 =10'b0;

   // m171_10 = W*in
   wire signed [9:0] m171_10;
   assign m171_10 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_11 = W*in
   wire signed [9:0] m171_11;
   assign m171_11 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_12 = W*in
   wire signed [9:0] m171_12;
   assign m171_12 =10'b0;

   // m171_13 = W*in
   wire signed [9:0] m171_13;
   assign m171_13 =10'b0;

   // m171_14 = W*in
   wire signed [9:0] m171_14;
   assign m171_14 =10'b0;

   // m171_15 = W*in
   wire signed [9:0] m171_15;
   assign m171_15 =10'b0;

   // m171_16 = W*in
   wire signed [9:0] m171_16;
   assign m171_16 =10'b0;

   // m171_17 = W*in
   wire signed [9:0] m171_17;
   assign m171_17 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_18 = W*in
   wire signed [9:0] m171_18;
   assign m171_18 ={ {3{in171[5]}} , in171 , {1{1'b0}} };

   // m171_19 = W*in
   wire signed [9:0] m171_19;
   assign m171_19 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_20 = W*in
   wire signed [9:0] m171_20;
   assign m171_20 ={ {5{in171[5]}} , in171[5:1] };

   // m171_21 = W*in
   wire signed [9:0] m171_21;
   assign m171_21 ={ {5{neg171[5]}} , neg171[5:1] };

   // m171_22 = W*in
   wire signed [9:0] m171_22;
   assign m171_22 =10'b0;

   // m171_23 = W*in
   wire signed [9:0] m171_23;
   assign m171_23 =10'b0;

   // m171_24 = W*in
   wire signed [9:0] m171_24;
   assign m171_24 =10'b0;

   // m171_25 = W*in
   wire signed [9:0] m171_25;
   assign m171_25 =10'b0;

   // m171_26 = W*in
   wire signed [9:0] m171_26;
   assign m171_26 ={ {4{in171[5]}} , in171[5:0] };

   // m171_27 = W*in
   wire signed [9:0] m171_27;
   assign m171_27 =10'b0;

   // m171_28 = W*in
   wire signed [9:0] m171_28;
   assign m171_28 ={ {5{neg171[5]}} , neg171[5:1] };

   // m171_29 = W*in
   wire signed [9:0] m171_29;
   assign m171_29 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_30 = W*in
   wire signed [9:0] m171_30;
   assign m171_30 ={ {4{in171[5]}} , in171[5:0] };

   // m171_31 = W*in
   wire signed [9:0] m171_31;
   assign m171_31 =10'b0;

   // m171_32 = W*in
   wire signed [9:0] m171_32;
   assign m171_32 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_33 = W*in
   wire signed [9:0] m171_33;
   assign m171_33 ={ {4{in171[5]}} , in171[5:0] };

   // m171_34 = W*in
   wire signed [9:0] m171_34;
   assign m171_34 =10'b0;

   // m171_35 = W*in
   wire signed [9:0] m171_35;
   assign m171_35 ={ {5{in171[5]}} , in171[5:1] };

   // m171_36 = W*in
   wire signed [9:0] m171_36;
   assign m171_36 =10'b0;

   // m171_37 = W*in
   wire signed [9:0] m171_37;
   assign m171_37 =10'b0;

   // m171_38 = W*in
   wire signed [9:0] m171_38;
   assign m171_38 ={ {5{neg171[5]}} , neg171[5:1] };

   // m171_39 = W*in
   wire signed [9:0] m171_39;
   assign m171_39 =10'b0;

   // m171_40 = W*in
   wire signed [9:0] m171_40;
   assign m171_40 =10'b0;

   // m171_41 = W*in
   wire signed [9:0] m171_41;
   assign m171_41 ={ {4{in171[5]}} , in171[5:0] };

   // m171_42 = W*in
   wire signed [9:0] m171_42;
   assign m171_42 ={ {4{in171[5]}} , in171[5:0] };

   // m171_43 = W*in
   wire signed [9:0] m171_43;
   assign m171_43 ={ {4{in171[5]}} , in171[5:0] };

   // m171_44 = W*in
   wire signed [9:0] m171_44;
   assign m171_44 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_45 = W*in
   wire signed [9:0] m171_45;
   assign m171_45 =10'b0;

   // m171_46 = W*in
   wire signed [9:0] m171_46;
   assign m171_46 =10'b0;

   // m171_47 = W*in
   wire signed [9:0] m171_47;
   assign m171_47 =10'b0;

   // m171_48 = W*in
   wire signed [9:0] m171_48;
   assign m171_48 ={ {4{in171[5]}} , in171[5:0] };

   // m171_49 = W*in
   wire signed [9:0] m171_49;
   assign m171_49 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_50 = W*in
   wire signed [9:0] m171_50;
   assign m171_50 =10'b0;

   // m171_51 = W*in
   wire signed [9:0] m171_51;
   assign m171_51 =10'b0;

   // m171_52 = W*in
   wire signed [9:0] m171_52;
   assign m171_52 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_53 = W*in
   wire signed [9:0] m171_53;
   assign m171_53 ={ {3{neg171[5]}} , neg171 , {1{1'b0}} };

   // m171_54 = W*in
   wire signed [9:0] m171_54;
   assign m171_54 ={ {3{neg171[5]}} , neg171 , {1{1'b0}} };

   // m171_55 = W*in
   wire signed [9:0] m171_55;
   assign m171_55 ={ {4{in171[5]}} , in171[5:0] };

   // m171_56 = W*in
   wire signed [9:0] m171_56;
   assign m171_56 =10'b0;

   // m171_57 = W*in
   wire signed [9:0] m171_57;
   assign m171_57 =10'b0;

   // m171_58 = W*in
   wire signed [9:0] m171_58;
   assign m171_58 =10'b0;

   // m171_59 = W*in
   wire signed [9:0] m171_59;
   assign m171_59 ={ {5{neg171[5]}} , neg171[5:1] };

   // m171_60 = W*in
   wire signed [9:0] m171_60;
   assign m171_60 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_61 = W*in
   wire signed [9:0] m171_61;
   assign m171_61 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_62 = W*in
   wire signed [9:0] m171_62;
   assign m171_62 =10'b0;

   // m171_63 = W*in
   wire signed [9:0] m171_63;
   assign m171_63 =10'b0;

   // m171_64 = W*in
   wire signed [9:0] m171_64;
   assign m171_64 ={ {4{in171[5]}} , in171[5:0] };

   // m171_65 = W*in
   wire signed [9:0] m171_65;
   assign m171_65 =10'b0;

   // m171_66 = W*in
   wire signed [9:0] m171_66;
   assign m171_66 =10'b0;

   // m171_67 = W*in
   wire signed [9:0] m171_67;
   assign m171_67 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_68 = W*in
   wire signed [9:0] m171_68;
   assign m171_68 ={ {4{in171[5]}} , in171[5:0] };

   // m171_69 = W*in
   wire signed [9:0] m171_69;
   assign m171_69 =10'b0;

   // m171_70 = W*in
   wire signed [9:0] m171_70;
   assign m171_70 =10'b0;

   // m171_71 = W*in
   wire signed [9:0] m171_71;
   assign m171_71 ={ {5{in171[5]}} , in171[5:1] };

   // m171_72 = W*in
   wire signed [9:0] m171_72;
   assign m171_72 =10'b0;

   // m171_73 = W*in
   wire signed [9:0] m171_73;
   assign m171_73 =10'b0;

   // m171_74 = W*in
   wire signed [9:0] m171_74;
   assign m171_74 ={ {5{in171[5]}} , in171[5:1] };

   // m171_75 = W*in
   wire signed [9:0] m171_75;
   assign m171_75 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_76 = W*in
   wire signed [9:0] m171_76;
   assign m171_76 =10'b0;

   // m171_77 = W*in
   wire signed [9:0] m171_77;
   assign m171_77 =10'b0;

   // m171_78 = W*in
   wire signed [9:0] m171_78;
   assign m171_78 ={ {4{in171[5]}} , in171[5:0] };

   // m171_79 = W*in
   wire signed [9:0] m171_79;
   assign m171_79 =10'b0;

   // m171_80 = W*in
   wire signed [9:0] m171_80;
   assign m171_80 =10'b0;

   // m171_81 = W*in
   wire signed [9:0] m171_81;
   assign m171_81 =10'b0;

   // m171_82 = W*in
   wire signed [9:0] m171_82;
   assign m171_82 =10'b0;

   // m171_83 = W*in
   wire signed [9:0] m171_83;
   assign m171_83 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_84 = W*in
   wire signed [9:0] m171_84;
   assign m171_84 =10'b0;

   // m171_85 = W*in
   wire signed [9:0] m171_85;
   assign m171_85 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_86 = W*in
   wire signed [9:0] m171_86;
   assign m171_86 =10'b0;

   // m171_87 = W*in
   wire signed [9:0] m171_87;
   assign m171_87 =10'b0;

   // m171_88 = W*in
   wire signed [9:0] m171_88;
   assign m171_88 =10'b0;

   // m171_89 = W*in
   wire signed [9:0] m171_89;
   assign m171_89 =10'b0;

   // m171_90 = W*in
   wire signed [9:0] m171_90;
   assign m171_90 =10'b0;

   // m171_91 = W*in
   wire signed [9:0] m171_91;
   assign m171_91 =10'b0;

   // m171_92 = W*in
   wire signed [9:0] m171_92;
   assign m171_92 =10'b0;

   // m171_93 = W*in
   wire signed [9:0] m171_93;
   assign m171_93 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_94 = W*in
   wire signed [9:0] m171_94;
   assign m171_94 ={ {5{in171[5]}} , in171[5:1] };

   // m171_95 = W*in
   wire signed [9:0] m171_95;
   assign m171_95 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_96 = W*in
   wire signed [9:0] m171_96;
   assign m171_96 ={ {4{in171[5]}} , in171[5:0] };

   // m171_97 = W*in
   wire signed [9:0] m171_97;
   assign m171_97 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_98 = W*in
   wire signed [9:0] m171_98;
   assign m171_98 =10'b0;

   // m171_99 = W*in
   wire signed [9:0] m171_99;
   assign m171_99 =10'b0;

   // m171_100 = W*in
   wire signed [9:0] m171_100;
   assign m171_100 =10'b0;

   // m171_101 = W*in
   wire signed [9:0] m171_101;
   assign m171_101 =10'b0;

   // m171_102 = W*in
   wire signed [9:0] m171_102;
   assign m171_102 =10'b0;

   // m171_103 = W*in
   wire signed [9:0] m171_103;
   assign m171_103 =10'b0;

   // m171_104 = W*in
   wire signed [9:0] m171_104;
   assign m171_104 =10'b0;

   // m171_105 = W*in
   wire signed [9:0] m171_105;
   assign m171_105 =10'b0;

   // m171_106 = W*in
   wire signed [9:0] m171_106;
   assign m171_106 ={ {4{in171[5]}} , in171[5:0] };

   // m171_107 = W*in
   wire signed [9:0] m171_107;
   assign m171_107 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_108 = W*in
   wire signed [9:0] m171_108;
   assign m171_108 ={ {5{in171[5]}} , in171[5:1] };

   // m171_109 = W*in
   wire signed [9:0] m171_109;
   assign m171_109 ={ {4{in171[5]}} , in171[5:0] };

   // m171_110 = W*in
   wire signed [9:0] m171_110;
   assign m171_110 ={ {4{neg171[5]}} , neg171[5:0] };

   // m171_111 = W*in
   wire signed [9:0] m171_111;
   assign m171_111 =10'b0;

   // m171_112 = W*in
   wire signed [9:0] m171_112;
   assign m171_112 ={ {5{neg171[5]}} , neg171[5:1] };

   // m171_113 = W*in
   wire signed [9:0] m171_113;
   assign m171_113 ={ {4{in171[5]}} , in171[5:0] };

   // m171_114 = W*in
   wire signed [9:0] m171_114;
   assign m171_114 =10'b0;

   // m171_115 = W*in
   wire signed [9:0] m171_115;
   assign m171_115 ={ {4{in171[5]}} , in171[5:0] };

   // m171_116 = W*in
   wire signed [9:0] m171_116;
   assign m171_116 ={ {3{in171[5]}} , in171 , {1{1'b0}} };

   // m171_117 = W*in
   wire signed [9:0] m171_117;
   assign m171_117 =10'b0;

   // m172_1 = W*in
   wire signed [9:0] m172_1;
   assign m172_1 =10'b0;

   // m172_2 = W*in
   wire signed [9:0] m172_2;
   assign m172_2 =10'b0;

   // m172_3 = W*in
   wire signed [9:0] m172_3;
   assign m172_3 =10'b0;

   // m172_4 = W*in
   wire signed [9:0] m172_4;
   assign m172_4 =10'b0;

   // m172_5 = W*in
   wire signed [9:0] m172_5;
   assign m172_5 =10'b0;

   // m172_6 = W*in
   wire signed [9:0] m172_6;
   assign m172_6 ={ {5{neg172[5]}} , neg172[5:1] };

   // m172_7 = W*in
   wire signed [9:0] m172_7;
   assign m172_7 =10'b0;

   // m172_8 = W*in
   wire signed [9:0] m172_8;
   assign m172_8 =10'b0;

   // m172_9 = W*in
   wire signed [9:0] m172_9;
   assign m172_9 =10'b0;

   // m172_10 = W*in
   wire signed [9:0] m172_10;
   assign m172_10 =10'b0;

   // m172_11 = W*in
   wire signed [9:0] m172_11;
   assign m172_11 =10'b0;

   // m172_12 = W*in
   wire signed [9:0] m172_12;
   assign m172_12 =10'b0;

   // m172_13 = W*in
   wire signed [9:0] m172_13;
   assign m172_13 =10'b0;

   // m172_14 = W*in
   wire signed [9:0] m172_14;
   assign m172_14 =10'b0;

   // m172_15 = W*in
   wire signed [9:0] m172_15;
   assign m172_15 =10'b0;

   // m172_16 = W*in
   wire signed [9:0] m172_16;
   assign m172_16 =10'b0;

   // m172_17 = W*in
   wire signed [9:0] m172_17;
   assign m172_17 ={ {5{in172[5]}} , in172[5:1] };

   // m172_18 = W*in
   wire signed [9:0] m172_18;
   assign m172_18 ={ {5{neg172[5]}} , neg172[5:1] };

   // m172_19 = W*in
   wire signed [9:0] m172_19;
   assign m172_19 =10'b0;

   // m172_20 = W*in
   wire signed [9:0] m172_20;
   assign m172_20 =10'b0;

   // m172_21 = W*in
   wire signed [9:0] m172_21;
   assign m172_21 =10'b0;

   // m172_22 = W*in
   wire signed [9:0] m172_22;
   assign m172_22 =10'b0;

   // m172_23 = W*in
   wire signed [9:0] m172_23;
   assign m172_23 =10'b0;

   // m172_24 = W*in
   wire signed [9:0] m172_24;
   assign m172_24 =10'b0;

   // m172_25 = W*in
   wire signed [9:0] m172_25;
   assign m172_25 ={ {4{in172[5]}} , in172[5:0] };

   // m172_26 = W*in
   wire signed [9:0] m172_26;
   assign m172_26 =10'b0;

   // m172_27 = W*in
   wire signed [9:0] m172_27;
   assign m172_27 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_28 = W*in
   wire signed [9:0] m172_28;
   assign m172_28 =10'b0;

   // m172_29 = W*in
   wire signed [9:0] m172_29;
   assign m172_29 =10'b0;

   // m172_30 = W*in
   wire signed [9:0] m172_30;
   assign m172_30 ={ {4{in172[5]}} , in172[5:0] };

   // m172_31 = W*in
   wire signed [9:0] m172_31;
   assign m172_31 ={ {5{neg172[5]}} , neg172[5:1] };

   // m172_32 = W*in
   wire signed [9:0] m172_32;
   assign m172_32 =10'b0;

   // m172_33 = W*in
   wire signed [9:0] m172_33;
   assign m172_33 ={ {5{in172[5]}} , in172[5:1] };

   // m172_34 = W*in
   wire signed [9:0] m172_34;
   assign m172_34 =10'b0;

   // m172_35 = W*in
   wire signed [9:0] m172_35;
   assign m172_35 =10'b0;

   // m172_36 = W*in
   wire signed [9:0] m172_36;
   assign m172_36 =10'b0;

   // m172_37 = W*in
   wire signed [9:0] m172_37;
   assign m172_37 =10'b0;

   // m172_38 = W*in
   wire signed [9:0] m172_38;
   assign m172_38 =10'b0;

   // m172_39 = W*in
   wire signed [9:0] m172_39;
   assign m172_39 =10'b0;

   // m172_40 = W*in
   wire signed [9:0] m172_40;
   assign m172_40 =10'b0;

   // m172_41 = W*in
   wire signed [9:0] m172_41;
   assign m172_41 =10'b0;

   // m172_42 = W*in
   wire signed [9:0] m172_42;
   assign m172_42 =10'b0;

   // m172_43 = W*in
   wire signed [9:0] m172_43;
   assign m172_43 =10'b0;

   // m172_44 = W*in
   wire signed [9:0] m172_44;
   assign m172_44 =10'b0;

   // m172_45 = W*in
   wire signed [9:0] m172_45;
   assign m172_45 =10'b0;

   // m172_46 = W*in
   wire signed [9:0] m172_46;
   assign m172_46 =10'b0;

   // m172_47 = W*in
   wire signed [9:0] m172_47;
   assign m172_47 =10'b0;

   // m172_48 = W*in
   wire signed [9:0] m172_48;
   assign m172_48 =10'b0;

   // m172_49 = W*in
   wire signed [9:0] m172_49;
   assign m172_49 =10'b0;

   // m172_50 = W*in
   wire signed [9:0] m172_50;
   assign m172_50 ={ {4{in172[5]}} , in172[5:0] };

   // m172_51 = W*in
   wire signed [9:0] m172_51;
   assign m172_51 =10'b0;

   // m172_52 = W*in
   wire signed [9:0] m172_52;
   assign m172_52 =10'b0;

   // m172_53 = W*in
   wire signed [9:0] m172_53;
   assign m172_53 =10'b0;

   // m172_54 = W*in
   wire signed [9:0] m172_54;
   assign m172_54 =10'b0;

   // m172_55 = W*in
   wire signed [9:0] m172_55;
   assign m172_55 =10'b0;

   // m172_56 = W*in
   wire signed [9:0] m172_56;
   assign m172_56 ={ {4{in172[5]}} , in172[5:0] };

   // m172_57 = W*in
   wire signed [9:0] m172_57;
   assign m172_57 =10'b0;

   // m172_58 = W*in
   wire signed [9:0] m172_58;
   assign m172_58 =10'b0;

   // m172_59 = W*in
   wire signed [9:0] m172_59;
   assign m172_59 =10'b0;

   // m172_60 = W*in
   wire signed [9:0] m172_60;
   assign m172_60 =10'b0;

   // m172_61 = W*in
   wire signed [9:0] m172_61;
   assign m172_61 ={ {5{neg172[5]}} , neg172[5:1] };

   // m172_62 = W*in
   wire signed [9:0] m172_62;
   assign m172_62 =10'b0;

   // m172_63 = W*in
   wire signed [9:0] m172_63;
   assign m172_63 =10'b0;

   // m172_64 = W*in
   wire signed [9:0] m172_64;
   assign m172_64 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_65 = W*in
   wire signed [9:0] m172_65;
   assign m172_65 =10'b0;

   // m172_66 = W*in
   wire signed [9:0] m172_66;
   assign m172_66 ={ {5{neg172[5]}} , neg172[5:1] };

   // m172_67 = W*in
   wire signed [9:0] m172_67;
   assign m172_67 =10'b0;

   // m172_68 = W*in
   wire signed [9:0] m172_68;
   assign m172_68 =10'b0;

   // m172_69 = W*in
   wire signed [9:0] m172_69;
   assign m172_69 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_70 = W*in
   wire signed [9:0] m172_70;
   assign m172_70 =10'b0;

   // m172_71 = W*in
   wire signed [9:0] m172_71;
   assign m172_71 =10'b0;

   // m172_72 = W*in
   wire signed [9:0] m172_72;
   assign m172_72 =10'b0;

   // m172_73 = W*in
   wire signed [9:0] m172_73;
   assign m172_73 ={ {5{in172[5]}} , in172[5:1] };

   // m172_74 = W*in
   wire signed [9:0] m172_74;
   assign m172_74 =10'b0;

   // m172_75 = W*in
   wire signed [9:0] m172_75;
   assign m172_75 ={ {4{in172[5]}} , in172[5:0] };

   // m172_76 = W*in
   wire signed [9:0] m172_76;
   assign m172_76 ={ {4{in172[5]}} , in172[5:0] };

   // m172_77 = W*in
   wire signed [9:0] m172_77;
   assign m172_77 =10'b0;

   // m172_78 = W*in
   wire signed [9:0] m172_78;
   assign m172_78 =10'b0;

   // m172_79 = W*in
   wire signed [9:0] m172_79;
   assign m172_79 =10'b0;

   // m172_80 = W*in
   wire signed [9:0] m172_80;
   assign m172_80 =10'b0;

   // m172_81 = W*in
   wire signed [9:0] m172_81;
   assign m172_81 ={ {5{neg172[5]}} , neg172[5:1] };

   // m172_82 = W*in
   wire signed [9:0] m172_82;
   assign m172_82 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_83 = W*in
   wire signed [9:0] m172_83;
   assign m172_83 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_84 = W*in
   wire signed [9:0] m172_84;
   assign m172_84 =10'b0;

   // m172_85 = W*in
   wire signed [9:0] m172_85;
   assign m172_85 =10'b0;

   // m172_86 = W*in
   wire signed [9:0] m172_86;
   assign m172_86 =10'b0;

   // m172_87 = W*in
   wire signed [9:0] m172_87;
   assign m172_87 =10'b0;

   // m172_88 = W*in
   wire signed [9:0] m172_88;
   assign m172_88 =10'b0;

   // m172_89 = W*in
   wire signed [9:0] m172_89;
   assign m172_89 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_90 = W*in
   wire signed [9:0] m172_90;
   assign m172_90 =10'b0;

   // m172_91 = W*in
   wire signed [9:0] m172_91;
   assign m172_91 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_92 = W*in
   wire signed [9:0] m172_92;
   assign m172_92 =10'b0;

   // m172_93 = W*in
   wire signed [9:0] m172_93;
   assign m172_93 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_94 = W*in
   wire signed [9:0] m172_94;
   assign m172_94 =10'b0;

   // m172_95 = W*in
   wire signed [9:0] m172_95;
   assign m172_95 =10'b0;

   // m172_96 = W*in
   wire signed [9:0] m172_96;
   assign m172_96 =10'b0;

   // m172_97 = W*in
   wire signed [9:0] m172_97;
   assign m172_97 ={ {4{neg172[5]}} , neg172[5:0] };

   // m172_98 = W*in
   wire signed [9:0] m172_98;
   assign m172_98 =10'b0;

   // m172_99 = W*in
   wire signed [9:0] m172_99;
   assign m172_99 =10'b0;

   // m172_100 = W*in
   wire signed [9:0] m172_100;
   assign m172_100 ={ {4{in172[5]}} , in172[5:0] };

   // m172_101 = W*in
   wire signed [9:0] m172_101;
   assign m172_101 =10'b0;

   // m172_102 = W*in
   wire signed [9:0] m172_102;
   assign m172_102 ={ {4{in172[5]}} , in172[5:0] };

   // m172_103 = W*in
   wire signed [9:0] m172_103;
   assign m172_103 =10'b0;

   // m172_104 = W*in
   wire signed [9:0] m172_104;
   assign m172_104 =10'b0;

   // m172_105 = W*in
   wire signed [9:0] m172_105;
   assign m172_105 =10'b0;

   // m172_106 = W*in
   wire signed [9:0] m172_106;
   assign m172_106 ={ {4{in172[5]}} , in172[5:0] };

   // m172_107 = W*in
   wire signed [9:0] m172_107;
   assign m172_107 =10'b0;

   // m172_108 = W*in
   wire signed [9:0] m172_108;
   assign m172_108 =10'b0;

   // m172_109 = W*in
   wire signed [9:0] m172_109;
   assign m172_109 =10'b0;

   // m172_110 = W*in
   wire signed [9:0] m172_110;
   assign m172_110 =10'b0;

   // m172_111 = W*in
   wire signed [9:0] m172_111;
   assign m172_111 =10'b0;

   // m172_112 = W*in
   wire signed [9:0] m172_112;
   assign m172_112 =10'b0;

   // m172_113 = W*in
   wire signed [9:0] m172_113;
   assign m172_113 =10'b0;

   // m172_114 = W*in
   wire signed [9:0] m172_114;
   assign m172_114 =10'b0;

   // m172_115 = W*in
   wire signed [9:0] m172_115;
   assign m172_115 =10'b0;

   // m172_116 = W*in
   wire signed [9:0] m172_116;
   assign m172_116 ={ {4{in172[5]}} , in172[5:0] };

   // m172_117 = W*in
   wire signed [9:0] m172_117;
   assign m172_117 ={ {4{neg172[5]}} , neg172[5:0] };

   // m173_1 = W*in
   wire signed [9:0] m173_1;
   assign m173_1 ={ {4{in173[5]}} , in173[5:0] };

   // m173_2 = W*in
   wire signed [9:0] m173_2;
   assign m173_2 =10'b0;

   // m173_3 = W*in
   wire signed [9:0] m173_3;
   assign m173_3 =10'b0;

   // m173_4 = W*in
   wire signed [9:0] m173_4;
   assign m173_4 =10'b0;

   // m173_5 = W*in
   wire signed [9:0] m173_5;
   assign m173_5 ={ {4{in173[5]}} , in173[5:0] };

   // m173_6 = W*in
   wire signed [9:0] m173_6;
   assign m173_6 =10'b0;

   // m173_7 = W*in
   wire signed [9:0] m173_7;
   assign m173_7 ={ {4{in173[5]}} , in173[5:0] };

   // m173_8 = W*in
   wire signed [9:0] m173_8;
   assign m173_8 =10'b0;

   // m173_9 = W*in
   wire signed [9:0] m173_9;
   assign m173_9 =10'b0;

   // m173_10 = W*in
   wire signed [9:0] m173_10;
   assign m173_10 =10'b0;

   // m173_11 = W*in
   wire signed [9:0] m173_11;
   assign m173_11 =10'b0;

   // m173_12 = W*in
   wire signed [9:0] m173_12;
   assign m173_12 =10'b0;

   // m173_13 = W*in
   wire signed [9:0] m173_13;
   assign m173_13 =10'b0;

   // m173_14 = W*in
   wire signed [9:0] m173_14;
   assign m173_14 =10'b0;

   // m173_15 = W*in
   wire signed [9:0] m173_15;
   assign m173_15 =10'b0;

   // m173_16 = W*in
   wire signed [9:0] m173_16;
   assign m173_16 =10'b0;

   // m173_17 = W*in
   wire signed [9:0] m173_17;
   assign m173_17 =10'b0;

   // m173_18 = W*in
   wire signed [9:0] m173_18;
   assign m173_18 =10'b0;

   // m173_19 = W*in
   wire signed [9:0] m173_19;
   assign m173_19 =10'b0;

   // m173_20 = W*in
   wire signed [9:0] m173_20;
   assign m173_20 ={ {5{neg173[5]}} , neg173[5:1] };

   // m173_21 = W*in
   wire signed [9:0] m173_21;
   assign m173_21 ={ {5{neg173[5]}} , neg173[5:1] };

   // m173_22 = W*in
   wire signed [9:0] m173_22;
   assign m173_22 ={ {4{in173[5]}} , in173[5:0] };

   // m173_23 = W*in
   wire signed [9:0] m173_23;
   assign m173_23 =10'b0;

   // m173_24 = W*in
   wire signed [9:0] m173_24;
   assign m173_24 =10'b0;

   // m173_25 = W*in
   wire signed [9:0] m173_25;
   assign m173_25 =10'b0;

   // m173_26 = W*in
   wire signed [9:0] m173_26;
   assign m173_26 =10'b0;

   // m173_27 = W*in
   wire signed [9:0] m173_27;
   assign m173_27 =10'b0;

   // m173_28 = W*in
   wire signed [9:0] m173_28;
   assign m173_28 ={ {4{in173[5]}} , in173[5:0] };

   // m173_29 = W*in
   wire signed [9:0] m173_29;
   assign m173_29 =10'b0;

   // m173_30 = W*in
   wire signed [9:0] m173_30;
   assign m173_30 =10'b0;

   // m173_31 = W*in
   wire signed [9:0] m173_31;
   assign m173_31 =10'b0;

   // m173_32 = W*in
   wire signed [9:0] m173_32;
   assign m173_32 =10'b0;

   // m173_33 = W*in
   wire signed [9:0] m173_33;
   assign m173_33 ={ {4{in173[5]}} , in173[5:0] };

   // m173_34 = W*in
   wire signed [9:0] m173_34;
   assign m173_34 =10'b0;

   // m173_35 = W*in
   wire signed [9:0] m173_35;
   assign m173_35 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_36 = W*in
   wire signed [9:0] m173_36;
   assign m173_36 =10'b0;

   // m173_37 = W*in
   wire signed [9:0] m173_37;
   assign m173_37 =10'b0;

   // m173_38 = W*in
   wire signed [9:0] m173_38;
   assign m173_38 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_39 = W*in
   wire signed [9:0] m173_39;
   assign m173_39 =10'b0;

   // m173_40 = W*in
   wire signed [9:0] m173_40;
   assign m173_40 =10'b0;

   // m173_41 = W*in
   wire signed [9:0] m173_41;
   assign m173_41 =10'b0;

   // m173_42 = W*in
   wire signed [9:0] m173_42;
   assign m173_42 =10'b0;

   // m173_43 = W*in
   wire signed [9:0] m173_43;
   assign m173_43 =10'b0;

   // m173_44 = W*in
   wire signed [9:0] m173_44;
   assign m173_44 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_45 = W*in
   wire signed [9:0] m173_45;
   assign m173_45 ={ {4{in173[5]}} , in173[5:0] };

   // m173_46 = W*in
   wire signed [9:0] m173_46;
   assign m173_46 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_47 = W*in
   wire signed [9:0] m173_47;
   assign m173_47 =10'b0;

   // m173_48 = W*in
   wire signed [9:0] m173_48;
   assign m173_48 =10'b0;

   // m173_49 = W*in
   wire signed [9:0] m173_49;
   assign m173_49 =10'b0;

   // m173_50 = W*in
   wire signed [9:0] m173_50;
   assign m173_50 =10'b0;

   // m173_51 = W*in
   wire signed [9:0] m173_51;
   assign m173_51 ={ {4{in173[5]}} , in173[5:0] };

   // m173_52 = W*in
   wire signed [9:0] m173_52;
   assign m173_52 =10'b0;

   // m173_53 = W*in
   wire signed [9:0] m173_53;
   assign m173_53 =10'b0;

   // m173_54 = W*in
   wire signed [9:0] m173_54;
   assign m173_54 =10'b0;

   // m173_55 = W*in
   wire signed [9:0] m173_55;
   assign m173_55 =10'b0;

   // m173_56 = W*in
   wire signed [9:0] m173_56;
   assign m173_56 =10'b0;

   // m173_57 = W*in
   wire signed [9:0] m173_57;
   assign m173_57 =10'b0;

   // m173_58 = W*in
   wire signed [9:0] m173_58;
   assign m173_58 =10'b0;

   // m173_59 = W*in
   wire signed [9:0] m173_59;
   assign m173_59 =10'b0;

   // m173_60 = W*in
   wire signed [9:0] m173_60;
   assign m173_60 =10'b0;

   // m173_61 = W*in
   wire signed [9:0] m173_61;
   assign m173_61 =10'b0;

   // m173_62 = W*in
   wire signed [9:0] m173_62;
   assign m173_62 =10'b0;

   // m173_63 = W*in
   wire signed [9:0] m173_63;
   assign m173_63 =10'b0;

   // m173_64 = W*in
   wire signed [9:0] m173_64;
   assign m173_64 =10'b0;

   // m173_65 = W*in
   wire signed [9:0] m173_65;
   assign m173_65 =10'b0;

   // m173_66 = W*in
   wire signed [9:0] m173_66;
   assign m173_66 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_67 = W*in
   wire signed [9:0] m173_67;
   assign m173_67 =10'b0;

   // m173_68 = W*in
   wire signed [9:0] m173_68;
   assign m173_68 =10'b0;

   // m173_69 = W*in
   wire signed [9:0] m173_69;
   assign m173_69 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_70 = W*in
   wire signed [9:0] m173_70;
   assign m173_70 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_71 = W*in
   wire signed [9:0] m173_71;
   assign m173_71 ={ {5{neg173[5]}} , neg173[5:1] };

   // m173_72 = W*in
   wire signed [9:0] m173_72;
   assign m173_72 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_73 = W*in
   wire signed [9:0] m173_73;
   assign m173_73 ={ {4{in173[5]}} , in173[5:0] };

   // m173_74 = W*in
   wire signed [9:0] m173_74;
   assign m173_74 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_75 = W*in
   wire signed [9:0] m173_75;
   assign m173_75 =10'b0;

   // m173_76 = W*in
   wire signed [9:0] m173_76;
   assign m173_76 =10'b0;

   // m173_77 = W*in
   wire signed [9:0] m173_77;
   assign m173_77 =10'b0;

   // m173_78 = W*in
   wire signed [9:0] m173_78;
   assign m173_78 ={ {4{in173[5]}} , in173[5:0] };

   // m173_79 = W*in
   wire signed [9:0] m173_79;
   assign m173_79 =10'b0;

   // m173_80 = W*in
   wire signed [9:0] m173_80;
   assign m173_80 =10'b0;

   // m173_81 = W*in
   wire signed [9:0] m173_81;
   assign m173_81 =10'b0;

   // m173_82 = W*in
   wire signed [9:0] m173_82;
   assign m173_82 ={ {5{neg173[5]}} , neg173[5:1] };

   // m173_83 = W*in
   wire signed [9:0] m173_83;
   assign m173_83 ={ {5{in173[5]}} , in173[5:1] };

   // m173_84 = W*in
   wire signed [9:0] m173_84;
   assign m173_84 =10'b0;

   // m173_85 = W*in
   wire signed [9:0] m173_85;
   assign m173_85 =10'b0;

   // m173_86 = W*in
   wire signed [9:0] m173_86;
   assign m173_86 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_87 = W*in
   wire signed [9:0] m173_87;
   assign m173_87 =10'b0;

   // m173_88 = W*in
   wire signed [9:0] m173_88;
   assign m173_88 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_89 = W*in
   wire signed [9:0] m173_89;
   assign m173_89 =10'b0;

   // m173_90 = W*in
   wire signed [9:0] m173_90;
   assign m173_90 ={ {4{in173[5]}} , in173[5:0] };

   // m173_91 = W*in
   wire signed [9:0] m173_91;
   assign m173_91 =10'b0;

   // m173_92 = W*in
   wire signed [9:0] m173_92;
   assign m173_92 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_93 = W*in
   wire signed [9:0] m173_93;
   assign m173_93 =10'b0;

   // m173_94 = W*in
   wire signed [9:0] m173_94;
   assign m173_94 =10'b0;

   // m173_95 = W*in
   wire signed [9:0] m173_95;
   assign m173_95 =10'b0;

   // m173_96 = W*in
   wire signed [9:0] m173_96;
   assign m173_96 =10'b0;

   // m173_97 = W*in
   wire signed [9:0] m173_97;
   assign m173_97 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_98 = W*in
   wire signed [9:0] m173_98;
   assign m173_98 =10'b0;

   // m173_99 = W*in
   wire signed [9:0] m173_99;
   assign m173_99 =10'b0;

   // m173_100 = W*in
   wire signed [9:0] m173_100;
   assign m173_100 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_101 = W*in
   wire signed [9:0] m173_101;
   assign m173_101 =10'b0;

   // m173_102 = W*in
   wire signed [9:0] m173_102;
   assign m173_102 =10'b0;

   // m173_103 = W*in
   wire signed [9:0] m173_103;
   assign m173_103 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_104 = W*in
   wire signed [9:0] m173_104;
   assign m173_104 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_105 = W*in
   wire signed [9:0] m173_105;
   assign m173_105 =10'b0;

   // m173_106 = W*in
   wire signed [9:0] m173_106;
   assign m173_106 =10'b0;

   // m173_107 = W*in
   wire signed [9:0] m173_107;
   assign m173_107 =10'b0;

   // m173_108 = W*in
   wire signed [9:0] m173_108;
   assign m173_108 ={ {5{neg173[5]}} , neg173[5:1] };

   // m173_109 = W*in
   wire signed [9:0] m173_109;
   assign m173_109 ={ {5{neg173[5]}} , neg173[5:1] };

   // m173_110 = W*in
   wire signed [9:0] m173_110;
   assign m173_110 ={ {4{neg173[5]}} , neg173[5:0] };

   // m173_111 = W*in
   wire signed [9:0] m173_111;
   assign m173_111 =10'b0;

   // m173_112 = W*in
   wire signed [9:0] m173_112;
   assign m173_112 =10'b0;

   // m173_113 = W*in
   wire signed [9:0] m173_113;
   assign m173_113 =10'b0;

   // m173_114 = W*in
   wire signed [9:0] m173_114;
   assign m173_114 =10'b0;

   // m173_115 = W*in
   wire signed [9:0] m173_115;
   assign m173_115 =10'b0;

   // m173_116 = W*in
   wire signed [9:0] m173_116;
   assign m173_116 =10'b0;

   // m173_117 = W*in
   wire signed [9:0] m173_117;
   assign m173_117 ={ {4{neg173[5]}} , neg173[5:0] };

   // m174_1 = W*in
   wire signed [9:0] m174_1;
   assign m174_1 =10'b0;

   // m174_2 = W*in
   wire signed [9:0] m174_2;
   assign m174_2 =10'b0;

   // m174_3 = W*in
   wire signed [9:0] m174_3;
   assign m174_3 =10'b0;

   // m174_4 = W*in
   wire signed [9:0] m174_4;
   assign m174_4 =10'b0;

   // m174_5 = W*in
   wire signed [9:0] m174_5;
   assign m174_5 =10'b0;

   // m174_6 = W*in
   wire signed [9:0] m174_6;
   assign m174_6 =10'b0;

   // m174_7 = W*in
   wire signed [9:0] m174_7;
   assign m174_7 ={ {4{in174[5]}} , in174[5:0] };

   // m174_8 = W*in
   wire signed [9:0] m174_8;
   assign m174_8 =10'b0;

   // m174_9 = W*in
   wire signed [9:0] m174_9;
   assign m174_9 =10'b0;

   // m174_10 = W*in
   wire signed [9:0] m174_10;
   assign m174_10 =10'b0;

   // m174_11 = W*in
   wire signed [9:0] m174_11;
   assign m174_11 =10'b0;

   // m174_12 = W*in
   wire signed [9:0] m174_12;
   assign m174_12 =10'b0;

   // m174_13 = W*in
   wire signed [9:0] m174_13;
   assign m174_13 =10'b0;

   // m174_14 = W*in
   wire signed [9:0] m174_14;
   assign m174_14 =10'b0;

   // m174_15 = W*in
   wire signed [9:0] m174_15;
   assign m174_15 =10'b0;

   // m174_16 = W*in
   wire signed [9:0] m174_16;
   assign m174_16 =10'b0;

   // m174_17 = W*in
   wire signed [9:0] m174_17;
   assign m174_17 =10'b0;

   // m174_18 = W*in
   wire signed [9:0] m174_18;
   assign m174_18 =10'b0;

   // m174_19 = W*in
   wire signed [9:0] m174_19;
   assign m174_19 =10'b0;

   // m174_20 = W*in
   wire signed [9:0] m174_20;
   assign m174_20 =10'b0;

   // m174_21 = W*in
   wire signed [9:0] m174_21;
   assign m174_21 ={ {5{neg174[5]}} , neg174[5:1] };

   // m174_22 = W*in
   wire signed [9:0] m174_22;
   assign m174_22 =10'b0;

   // m174_23 = W*in
   wire signed [9:0] m174_23;
   assign m174_23 =10'b0;

   // m174_24 = W*in
   wire signed [9:0] m174_24;
   assign m174_24 =10'b0;

   // m174_25 = W*in
   wire signed [9:0] m174_25;
   assign m174_25 =10'b0;

   // m174_26 = W*in
   wire signed [9:0] m174_26;
   assign m174_26 =10'b0;

   // m174_27 = W*in
   wire signed [9:0] m174_27;
   assign m174_27 ={ {5{in174[5]}} , in174[5:1] };

   // m174_28 = W*in
   wire signed [9:0] m174_28;
   assign m174_28 =10'b0;

   // m174_29 = W*in
   wire signed [9:0] m174_29;
   assign m174_29 =10'b0;

   // m174_30 = W*in
   wire signed [9:0] m174_30;
   assign m174_30 =10'b0;

   // m174_31 = W*in
   wire signed [9:0] m174_31;
   assign m174_31 =10'b0;

   // m174_32 = W*in
   wire signed [9:0] m174_32;
   assign m174_32 =10'b0;

   // m174_33 = W*in
   wire signed [9:0] m174_33;
   assign m174_33 =10'b0;

   // m174_34 = W*in
   wire signed [9:0] m174_34;
   assign m174_34 =10'b0;

   // m174_35 = W*in
   wire signed [9:0] m174_35;
   assign m174_35 =10'b0;

   // m174_36 = W*in
   wire signed [9:0] m174_36;
   assign m174_36 ={ {5{in174[5]}} , in174[5:1] };

   // m174_37 = W*in
   wire signed [9:0] m174_37;
   assign m174_37 =10'b0;

   // m174_38 = W*in
   wire signed [9:0] m174_38;
   assign m174_38 =10'b0;

   // m174_39 = W*in
   wire signed [9:0] m174_39;
   assign m174_39 =10'b0;

   // m174_40 = W*in
   wire signed [9:0] m174_40;
   assign m174_40 =10'b0;

   // m174_41 = W*in
   wire signed [9:0] m174_41;
   assign m174_41 =10'b0;

   // m174_42 = W*in
   wire signed [9:0] m174_42;
   assign m174_42 =10'b0;

   // m174_43 = W*in
   wire signed [9:0] m174_43;
   assign m174_43 =10'b0;

   // m174_44 = W*in
   wire signed [9:0] m174_44;
   assign m174_44 =10'b0;

   // m174_45 = W*in
   wire signed [9:0] m174_45;
   assign m174_45 =10'b0;

   // m174_46 = W*in
   wire signed [9:0] m174_46;
   assign m174_46 =10'b0;

   // m174_47 = W*in
   wire signed [9:0] m174_47;
   assign m174_47 =10'b0;

   // m174_48 = W*in
   wire signed [9:0] m174_48;
   assign m174_48 =10'b0;

   // m174_49 = W*in
   wire signed [9:0] m174_49;
   assign m174_49 =10'b0;

   // m174_50 = W*in
   wire signed [9:0] m174_50;
   assign m174_50 =10'b0;

   // m174_51 = W*in
   wire signed [9:0] m174_51;
   assign m174_51 =10'b0;

   // m174_52 = W*in
   wire signed [9:0] m174_52;
   assign m174_52 =10'b0;

   // m174_53 = W*in
   wire signed [9:0] m174_53;
   assign m174_53 =10'b0;

   // m174_54 = W*in
   wire signed [9:0] m174_54;
   assign m174_54 =10'b0;

   // m174_55 = W*in
   wire signed [9:0] m174_55;
   assign m174_55 =10'b0;

   // m174_56 = W*in
   wire signed [9:0] m174_56;
   assign m174_56 =10'b0;

   // m174_57 = W*in
   wire signed [9:0] m174_57;
   assign m174_57 =10'b0;

   // m174_58 = W*in
   wire signed [9:0] m174_58;
   assign m174_58 =10'b0;

   // m174_59 = W*in
   wire signed [9:0] m174_59;
   assign m174_59 =10'b0;

   // m174_60 = W*in
   wire signed [9:0] m174_60;
   assign m174_60 =10'b0;

   // m174_61 = W*in
   wire signed [9:0] m174_61;
   assign m174_61 =10'b0;

   // m174_62 = W*in
   wire signed [9:0] m174_62;
   assign m174_62 =10'b0;

   // m174_63 = W*in
   wire signed [9:0] m174_63;
   assign m174_63 =10'b0;

   // m174_64 = W*in
   wire signed [9:0] m174_64;
   assign m174_64 =10'b0;

   // m174_65 = W*in
   wire signed [9:0] m174_65;
   assign m174_65 =10'b0;

   // m174_66 = W*in
   wire signed [9:0] m174_66;
   assign m174_66 =10'b0;

   // m174_67 = W*in
   wire signed [9:0] m174_67;
   assign m174_67 =10'b0;

   // m174_68 = W*in
   wire signed [9:0] m174_68;
   assign m174_68 =10'b0;

   // m174_69 = W*in
   wire signed [9:0] m174_69;
   assign m174_69 =10'b0;

   // m174_70 = W*in
   wire signed [9:0] m174_70;
   assign m174_70 ={ {5{neg174[5]}} , neg174[5:1] };

   // m174_71 = W*in
   wire signed [9:0] m174_71;
   assign m174_71 =10'b0;

   // m174_72 = W*in
   wire signed [9:0] m174_72;
   assign m174_72 ={ {5{neg174[5]}} , neg174[5:1] };

   // m174_73 = W*in
   wire signed [9:0] m174_73;
   assign m174_73 ={ {5{in174[5]}} , in174[5:1] };

   // m174_74 = W*in
   wire signed [9:0] m174_74;
   assign m174_74 ={ {5{neg174[5]}} , neg174[5:1] };

   // m174_75 = W*in
   wire signed [9:0] m174_75;
   assign m174_75 =10'b0;

   // m174_76 = W*in
   wire signed [9:0] m174_76;
   assign m174_76 =10'b0;

   // m174_77 = W*in
   wire signed [9:0] m174_77;
   assign m174_77 =10'b0;

   // m174_78 = W*in
   wire signed [9:0] m174_78;
   assign m174_78 =10'b0;

   // m174_79 = W*in
   wire signed [9:0] m174_79;
   assign m174_79 =10'b0;

   // m174_80 = W*in
   wire signed [9:0] m174_80;
   assign m174_80 =10'b0;

   // m174_81 = W*in
   wire signed [9:0] m174_81;
   assign m174_81 =10'b0;

   // m174_82 = W*in
   wire signed [9:0] m174_82;
   assign m174_82 =10'b0;

   // m174_83 = W*in
   wire signed [9:0] m174_83;
   assign m174_83 =10'b0;

   // m174_84 = W*in
   wire signed [9:0] m174_84;
   assign m174_84 =10'b0;

   // m174_85 = W*in
   wire signed [9:0] m174_85;
   assign m174_85 =10'b0;

   // m174_86 = W*in
   wire signed [9:0] m174_86;
   assign m174_86 =10'b0;

   // m174_87 = W*in
   wire signed [9:0] m174_87;
   assign m174_87 =10'b0;

   // m174_88 = W*in
   wire signed [9:0] m174_88;
   assign m174_88 =10'b0;

   // m174_89 = W*in
   wire signed [9:0] m174_89;
   assign m174_89 =10'b0;

   // m174_90 = W*in
   wire signed [9:0] m174_90;
   assign m174_90 =10'b0;

   // m174_91 = W*in
   wire signed [9:0] m174_91;
   assign m174_91 =10'b0;

   // m174_92 = W*in
   wire signed [9:0] m174_92;
   assign m174_92 =10'b0;

   // m174_93 = W*in
   wire signed [9:0] m174_93;
   assign m174_93 =10'b0;

   // m174_94 = W*in
   wire signed [9:0] m174_94;
   assign m174_94 =10'b0;

   // m174_95 = W*in
   wire signed [9:0] m174_95;
   assign m174_95 =10'b0;

   // m174_96 = W*in
   wire signed [9:0] m174_96;
   assign m174_96 =10'b0;

   // m174_97 = W*in
   wire signed [9:0] m174_97;
   assign m174_97 =10'b0;

   // m174_98 = W*in
   wire signed [9:0] m174_98;
   assign m174_98 =10'b0;

   // m174_99 = W*in
   wire signed [9:0] m174_99;
   assign m174_99 =10'b0;

   // m174_100 = W*in
   wire signed [9:0] m174_100;
   assign m174_100 =10'b0;

   // m174_101 = W*in
   wire signed [9:0] m174_101;
   assign m174_101 =10'b0;

   // m174_102 = W*in
   wire signed [9:0] m174_102;
   assign m174_102 =10'b0;

   // m174_103 = W*in
   wire signed [9:0] m174_103;
   assign m174_103 =10'b0;

   // m174_104 = W*in
   wire signed [9:0] m174_104;
   assign m174_104 =10'b0;

   // m174_105 = W*in
   wire signed [9:0] m174_105;
   assign m174_105 =10'b0;

   // m174_106 = W*in
   wire signed [9:0] m174_106;
   assign m174_106 =10'b0;

   // m174_107 = W*in
   wire signed [9:0] m174_107;
   assign m174_107 =10'b0;

   // m174_108 = W*in
   wire signed [9:0] m174_108;
   assign m174_108 =10'b0;

   // m174_109 = W*in
   wire signed [9:0] m174_109;
   assign m174_109 =10'b0;

   // m174_110 = W*in
   wire signed [9:0] m174_110;
   assign m174_110 =10'b0;

   // m174_111 = W*in
   wire signed [9:0] m174_111;
   assign m174_111 =10'b0;

   // m174_112 = W*in
   wire signed [9:0] m174_112;
   assign m174_112 =10'b0;

   // m174_113 = W*in
   wire signed [9:0] m174_113;
   assign m174_113 =10'b0;

   // m174_114 = W*in
   wire signed [9:0] m174_114;
   assign m174_114 =10'b0;

   // m174_115 = W*in
   wire signed [9:0] m174_115;
   assign m174_115 =10'b0;

   // m174_116 = W*in
   wire signed [9:0] m174_116;
   assign m174_116 =10'b0;

   // m174_117 = W*in
   wire signed [9:0] m174_117;
   assign m174_117 =10'b0;

   // m175_1 = W*in
   wire signed [9:0] m175_1;
   assign m175_1 =10'b0;

   // m175_2 = W*in
   wire signed [9:0] m175_2;
   assign m175_2 =10'b0;

   // m175_3 = W*in
   wire signed [9:0] m175_3;
   assign m175_3 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_4 = W*in
   wire signed [9:0] m175_4;
   assign m175_4 =10'b0;

   // m175_5 = W*in
   wire signed [9:0] m175_5;
   assign m175_5 =10'b0;

   // m175_6 = W*in
   wire signed [9:0] m175_6;
   assign m175_6 ={ {4{in175[5]}} , in175[5:0] };

   // m175_7 = W*in
   wire signed [9:0] m175_7;
   assign m175_7 =10'b0;

   // m175_8 = W*in
   wire signed [9:0] m175_8;
   assign m175_8 =10'b0;

   // m175_9 = W*in
   wire signed [9:0] m175_9;
   assign m175_9 =10'b0;

   // m175_10 = W*in
   wire signed [9:0] m175_10;
   assign m175_10 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_11 = W*in
   wire signed [9:0] m175_11;
   assign m175_11 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_12 = W*in
   wire signed [9:0] m175_12;
   assign m175_12 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_13 = W*in
   wire signed [9:0] m175_13;
   assign m175_13 =10'b0;

   // m175_14 = W*in
   wire signed [9:0] m175_14;
   assign m175_14 =10'b0;

   // m175_15 = W*in
   wire signed [9:0] m175_15;
   assign m175_15 =10'b0;

   // m175_16 = W*in
   wire signed [9:0] m175_16;
   assign m175_16 ={ {4{in175[5]}} , in175[5:0] };

   // m175_17 = W*in
   wire signed [9:0] m175_17;
   assign m175_17 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_18 = W*in
   wire signed [9:0] m175_18;
   assign m175_18 ={ {4{in175[5]}} , in175[5:0] };

   // m175_19 = W*in
   wire signed [9:0] m175_19;
   assign m175_19 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_20 = W*in
   wire signed [9:0] m175_20;
   assign m175_20 ={ {4{in175[5]}} , in175[5:0] };

   // m175_21 = W*in
   wire signed [9:0] m175_21;
   assign m175_21 =10'b0;

   // m175_22 = W*in
   wire signed [9:0] m175_22;
   assign m175_22 =10'b0;

   // m175_23 = W*in
   wire signed [9:0] m175_23;
   assign m175_23 =10'b0;

   // m175_24 = W*in
   wire signed [9:0] m175_24;
   assign m175_24 =10'b0;

   // m175_25 = W*in
   wire signed [9:0] m175_25;
   assign m175_25 =10'b0;

   // m175_26 = W*in
   wire signed [9:0] m175_26;
   assign m175_26 =10'b0;

   // m175_27 = W*in
   wire signed [9:0] m175_27;
   assign m175_27 =10'b0;

   // m175_28 = W*in
   wire signed [9:0] m175_28;
   assign m175_28 =10'b0;

   // m175_29 = W*in
   wire signed [9:0] m175_29;
   assign m175_29 =10'b0;

   // m175_30 = W*in
   wire signed [9:0] m175_30;
   assign m175_30 ={ {4{in175[5]}} , in175[5:0] };

   // m175_31 = W*in
   wire signed [9:0] m175_31;
   assign m175_31 =10'b0;

   // m175_32 = W*in
   wire signed [9:0] m175_32;
   assign m175_32 =10'b0;

   // m175_33 = W*in
   wire signed [9:0] m175_33;
   assign m175_33 =10'b0;

   // m175_34 = W*in
   wire signed [9:0] m175_34;
   assign m175_34 ={ {4{in175[5]}} , in175[5:0] };

   // m175_35 = W*in
   wire signed [9:0] m175_35;
   assign m175_35 =10'b0;

   // m175_36 = W*in
   wire signed [9:0] m175_36;
   assign m175_36 =10'b0;

   // m175_37 = W*in
   wire signed [9:0] m175_37;
   assign m175_37 =10'b0;

   // m175_38 = W*in
   wire signed [9:0] m175_38;
   assign m175_38 =10'b0;

   // m175_39 = W*in
   wire signed [9:0] m175_39;
   assign m175_39 =10'b0;

   // m175_40 = W*in
   wire signed [9:0] m175_40;
   assign m175_40 =10'b0;

   // m175_41 = W*in
   wire signed [9:0] m175_41;
   assign m175_41 =10'b0;

   // m175_42 = W*in
   wire signed [9:0] m175_42;
   assign m175_42 ={ {4{in175[5]}} , in175[5:0] };

   // m175_43 = W*in
   wire signed [9:0] m175_43;
   assign m175_43 ={ {5{in175[5]}} , in175[5:1] };

   // m175_44 = W*in
   wire signed [9:0] m175_44;
   assign m175_44 =10'b0;

   // m175_45 = W*in
   wire signed [9:0] m175_45;
   assign m175_45 =10'b0;

   // m175_46 = W*in
   wire signed [9:0] m175_46;
   assign m175_46 =10'b0;

   // m175_47 = W*in
   wire signed [9:0] m175_47;
   assign m175_47 =10'b0;

   // m175_48 = W*in
   wire signed [9:0] m175_48;
   assign m175_48 =10'b0;

   // m175_49 = W*in
   wire signed [9:0] m175_49;
   assign m175_49 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_50 = W*in
   wire signed [9:0] m175_50;
   assign m175_50 =10'b0;

   // m175_51 = W*in
   wire signed [9:0] m175_51;
   assign m175_51 =10'b0;

   // m175_52 = W*in
   wire signed [9:0] m175_52;
   assign m175_52 =10'b0;

   // m175_53 = W*in
   wire signed [9:0] m175_53;
   assign m175_53 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_54 = W*in
   wire signed [9:0] m175_54;
   assign m175_54 =10'b0;

   // m175_55 = W*in
   wire signed [9:0] m175_55;
   assign m175_55 ={ {4{in175[5]}} , in175[5:0] };

   // m175_56 = W*in
   wire signed [9:0] m175_56;
   assign m175_56 ={ {4{in175[5]}} , in175[5:0] };

   // m175_57 = W*in
   wire signed [9:0] m175_57;
   assign m175_57 =10'b0;

   // m175_58 = W*in
   wire signed [9:0] m175_58;
   assign m175_58 =10'b0;

   // m175_59 = W*in
   wire signed [9:0] m175_59;
   assign m175_59 =10'b0;

   // m175_60 = W*in
   wire signed [9:0] m175_60;
   assign m175_60 =10'b0;

   // m175_61 = W*in
   wire signed [9:0] m175_61;
   assign m175_61 =10'b0;

   // m175_62 = W*in
   wire signed [9:0] m175_62;
   assign m175_62 =10'b0;

   // m175_63 = W*in
   wire signed [9:0] m175_63;
   assign m175_63 =10'b0;

   // m175_64 = W*in
   wire signed [9:0] m175_64;
   assign m175_64 ={ {4{in175[5]}} , in175[5:0] };

   // m175_65 = W*in
   wire signed [9:0] m175_65;
   assign m175_65 =10'b0;

   // m175_66 = W*in
   wire signed [9:0] m175_66;
   assign m175_66 ={ {5{neg175[5]}} , neg175[5:1] };

   // m175_67 = W*in
   wire signed [9:0] m175_67;
   assign m175_67 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_68 = W*in
   wire signed [9:0] m175_68;
   assign m175_68 =10'b0;

   // m175_69 = W*in
   wire signed [9:0] m175_69;
   assign m175_69 =10'b0;

   // m175_70 = W*in
   wire signed [9:0] m175_70;
   assign m175_70 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_71 = W*in
   wire signed [9:0] m175_71;
   assign m175_71 =10'b0;

   // m175_72 = W*in
   wire signed [9:0] m175_72;
   assign m175_72 =10'b0;

   // m175_73 = W*in
   wire signed [9:0] m175_73;
   assign m175_73 =10'b0;

   // m175_74 = W*in
   wire signed [9:0] m175_74;
   assign m175_74 =10'b0;

   // m175_75 = W*in
   wire signed [9:0] m175_75;
   assign m175_75 =10'b0;

   // m175_76 = W*in
   wire signed [9:0] m175_76;
   assign m175_76 ={ {4{in175[5]}} , in175[5:0] };

   // m175_77 = W*in
   wire signed [9:0] m175_77;
   assign m175_77 =10'b0;

   // m175_78 = W*in
   wire signed [9:0] m175_78;
   assign m175_78 =10'b0;

   // m175_79 = W*in
   wire signed [9:0] m175_79;
   assign m175_79 =10'b0;

   // m175_80 = W*in
   wire signed [9:0] m175_80;
   assign m175_80 =10'b0;

   // m175_81 = W*in
   wire signed [9:0] m175_81;
   assign m175_81 ={ {4{in175[5]}} , in175[5:0] };

   // m175_82 = W*in
   wire signed [9:0] m175_82;
   assign m175_82 =10'b0;

   // m175_83 = W*in
   wire signed [9:0] m175_83;
   assign m175_83 ={ {5{neg175[5]}} , neg175[5:1] };

   // m175_84 = W*in
   wire signed [9:0] m175_84;
   assign m175_84 =10'b0;

   // m175_85 = W*in
   wire signed [9:0] m175_85;
   assign m175_85 =10'b0;

   // m175_86 = W*in
   wire signed [9:0] m175_86;
   assign m175_86 =10'b0;

   // m175_87 = W*in
   wire signed [9:0] m175_87;
   assign m175_87 ={ {4{in175[5]}} , in175[5:0] };

   // m175_88 = W*in
   wire signed [9:0] m175_88;
   assign m175_88 =10'b0;

   // m175_89 = W*in
   wire signed [9:0] m175_89;
   assign m175_89 ={ {4{in175[5]}} , in175[5:0] };

   // m175_90 = W*in
   wire signed [9:0] m175_90;
   assign m175_90 =10'b0;

   // m175_91 = W*in
   wire signed [9:0] m175_91;
   assign m175_91 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_92 = W*in
   wire signed [9:0] m175_92;
   assign m175_92 =10'b0;

   // m175_93 = W*in
   wire signed [9:0] m175_93;
   assign m175_93 =10'b0;

   // m175_94 = W*in
   wire signed [9:0] m175_94;
   assign m175_94 ={ {4{in175[5]}} , in175[5:0] };

   // m175_95 = W*in
   wire signed [9:0] m175_95;
   assign m175_95 =10'b0;

   // m175_96 = W*in
   wire signed [9:0] m175_96;
   assign m175_96 =10'b0;

   // m175_97 = W*in
   wire signed [9:0] m175_97;
   assign m175_97 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_98 = W*in
   wire signed [9:0] m175_98;
   assign m175_98 =10'b0;

   // m175_99 = W*in
   wire signed [9:0] m175_99;
   assign m175_99 ={ {4{in175[5]}} , in175[5:0] };

   // m175_100 = W*in
   wire signed [9:0] m175_100;
   assign m175_100 =10'b0;

   // m175_101 = W*in
   wire signed [9:0] m175_101;
   assign m175_101 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_102 = W*in
   wire signed [9:0] m175_102;
   assign m175_102 =10'b0;

   // m175_103 = W*in
   wire signed [9:0] m175_103;
   assign m175_103 =10'b0;

   // m175_104 = W*in
   wire signed [9:0] m175_104;
   assign m175_104 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_105 = W*in
   wire signed [9:0] m175_105;
   assign m175_105 =10'b0;

   // m175_106 = W*in
   wire signed [9:0] m175_106;
   assign m175_106 ={ {4{in175[5]}} , in175[5:0] };

   // m175_107 = W*in
   wire signed [9:0] m175_107;
   assign m175_107 ={ {4{neg175[5]}} , neg175[5:0] };

   // m175_108 = W*in
   wire signed [9:0] m175_108;
   assign m175_108 ={ {4{in175[5]}} , in175[5:0] };

   // m175_109 = W*in
   wire signed [9:0] m175_109;
   assign m175_109 =10'b0;

   // m175_110 = W*in
   wire signed [9:0] m175_110;
   assign m175_110 =10'b0;

   // m175_111 = W*in
   wire signed [9:0] m175_111;
   assign m175_111 ={ {4{in175[5]}} , in175[5:0] };

   // m175_112 = W*in
   wire signed [9:0] m175_112;
   assign m175_112 =10'b0;

   // m175_113 = W*in
   wire signed [9:0] m175_113;
   assign m175_113 ={ {4{in175[5]}} , in175[5:0] };

   // m175_114 = W*in
   wire signed [9:0] m175_114;
   assign m175_114 ={ {4{in175[5]}} , in175[5:0] };

   // m175_115 = W*in
   wire signed [9:0] m175_115;
   assign m175_115 ={ {4{in175[5]}} , in175[5:0] };

   // m175_116 = W*in
   wire signed [9:0] m175_116;
   assign m175_116 =10'b0;

   // m175_117 = W*in
   wire signed [9:0] m175_117;
   assign m175_117 =10'b0;

   // m176_1 = W*in
   wire signed [9:0] m176_1;
   assign m176_1 =10'b0;

   // m176_2 = W*in
   wire signed [9:0] m176_2;
   assign m176_2 =10'b0;

   // m176_3 = W*in
   wire signed [9:0] m176_3;
   assign m176_3 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_4 = W*in
   wire signed [9:0] m176_4;
   assign m176_4 =10'b0;

   // m176_5 = W*in
   wire signed [9:0] m176_5;
   assign m176_5 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_6 = W*in
   wire signed [9:0] m176_6;
   assign m176_6 =10'b0;

   // m176_7 = W*in
   wire signed [9:0] m176_7;
   assign m176_7 ={ {5{in176[5]}} , in176[5:1] };

   // m176_8 = W*in
   wire signed [9:0] m176_8;
   assign m176_8 =10'b0;

   // m176_9 = W*in
   wire signed [9:0] m176_9;
   assign m176_9 =10'b0;

   // m176_10 = W*in
   wire signed [9:0] m176_10;
   assign m176_10 =10'b0;

   // m176_11 = W*in
   wire signed [9:0] m176_11;
   assign m176_11 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_12 = W*in
   wire signed [9:0] m176_12;
   assign m176_12 =10'b0;

   // m176_13 = W*in
   wire signed [9:0] m176_13;
   assign m176_13 =10'b0;

   // m176_14 = W*in
   wire signed [9:0] m176_14;
   assign m176_14 ={ {4{in176[5]}} , in176[5:0] };

   // m176_15 = W*in
   wire signed [9:0] m176_15;
   assign m176_15 =10'b0;

   // m176_16 = W*in
   wire signed [9:0] m176_16;
   assign m176_16 =10'b0;

   // m176_17 = W*in
   wire signed [9:0] m176_17;
   assign m176_17 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_18 = W*in
   wire signed [9:0] m176_18;
   assign m176_18 ={ {3{in176[5]}} , in176 , {1{1'b0}} };

   // m176_19 = W*in
   wire signed [9:0] m176_19;
   assign m176_19 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_20 = W*in
   wire signed [9:0] m176_20;
   assign m176_20 =10'b0;

   // m176_21 = W*in
   wire signed [9:0] m176_21;
   assign m176_21 =10'b0;

   // m176_22 = W*in
   wire signed [9:0] m176_22;
   assign m176_22 =10'b0;

   // m176_23 = W*in
   wire signed [9:0] m176_23;
   assign m176_23 =10'b0;

   // m176_24 = W*in
   wire signed [9:0] m176_24;
   assign m176_24 =10'b0;

   // m176_25 = W*in
   wire signed [9:0] m176_25;
   assign m176_25 =10'b0;

   // m176_26 = W*in
   wire signed [9:0] m176_26;
   assign m176_26 ={ {4{in176[5]}} , in176[5:0] };

   // m176_27 = W*in
   wire signed [9:0] m176_27;
   assign m176_27 =10'b0;

   // m176_28 = W*in
   wire signed [9:0] m176_28;
   assign m176_28 =10'b0;

   // m176_29 = W*in
   wire signed [9:0] m176_29;
   assign m176_29 =10'b0;

   // m176_30 = W*in
   wire signed [9:0] m176_30;
   assign m176_30 =10'b0;

   // m176_31 = W*in
   wire signed [9:0] m176_31;
   assign m176_31 =10'b0;

   // m176_32 = W*in
   wire signed [9:0] m176_32;
   assign m176_32 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_33 = W*in
   wire signed [9:0] m176_33;
   assign m176_33 ={ {4{in176[5]}} , in176[5:0] };

   // m176_34 = W*in
   wire signed [9:0] m176_34;
   assign m176_34 =10'b0;

   // m176_35 = W*in
   wire signed [9:0] m176_35;
   assign m176_35 =10'b0;

   // m176_36 = W*in
   wire signed [9:0] m176_36;
   assign m176_36 =10'b0;

   // m176_37 = W*in
   wire signed [9:0] m176_37;
   assign m176_37 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_38 = W*in
   wire signed [9:0] m176_38;
   assign m176_38 ={ {4{in176[5]}} , in176[5:0] };

   // m176_39 = W*in
   wire signed [9:0] m176_39;
   assign m176_39 =10'b0;

   // m176_40 = W*in
   wire signed [9:0] m176_40;
   assign m176_40 =10'b0;

   // m176_41 = W*in
   wire signed [9:0] m176_41;
   assign m176_41 =10'b0;

   // m176_42 = W*in
   wire signed [9:0] m176_42;
   assign m176_42 =10'b0;

   // m176_43 = W*in
   wire signed [9:0] m176_43;
   assign m176_43 =10'b0;

   // m176_44 = W*in
   wire signed [9:0] m176_44;
   assign m176_44 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_45 = W*in
   wire signed [9:0] m176_45;
   assign m176_45 =10'b0;

   // m176_46 = W*in
   wire signed [9:0] m176_46;
   assign m176_46 =10'b0;

   // m176_47 = W*in
   wire signed [9:0] m176_47;
   assign m176_47 ={ {4{in176[5]}} , in176[5:0] };

   // m176_48 = W*in
   wire signed [9:0] m176_48;
   assign m176_48 ={ {4{in176[5]}} , in176[5:0] };

   // m176_49 = W*in
   wire signed [9:0] m176_49;
   assign m176_49 =10'b0;

   // m176_50 = W*in
   wire signed [9:0] m176_50;
   assign m176_50 =10'b0;

   // m176_51 = W*in
   wire signed [9:0] m176_51;
   assign m176_51 =10'b0;

   // m176_52 = W*in
   wire signed [9:0] m176_52;
   assign m176_52 =10'b0;

   // m176_53 = W*in
   wire signed [9:0] m176_53;
   assign m176_53 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_54 = W*in
   wire signed [9:0] m176_54;
   assign m176_54 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_55 = W*in
   wire signed [9:0] m176_55;
   assign m176_55 ={ {4{in176[5]}} , in176[5:0] };

   // m176_56 = W*in
   wire signed [9:0] m176_56;
   assign m176_56 =10'b0;

   // m176_57 = W*in
   wire signed [9:0] m176_57;
   assign m176_57 =10'b0;

   // m176_58 = W*in
   wire signed [9:0] m176_58;
   assign m176_58 =10'b0;

   // m176_59 = W*in
   wire signed [9:0] m176_59;
   assign m176_59 =10'b0;

   // m176_60 = W*in
   wire signed [9:0] m176_60;
   assign m176_60 =10'b0;

   // m176_61 = W*in
   wire signed [9:0] m176_61;
   assign m176_61 ={ {5{neg176[5]}} , neg176[5:1] };

   // m176_62 = W*in
   wire signed [9:0] m176_62;
   assign m176_62 =10'b0;

   // m176_63 = W*in
   wire signed [9:0] m176_63;
   assign m176_63 =10'b0;

   // m176_64 = W*in
   wire signed [9:0] m176_64;
   assign m176_64 =10'b0;

   // m176_65 = W*in
   wire signed [9:0] m176_65;
   assign m176_65 =10'b0;

   // m176_66 = W*in
   wire signed [9:0] m176_66;
   assign m176_66 ={ {5{in176[5]}} , in176[5:1] };

   // m176_67 = W*in
   wire signed [9:0] m176_67;
   assign m176_67 ={ {3{neg176[5]}} , neg176 , {1{1'b0}} };

   // m176_68 = W*in
   wire signed [9:0] m176_68;
   assign m176_68 =10'b0;

   // m176_69 = W*in
   wire signed [9:0] m176_69;
   assign m176_69 ={ {4{in176[5]}} , in176[5:0] };

   // m176_70 = W*in
   wire signed [9:0] m176_70;
   assign m176_70 ={ {4{in176[5]}} , in176[5:0] };

   // m176_71 = W*in
   wire signed [9:0] m176_71;
   assign m176_71 ={ {4{in176[5]}} , in176[5:0] };

   // m176_72 = W*in
   wire signed [9:0] m176_72;
   assign m176_72 =10'b0;

   // m176_73 = W*in
   wire signed [9:0] m176_73;
   assign m176_73 ={ {5{neg176[5]}} , neg176[5:1] };

   // m176_74 = W*in
   wire signed [9:0] m176_74;
   assign m176_74 ={ {4{in176[5]}} , in176[5:0] };

   // m176_75 = W*in
   wire signed [9:0] m176_75;
   assign m176_75 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_76 = W*in
   wire signed [9:0] m176_76;
   assign m176_76 ={ {5{in176[5]}} , in176[5:1] };

   // m176_77 = W*in
   wire signed [9:0] m176_77;
   assign m176_77 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_78 = W*in
   wire signed [9:0] m176_78;
   assign m176_78 ={ {3{in176[5]}} , in176 , {1{1'b0}} };

   // m176_79 = W*in
   wire signed [9:0] m176_79;
   assign m176_79 =10'b0;

   // m176_80 = W*in
   wire signed [9:0] m176_80;
   assign m176_80 =10'b0;

   // m176_81 = W*in
   wire signed [9:0] m176_81;
   assign m176_81 =10'b0;

   // m176_82 = W*in
   wire signed [9:0] m176_82;
   assign m176_82 ={ {4{in176[5]}} , in176[5:0] };

   // m176_83 = W*in
   wire signed [9:0] m176_83;
   assign m176_83 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_84 = W*in
   wire signed [9:0] m176_84;
   assign m176_84 =10'b0;

   // m176_85 = W*in
   wire signed [9:0] m176_85;
   assign m176_85 =10'b0;

   // m176_86 = W*in
   wire signed [9:0] m176_86;
   assign m176_86 ={ {4{in176[5]}} , in176[5:0] };

   // m176_87 = W*in
   wire signed [9:0] m176_87;
   assign m176_87 ={ {4{in176[5]}} , in176[5:0] };

   // m176_88 = W*in
   wire signed [9:0] m176_88;
   assign m176_88 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_89 = W*in
   wire signed [9:0] m176_89;
   assign m176_89 =10'b0;

   // m176_90 = W*in
   wire signed [9:0] m176_90;
   assign m176_90 =10'b0;

   // m176_91 = W*in
   wire signed [9:0] m176_91;
   assign m176_91 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_92 = W*in
   wire signed [9:0] m176_92;
   assign m176_92 =10'b0;

   // m176_93 = W*in
   wire signed [9:0] m176_93;
   assign m176_93 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_94 = W*in
   wire signed [9:0] m176_94;
   assign m176_94 =10'b0;

   // m176_95 = W*in
   wire signed [9:0] m176_95;
   assign m176_95 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_96 = W*in
   wire signed [9:0] m176_96;
   assign m176_96 ={ {4{in176[5]}} , in176[5:0] };

   // m176_97 = W*in
   wire signed [9:0] m176_97;
   assign m176_97 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_98 = W*in
   wire signed [9:0] m176_98;
   assign m176_98 =10'b0;

   // m176_99 = W*in
   wire signed [9:0] m176_99;
   assign m176_99 ={ {4{in176[5]}} , in176[5:0] };

   // m176_100 = W*in
   wire signed [9:0] m176_100;
   assign m176_100 =10'b0;

   // m176_101 = W*in
   wire signed [9:0] m176_101;
   assign m176_101 =10'b0;

   // m176_102 = W*in
   wire signed [9:0] m176_102;
   assign m176_102 =10'b0;

   // m176_103 = W*in
   wire signed [9:0] m176_103;
   assign m176_103 =10'b0;

   // m176_104 = W*in
   wire signed [9:0] m176_104;
   assign m176_104 =10'b0;

   // m176_105 = W*in
   wire signed [9:0] m176_105;
   assign m176_105 =10'b0;

   // m176_106 = W*in
   wire signed [9:0] m176_106;
   assign m176_106 ={ {4{in176[5]}} , in176[5:0] };

   // m176_107 = W*in
   wire signed [9:0] m176_107;
   assign m176_107 ={ {4{neg176[5]}} , neg176[5:0] };

   // m176_108 = W*in
   wire signed [9:0] m176_108;
   assign m176_108 ={ {5{neg176[5]}} , neg176[5:1] };

   // m176_109 = W*in
   wire signed [9:0] m176_109;
   assign m176_109 ={ {5{in176[5]}} , in176[5:1] };

   // m176_110 = W*in
   wire signed [9:0] m176_110;
   assign m176_110 ={ {4{in176[5]}} , in176[5:0] };

   // m176_111 = W*in
   wire signed [9:0] m176_111;
   assign m176_111 =10'b0;

   // m176_112 = W*in
   wire signed [9:0] m176_112;
   assign m176_112 =10'b0;

   // m176_113 = W*in
   wire signed [9:0] m176_113;
   assign m176_113 =10'b0;

   // m176_114 = W*in
   wire signed [9:0] m176_114;
   assign m176_114 =10'b0;

   // m176_115 = W*in
   wire signed [9:0] m176_115;
   assign m176_115 =10'b0;

   // m176_116 = W*in
   wire signed [9:0] m176_116;
   assign m176_116 =10'b0;

   // m176_117 = W*in
   wire signed [9:0] m176_117;
   assign m176_117 =10'b0;

   // m177_1 = W*in
   wire signed [9:0] m177_1;
   assign m177_1 =10'b0;

   // m177_2 = W*in
   wire signed [9:0] m177_2;
   assign m177_2 ={ {4{in177[5]}} , in177[5:0] };

   // m177_3 = W*in
   wire signed [9:0] m177_3;
   assign m177_3 =10'b0;

   // m177_4 = W*in
   wire signed [9:0] m177_4;
   assign m177_4 =10'b0;

   // m177_5 = W*in
   wire signed [9:0] m177_5;
   assign m177_5 =10'b0;

   // m177_6 = W*in
   wire signed [9:0] m177_6;
   assign m177_6 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_7 = W*in
   wire signed [9:0] m177_7;
   assign m177_7 =10'b0;

   // m177_8 = W*in
   wire signed [9:0] m177_8;
   assign m177_8 ={ {4{in177[5]}} , in177[5:0] };

   // m177_9 = W*in
   wire signed [9:0] m177_9;
   assign m177_9 ={ {4{in177[5]}} , in177[5:0] };

   // m177_10 = W*in
   wire signed [9:0] m177_10;
   assign m177_10 ={ {4{in177[5]}} , in177[5:0] };

   // m177_11 = W*in
   wire signed [9:0] m177_11;
   assign m177_11 =10'b0;

   // m177_12 = W*in
   wire signed [9:0] m177_12;
   assign m177_12 ={ {4{in177[5]}} , in177[5:0] };

   // m177_13 = W*in
   wire signed [9:0] m177_13;
   assign m177_13 =10'b0;

   // m177_14 = W*in
   wire signed [9:0] m177_14;
   assign m177_14 ={ {4{in177[5]}} , in177[5:0] };

   // m177_15 = W*in
   wire signed [9:0] m177_15;
   assign m177_15 =10'b0;

   // m177_16 = W*in
   wire signed [9:0] m177_16;
   assign m177_16 ={ {4{in177[5]}} , in177[5:0] };

   // m177_17 = W*in
   wire signed [9:0] m177_17;
   assign m177_17 ={ {5{in177[5]}} , in177[5:1] };

   // m177_18 = W*in
   wire signed [9:0] m177_18;
   assign m177_18 ={ {4{in177[5]}} , in177[5:0] };

   // m177_19 = W*in
   wire signed [9:0] m177_19;
   assign m177_19 =10'b0;

   // m177_20 = W*in
   wire signed [9:0] m177_20;
   assign m177_20 ={ {5{neg177[5]}} , neg177[5:1] };

   // m177_21 = W*in
   wire signed [9:0] m177_21;
   assign m177_21 ={ {5{neg177[5]}} , neg177[5:1] };

   // m177_22 = W*in
   wire signed [9:0] m177_22;
   assign m177_22 =10'b0;

   // m177_23 = W*in
   wire signed [9:0] m177_23;
   assign m177_23 ={ {5{neg177[5]}} , neg177[5:1] };

   // m177_24 = W*in
   wire signed [9:0] m177_24;
   assign m177_24 =10'b0;

   // m177_25 = W*in
   wire signed [9:0] m177_25;
   assign m177_25 ={ {4{in177[5]}} , in177[5:0] };

   // m177_26 = W*in
   wire signed [9:0] m177_26;
   assign m177_26 =10'b0;

   // m177_27 = W*in
   wire signed [9:0] m177_27;
   assign m177_27 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_28 = W*in
   wire signed [9:0] m177_28;
   assign m177_28 =10'b0;

   // m177_29 = W*in
   wire signed [9:0] m177_29;
   assign m177_29 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_30 = W*in
   wire signed [9:0] m177_30;
   assign m177_30 =10'b0;

   // m177_31 = W*in
   wire signed [9:0] m177_31;
   assign m177_31 =10'b0;

   // m177_32 = W*in
   wire signed [9:0] m177_32;
   assign m177_32 =10'b0;

   // m177_33 = W*in
   wire signed [9:0] m177_33;
   assign m177_33 =10'b0;

   // m177_34 = W*in
   wire signed [9:0] m177_34;
   assign m177_34 =10'b0;

   // m177_35 = W*in
   wire signed [9:0] m177_35;
   assign m177_35 =10'b0;

   // m177_36 = W*in
   wire signed [9:0] m177_36;
   assign m177_36 =10'b0;

   // m177_37 = W*in
   wire signed [9:0] m177_37;
   assign m177_37 =10'b0;

   // m177_38 = W*in
   wire signed [9:0] m177_38;
   assign m177_38 =10'b0;

   // m177_39 = W*in
   wire signed [9:0] m177_39;
   assign m177_39 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_40 = W*in
   wire signed [9:0] m177_40;
   assign m177_40 =10'b0;

   // m177_41 = W*in
   wire signed [9:0] m177_41;
   assign m177_41 =10'b0;

   // m177_42 = W*in
   wire signed [9:0] m177_42;
   assign m177_42 ={ {4{in177[5]}} , in177[5:0] };

   // m177_43 = W*in
   wire signed [9:0] m177_43;
   assign m177_43 =10'b0;

   // m177_44 = W*in
   wire signed [9:0] m177_44;
   assign m177_44 =10'b0;

   // m177_45 = W*in
   wire signed [9:0] m177_45;
   assign m177_45 =10'b0;

   // m177_46 = W*in
   wire signed [9:0] m177_46;
   assign m177_46 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_47 = W*in
   wire signed [9:0] m177_47;
   assign m177_47 =10'b0;

   // m177_48 = W*in
   wire signed [9:0] m177_48;
   assign m177_48 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_49 = W*in
   wire signed [9:0] m177_49;
   assign m177_49 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_50 = W*in
   wire signed [9:0] m177_50;
   assign m177_50 =10'b0;

   // m177_51 = W*in
   wire signed [9:0] m177_51;
   assign m177_51 ={ {4{in177[5]}} , in177[5:0] };

   // m177_52 = W*in
   wire signed [9:0] m177_52;
   assign m177_52 ={ {4{in177[5]}} , in177[5:0] };

   // m177_53 = W*in
   wire signed [9:0] m177_53;
   assign m177_53 =10'b0;

   // m177_54 = W*in
   wire signed [9:0] m177_54;
   assign m177_54 =10'b0;

   // m177_55 = W*in
   wire signed [9:0] m177_55;
   assign m177_55 =10'b0;

   // m177_56 = W*in
   wire signed [9:0] m177_56;
   assign m177_56 ={ {4{in177[5]}} , in177[5:0] };

   // m177_57 = W*in
   wire signed [9:0] m177_57;
   assign m177_57 =10'b0;

   // m177_58 = W*in
   wire signed [9:0] m177_58;
   assign m177_58 =10'b0;

   // m177_59 = W*in
   wire signed [9:0] m177_59;
   assign m177_59 =10'b0;

   // m177_60 = W*in
   wire signed [9:0] m177_60;
   assign m177_60 =10'b0;

   // m177_61 = W*in
   wire signed [9:0] m177_61;
   assign m177_61 ={ {5{in177[5]}} , in177[5:1] };

   // m177_62 = W*in
   wire signed [9:0] m177_62;
   assign m177_62 =10'b0;

   // m177_63 = W*in
   wire signed [9:0] m177_63;
   assign m177_63 =10'b0;

   // m177_64 = W*in
   wire signed [9:0] m177_64;
   assign m177_64 ={ {4{in177[5]}} , in177[5:0] };

   // m177_65 = W*in
   wire signed [9:0] m177_65;
   assign m177_65 ={ {5{in177[5]}} , in177[5:1] };

   // m177_66 = W*in
   wire signed [9:0] m177_66;
   assign m177_66 =10'b0;

   // m177_67 = W*in
   wire signed [9:0] m177_67;
   assign m177_67 =10'b0;

   // m177_68 = W*in
   wire signed [9:0] m177_68;
   assign m177_68 ={ {4{in177[5]}} , in177[5:0] };

   // m177_69 = W*in
   wire signed [9:0] m177_69;
   assign m177_69 ={ {5{neg177[5]}} , neg177[5:1] };

   // m177_70 = W*in
   wire signed [9:0] m177_70;
   assign m177_70 =10'b0;

   // m177_71 = W*in
   wire signed [9:0] m177_71;
   assign m177_71 =10'b0;

   // m177_72 = W*in
   wire signed [9:0] m177_72;
   assign m177_72 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_73 = W*in
   wire signed [9:0] m177_73;
   assign m177_73 =10'b0;

   // m177_74 = W*in
   wire signed [9:0] m177_74;
   assign m177_74 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_75 = W*in
   wire signed [9:0] m177_75;
   assign m177_75 ={ {4{in177[5]}} , in177[5:0] };

   // m177_76 = W*in
   wire signed [9:0] m177_76;
   assign m177_76 =10'b0;

   // m177_77 = W*in
   wire signed [9:0] m177_77;
   assign m177_77 ={ {4{in177[5]}} , in177[5:0] };

   // m177_78 = W*in
   wire signed [9:0] m177_78;
   assign m177_78 =10'b0;

   // m177_79 = W*in
   wire signed [9:0] m177_79;
   assign m177_79 =10'b0;

   // m177_80 = W*in
   wire signed [9:0] m177_80;
   assign m177_80 ={ {4{in177[5]}} , in177[5:0] };

   // m177_81 = W*in
   wire signed [9:0] m177_81;
   assign m177_81 =10'b0;

   // m177_82 = W*in
   wire signed [9:0] m177_82;
   assign m177_82 =10'b0;

   // m177_83 = W*in
   wire signed [9:0] m177_83;
   assign m177_83 =10'b0;

   // m177_84 = W*in
   wire signed [9:0] m177_84;
   assign m177_84 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_85 = W*in
   wire signed [9:0] m177_85;
   assign m177_85 =10'b0;

   // m177_86 = W*in
   wire signed [9:0] m177_86;
   assign m177_86 =10'b0;

   // m177_87 = W*in
   wire signed [9:0] m177_87;
   assign m177_87 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_88 = W*in
   wire signed [9:0] m177_88;
   assign m177_88 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_89 = W*in
   wire signed [9:0] m177_89;
   assign m177_89 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_90 = W*in
   wire signed [9:0] m177_90;
   assign m177_90 =10'b0;

   // m177_91 = W*in
   wire signed [9:0] m177_91;
   assign m177_91 =10'b0;

   // m177_92 = W*in
   wire signed [9:0] m177_92;
   assign m177_92 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_93 = W*in
   wire signed [9:0] m177_93;
   assign m177_93 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_94 = W*in
   wire signed [9:0] m177_94;
   assign m177_94 ={ {4{in177[5]}} , in177[5:0] };

   // m177_95 = W*in
   wire signed [9:0] m177_95;
   assign m177_95 =10'b0;

   // m177_96 = W*in
   wire signed [9:0] m177_96;
   assign m177_96 =10'b0;

   // m177_97 = W*in
   wire signed [9:0] m177_97;
   assign m177_97 ={ {5{in177[5]}} , in177[5:1] };

   // m177_98 = W*in
   wire signed [9:0] m177_98;
   assign m177_98 =10'b0;

   // m177_99 = W*in
   wire signed [9:0] m177_99;
   assign m177_99 =10'b0;

   // m177_100 = W*in
   wire signed [9:0] m177_100;
   assign m177_100 ={ {4{in177[5]}} , in177[5:0] };

   // m177_101 = W*in
   wire signed [9:0] m177_101;
   assign m177_101 =10'b0;

   // m177_102 = W*in
   wire signed [9:0] m177_102;
   assign m177_102 =10'b0;

   // m177_103 = W*in
   wire signed [9:0] m177_103;
   assign m177_103 =10'b0;

   // m177_104 = W*in
   wire signed [9:0] m177_104;
   assign m177_104 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_105 = W*in
   wire signed [9:0] m177_105;
   assign m177_105 =10'b0;

   // m177_106 = W*in
   wire signed [9:0] m177_106;
   assign m177_106 =10'b0;

   // m177_107 = W*in
   wire signed [9:0] m177_107;
   assign m177_107 ={ {4{in177[5]}} , in177[5:0] };

   // m177_108 = W*in
   wire signed [9:0] m177_108;
   assign m177_108 =10'b0;

   // m177_109 = W*in
   wire signed [9:0] m177_109;
   assign m177_109 ={ {5{neg177[5]}} , neg177[5:1] };

   // m177_110 = W*in
   wire signed [9:0] m177_110;
   assign m177_110 ={ {4{neg177[5]}} , neg177[5:0] };

   // m177_111 = W*in
   wire signed [9:0] m177_111;
   assign m177_111 =10'b0;

   // m177_112 = W*in
   wire signed [9:0] m177_112;
   assign m177_112 ={ {4{in177[5]}} , in177[5:0] };

   // m177_113 = W*in
   wire signed [9:0] m177_113;
   assign m177_113 =10'b0;

   // m177_114 = W*in
   wire signed [9:0] m177_114;
   assign m177_114 ={ {5{neg177[5]}} , neg177[5:1] };

   // m177_115 = W*in
   wire signed [9:0] m177_115;
   assign m177_115 =10'b0;

   // m177_116 = W*in
   wire signed [9:0] m177_116;
   assign m177_116 =10'b0;

   // m177_117 = W*in
   wire signed [9:0] m177_117;
   assign m177_117 =10'b0;

   // m178_1 = W*in
   wire signed [9:0] m178_1;
   assign m178_1 =10'b0;

   // m178_2 = W*in
   wire signed [9:0] m178_2;
   assign m178_2 =10'b0;

   // m178_3 = W*in
   wire signed [9:0] m178_3;
   assign m178_3 =10'b0;

   // m178_4 = W*in
   wire signed [9:0] m178_4;
   assign m178_4 =10'b0;

   // m178_5 = W*in
   wire signed [9:0] m178_5;
   assign m178_5 =10'b0;

   // m178_6 = W*in
   wire signed [9:0] m178_6;
   assign m178_6 =10'b0;

   // m178_7 = W*in
   wire signed [9:0] m178_7;
   assign m178_7 ={ {4{in178[5]}} , in178[5:0] };

   // m178_8 = W*in
   wire signed [9:0] m178_8;
   assign m178_8 ={ {4{in178[5]}} , in178[5:0] };

   // m178_9 = W*in
   wire signed [9:0] m178_9;
   assign m178_9 =10'b0;

   // m178_10 = W*in
   wire signed [9:0] m178_10;
   assign m178_10 =10'b0;

   // m178_11 = W*in
   wire signed [9:0] m178_11;
   assign m178_11 =10'b0;

   // m178_12 = W*in
   wire signed [9:0] m178_12;
   assign m178_12 ={ {4{in178[5]}} , in178[5:0] };

   // m178_13 = W*in
   wire signed [9:0] m178_13;
   assign m178_13 =10'b0;

   // m178_14 = W*in
   wire signed [9:0] m178_14;
   assign m178_14 =10'b0;

   // m178_15 = W*in
   wire signed [9:0] m178_15;
   assign m178_15 =10'b0;

   // m178_16 = W*in
   wire signed [9:0] m178_16;
   assign m178_16 =10'b0;

   // m178_17 = W*in
   wire signed [9:0] m178_17;
   assign m178_17 =10'b0;

   // m178_18 = W*in
   wire signed [9:0] m178_18;
   assign m178_18 =10'b0;

   // m178_19 = W*in
   wire signed [9:0] m178_19;
   assign m178_19 =10'b0;

   // m178_20 = W*in
   wire signed [9:0] m178_20;
   assign m178_20 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_21 = W*in
   wire signed [9:0] m178_21;
   assign m178_21 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_22 = W*in
   wire signed [9:0] m178_22;
   assign m178_22 =10'b0;

   // m178_23 = W*in
   wire signed [9:0] m178_23;
   assign m178_23 =10'b0;

   // m178_24 = W*in
   wire signed [9:0] m178_24;
   assign m178_24 =10'b0;

   // m178_25 = W*in
   wire signed [9:0] m178_25;
   assign m178_25 ={ {4{in178[5]}} , in178[5:0] };

   // m178_26 = W*in
   wire signed [9:0] m178_26;
   assign m178_26 =10'b0;

   // m178_27 = W*in
   wire signed [9:0] m178_27;
   assign m178_27 =10'b0;

   // m178_28 = W*in
   wire signed [9:0] m178_28;
   assign m178_28 ={ {4{in178[5]}} , in178[5:0] };

   // m178_29 = W*in
   wire signed [9:0] m178_29;
   assign m178_29 =10'b0;

   // m178_30 = W*in
   wire signed [9:0] m178_30;
   assign m178_30 =10'b0;

   // m178_31 = W*in
   wire signed [9:0] m178_31;
   assign m178_31 ={ {5{in178[5]}} , in178[5:1] };

   // m178_32 = W*in
   wire signed [9:0] m178_32;
   assign m178_32 =10'b0;

   // m178_33 = W*in
   wire signed [9:0] m178_33;
   assign m178_33 ={ {4{in178[5]}} , in178[5:0] };

   // m178_34 = W*in
   wire signed [9:0] m178_34;
   assign m178_34 =10'b0;

   // m178_35 = W*in
   wire signed [9:0] m178_35;
   assign m178_35 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_36 = W*in
   wire signed [9:0] m178_36;
   assign m178_36 =10'b0;

   // m178_37 = W*in
   wire signed [9:0] m178_37;
   assign m178_37 =10'b0;

   // m178_38 = W*in
   wire signed [9:0] m178_38;
   assign m178_38 =10'b0;

   // m178_39 = W*in
   wire signed [9:0] m178_39;
   assign m178_39 =10'b0;

   // m178_40 = W*in
   wire signed [9:0] m178_40;
   assign m178_40 =10'b0;

   // m178_41 = W*in
   wire signed [9:0] m178_41;
   assign m178_41 =10'b0;

   // m178_42 = W*in
   wire signed [9:0] m178_42;
   assign m178_42 =10'b0;

   // m178_43 = W*in
   wire signed [9:0] m178_43;
   assign m178_43 =10'b0;

   // m178_44 = W*in
   wire signed [9:0] m178_44;
   assign m178_44 =10'b0;

   // m178_45 = W*in
   wire signed [9:0] m178_45;
   assign m178_45 =10'b0;

   // m178_46 = W*in
   wire signed [9:0] m178_46;
   assign m178_46 =10'b0;

   // m178_47 = W*in
   wire signed [9:0] m178_47;
   assign m178_47 =10'b0;

   // m178_48 = W*in
   wire signed [9:0] m178_48;
   assign m178_48 =10'b0;

   // m178_49 = W*in
   wire signed [9:0] m178_49;
   assign m178_49 =10'b0;

   // m178_50 = W*in
   wire signed [9:0] m178_50;
   assign m178_50 =10'b0;

   // m178_51 = W*in
   wire signed [9:0] m178_51;
   assign m178_51 ={ {4{in178[5]}} , in178[5:0] };

   // m178_52 = W*in
   wire signed [9:0] m178_52;
   assign m178_52 ={ {4{in178[5]}} , in178[5:0] };

   // m178_53 = W*in
   wire signed [9:0] m178_53;
   assign m178_53 =10'b0;

   // m178_54 = W*in
   wire signed [9:0] m178_54;
   assign m178_54 =10'b0;

   // m178_55 = W*in
   wire signed [9:0] m178_55;
   assign m178_55 =10'b0;

   // m178_56 = W*in
   wire signed [9:0] m178_56;
   assign m178_56 =10'b0;

   // m178_57 = W*in
   wire signed [9:0] m178_57;
   assign m178_57 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_58 = W*in
   wire signed [9:0] m178_58;
   assign m178_58 =10'b0;

   // m178_59 = W*in
   wire signed [9:0] m178_59;
   assign m178_59 ={ {4{in178[5]}} , in178[5:0] };

   // m178_60 = W*in
   wire signed [9:0] m178_60;
   assign m178_60 =10'b0;

   // m178_61 = W*in
   wire signed [9:0] m178_61;
   assign m178_61 =10'b0;

   // m178_62 = W*in
   wire signed [9:0] m178_62;
   assign m178_62 =10'b0;

   // m178_63 = W*in
   wire signed [9:0] m178_63;
   assign m178_63 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_64 = W*in
   wire signed [9:0] m178_64;
   assign m178_64 =10'b0;

   // m178_65 = W*in
   wire signed [9:0] m178_65;
   assign m178_65 =10'b0;

   // m178_66 = W*in
   wire signed [9:0] m178_66;
   assign m178_66 =10'b0;

   // m178_67 = W*in
   wire signed [9:0] m178_67;
   assign m178_67 =10'b0;

   // m178_68 = W*in
   wire signed [9:0] m178_68;
   assign m178_68 ={ {4{in178[5]}} , in178[5:0] };

   // m178_69 = W*in
   wire signed [9:0] m178_69;
   assign m178_69 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_70 = W*in
   wire signed [9:0] m178_70;
   assign m178_70 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_71 = W*in
   wire signed [9:0] m178_71;
   assign m178_71 =10'b0;

   // m178_72 = W*in
   wire signed [9:0] m178_72;
   assign m178_72 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_73 = W*in
   wire signed [9:0] m178_73;
   assign m178_73 ={ {4{in178[5]}} , in178[5:0] };

   // m178_74 = W*in
   wire signed [9:0] m178_74;
   assign m178_74 =10'b0;

   // m178_75 = W*in
   wire signed [9:0] m178_75;
   assign m178_75 ={ {5{neg178[5]}} , neg178[5:1] };

   // m178_76 = W*in
   wire signed [9:0] m178_76;
   assign m178_76 =10'b0;

   // m178_77 = W*in
   wire signed [9:0] m178_77;
   assign m178_77 =10'b0;

   // m178_78 = W*in
   wire signed [9:0] m178_78;
   assign m178_78 ={ {4{in178[5]}} , in178[5:0] };

   // m178_79 = W*in
   wire signed [9:0] m178_79;
   assign m178_79 =10'b0;

   // m178_80 = W*in
   wire signed [9:0] m178_80;
   assign m178_80 =10'b0;

   // m178_81 = W*in
   wire signed [9:0] m178_81;
   assign m178_81 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_82 = W*in
   wire signed [9:0] m178_82;
   assign m178_82 ={ {5{neg178[5]}} , neg178[5:1] };

   // m178_83 = W*in
   wire signed [9:0] m178_83;
   assign m178_83 ={ {5{neg178[5]}} , neg178[5:1] };

   // m178_84 = W*in
   wire signed [9:0] m178_84;
   assign m178_84 =10'b0;

   // m178_85 = W*in
   wire signed [9:0] m178_85;
   assign m178_85 =10'b0;

   // m178_86 = W*in
   wire signed [9:0] m178_86;
   assign m178_86 =10'b0;

   // m178_87 = W*in
   wire signed [9:0] m178_87;
   assign m178_87 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_88 = W*in
   wire signed [9:0] m178_88;
   assign m178_88 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_89 = W*in
   wire signed [9:0] m178_89;
   assign m178_89 =10'b0;

   // m178_90 = W*in
   wire signed [9:0] m178_90;
   assign m178_90 =10'b0;

   // m178_91 = W*in
   wire signed [9:0] m178_91;
   assign m178_91 =10'b0;

   // m178_92 = W*in
   wire signed [9:0] m178_92;
   assign m178_92 =10'b0;

   // m178_93 = W*in
   wire signed [9:0] m178_93;
   assign m178_93 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_94 = W*in
   wire signed [9:0] m178_94;
   assign m178_94 =10'b0;

   // m178_95 = W*in
   wire signed [9:0] m178_95;
   assign m178_95 =10'b0;

   // m178_96 = W*in
   wire signed [9:0] m178_96;
   assign m178_96 =10'b0;

   // m178_97 = W*in
   wire signed [9:0] m178_97;
   assign m178_97 =10'b0;

   // m178_98 = W*in
   wire signed [9:0] m178_98;
   assign m178_98 =10'b0;

   // m178_99 = W*in
   wire signed [9:0] m178_99;
   assign m178_99 =10'b0;

   // m178_100 = W*in
   wire signed [9:0] m178_100;
   assign m178_100 =10'b0;

   // m178_101 = W*in
   wire signed [9:0] m178_101;
   assign m178_101 =10'b0;

   // m178_102 = W*in
   wire signed [9:0] m178_102;
   assign m178_102 =10'b0;

   // m178_103 = W*in
   wire signed [9:0] m178_103;
   assign m178_103 =10'b0;

   // m178_104 = W*in
   wire signed [9:0] m178_104;
   assign m178_104 ={ {4{in178[5]}} , in178[5:0] };

   // m178_105 = W*in
   wire signed [9:0] m178_105;
   assign m178_105 =10'b0;

   // m178_106 = W*in
   wire signed [9:0] m178_106;
   assign m178_106 =10'b0;

   // m178_107 = W*in
   wire signed [9:0] m178_107;
   assign m178_107 =10'b0;

   // m178_108 = W*in
   wire signed [9:0] m178_108;
   assign m178_108 ={ {4{neg178[5]}} , neg178[5:0] };

   // m178_109 = W*in
   wire signed [9:0] m178_109;
   assign m178_109 =10'b0;

   // m178_110 = W*in
   wire signed [9:0] m178_110;
   assign m178_110 =10'b0;

   // m178_111 = W*in
   wire signed [9:0] m178_111;
   assign m178_111 =10'b0;

   // m178_112 = W*in
   wire signed [9:0] m178_112;
   assign m178_112 =10'b0;

   // m178_113 = W*in
   wire signed [9:0] m178_113;
   assign m178_113 =10'b0;

   // m178_114 = W*in
   wire signed [9:0] m178_114;
   assign m178_114 ={ {5{neg178[5]}} , neg178[5:1] };

   // m178_115 = W*in
   wire signed [9:0] m178_115;
   assign m178_115 =10'b0;

   // m178_116 = W*in
   wire signed [9:0] m178_116;
   assign m178_116 =10'b0;

   // m178_117 = W*in
   wire signed [9:0] m178_117;
   assign m178_117 =10'b0;

   // m179_1 = W*in
   wire signed [9:0] m179_1;
   assign m179_1 =10'b0;

   // m179_2 = W*in
   wire signed [9:0] m179_2;
   assign m179_2 =10'b0;

   // m179_3 = W*in
   wire signed [9:0] m179_3;
   assign m179_3 =10'b0;

   // m179_4 = W*in
   wire signed [9:0] m179_4;
   assign m179_4 =10'b0;

   // m179_5 = W*in
   wire signed [9:0] m179_5;
   assign m179_5 =10'b0;

   // m179_6 = W*in
   wire signed [9:0] m179_6;
   assign m179_6 =10'b0;

   // m179_7 = W*in
   wire signed [9:0] m179_7;
   assign m179_7 =10'b0;

   // m179_8 = W*in
   wire signed [9:0] m179_8;
   assign m179_8 =10'b0;

   // m179_9 = W*in
   wire signed [9:0] m179_9;
   assign m179_9 =10'b0;

   // m179_10 = W*in
   wire signed [9:0] m179_10;
   assign m179_10 =10'b0;

   // m179_11 = W*in
   wire signed [9:0] m179_11;
   assign m179_11 =10'b0;

   // m179_12 = W*in
   wire signed [9:0] m179_12;
   assign m179_12 =10'b0;

   // m179_13 = W*in
   wire signed [9:0] m179_13;
   assign m179_13 =10'b0;

   // m179_14 = W*in
   wire signed [9:0] m179_14;
   assign m179_14 =10'b0;

   // m179_15 = W*in
   wire signed [9:0] m179_15;
   assign m179_15 =10'b0;

   // m179_16 = W*in
   wire signed [9:0] m179_16;
   assign m179_16 =10'b0;

   // m179_17 = W*in
   wire signed [9:0] m179_17;
   assign m179_17 =10'b0;

   // m179_18 = W*in
   wire signed [9:0] m179_18;
   assign m179_18 =10'b0;

   // m179_19 = W*in
   wire signed [9:0] m179_19;
   assign m179_19 =10'b0;

   // m179_20 = W*in
   wire signed [9:0] m179_20;
   assign m179_20 =10'b0;

   // m179_21 = W*in
   wire signed [9:0] m179_21;
   assign m179_21 =10'b0;

   // m179_22 = W*in
   wire signed [9:0] m179_22;
   assign m179_22 ={ {5{in179[5]}} , in179[5:1] };

   // m179_23 = W*in
   wire signed [9:0] m179_23;
   assign m179_23 ={ {5{in179[5]}} , in179[5:1] };

   // m179_24 = W*in
   wire signed [9:0] m179_24;
   assign m179_24 =10'b0;

   // m179_25 = W*in
   wire signed [9:0] m179_25;
   assign m179_25 =10'b0;

   // m179_26 = W*in
   wire signed [9:0] m179_26;
   assign m179_26 =10'b0;

   // m179_27 = W*in
   wire signed [9:0] m179_27;
   assign m179_27 ={ {5{in179[5]}} , in179[5:1] };

   // m179_28 = W*in
   wire signed [9:0] m179_28;
   assign m179_28 =10'b0;

   // m179_29 = W*in
   wire signed [9:0] m179_29;
   assign m179_29 =10'b0;

   // m179_30 = W*in
   wire signed [9:0] m179_30;
   assign m179_30 =10'b0;

   // m179_31 = W*in
   wire signed [9:0] m179_31;
   assign m179_31 ={ {5{in179[5]}} , in179[5:1] };

   // m179_32 = W*in
   wire signed [9:0] m179_32;
   assign m179_32 =10'b0;

   // m179_33 = W*in
   wire signed [9:0] m179_33;
   assign m179_33 =10'b0;

   // m179_34 = W*in
   wire signed [9:0] m179_34;
   assign m179_34 =10'b0;

   // m179_35 = W*in
   wire signed [9:0] m179_35;
   assign m179_35 =10'b0;

   // m179_36 = W*in
   wire signed [9:0] m179_36;
   assign m179_36 ={ {5{in179[5]}} , in179[5:1] };

   // m179_37 = W*in
   wire signed [9:0] m179_37;
   assign m179_37 =10'b0;

   // m179_38 = W*in
   wire signed [9:0] m179_38;
   assign m179_38 =10'b0;

   // m179_39 = W*in
   wire signed [9:0] m179_39;
   assign m179_39 =10'b0;

   // m179_40 = W*in
   wire signed [9:0] m179_40;
   assign m179_40 =10'b0;

   // m179_41 = W*in
   wire signed [9:0] m179_41;
   assign m179_41 =10'b0;

   // m179_42 = W*in
   wire signed [9:0] m179_42;
   assign m179_42 =10'b0;

   // m179_43 = W*in
   wire signed [9:0] m179_43;
   assign m179_43 =10'b0;

   // m179_44 = W*in
   wire signed [9:0] m179_44;
   assign m179_44 =10'b0;

   // m179_45 = W*in
   wire signed [9:0] m179_45;
   assign m179_45 =10'b0;

   // m179_46 = W*in
   wire signed [9:0] m179_46;
   assign m179_46 =10'b0;

   // m179_47 = W*in
   wire signed [9:0] m179_47;
   assign m179_47 =10'b0;

   // m179_48 = W*in
   wire signed [9:0] m179_48;
   assign m179_48 =10'b0;

   // m179_49 = W*in
   wire signed [9:0] m179_49;
   assign m179_49 =10'b0;

   // m179_50 = W*in
   wire signed [9:0] m179_50;
   assign m179_50 =10'b0;

   // m179_51 = W*in
   wire signed [9:0] m179_51;
   assign m179_51 =10'b0;

   // m179_52 = W*in
   wire signed [9:0] m179_52;
   assign m179_52 =10'b0;

   // m179_53 = W*in
   wire signed [9:0] m179_53;
   assign m179_53 =10'b0;

   // m179_54 = W*in
   wire signed [9:0] m179_54;
   assign m179_54 =10'b0;

   // m179_55 = W*in
   wire signed [9:0] m179_55;
   assign m179_55 =10'b0;

   // m179_56 = W*in
   wire signed [9:0] m179_56;
   assign m179_56 =10'b0;

   // m179_57 = W*in
   wire signed [9:0] m179_57;
   assign m179_57 =10'b0;

   // m179_58 = W*in
   wire signed [9:0] m179_58;
   assign m179_58 =10'b0;

   // m179_59 = W*in
   wire signed [9:0] m179_59;
   assign m179_59 =10'b0;

   // m179_60 = W*in
   wire signed [9:0] m179_60;
   assign m179_60 =10'b0;

   // m179_61 = W*in
   wire signed [9:0] m179_61;
   assign m179_61 =10'b0;

   // m179_62 = W*in
   wire signed [9:0] m179_62;
   assign m179_62 =10'b0;

   // m179_63 = W*in
   wire signed [9:0] m179_63;
   assign m179_63 =10'b0;

   // m179_64 = W*in
   wire signed [9:0] m179_64;
   assign m179_64 =10'b0;

   // m179_65 = W*in
   wire signed [9:0] m179_65;
   assign m179_65 =10'b0;

   // m179_66 = W*in
   wire signed [9:0] m179_66;
   assign m179_66 =10'b0;

   // m179_67 = W*in
   wire signed [9:0] m179_67;
   assign m179_67 =10'b0;

   // m179_68 = W*in
   wire signed [9:0] m179_68;
   assign m179_68 =10'b0;

   // m179_69 = W*in
   wire signed [9:0] m179_69;
   assign m179_69 =10'b0;

   // m179_70 = W*in
   wire signed [9:0] m179_70;
   assign m179_70 =10'b0;

   // m179_71 = W*in
   wire signed [9:0] m179_71;
   assign m179_71 =10'b0;

   // m179_72 = W*in
   wire signed [9:0] m179_72;
   assign m179_72 =10'b0;

   // m179_73 = W*in
   wire signed [9:0] m179_73;
   assign m179_73 =10'b0;

   // m179_74 = W*in
   wire signed [9:0] m179_74;
   assign m179_74 =10'b0;

   // m179_75 = W*in
   wire signed [9:0] m179_75;
   assign m179_75 =10'b0;

   // m179_76 = W*in
   wire signed [9:0] m179_76;
   assign m179_76 =10'b0;

   // m179_77 = W*in
   wire signed [9:0] m179_77;
   assign m179_77 =10'b0;

   // m179_78 = W*in
   wire signed [9:0] m179_78;
   assign m179_78 =10'b0;

   // m179_79 = W*in
   wire signed [9:0] m179_79;
   assign m179_79 =10'b0;

   // m179_80 = W*in
   wire signed [9:0] m179_80;
   assign m179_80 =10'b0;

   // m179_81 = W*in
   wire signed [9:0] m179_81;
   assign m179_81 =10'b0;

   // m179_82 = W*in
   wire signed [9:0] m179_82;
   assign m179_82 =10'b0;

   // m179_83 = W*in
   wire signed [9:0] m179_83;
   assign m179_83 =10'b0;

   // m179_84 = W*in
   wire signed [9:0] m179_84;
   assign m179_84 =10'b0;

   // m179_85 = W*in
   wire signed [9:0] m179_85;
   assign m179_85 =10'b0;

   // m179_86 = W*in
   wire signed [9:0] m179_86;
   assign m179_86 =10'b0;

   // m179_87 = W*in
   wire signed [9:0] m179_87;
   assign m179_87 =10'b0;

   // m179_88 = W*in
   wire signed [9:0] m179_88;
   assign m179_88 =10'b0;

   // m179_89 = W*in
   wire signed [9:0] m179_89;
   assign m179_89 =10'b0;

   // m179_90 = W*in
   wire signed [9:0] m179_90;
   assign m179_90 =10'b0;

   // m179_91 = W*in
   wire signed [9:0] m179_91;
   assign m179_91 =10'b0;

   // m179_92 = W*in
   wire signed [9:0] m179_92;
   assign m179_92 =10'b0;

   // m179_93 = W*in
   wire signed [9:0] m179_93;
   assign m179_93 =10'b0;

   // m179_94 = W*in
   wire signed [9:0] m179_94;
   assign m179_94 =10'b0;

   // m179_95 = W*in
   wire signed [9:0] m179_95;
   assign m179_95 =10'b0;

   // m179_96 = W*in
   wire signed [9:0] m179_96;
   assign m179_96 =10'b0;

   // m179_97 = W*in
   wire signed [9:0] m179_97;
   assign m179_97 =10'b0;

   // m179_98 = W*in
   wire signed [9:0] m179_98;
   assign m179_98 =10'b0;

   // m179_99 = W*in
   wire signed [9:0] m179_99;
   assign m179_99 =10'b0;

   // m179_100 = W*in
   wire signed [9:0] m179_100;
   assign m179_100 =10'b0;

   // m179_101 = W*in
   wire signed [9:0] m179_101;
   assign m179_101 =10'b0;

   // m179_102 = W*in
   wire signed [9:0] m179_102;
   assign m179_102 =10'b0;

   // m179_103 = W*in
   wire signed [9:0] m179_103;
   assign m179_103 =10'b0;

   // m179_104 = W*in
   wire signed [9:0] m179_104;
   assign m179_104 =10'b0;

   // m179_105 = W*in
   wire signed [9:0] m179_105;
   assign m179_105 =10'b0;

   // m179_106 = W*in
   wire signed [9:0] m179_106;
   assign m179_106 =10'b0;

   // m179_107 = W*in
   wire signed [9:0] m179_107;
   assign m179_107 =10'b0;

   // m179_108 = W*in
   wire signed [9:0] m179_108;
   assign m179_108 =10'b0;

   // m179_109 = W*in
   wire signed [9:0] m179_109;
   assign m179_109 ={ {5{in179[5]}} , in179[5:1] };

   // m179_110 = W*in
   wire signed [9:0] m179_110;
   assign m179_110 =10'b0;

   // m179_111 = W*in
   wire signed [9:0] m179_111;
   assign m179_111 =10'b0;

   // m179_112 = W*in
   wire signed [9:0] m179_112;
   assign m179_112 =10'b0;

   // m179_113 = W*in
   wire signed [9:0] m179_113;
   assign m179_113 =10'b0;

   // m179_114 = W*in
   wire signed [9:0] m179_114;
   assign m179_114 =10'b0;

   // m179_115 = W*in
   wire signed [9:0] m179_115;
   assign m179_115 =10'b0;

   // m179_116 = W*in
   wire signed [9:0] m179_116;
   assign m179_116 =10'b0;

   // m179_117 = W*in
   wire signed [9:0] m179_117;
   assign m179_117 =10'b0;

   // m180_1 = W*in
   wire signed [9:0] m180_1;
   assign m180_1 =10'b0;

   // m180_2 = W*in
   wire signed [9:0] m180_2;
   assign m180_2 =10'b0;

   // m180_3 = W*in
   wire signed [9:0] m180_3;
   assign m180_3 =10'b0;

   // m180_4 = W*in
   wire signed [9:0] m180_4;
   assign m180_4 =10'b0;

   // m180_5 = W*in
   wire signed [9:0] m180_5;
   assign m180_5 =10'b0;

   // m180_6 = W*in
   wire signed [9:0] m180_6;
   assign m180_6 =10'b0;

   // m180_7 = W*in
   wire signed [9:0] m180_7;
   assign m180_7 =10'b0;

   // m180_8 = W*in
   wire signed [9:0] m180_8;
   assign m180_8 =10'b0;

   // m180_9 = W*in
   wire signed [9:0] m180_9;
   assign m180_9 =10'b0;

   // m180_10 = W*in
   wire signed [9:0] m180_10;
   assign m180_10 =10'b0;

   // m180_11 = W*in
   wire signed [9:0] m180_11;
   assign m180_11 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_12 = W*in
   wire signed [9:0] m180_12;
   assign m180_12 =10'b0;

   // m180_13 = W*in
   wire signed [9:0] m180_13;
   assign m180_13 =10'b0;

   // m180_14 = W*in
   wire signed [9:0] m180_14;
   assign m180_14 =10'b0;

   // m180_15 = W*in
   wire signed [9:0] m180_15;
   assign m180_15 =10'b0;

   // m180_16 = W*in
   wire signed [9:0] m180_16;
   assign m180_16 =10'b0;

   // m180_17 = W*in
   wire signed [9:0] m180_17;
   assign m180_17 =10'b0;

   // m180_18 = W*in
   wire signed [9:0] m180_18;
   assign m180_18 =10'b0;

   // m180_19 = W*in
   wire signed [9:0] m180_19;
   assign m180_19 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_20 = W*in
   wire signed [9:0] m180_20;
   assign m180_20 ={ {5{in180[5]}} , in180[5:1] };

   // m180_21 = W*in
   wire signed [9:0] m180_21;
   assign m180_21 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_22 = W*in
   wire signed [9:0] m180_22;
   assign m180_22 =10'b0;

   // m180_23 = W*in
   wire signed [9:0] m180_23;
   assign m180_23 ={ {4{in180[5]}} , in180[5:0] };

   // m180_24 = W*in
   wire signed [9:0] m180_24;
   assign m180_24 =10'b0;

   // m180_25 = W*in
   wire signed [9:0] m180_25;
   assign m180_25 ={ {4{in180[5]}} , in180[5:0] };

   // m180_26 = W*in
   wire signed [9:0] m180_26;
   assign m180_26 ={ {5{in180[5]}} , in180[5:1] };

   // m180_27 = W*in
   wire signed [9:0] m180_27;
   assign m180_27 ={ {4{in180[5]}} , in180[5:0] };

   // m180_28 = W*in
   wire signed [9:0] m180_28;
   assign m180_28 ={ {4{in180[5]}} , in180[5:0] };

   // m180_29 = W*in
   wire signed [9:0] m180_29;
   assign m180_29 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_30 = W*in
   wire signed [9:0] m180_30;
   assign m180_30 =10'b0;

   // m180_31 = W*in
   wire signed [9:0] m180_31;
   assign m180_31 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_32 = W*in
   wire signed [9:0] m180_32;
   assign m180_32 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_33 = W*in
   wire signed [9:0] m180_33;
   assign m180_33 =10'b0;

   // m180_34 = W*in
   wire signed [9:0] m180_34;
   assign m180_34 =10'b0;

   // m180_35 = W*in
   wire signed [9:0] m180_35;
   assign m180_35 =10'b0;

   // m180_36 = W*in
   wire signed [9:0] m180_36;
   assign m180_36 ={ {5{in180[5]}} , in180[5:1] };

   // m180_37 = W*in
   wire signed [9:0] m180_37;
   assign m180_37 =10'b0;

   // m180_38 = W*in
   wire signed [9:0] m180_38;
   assign m180_38 ={ {5{in180[5]}} , in180[5:1] };

   // m180_39 = W*in
   wire signed [9:0] m180_39;
   assign m180_39 =10'b0;

   // m180_40 = W*in
   wire signed [9:0] m180_40;
   assign m180_40 =10'b0;

   // m180_41 = W*in
   wire signed [9:0] m180_41;
   assign m180_41 =10'b0;

   // m180_42 = W*in
   wire signed [9:0] m180_42;
   assign m180_42 =10'b0;

   // m180_43 = W*in
   wire signed [9:0] m180_43;
   assign m180_43 =10'b0;

   // m180_44 = W*in
   wire signed [9:0] m180_44;
   assign m180_44 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_45 = W*in
   wire signed [9:0] m180_45;
   assign m180_45 =10'b0;

   // m180_46 = W*in
   wire signed [9:0] m180_46;
   assign m180_46 =10'b0;

   // m180_47 = W*in
   wire signed [9:0] m180_47;
   assign m180_47 ={ {4{in180[5]}} , in180[5:0] };

   // m180_48 = W*in
   wire signed [9:0] m180_48;
   assign m180_48 =10'b0;

   // m180_49 = W*in
   wire signed [9:0] m180_49;
   assign m180_49 =10'b0;

   // m180_50 = W*in
   wire signed [9:0] m180_50;
   assign m180_50 =10'b0;

   // m180_51 = W*in
   wire signed [9:0] m180_51;
   assign m180_51 =10'b0;

   // m180_52 = W*in
   wire signed [9:0] m180_52;
   assign m180_52 =10'b0;

   // m180_53 = W*in
   wire signed [9:0] m180_53;
   assign m180_53 =10'b0;

   // m180_54 = W*in
   wire signed [9:0] m180_54;
   assign m180_54 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_55 = W*in
   wire signed [9:0] m180_55;
   assign m180_55 =10'b0;

   // m180_56 = W*in
   wire signed [9:0] m180_56;
   assign m180_56 =10'b0;

   // m180_57 = W*in
   wire signed [9:0] m180_57;
   assign m180_57 =10'b0;

   // m180_58 = W*in
   wire signed [9:0] m180_58;
   assign m180_58 =10'b0;

   // m180_59 = W*in
   wire signed [9:0] m180_59;
   assign m180_59 ={ {4{in180[5]}} , in180[5:0] };

   // m180_60 = W*in
   wire signed [9:0] m180_60;
   assign m180_60 ={ {4{in180[5]}} , in180[5:0] };

   // m180_61 = W*in
   wire signed [9:0] m180_61;
   assign m180_61 =10'b0;

   // m180_62 = W*in
   wire signed [9:0] m180_62;
   assign m180_62 =10'b0;

   // m180_63 = W*in
   wire signed [9:0] m180_63;
   assign m180_63 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_64 = W*in
   wire signed [9:0] m180_64;
   assign m180_64 =10'b0;

   // m180_65 = W*in
   wire signed [9:0] m180_65;
   assign m180_65 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_66 = W*in
   wire signed [9:0] m180_66;
   assign m180_66 =10'b0;

   // m180_67 = W*in
   wire signed [9:0] m180_67;
   assign m180_67 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_68 = W*in
   wire signed [9:0] m180_68;
   assign m180_68 =10'b0;

   // m180_69 = W*in
   wire signed [9:0] m180_69;
   assign m180_69 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_70 = W*in
   wire signed [9:0] m180_70;
   assign m180_70 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_71 = W*in
   wire signed [9:0] m180_71;
   assign m180_71 ={ {5{in180[5]}} , in180[5:1] };

   // m180_72 = W*in
   wire signed [9:0] m180_72;
   assign m180_72 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_73 = W*in
   wire signed [9:0] m180_73;
   assign m180_73 =10'b0;

   // m180_74 = W*in
   wire signed [9:0] m180_74;
   assign m180_74 =10'b0;

   // m180_75 = W*in
   wire signed [9:0] m180_75;
   assign m180_75 =10'b0;

   // m180_76 = W*in
   wire signed [9:0] m180_76;
   assign m180_76 =10'b0;

   // m180_77 = W*in
   wire signed [9:0] m180_77;
   assign m180_77 ={ {4{in180[5]}} , in180[5:0] };

   // m180_78 = W*in
   wire signed [9:0] m180_78;
   assign m180_78 =10'b0;

   // m180_79 = W*in
   wire signed [9:0] m180_79;
   assign m180_79 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_80 = W*in
   wire signed [9:0] m180_80;
   assign m180_80 =10'b0;

   // m180_81 = W*in
   wire signed [9:0] m180_81;
   assign m180_81 ={ {4{in180[5]}} , in180[5:0] };

   // m180_82 = W*in
   wire signed [9:0] m180_82;
   assign m180_82 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_83 = W*in
   wire signed [9:0] m180_83;
   assign m180_83 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_84 = W*in
   wire signed [9:0] m180_84;
   assign m180_84 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_85 = W*in
   wire signed [9:0] m180_85;
   assign m180_85 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_86 = W*in
   wire signed [9:0] m180_86;
   assign m180_86 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_87 = W*in
   wire signed [9:0] m180_87;
   assign m180_87 ={ {4{in180[5]}} , in180[5:0] };

   // m180_88 = W*in
   wire signed [9:0] m180_88;
   assign m180_88 =10'b0;

   // m180_89 = W*in
   wire signed [9:0] m180_89;
   assign m180_89 =10'b0;

   // m180_90 = W*in
   wire signed [9:0] m180_90;
   assign m180_90 =10'b0;

   // m180_91 = W*in
   wire signed [9:0] m180_91;
   assign m180_91 =10'b0;

   // m180_92 = W*in
   wire signed [9:0] m180_92;
   assign m180_92 =10'b0;

   // m180_93 = W*in
   wire signed [9:0] m180_93;
   assign m180_93 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_94 = W*in
   wire signed [9:0] m180_94;
   assign m180_94 =10'b0;

   // m180_95 = W*in
   wire signed [9:0] m180_95;
   assign m180_95 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_96 = W*in
   wire signed [9:0] m180_96;
   assign m180_96 =10'b0;

   // m180_97 = W*in
   wire signed [9:0] m180_97;
   assign m180_97 ={ {4{in180[5]}} , in180[5:0] };

   // m180_98 = W*in
   wire signed [9:0] m180_98;
   assign m180_98 =10'b0;

   // m180_99 = W*in
   wire signed [9:0] m180_99;
   assign m180_99 ={ {4{in180[5]}} , in180[5:0] };

   // m180_100 = W*in
   wire signed [9:0] m180_100;
   assign m180_100 =10'b0;

   // m180_101 = W*in
   wire signed [9:0] m180_101;
   assign m180_101 =10'b0;

   // m180_102 = W*in
   wire signed [9:0] m180_102;
   assign m180_102 =10'b0;

   // m180_103 = W*in
   wire signed [9:0] m180_103;
   assign m180_103 =10'b0;

   // m180_104 = W*in
   wire signed [9:0] m180_104;
   assign m180_104 =10'b0;

   // m180_105 = W*in
   wire signed [9:0] m180_105;
   assign m180_105 =10'b0;

   // m180_106 = W*in
   wire signed [9:0] m180_106;
   assign m180_106 =10'b0;

   // m180_107 = W*in
   wire signed [9:0] m180_107;
   assign m180_107 =10'b0;

   // m180_108 = W*in
   wire signed [9:0] m180_108;
   assign m180_108 ={ {5{neg180[5]}} , neg180[5:1] };

   // m180_109 = W*in
   wire signed [9:0] m180_109;
   assign m180_109 =10'b0;

   // m180_110 = W*in
   wire signed [9:0] m180_110;
   assign m180_110 ={ {4{in180[5]}} , in180[5:0] };

   // m180_111 = W*in
   wire signed [9:0] m180_111;
   assign m180_111 =10'b0;

   // m180_112 = W*in
   wire signed [9:0] m180_112;
   assign m180_112 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_113 = W*in
   wire signed [9:0] m180_113;
   assign m180_113 =10'b0;

   // m180_114 = W*in
   wire signed [9:0] m180_114;
   assign m180_114 ={ {4{in180[5]}} , in180[5:0] };

   // m180_115 = W*in
   wire signed [9:0] m180_115;
   assign m180_115 =10'b0;

   // m180_116 = W*in
   wire signed [9:0] m180_116;
   assign m180_116 ={ {4{neg180[5]}} , neg180[5:0] };

   // m180_117 = W*in
   wire signed [9:0] m180_117;
   assign m180_117 ={ {5{in180[5]}} , in180[5:1] };

   // m181_1 = W*in
   wire signed [9:0] m181_1;
   assign m181_1 =10'b0;

   // m181_2 = W*in
   wire signed [9:0] m181_2;
   assign m181_2 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_3 = W*in
   wire signed [9:0] m181_3;
   assign m181_3 =10'b0;

   // m181_4 = W*in
   wire signed [9:0] m181_4;
   assign m181_4 =10'b0;

   // m181_5 = W*in
   wire signed [9:0] m181_5;
   assign m181_5 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_6 = W*in
   wire signed [9:0] m181_6;
   assign m181_6 =10'b0;

   // m181_7 = W*in
   wire signed [9:0] m181_7;
   assign m181_7 =10'b0;

   // m181_8 = W*in
   wire signed [9:0] m181_8;
   assign m181_8 =10'b0;

   // m181_9 = W*in
   wire signed [9:0] m181_9;
   assign m181_9 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_10 = W*in
   wire signed [9:0] m181_10;
   assign m181_10 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_11 = W*in
   wire signed [9:0] m181_11;
   assign m181_11 =10'b0;

   // m181_12 = W*in
   wire signed [9:0] m181_12;
   assign m181_12 ={ {4{in181[5]}} , in181[5:0] };

   // m181_13 = W*in
   wire signed [9:0] m181_13;
   assign m181_13 =10'b0;

   // m181_14 = W*in
   wire signed [9:0] m181_14;
   assign m181_14 =10'b0;

   // m181_15 = W*in
   wire signed [9:0] m181_15;
   assign m181_15 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_16 = W*in
   wire signed [9:0] m181_16;
   assign m181_16 =10'b0;

   // m181_17 = W*in
   wire signed [9:0] m181_17;
   assign m181_17 ={ {4{in181[5]}} , in181[5:0] };

   // m181_18 = W*in
   wire signed [9:0] m181_18;
   assign m181_18 =10'b0;

   // m181_19 = W*in
   wire signed [9:0] m181_19;
   assign m181_19 =10'b0;

   // m181_20 = W*in
   wire signed [9:0] m181_20;
   assign m181_20 =10'b0;

   // m181_21 = W*in
   wire signed [9:0] m181_21;
   assign m181_21 =10'b0;

   // m181_22 = W*in
   wire signed [9:0] m181_22;
   assign m181_22 ={ {5{in181[5]}} , in181[5:1] };

   // m181_23 = W*in
   wire signed [9:0] m181_23;
   assign m181_23 ={ {5{in181[5]}} , in181[5:1] };

   // m181_24 = W*in
   wire signed [9:0] m181_24;
   assign m181_24 ={ {5{in181[5]}} , in181[5:1] };

   // m181_25 = W*in
   wire signed [9:0] m181_25;
   assign m181_25 =10'b0;

   // m181_26 = W*in
   wire signed [9:0] m181_26;
   assign m181_26 ={ {4{in181[5]}} , in181[5:0] };

   // m181_27 = W*in
   wire signed [9:0] m181_27;
   assign m181_27 ={ {4{in181[5]}} , in181[5:0] };

   // m181_28 = W*in
   wire signed [9:0] m181_28;
   assign m181_28 ={ {4{in181[5]}} , in181[5:0] };

   // m181_29 = W*in
   wire signed [9:0] m181_29;
   assign m181_29 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_30 = W*in
   wire signed [9:0] m181_30;
   assign m181_30 =10'b0;

   // m181_31 = W*in
   wire signed [9:0] m181_31;
   assign m181_31 =10'b0;

   // m181_32 = W*in
   wire signed [9:0] m181_32;
   assign m181_32 ={ {3{neg181[5]}} , neg181 , {1{1'b0}} };

   // m181_33 = W*in
   wire signed [9:0] m181_33;
   assign m181_33 =10'b0;

   // m181_34 = W*in
   wire signed [9:0] m181_34;
   assign m181_34 ={ {4{in181[5]}} , in181[5:0] };

   // m181_35 = W*in
   wire signed [9:0] m181_35;
   assign m181_35 =10'b0;

   // m181_36 = W*in
   wire signed [9:0] m181_36;
   assign m181_36 =10'b0;

   // m181_37 = W*in
   wire signed [9:0] m181_37;
   assign m181_37 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_38 = W*in
   wire signed [9:0] m181_38;
   assign m181_38 ={ {3{in181[5]}} , in181 , {1{1'b0}} };

   // m181_39 = W*in
   wire signed [9:0] m181_39;
   assign m181_39 ={ {4{in181[5]}} , in181[5:0] };

   // m181_40 = W*in
   wire signed [9:0] m181_40;
   assign m181_40 =10'b0;

   // m181_41 = W*in
   wire signed [9:0] m181_41;
   assign m181_41 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_42 = W*in
   wire signed [9:0] m181_42;
   assign m181_42 ={ {3{in181[5]}} , in181 , {1{1'b0}} };

   // m181_43 = W*in
   wire signed [9:0] m181_43;
   assign m181_43 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_44 = W*in
   wire signed [9:0] m181_44;
   assign m181_44 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_45 = W*in
   wire signed [9:0] m181_45;
   assign m181_45 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_46 = W*in
   wire signed [9:0] m181_46;
   assign m181_46 ={ {4{in181[5]}} , in181[5:0] };

   // m181_47 = W*in
   wire signed [9:0] m181_47;
   assign m181_47 ={ {4{in181[5]}} , in181[5:0] };

   // m181_48 = W*in
   wire signed [9:0] m181_48;
   assign m181_48 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_49 = W*in
   wire signed [9:0] m181_49;
   assign m181_49 ={ {5{in181[5]}} , in181[5:1] };

   // m181_50 = W*in
   wire signed [9:0] m181_50;
   assign m181_50 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_51 = W*in
   wire signed [9:0] m181_51;
   assign m181_51 =10'b0;

   // m181_52 = W*in
   wire signed [9:0] m181_52;
   assign m181_52 =10'b0;

   // m181_53 = W*in
   wire signed [9:0] m181_53;
   assign m181_53 =10'b0;

   // m181_54 = W*in
   wire signed [9:0] m181_54;
   assign m181_54 =10'b0;

   // m181_55 = W*in
   wire signed [9:0] m181_55;
   assign m181_55 =10'b0;

   // m181_56 = W*in
   wire signed [9:0] m181_56;
   assign m181_56 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_57 = W*in
   wire signed [9:0] m181_57;
   assign m181_57 =10'b0;

   // m181_58 = W*in
   wire signed [9:0] m181_58;
   assign m181_58 ={ {5{neg181[5]}} , neg181[5:1] };

   // m181_59 = W*in
   wire signed [9:0] m181_59;
   assign m181_59 =10'b0;

   // m181_60 = W*in
   wire signed [9:0] m181_60;
   assign m181_60 ={ {4{in181[5]}} , in181[5:0] };

   // m181_61 = W*in
   wire signed [9:0] m181_61;
   assign m181_61 =10'b0;

   // m181_62 = W*in
   wire signed [9:0] m181_62;
   assign m181_62 =10'b0;

   // m181_63 = W*in
   wire signed [9:0] m181_63;
   assign m181_63 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_64 = W*in
   wire signed [9:0] m181_64;
   assign m181_64 ={ {3{in181[5]}} , in181 , {1{1'b0}} };

   // m181_65 = W*in
   wire signed [9:0] m181_65;
   assign m181_65 ={ {4{in181[5]}} , in181[5:0] };

   // m181_66 = W*in
   wire signed [9:0] m181_66;
   assign m181_66 ={ {4{in181[5]}} , in181[5:0] };

   // m181_67 = W*in
   wire signed [9:0] m181_67;
   assign m181_67 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_68 = W*in
   wire signed [9:0] m181_68;
   assign m181_68 =10'b0;

   // m181_69 = W*in
   wire signed [9:0] m181_69;
   assign m181_69 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_70 = W*in
   wire signed [9:0] m181_70;
   assign m181_70 =10'b0;

   // m181_71 = W*in
   wire signed [9:0] m181_71;
   assign m181_71 ={ {4{in181[5]}} , in181[5:0] };

   // m181_72 = W*in
   wire signed [9:0] m181_72;
   assign m181_72 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_73 = W*in
   wire signed [9:0] m181_73;
   assign m181_73 =10'b0;

   // m181_74 = W*in
   wire signed [9:0] m181_74;
   assign m181_74 ={ {4{in181[5]}} , in181[5:0] };

   // m181_75 = W*in
   wire signed [9:0] m181_75;
   assign m181_75 ={ {4{in181[5]}} , in181[5:0] };

   // m181_76 = W*in
   wire signed [9:0] m181_76;
   assign m181_76 =10'b0;

   // m181_77 = W*in
   wire signed [9:0] m181_77;
   assign m181_77 =10'b0;

   // m181_78 = W*in
   wire signed [9:0] m181_78;
   assign m181_78 =10'b0;

   // m181_79 = W*in
   wire signed [9:0] m181_79;
   assign m181_79 ={ {5{neg181[5]}} , neg181[5:1] };

   // m181_80 = W*in
   wire signed [9:0] m181_80;
   assign m181_80 =10'b0;

   // m181_81 = W*in
   wire signed [9:0] m181_81;
   assign m181_81 ={ {4{in181[5]}} , in181[5:0] };

   // m181_82 = W*in
   wire signed [9:0] m181_82;
   assign m181_82 =10'b0;

   // m181_83 = W*in
   wire signed [9:0] m181_83;
   assign m181_83 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_84 = W*in
   wire signed [9:0] m181_84;
   assign m181_84 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_85 = W*in
   wire signed [9:0] m181_85;
   assign m181_85 ={ {3{neg181[5]}} , neg181 , {1{1'b0}} };

   // m181_86 = W*in
   wire signed [9:0] m181_86;
   assign m181_86 ={ {4{in181[5]}} , in181[5:0] };

   // m181_87 = W*in
   wire signed [9:0] m181_87;
   assign m181_87 =10'b0;

   // m181_88 = W*in
   wire signed [9:0] m181_88;
   assign m181_88 =10'b0;

   // m181_89 = W*in
   wire signed [9:0] m181_89;
   assign m181_89 =10'b0;

   // m181_90 = W*in
   wire signed [9:0] m181_90;
   assign m181_90 =10'b0;

   // m181_91 = W*in
   wire signed [9:0] m181_91;
   assign m181_91 ={ {3{in181[5]}} , in181 , {1{1'b0}} };

   // m181_92 = W*in
   wire signed [9:0] m181_92;
   assign m181_92 =10'b0;

   // m181_93 = W*in
   wire signed [9:0] m181_93;
   assign m181_93 =10'b0;

   // m181_94 = W*in
   wire signed [9:0] m181_94;
   assign m181_94 ={ {4{in181[5]}} , in181[5:0] };

   // m181_95 = W*in
   wire signed [9:0] m181_95;
   assign m181_95 =10'b0;

   // m181_96 = W*in
   wire signed [9:0] m181_96;
   assign m181_96 =10'b0;

   // m181_97 = W*in
   wire signed [9:0] m181_97;
   assign m181_97 ={ {5{in181[5]}} , in181[5:1] };

   // m181_98 = W*in
   wire signed [9:0] m181_98;
   assign m181_98 =10'b0;

   // m181_99 = W*in
   wire signed [9:0] m181_99;
   assign m181_99 ={ {4{in181[5]}} , in181[5:0] };

   // m181_100 = W*in
   wire signed [9:0] m181_100;
   assign m181_100 ={ {4{in181[5]}} , in181[5:0] };

   // m181_101 = W*in
   wire signed [9:0] m181_101;
   assign m181_101 =10'b0;

   // m181_102 = W*in
   wire signed [9:0] m181_102;
   assign m181_102 =10'b0;

   // m181_103 = W*in
   wire signed [9:0] m181_103;
   assign m181_103 ={ {4{in181[5]}} , in181[5:0] };

   // m181_104 = W*in
   wire signed [9:0] m181_104;
   assign m181_104 ={ {4{in181[5]}} , in181[5:0] };

   // m181_105 = W*in
   wire signed [9:0] m181_105;
   assign m181_105 =10'b0;

   // m181_106 = W*in
   wire signed [9:0] m181_106;
   assign m181_106 =10'b0;

   // m181_107 = W*in
   wire signed [9:0] m181_107;
   assign m181_107 =10'b0;

   // m181_108 = W*in
   wire signed [9:0] m181_108;
   assign m181_108 =10'b0;

   // m181_109 = W*in
   wire signed [9:0] m181_109;
   assign m181_109 =10'b0;

   // m181_110 = W*in
   wire signed [9:0] m181_110;
   assign m181_110 ={ {4{in181[5]}} , in181[5:0] };

   // m181_111 = W*in
   wire signed [9:0] m181_111;
   assign m181_111 =10'b0;

   // m181_112 = W*in
   wire signed [9:0] m181_112;
   assign m181_112 ={ {4{in181[5]}} , in181[5:0] };

   // m181_113 = W*in
   wire signed [9:0] m181_113;
   assign m181_113 ={ {4{neg181[5]}} , neg181[5:0] };

   // m181_114 = W*in
   wire signed [9:0] m181_114;
   assign m181_114 =10'b0;

   // m181_115 = W*in
   wire signed [9:0] m181_115;
   assign m181_115 =10'b0;

   // m181_116 = W*in
   wire signed [9:0] m181_116;
   assign m181_116 =10'b0;

   // m181_117 = W*in
   wire signed [9:0] m181_117;
   assign m181_117 ={ {4{in181[5]}} , in181[5:0] };

   // m182_1 = W*in
   wire signed [9:0] m182_1;
   assign m182_1 =10'b0;

   // m182_2 = W*in
   wire signed [9:0] m182_2;
   assign m182_2 ={ {5{neg182[5]}} , neg182[5:1] };

   // m182_3 = W*in
   wire signed [9:0] m182_3;
   assign m182_3 =10'b0;

   // m182_4 = W*in
   wire signed [9:0] m182_4;
   assign m182_4 =10'b0;

   // m182_5 = W*in
   wire signed [9:0] m182_5;
   assign m182_5 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_6 = W*in
   wire signed [9:0] m182_6;
   assign m182_6 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_7 = W*in
   wire signed [9:0] m182_7;
   assign m182_7 =10'b0;

   // m182_8 = W*in
   wire signed [9:0] m182_8;
   assign m182_8 =10'b0;

   // m182_9 = W*in
   wire signed [9:0] m182_9;
   assign m182_9 =10'b0;

   // m182_10 = W*in
   wire signed [9:0] m182_10;
   assign m182_10 ={ {4{in182[5]}} , in182[5:0] };

   // m182_11 = W*in
   wire signed [9:0] m182_11;
   assign m182_11 =10'b0;

   // m182_12 = W*in
   wire signed [9:0] m182_12;
   assign m182_12 ={ {5{in182[5]}} , in182[5:1] };

   // m182_13 = W*in
   wire signed [9:0] m182_13;
   assign m182_13 =10'b0;

   // m182_14 = W*in
   wire signed [9:0] m182_14;
   assign m182_14 =10'b0;

   // m182_15 = W*in
   wire signed [9:0] m182_15;
   assign m182_15 =10'b0;

   // m182_16 = W*in
   wire signed [9:0] m182_16;
   assign m182_16 =10'b0;

   // m182_17 = W*in
   wire signed [9:0] m182_17;
   assign m182_17 =10'b0;

   // m182_18 = W*in
   wire signed [9:0] m182_18;
   assign m182_18 ={ {4{in182[5]}} , in182[5:0] };

   // m182_19 = W*in
   wire signed [9:0] m182_19;
   assign m182_19 =10'b0;

   // m182_20 = W*in
   wire signed [9:0] m182_20;
   assign m182_20 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_21 = W*in
   wire signed [9:0] m182_21;
   assign m182_21 ={ {5{neg182[5]}} , neg182[5:1] };

   // m182_22 = W*in
   wire signed [9:0] m182_22;
   assign m182_22 =10'b0;

   // m182_23 = W*in
   wire signed [9:0] m182_23;
   assign m182_23 ={ {5{neg182[5]}} , neg182[5:1] };

   // m182_24 = W*in
   wire signed [9:0] m182_24;
   assign m182_24 =10'b0;

   // m182_25 = W*in
   wire signed [9:0] m182_25;
   assign m182_25 =10'b0;

   // m182_26 = W*in
   wire signed [9:0] m182_26;
   assign m182_26 ={ {4{in182[5]}} , in182[5:0] };

   // m182_27 = W*in
   wire signed [9:0] m182_27;
   assign m182_27 =10'b0;

   // m182_28 = W*in
   wire signed [9:0] m182_28;
   assign m182_28 =10'b0;

   // m182_29 = W*in
   wire signed [9:0] m182_29;
   assign m182_29 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_30 = W*in
   wire signed [9:0] m182_30;
   assign m182_30 =10'b0;

   // m182_31 = W*in
   wire signed [9:0] m182_31;
   assign m182_31 =10'b0;

   // m182_32 = W*in
   wire signed [9:0] m182_32;
   assign m182_32 =10'b0;

   // m182_33 = W*in
   wire signed [9:0] m182_33;
   assign m182_33 =10'b0;

   // m182_34 = W*in
   wire signed [9:0] m182_34;
   assign m182_34 ={ {3{neg182[5]}} , neg182 , {1{1'b0}} };

   // m182_35 = W*in
   wire signed [9:0] m182_35;
   assign m182_35 ={ {5{neg182[5]}} , neg182[5:1] };

   // m182_36 = W*in
   wire signed [9:0] m182_36;
   assign m182_36 ={ {5{in182[5]}} , in182[5:1] };

   // m182_37 = W*in
   wire signed [9:0] m182_37;
   assign m182_37 =10'b0;

   // m182_38 = W*in
   wire signed [9:0] m182_38;
   assign m182_38 =10'b0;

   // m182_39 = W*in
   wire signed [9:0] m182_39;
   assign m182_39 =10'b0;

   // m182_40 = W*in
   wire signed [9:0] m182_40;
   assign m182_40 =10'b0;

   // m182_41 = W*in
   wire signed [9:0] m182_41;
   assign m182_41 =10'b0;

   // m182_42 = W*in
   wire signed [9:0] m182_42;
   assign m182_42 ={ {4{in182[5]}} , in182[5:0] };

   // m182_43 = W*in
   wire signed [9:0] m182_43;
   assign m182_43 =10'b0;

   // m182_44 = W*in
   wire signed [9:0] m182_44;
   assign m182_44 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_45 = W*in
   wire signed [9:0] m182_45;
   assign m182_45 =10'b0;

   // m182_46 = W*in
   wire signed [9:0] m182_46;
   assign m182_46 =10'b0;

   // m182_47 = W*in
   wire signed [9:0] m182_47;
   assign m182_47 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_48 = W*in
   wire signed [9:0] m182_48;
   assign m182_48 =10'b0;

   // m182_49 = W*in
   wire signed [9:0] m182_49;
   assign m182_49 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_50 = W*in
   wire signed [9:0] m182_50;
   assign m182_50 =10'b0;

   // m182_51 = W*in
   wire signed [9:0] m182_51;
   assign m182_51 =10'b0;

   // m182_52 = W*in
   wire signed [9:0] m182_52;
   assign m182_52 ={ {5{in182[5]}} , in182[5:1] };

   // m182_53 = W*in
   wire signed [9:0] m182_53;
   assign m182_53 =10'b0;

   // m182_54 = W*in
   wire signed [9:0] m182_54;
   assign m182_54 =10'b0;

   // m182_55 = W*in
   wire signed [9:0] m182_55;
   assign m182_55 ={ {4{in182[5]}} , in182[5:0] };

   // m182_56 = W*in
   wire signed [9:0] m182_56;
   assign m182_56 =10'b0;

   // m182_57 = W*in
   wire signed [9:0] m182_57;
   assign m182_57 =10'b0;

   // m182_58 = W*in
   wire signed [9:0] m182_58;
   assign m182_58 =10'b0;

   // m182_59 = W*in
   wire signed [9:0] m182_59;
   assign m182_59 ={ {5{in182[5]}} , in182[5:1] };

   // m182_60 = W*in
   wire signed [9:0] m182_60;
   assign m182_60 =10'b0;

   // m182_61 = W*in
   wire signed [9:0] m182_61;
   assign m182_61 =10'b0;

   // m182_62 = W*in
   wire signed [9:0] m182_62;
   assign m182_62 =10'b0;

   // m182_63 = W*in
   wire signed [9:0] m182_63;
   assign m182_63 =10'b0;

   // m182_64 = W*in
   wire signed [9:0] m182_64;
   assign m182_64 =10'b0;

   // m182_65 = W*in
   wire signed [9:0] m182_65;
   assign m182_65 ={ {4{in182[5]}} , in182[5:0] };

   // m182_66 = W*in
   wire signed [9:0] m182_66;
   assign m182_66 =10'b0;

   // m182_67 = W*in
   wire signed [9:0] m182_67;
   assign m182_67 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_68 = W*in
   wire signed [9:0] m182_68;
   assign m182_68 =10'b0;

   // m182_69 = W*in
   wire signed [9:0] m182_69;
   assign m182_69 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_70 = W*in
   wire signed [9:0] m182_70;
   assign m182_70 =10'b0;

   // m182_71 = W*in
   wire signed [9:0] m182_71;
   assign m182_71 =10'b0;

   // m182_72 = W*in
   wire signed [9:0] m182_72;
   assign m182_72 =10'b0;

   // m182_73 = W*in
   wire signed [9:0] m182_73;
   assign m182_73 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_74 = W*in
   wire signed [9:0] m182_74;
   assign m182_74 =10'b0;

   // m182_75 = W*in
   wire signed [9:0] m182_75;
   assign m182_75 =10'b0;

   // m182_76 = W*in
   wire signed [9:0] m182_76;
   assign m182_76 =10'b0;

   // m182_77 = W*in
   wire signed [9:0] m182_77;
   assign m182_77 =10'b0;

   // m182_78 = W*in
   wire signed [9:0] m182_78;
   assign m182_78 =10'b0;

   // m182_79 = W*in
   wire signed [9:0] m182_79;
   assign m182_79 =10'b0;

   // m182_80 = W*in
   wire signed [9:0] m182_80;
   assign m182_80 =10'b0;

   // m182_81 = W*in
   wire signed [9:0] m182_81;
   assign m182_81 =10'b0;

   // m182_82 = W*in
   wire signed [9:0] m182_82;
   assign m182_82 =10'b0;

   // m182_83 = W*in
   wire signed [9:0] m182_83;
   assign m182_83 =10'b0;

   // m182_84 = W*in
   wire signed [9:0] m182_84;
   assign m182_84 =10'b0;

   // m182_85 = W*in
   wire signed [9:0] m182_85;
   assign m182_85 =10'b0;

   // m182_86 = W*in
   wire signed [9:0] m182_86;
   assign m182_86 ={ {4{in182[5]}} , in182[5:0] };

   // m182_87 = W*in
   wire signed [9:0] m182_87;
   assign m182_87 =10'b0;

   // m182_88 = W*in
   wire signed [9:0] m182_88;
   assign m182_88 =10'b0;

   // m182_89 = W*in
   wire signed [9:0] m182_89;
   assign m182_89 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_90 = W*in
   wire signed [9:0] m182_90;
   assign m182_90 =10'b0;

   // m182_91 = W*in
   wire signed [9:0] m182_91;
   assign m182_91 ={ {4{in182[5]}} , in182[5:0] };

   // m182_92 = W*in
   wire signed [9:0] m182_92;
   assign m182_92 =10'b0;

   // m182_93 = W*in
   wire signed [9:0] m182_93;
   assign m182_93 ={ {4{neg182[5]}} , neg182[5:0] };

   // m182_94 = W*in
   wire signed [9:0] m182_94;
   assign m182_94 ={ {4{in182[5]}} , in182[5:0] };

   // m182_95 = W*in
   wire signed [9:0] m182_95;
   assign m182_95 =10'b0;

   // m182_96 = W*in
   wire signed [9:0] m182_96;
   assign m182_96 =10'b0;

   // m182_97 = W*in
   wire signed [9:0] m182_97;
   assign m182_97 =10'b0;

   // m182_98 = W*in
   wire signed [9:0] m182_98;
   assign m182_98 =10'b0;

   // m182_99 = W*in
   wire signed [9:0] m182_99;
   assign m182_99 =10'b0;

   // m182_100 = W*in
   wire signed [9:0] m182_100;
   assign m182_100 =10'b0;

   // m182_101 = W*in
   wire signed [9:0] m182_101;
   assign m182_101 =10'b0;

   // m182_102 = W*in
   wire signed [9:0] m182_102;
   assign m182_102 =10'b0;

   // m182_103 = W*in
   wire signed [9:0] m182_103;
   assign m182_103 =10'b0;

   // m182_104 = W*in
   wire signed [9:0] m182_104;
   assign m182_104 =10'b0;

   // m182_105 = W*in
   wire signed [9:0] m182_105;
   assign m182_105 =10'b0;

   // m182_106 = W*in
   wire signed [9:0] m182_106;
   assign m182_106 =10'b0;

   // m182_107 = W*in
   wire signed [9:0] m182_107;
   assign m182_107 ={ {5{in182[5]}} , in182[5:1] };

   // m182_108 = W*in
   wire signed [9:0] m182_108;
   assign m182_108 =10'b0;

   // m182_109 = W*in
   wire signed [9:0] m182_109;
   assign m182_109 =10'b0;

   // m182_110 = W*in
   wire signed [9:0] m182_110;
   assign m182_110 =10'b0;

   // m182_111 = W*in
   wire signed [9:0] m182_111;
   assign m182_111 =10'b0;

   // m182_112 = W*in
   wire signed [9:0] m182_112;
   assign m182_112 ={ {4{in182[5]}} , in182[5:0] };

   // m182_113 = W*in
   wire signed [9:0] m182_113;
   assign m182_113 =10'b0;

   // m182_114 = W*in
   wire signed [9:0] m182_114;
   assign m182_114 ={ {5{neg182[5]}} , neg182[5:1] };

   // m182_115 = W*in
   wire signed [9:0] m182_115;
   assign m182_115 ={ {5{neg182[5]}} , neg182[5:1] };

   // m182_116 = W*in
   wire signed [9:0] m182_116;
   assign m182_116 =10'b0;

   // m182_117 = W*in
   wire signed [9:0] m182_117;
   assign m182_117 =10'b0;

   // m183_1 = W*in
   wire signed [9:0] m183_1;
   assign m183_1 =10'b0;

   // m183_2 = W*in
   wire signed [9:0] m183_2;
   assign m183_2 =10'b0;

   // m183_3 = W*in
   wire signed [9:0] m183_3;
   assign m183_3 =10'b0;

   // m183_4 = W*in
   wire signed [9:0] m183_4;
   assign m183_4 =10'b0;

   // m183_5 = W*in
   wire signed [9:0] m183_5;
   assign m183_5 ={ {4{in183[5]}} , in183[5:0] };

   // m183_6 = W*in
   wire signed [9:0] m183_6;
   assign m183_6 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_7 = W*in
   wire signed [9:0] m183_7;
   assign m183_7 ={ {4{in183[5]}} , in183[5:0] };

   // m183_8 = W*in
   wire signed [9:0] m183_8;
   assign m183_8 =10'b0;

   // m183_9 = W*in
   wire signed [9:0] m183_9;
   assign m183_9 =10'b0;

   // m183_10 = W*in
   wire signed [9:0] m183_10;
   assign m183_10 =10'b0;

   // m183_11 = W*in
   wire signed [9:0] m183_11;
   assign m183_11 =10'b0;

   // m183_12 = W*in
   wire signed [9:0] m183_12;
   assign m183_12 =10'b0;

   // m183_13 = W*in
   wire signed [9:0] m183_13;
   assign m183_13 ={ {4{in183[5]}} , in183[5:0] };

   // m183_14 = W*in
   wire signed [9:0] m183_14;
   assign m183_14 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_15 = W*in
   wire signed [9:0] m183_15;
   assign m183_15 =10'b0;

   // m183_16 = W*in
   wire signed [9:0] m183_16;
   assign m183_16 ={ {5{neg183[5]}} , neg183[5:1] };

   // m183_17 = W*in
   wire signed [9:0] m183_17;
   assign m183_17 =10'b0;

   // m183_18 = W*in
   wire signed [9:0] m183_18;
   assign m183_18 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_19 = W*in
   wire signed [9:0] m183_19;
   assign m183_19 =10'b0;

   // m183_20 = W*in
   wire signed [9:0] m183_20;
   assign m183_20 =10'b0;

   // m183_21 = W*in
   wire signed [9:0] m183_21;
   assign m183_21 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_22 = W*in
   wire signed [9:0] m183_22;
   assign m183_22 ={ {4{in183[5]}} , in183[5:0] };

   // m183_23 = W*in
   wire signed [9:0] m183_23;
   assign m183_23 =10'b0;

   // m183_24 = W*in
   wire signed [9:0] m183_24;
   assign m183_24 ={ {4{in183[5]}} , in183[5:0] };

   // m183_25 = W*in
   wire signed [9:0] m183_25;
   assign m183_25 ={ {4{in183[5]}} , in183[5:0] };

   // m183_26 = W*in
   wire signed [9:0] m183_26;
   assign m183_26 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_27 = W*in
   wire signed [9:0] m183_27;
   assign m183_27 ={ {4{in183[5]}} , in183[5:0] };

   // m183_28 = W*in
   wire signed [9:0] m183_28;
   assign m183_28 ={ {4{in183[5]}} , in183[5:0] };

   // m183_29 = W*in
   wire signed [9:0] m183_29;
   assign m183_29 =10'b0;

   // m183_30 = W*in
   wire signed [9:0] m183_30;
   assign m183_30 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_31 = W*in
   wire signed [9:0] m183_31;
   assign m183_31 =10'b0;

   // m183_32 = W*in
   wire signed [9:0] m183_32;
   assign m183_32 =10'b0;

   // m183_33 = W*in
   wire signed [9:0] m183_33;
   assign m183_33 ={ {4{in183[5]}} , in183[5:0] };

   // m183_34 = W*in
   wire signed [9:0] m183_34;
   assign m183_34 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_35 = W*in
   wire signed [9:0] m183_35;
   assign m183_35 =10'b0;

   // m183_36 = W*in
   wire signed [9:0] m183_36;
   assign m183_36 =10'b0;

   // m183_37 = W*in
   wire signed [9:0] m183_37;
   assign m183_37 =10'b0;

   // m183_38 = W*in
   wire signed [9:0] m183_38;
   assign m183_38 =10'b0;

   // m183_39 = W*in
   wire signed [9:0] m183_39;
   assign m183_39 ={ {4{in183[5]}} , in183[5:0] };

   // m183_40 = W*in
   wire signed [9:0] m183_40;
   assign m183_40 =10'b0;

   // m183_41 = W*in
   wire signed [9:0] m183_41;
   assign m183_41 =10'b0;

   // m183_42 = W*in
   wire signed [9:0] m183_42;
   assign m183_42 ={ {3{neg183[5]}} , neg183 , {1{1'b0}} };

   // m183_43 = W*in
   wire signed [9:0] m183_43;
   assign m183_43 =10'b0;

   // m183_44 = W*in
   wire signed [9:0] m183_44;
   assign m183_44 =10'b0;

   // m183_45 = W*in
   wire signed [9:0] m183_45;
   assign m183_45 =10'b0;

   // m183_46 = W*in
   wire signed [9:0] m183_46;
   assign m183_46 ={ {4{in183[5]}} , in183[5:0] };

   // m183_47 = W*in
   wire signed [9:0] m183_47;
   assign m183_47 =10'b0;

   // m183_48 = W*in
   wire signed [9:0] m183_48;
   assign m183_48 ={ {4{in183[5]}} , in183[5:0] };

   // m183_49 = W*in
   wire signed [9:0] m183_49;
   assign m183_49 =10'b0;

   // m183_50 = W*in
   wire signed [9:0] m183_50;
   assign m183_50 =10'b0;

   // m183_51 = W*in
   wire signed [9:0] m183_51;
   assign m183_51 ={ {4{in183[5]}} , in183[5:0] };

   // m183_52 = W*in
   wire signed [9:0] m183_52;
   assign m183_52 =10'b0;

   // m183_53 = W*in
   wire signed [9:0] m183_53;
   assign m183_53 =10'b0;

   // m183_54 = W*in
   wire signed [9:0] m183_54;
   assign m183_54 =10'b0;

   // m183_55 = W*in
   wire signed [9:0] m183_55;
   assign m183_55 =10'b0;

   // m183_56 = W*in
   wire signed [9:0] m183_56;
   assign m183_56 =10'b0;

   // m183_57 = W*in
   wire signed [9:0] m183_57;
   assign m183_57 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_58 = W*in
   wire signed [9:0] m183_58;
   assign m183_58 =10'b0;

   // m183_59 = W*in
   wire signed [9:0] m183_59;
   assign m183_59 ={ {4{in183[5]}} , in183[5:0] };

   // m183_60 = W*in
   wire signed [9:0] m183_60;
   assign m183_60 =10'b0;

   // m183_61 = W*in
   wire signed [9:0] m183_61;
   assign m183_61 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_62 = W*in
   wire signed [9:0] m183_62;
   assign m183_62 =10'b0;

   // m183_63 = W*in
   wire signed [9:0] m183_63;
   assign m183_63 =10'b0;

   // m183_64 = W*in
   wire signed [9:0] m183_64;
   assign m183_64 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_65 = W*in
   wire signed [9:0] m183_65;
   assign m183_65 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_66 = W*in
   wire signed [9:0] m183_66;
   assign m183_66 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_67 = W*in
   wire signed [9:0] m183_67;
   assign m183_67 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_68 = W*in
   wire signed [9:0] m183_68;
   assign m183_68 ={ {4{in183[5]}} , in183[5:0] };

   // m183_69 = W*in
   wire signed [9:0] m183_69;
   assign m183_69 =10'b0;

   // m183_70 = W*in
   wire signed [9:0] m183_70;
   assign m183_70 =10'b0;

   // m183_71 = W*in
   wire signed [9:0] m183_71;
   assign m183_71 ={ {5{in183[5]}} , in183[5:1] };

   // m183_72 = W*in
   wire signed [9:0] m183_72;
   assign m183_72 ={ {5{in183[5]}} , in183[5:1] };

   // m183_73 = W*in
   wire signed [9:0] m183_73;
   assign m183_73 ={ {4{in183[5]}} , in183[5:0] };

   // m183_74 = W*in
   wire signed [9:0] m183_74;
   assign m183_74 =10'b0;

   // m183_75 = W*in
   wire signed [9:0] m183_75;
   assign m183_75 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_76 = W*in
   wire signed [9:0] m183_76;
   assign m183_76 =10'b0;

   // m183_77 = W*in
   wire signed [9:0] m183_77;
   assign m183_77 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_78 = W*in
   wire signed [9:0] m183_78;
   assign m183_78 =10'b0;

   // m183_79 = W*in
   wire signed [9:0] m183_79;
   assign m183_79 =10'b0;

   // m183_80 = W*in
   wire signed [9:0] m183_80;
   assign m183_80 =10'b0;

   // m183_81 = W*in
   wire signed [9:0] m183_81;
   assign m183_81 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_82 = W*in
   wire signed [9:0] m183_82;
   assign m183_82 =10'b0;

   // m183_83 = W*in
   wire signed [9:0] m183_83;
   assign m183_83 =10'b0;

   // m183_84 = W*in
   wire signed [9:0] m183_84;
   assign m183_84 =10'b0;

   // m183_85 = W*in
   wire signed [9:0] m183_85;
   assign m183_85 =10'b0;

   // m183_86 = W*in
   wire signed [9:0] m183_86;
   assign m183_86 =10'b0;

   // m183_87 = W*in
   wire signed [9:0] m183_87;
   assign m183_87 =10'b0;

   // m183_88 = W*in
   wire signed [9:0] m183_88;
   assign m183_88 =10'b0;

   // m183_89 = W*in
   wire signed [9:0] m183_89;
   assign m183_89 =10'b0;

   // m183_90 = W*in
   wire signed [9:0] m183_90;
   assign m183_90 =10'b0;

   // m183_91 = W*in
   wire signed [9:0] m183_91;
   assign m183_91 =10'b0;

   // m183_92 = W*in
   wire signed [9:0] m183_92;
   assign m183_92 =10'b0;

   // m183_93 = W*in
   wire signed [9:0] m183_93;
   assign m183_93 =10'b0;

   // m183_94 = W*in
   wire signed [9:0] m183_94;
   assign m183_94 ={ {3{neg183[5]}} , neg183 , {1{1'b0}} };

   // m183_95 = W*in
   wire signed [9:0] m183_95;
   assign m183_95 =10'b0;

   // m183_96 = W*in
   wire signed [9:0] m183_96;
   assign m183_96 =10'b0;

   // m183_97 = W*in
   wire signed [9:0] m183_97;
   assign m183_97 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_98 = W*in
   wire signed [9:0] m183_98;
   assign m183_98 =10'b0;

   // m183_99 = W*in
   wire signed [9:0] m183_99;
   assign m183_99 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_100 = W*in
   wire signed [9:0] m183_100;
   assign m183_100 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_101 = W*in
   wire signed [9:0] m183_101;
   assign m183_101 =10'b0;

   // m183_102 = W*in
   wire signed [9:0] m183_102;
   assign m183_102 =10'b0;

   // m183_103 = W*in
   wire signed [9:0] m183_103;
   assign m183_103 ={ {4{in183[5]}} , in183[5:0] };

   // m183_104 = W*in
   wire signed [9:0] m183_104;
   assign m183_104 ={ {4{in183[5]}} , in183[5:0] };

   // m183_105 = W*in
   wire signed [9:0] m183_105;
   assign m183_105 =10'b0;

   // m183_106 = W*in
   wire signed [9:0] m183_106;
   assign m183_106 =10'b0;

   // m183_107 = W*in
   wire signed [9:0] m183_107;
   assign m183_107 =10'b0;

   // m183_108 = W*in
   wire signed [9:0] m183_108;
   assign m183_108 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_109 = W*in
   wire signed [9:0] m183_109;
   assign m183_109 ={ {5{in183[5]}} , in183[5:1] };

   // m183_110 = W*in
   wire signed [9:0] m183_110;
   assign m183_110 =10'b0;

   // m183_111 = W*in
   wire signed [9:0] m183_111;
   assign m183_111 ={ {4{in183[5]}} , in183[5:0] };

   // m183_112 = W*in
   wire signed [9:0] m183_112;
   assign m183_112 ={ {4{neg183[5]}} , neg183[5:0] };

   // m183_113 = W*in
   wire signed [9:0] m183_113;
   assign m183_113 =10'b0;

   // m183_114 = W*in
   wire signed [9:0] m183_114;
   assign m183_114 =10'b0;

   // m183_115 = W*in
   wire signed [9:0] m183_115;
   assign m183_115 =10'b0;

   // m183_116 = W*in
   wire signed [9:0] m183_116;
   assign m183_116 =10'b0;

   // m183_117 = W*in
   wire signed [9:0] m183_117;
   assign m183_117 =10'b0;

   // m184_1 = W*in
   wire signed [9:0] m184_1;
   assign m184_1 =10'b0;

   // m184_2 = W*in
   wire signed [9:0] m184_2;
   assign m184_2 =10'b0;

   // m184_3 = W*in
   wire signed [9:0] m184_3;
   assign m184_3 =10'b0;

   // m184_4 = W*in
   wire signed [9:0] m184_4;
   assign m184_4 =10'b0;

   // m184_5 = W*in
   wire signed [9:0] m184_5;
   assign m184_5 =10'b0;

   // m184_6 = W*in
   wire signed [9:0] m184_6;
   assign m184_6 =10'b0;

   // m184_7 = W*in
   wire signed [9:0] m184_7;
   assign m184_7 =10'b0;

   // m184_8 = W*in
   wire signed [9:0] m184_8;
   assign m184_8 =10'b0;

   // m184_9 = W*in
   wire signed [9:0] m184_9;
   assign m184_9 =10'b0;

   // m184_10 = W*in
   wire signed [9:0] m184_10;
   assign m184_10 =10'b0;

   // m184_11 = W*in
   wire signed [9:0] m184_11;
   assign m184_11 =10'b0;

   // m184_12 = W*in
   wire signed [9:0] m184_12;
   assign m184_12 =10'b0;

   // m184_13 = W*in
   wire signed [9:0] m184_13;
   assign m184_13 =10'b0;

   // m184_14 = W*in
   wire signed [9:0] m184_14;
   assign m184_14 =10'b0;

   // m184_15 = W*in
   wire signed [9:0] m184_15;
   assign m184_15 =10'b0;

   // m184_16 = W*in
   wire signed [9:0] m184_16;
   assign m184_16 =10'b0;

   // m184_17 = W*in
   wire signed [9:0] m184_17;
   assign m184_17 =10'b0;

   // m184_18 = W*in
   wire signed [9:0] m184_18;
   assign m184_18 =10'b0;

   // m184_19 = W*in
   wire signed [9:0] m184_19;
   assign m184_19 =10'b0;

   // m184_20 = W*in
   wire signed [9:0] m184_20;
   assign m184_20 =10'b0;

   // m184_21 = W*in
   wire signed [9:0] m184_21;
   assign m184_21 =10'b0;

   // m184_22 = W*in
   wire signed [9:0] m184_22;
   assign m184_22 =10'b0;

   // m184_23 = W*in
   wire signed [9:0] m184_23;
   assign m184_23 =10'b0;

   // m184_24 = W*in
   wire signed [9:0] m184_24;
   assign m184_24 =10'b0;

   // m184_25 = W*in
   wire signed [9:0] m184_25;
   assign m184_25 ={ {5{in184[5]}} , in184[5:1] };

   // m184_26 = W*in
   wire signed [9:0] m184_26;
   assign m184_26 =10'b0;

   // m184_27 = W*in
   wire signed [9:0] m184_27;
   assign m184_27 =10'b0;

   // m184_28 = W*in
   wire signed [9:0] m184_28;
   assign m184_28 =10'b0;

   // m184_29 = W*in
   wire signed [9:0] m184_29;
   assign m184_29 =10'b0;

   // m184_30 = W*in
   wire signed [9:0] m184_30;
   assign m184_30 =10'b0;

   // m184_31 = W*in
   wire signed [9:0] m184_31;
   assign m184_31 =10'b0;

   // m184_32 = W*in
   wire signed [9:0] m184_32;
   assign m184_32 =10'b0;

   // m184_33 = W*in
   wire signed [9:0] m184_33;
   assign m184_33 =10'b0;

   // m184_34 = W*in
   wire signed [9:0] m184_34;
   assign m184_34 =10'b0;

   // m184_35 = W*in
   wire signed [9:0] m184_35;
   assign m184_35 =10'b0;

   // m184_36 = W*in
   wire signed [9:0] m184_36;
   assign m184_36 =10'b0;

   // m184_37 = W*in
   wire signed [9:0] m184_37;
   assign m184_37 =10'b0;

   // m184_38 = W*in
   wire signed [9:0] m184_38;
   assign m184_38 =10'b0;

   // m184_39 = W*in
   wire signed [9:0] m184_39;
   assign m184_39 =10'b0;

   // m184_40 = W*in
   wire signed [9:0] m184_40;
   assign m184_40 =10'b0;

   // m184_41 = W*in
   wire signed [9:0] m184_41;
   assign m184_41 =10'b0;

   // m184_42 = W*in
   wire signed [9:0] m184_42;
   assign m184_42 =10'b0;

   // m184_43 = W*in
   wire signed [9:0] m184_43;
   assign m184_43 =10'b0;

   // m184_44 = W*in
   wire signed [9:0] m184_44;
   assign m184_44 =10'b0;

   // m184_45 = W*in
   wire signed [9:0] m184_45;
   assign m184_45 =10'b0;

   // m184_46 = W*in
   wire signed [9:0] m184_46;
   assign m184_46 =10'b0;

   // m184_47 = W*in
   wire signed [9:0] m184_47;
   assign m184_47 =10'b0;

   // m184_48 = W*in
   wire signed [9:0] m184_48;
   assign m184_48 =10'b0;

   // m184_49 = W*in
   wire signed [9:0] m184_49;
   assign m184_49 =10'b0;

   // m184_50 = W*in
   wire signed [9:0] m184_50;
   assign m184_50 =10'b0;

   // m184_51 = W*in
   wire signed [9:0] m184_51;
   assign m184_51 =10'b0;

   // m184_52 = W*in
   wire signed [9:0] m184_52;
   assign m184_52 =10'b0;

   // m184_53 = W*in
   wire signed [9:0] m184_53;
   assign m184_53 =10'b0;

   // m184_54 = W*in
   wire signed [9:0] m184_54;
   assign m184_54 =10'b0;

   // m184_55 = W*in
   wire signed [9:0] m184_55;
   assign m184_55 =10'b0;

   // m184_56 = W*in
   wire signed [9:0] m184_56;
   assign m184_56 =10'b0;

   // m184_57 = W*in
   wire signed [9:0] m184_57;
   assign m184_57 =10'b0;

   // m184_58 = W*in
   wire signed [9:0] m184_58;
   assign m184_58 =10'b0;

   // m184_59 = W*in
   wire signed [9:0] m184_59;
   assign m184_59 =10'b0;

   // m184_60 = W*in
   wire signed [9:0] m184_60;
   assign m184_60 =10'b0;

   // m184_61 = W*in
   wire signed [9:0] m184_61;
   assign m184_61 =10'b0;

   // m184_62 = W*in
   wire signed [9:0] m184_62;
   assign m184_62 =10'b0;

   // m184_63 = W*in
   wire signed [9:0] m184_63;
   assign m184_63 =10'b0;

   // m184_64 = W*in
   wire signed [9:0] m184_64;
   assign m184_64 =10'b0;

   // m184_65 = W*in
   wire signed [9:0] m184_65;
   assign m184_65 =10'b0;

   // m184_66 = W*in
   wire signed [9:0] m184_66;
   assign m184_66 ={ {5{neg184[5]}} , neg184[5:1] };

   // m184_67 = W*in
   wire signed [9:0] m184_67;
   assign m184_67 =10'b0;

   // m184_68 = W*in
   wire signed [9:0] m184_68;
   assign m184_68 =10'b0;

   // m184_69 = W*in
   wire signed [9:0] m184_69;
   assign m184_69 =10'b0;

   // m184_70 = W*in
   wire signed [9:0] m184_70;
   assign m184_70 =10'b0;

   // m184_71 = W*in
   wire signed [9:0] m184_71;
   assign m184_71 =10'b0;

   // m184_72 = W*in
   wire signed [9:0] m184_72;
   assign m184_72 =10'b0;

   // m184_73 = W*in
   wire signed [9:0] m184_73;
   assign m184_73 =10'b0;

   // m184_74 = W*in
   wire signed [9:0] m184_74;
   assign m184_74 =10'b0;

   // m184_75 = W*in
   wire signed [9:0] m184_75;
   assign m184_75 =10'b0;

   // m184_76 = W*in
   wire signed [9:0] m184_76;
   assign m184_76 =10'b0;

   // m184_77 = W*in
   wire signed [9:0] m184_77;
   assign m184_77 =10'b0;

   // m184_78 = W*in
   wire signed [9:0] m184_78;
   assign m184_78 ={ {5{in184[5]}} , in184[5:1] };

   // m184_79 = W*in
   wire signed [9:0] m184_79;
   assign m184_79 =10'b0;

   // m184_80 = W*in
   wire signed [9:0] m184_80;
   assign m184_80 =10'b0;

   // m184_81 = W*in
   wire signed [9:0] m184_81;
   assign m184_81 =10'b0;

   // m184_82 = W*in
   wire signed [9:0] m184_82;
   assign m184_82 =10'b0;

   // m184_83 = W*in
   wire signed [9:0] m184_83;
   assign m184_83 =10'b0;

   // m184_84 = W*in
   wire signed [9:0] m184_84;
   assign m184_84 =10'b0;

   // m184_85 = W*in
   wire signed [9:0] m184_85;
   assign m184_85 =10'b0;

   // m184_86 = W*in
   wire signed [9:0] m184_86;
   assign m184_86 =10'b0;

   // m184_87 = W*in
   wire signed [9:0] m184_87;
   assign m184_87 =10'b0;

   // m184_88 = W*in
   wire signed [9:0] m184_88;
   assign m184_88 =10'b0;

   // m184_89 = W*in
   wire signed [9:0] m184_89;
   assign m184_89 =10'b0;

   // m184_90 = W*in
   wire signed [9:0] m184_90;
   assign m184_90 =10'b0;

   // m184_91 = W*in
   wire signed [9:0] m184_91;
   assign m184_91 =10'b0;

   // m184_92 = W*in
   wire signed [9:0] m184_92;
   assign m184_92 =10'b0;

   // m184_93 = W*in
   wire signed [9:0] m184_93;
   assign m184_93 =10'b0;

   // m184_94 = W*in
   wire signed [9:0] m184_94;
   assign m184_94 =10'b0;

   // m184_95 = W*in
   wire signed [9:0] m184_95;
   assign m184_95 =10'b0;

   // m184_96 = W*in
   wire signed [9:0] m184_96;
   assign m184_96 =10'b0;

   // m184_97 = W*in
   wire signed [9:0] m184_97;
   assign m184_97 =10'b0;

   // m184_98 = W*in
   wire signed [9:0] m184_98;
   assign m184_98 =10'b0;

   // m184_99 = W*in
   wire signed [9:0] m184_99;
   assign m184_99 =10'b0;

   // m184_100 = W*in
   wire signed [9:0] m184_100;
   assign m184_100 =10'b0;

   // m184_101 = W*in
   wire signed [9:0] m184_101;
   assign m184_101 =10'b0;

   // m184_102 = W*in
   wire signed [9:0] m184_102;
   assign m184_102 =10'b0;

   // m184_103 = W*in
   wire signed [9:0] m184_103;
   assign m184_103 =10'b0;

   // m184_104 = W*in
   wire signed [9:0] m184_104;
   assign m184_104 =10'b0;

   // m184_105 = W*in
   wire signed [9:0] m184_105;
   assign m184_105 =10'b0;

   // m184_106 = W*in
   wire signed [9:0] m184_106;
   assign m184_106 =10'b0;

   // m184_107 = W*in
   wire signed [9:0] m184_107;
   assign m184_107 =10'b0;

   // m184_108 = W*in
   wire signed [9:0] m184_108;
   assign m184_108 =10'b0;

   // m184_109 = W*in
   wire signed [9:0] m184_109;
   assign m184_109 ={ {5{in184[5]}} , in184[5:1] };

   // m184_110 = W*in
   wire signed [9:0] m184_110;
   assign m184_110 =10'b0;

   // m184_111 = W*in
   wire signed [9:0] m184_111;
   assign m184_111 =10'b0;

   // m184_112 = W*in
   wire signed [9:0] m184_112;
   assign m184_112 =10'b0;

   // m184_113 = W*in
   wire signed [9:0] m184_113;
   assign m184_113 =10'b0;

   // m184_114 = W*in
   wire signed [9:0] m184_114;
   assign m184_114 =10'b0;

   // m184_115 = W*in
   wire signed [9:0] m184_115;
   assign m184_115 =10'b0;

   // m184_116 = W*in
   wire signed [9:0] m184_116;
   assign m184_116 =10'b0;

   // m184_117 = W*in
   wire signed [9:0] m184_117;
   assign m184_117 =10'b0;

   // m185_1 = W*in
   wire signed [9:0] m185_1;
   assign m185_1 =10'b0;

   // m185_2 = W*in
   wire signed [9:0] m185_2;
   assign m185_2 =10'b0;

   // m185_3 = W*in
   wire signed [9:0] m185_3;
   assign m185_3 =10'b0;

   // m185_4 = W*in
   wire signed [9:0] m185_4;
   assign m185_4 =10'b0;

   // m185_5 = W*in
   wire signed [9:0] m185_5;
   assign m185_5 =10'b0;

   // m185_6 = W*in
   wire signed [9:0] m185_6;
   assign m185_6 =10'b0;

   // m185_7 = W*in
   wire signed [9:0] m185_7;
   assign m185_7 =10'b0;

   // m185_8 = W*in
   wire signed [9:0] m185_8;
   assign m185_8 =10'b0;

   // m185_9 = W*in
   wire signed [9:0] m185_9;
   assign m185_9 =10'b0;

   // m185_10 = W*in
   wire signed [9:0] m185_10;
   assign m185_10 =10'b0;

   // m185_11 = W*in
   wire signed [9:0] m185_11;
   assign m185_11 =10'b0;

   // m185_12 = W*in
   wire signed [9:0] m185_12;
   assign m185_12 =10'b0;

   // m185_13 = W*in
   wire signed [9:0] m185_13;
   assign m185_13 =10'b0;

   // m185_14 = W*in
   wire signed [9:0] m185_14;
   assign m185_14 =10'b0;

   // m185_15 = W*in
   wire signed [9:0] m185_15;
   assign m185_15 =10'b0;

   // m185_16 = W*in
   wire signed [9:0] m185_16;
   assign m185_16 ={ {5{neg185[5]}} , neg185[5:1] };

   // m185_17 = W*in
   wire signed [9:0] m185_17;
   assign m185_17 ={ {5{in185[5]}} , in185[5:1] };

   // m185_18 = W*in
   wire signed [9:0] m185_18;
   assign m185_18 =10'b0;

   // m185_19 = W*in
   wire signed [9:0] m185_19;
   assign m185_19 =10'b0;

   // m185_20 = W*in
   wire signed [9:0] m185_20;
   assign m185_20 =10'b0;

   // m185_21 = W*in
   wire signed [9:0] m185_21;
   assign m185_21 =10'b0;

   // m185_22 = W*in
   wire signed [9:0] m185_22;
   assign m185_22 ={ {5{in185[5]}} , in185[5:1] };

   // m185_23 = W*in
   wire signed [9:0] m185_23;
   assign m185_23 =10'b0;

   // m185_24 = W*in
   wire signed [9:0] m185_24;
   assign m185_24 =10'b0;

   // m185_25 = W*in
   wire signed [9:0] m185_25;
   assign m185_25 =10'b0;

   // m185_26 = W*in
   wire signed [9:0] m185_26;
   assign m185_26 =10'b0;

   // m185_27 = W*in
   wire signed [9:0] m185_27;
   assign m185_27 ={ {5{in185[5]}} , in185[5:1] };

   // m185_28 = W*in
   wire signed [9:0] m185_28;
   assign m185_28 ={ {5{neg185[5]}} , neg185[5:1] };

   // m185_29 = W*in
   wire signed [9:0] m185_29;
   assign m185_29 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_30 = W*in
   wire signed [9:0] m185_30;
   assign m185_30 =10'b0;

   // m185_31 = W*in
   wire signed [9:0] m185_31;
   assign m185_31 =10'b0;

   // m185_32 = W*in
   wire signed [9:0] m185_32;
   assign m185_32 =10'b0;

   // m185_33 = W*in
   wire signed [9:0] m185_33;
   assign m185_33 =10'b0;

   // m185_34 = W*in
   wire signed [9:0] m185_34;
   assign m185_34 =10'b0;

   // m185_35 = W*in
   wire signed [9:0] m185_35;
   assign m185_35 =10'b0;

   // m185_36 = W*in
   wire signed [9:0] m185_36;
   assign m185_36 =10'b0;

   // m185_37 = W*in
   wire signed [9:0] m185_37;
   assign m185_37 =10'b0;

   // m185_38 = W*in
   wire signed [9:0] m185_38;
   assign m185_38 =10'b0;

   // m185_39 = W*in
   wire signed [9:0] m185_39;
   assign m185_39 =10'b0;

   // m185_40 = W*in
   wire signed [9:0] m185_40;
   assign m185_40 =10'b0;

   // m185_41 = W*in
   wire signed [9:0] m185_41;
   assign m185_41 =10'b0;

   // m185_42 = W*in
   wire signed [9:0] m185_42;
   assign m185_42 =10'b0;

   // m185_43 = W*in
   wire signed [9:0] m185_43;
   assign m185_43 =10'b0;

   // m185_44 = W*in
   wire signed [9:0] m185_44;
   assign m185_44 =10'b0;

   // m185_45 = W*in
   wire signed [9:0] m185_45;
   assign m185_45 =10'b0;

   // m185_46 = W*in
   wire signed [9:0] m185_46;
   assign m185_46 ={ {4{in185[5]}} , in185[5:0] };

   // m185_47 = W*in
   wire signed [9:0] m185_47;
   assign m185_47 =10'b0;

   // m185_48 = W*in
   wire signed [9:0] m185_48;
   assign m185_48 =10'b0;

   // m185_49 = W*in
   wire signed [9:0] m185_49;
   assign m185_49 =10'b0;

   // m185_50 = W*in
   wire signed [9:0] m185_50;
   assign m185_50 =10'b0;

   // m185_51 = W*in
   wire signed [9:0] m185_51;
   assign m185_51 =10'b0;

   // m185_52 = W*in
   wire signed [9:0] m185_52;
   assign m185_52 =10'b0;

   // m185_53 = W*in
   wire signed [9:0] m185_53;
   assign m185_53 =10'b0;

   // m185_54 = W*in
   wire signed [9:0] m185_54;
   assign m185_54 =10'b0;

   // m185_55 = W*in
   wire signed [9:0] m185_55;
   assign m185_55 =10'b0;

   // m185_56 = W*in
   wire signed [9:0] m185_56;
   assign m185_56 =10'b0;

   // m185_57 = W*in
   wire signed [9:0] m185_57;
   assign m185_57 =10'b0;

   // m185_58 = W*in
   wire signed [9:0] m185_58;
   assign m185_58 =10'b0;

   // m185_59 = W*in
   wire signed [9:0] m185_59;
   assign m185_59 =10'b0;

   // m185_60 = W*in
   wire signed [9:0] m185_60;
   assign m185_60 =10'b0;

   // m185_61 = W*in
   wire signed [9:0] m185_61;
   assign m185_61 =10'b0;

   // m185_62 = W*in
   wire signed [9:0] m185_62;
   assign m185_62 =10'b0;

   // m185_63 = W*in
   wire signed [9:0] m185_63;
   assign m185_63 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_64 = W*in
   wire signed [9:0] m185_64;
   assign m185_64 ={ {4{in185[5]}} , in185[5:0] };

   // m185_65 = W*in
   wire signed [9:0] m185_65;
   assign m185_65 =10'b0;

   // m185_66 = W*in
   wire signed [9:0] m185_66;
   assign m185_66 =10'b0;

   // m185_67 = W*in
   wire signed [9:0] m185_67;
   assign m185_67 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_68 = W*in
   wire signed [9:0] m185_68;
   assign m185_68 =10'b0;

   // m185_69 = W*in
   wire signed [9:0] m185_69;
   assign m185_69 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_70 = W*in
   wire signed [9:0] m185_70;
   assign m185_70 ={ {5{neg185[5]}} , neg185[5:1] };

   // m185_71 = W*in
   wire signed [9:0] m185_71;
   assign m185_71 ={ {5{in185[5]}} , in185[5:1] };

   // m185_72 = W*in
   wire signed [9:0] m185_72;
   assign m185_72 =10'b0;

   // m185_73 = W*in
   wire signed [9:0] m185_73;
   assign m185_73 =10'b0;

   // m185_74 = W*in
   wire signed [9:0] m185_74;
   assign m185_74 =10'b0;

   // m185_75 = W*in
   wire signed [9:0] m185_75;
   assign m185_75 =10'b0;

   // m185_76 = W*in
   wire signed [9:0] m185_76;
   assign m185_76 =10'b0;

   // m185_77 = W*in
   wire signed [9:0] m185_77;
   assign m185_77 =10'b0;

   // m185_78 = W*in
   wire signed [9:0] m185_78;
   assign m185_78 =10'b0;

   // m185_79 = W*in
   wire signed [9:0] m185_79;
   assign m185_79 =10'b0;

   // m185_80 = W*in
   wire signed [9:0] m185_80;
   assign m185_80 =10'b0;

   // m185_81 = W*in
   wire signed [9:0] m185_81;
   assign m185_81 =10'b0;

   // m185_82 = W*in
   wire signed [9:0] m185_82;
   assign m185_82 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_83 = W*in
   wire signed [9:0] m185_83;
   assign m185_83 =10'b0;

   // m185_84 = W*in
   wire signed [9:0] m185_84;
   assign m185_84 =10'b0;

   // m185_85 = W*in
   wire signed [9:0] m185_85;
   assign m185_85 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_86 = W*in
   wire signed [9:0] m185_86;
   assign m185_86 =10'b0;

   // m185_87 = W*in
   wire signed [9:0] m185_87;
   assign m185_87 =10'b0;

   // m185_88 = W*in
   wire signed [9:0] m185_88;
   assign m185_88 =10'b0;

   // m185_89 = W*in
   wire signed [9:0] m185_89;
   assign m185_89 =10'b0;

   // m185_90 = W*in
   wire signed [9:0] m185_90;
   assign m185_90 =10'b0;

   // m185_91 = W*in
   wire signed [9:0] m185_91;
   assign m185_91 =10'b0;

   // m185_92 = W*in
   wire signed [9:0] m185_92;
   assign m185_92 =10'b0;

   // m185_93 = W*in
   wire signed [9:0] m185_93;
   assign m185_93 ={ {4{neg185[5]}} , neg185[5:0] };

   // m185_94 = W*in
   wire signed [9:0] m185_94;
   assign m185_94 =10'b0;

   // m185_95 = W*in
   wire signed [9:0] m185_95;
   assign m185_95 =10'b0;

   // m185_96 = W*in
   wire signed [9:0] m185_96;
   assign m185_96 =10'b0;

   // m185_97 = W*in
   wire signed [9:0] m185_97;
   assign m185_97 =10'b0;

   // m185_98 = W*in
   wire signed [9:0] m185_98;
   assign m185_98 =10'b0;

   // m185_99 = W*in
   wire signed [9:0] m185_99;
   assign m185_99 =10'b0;

   // m185_100 = W*in
   wire signed [9:0] m185_100;
   assign m185_100 =10'b0;

   // m185_101 = W*in
   wire signed [9:0] m185_101;
   assign m185_101 =10'b0;

   // m185_102 = W*in
   wire signed [9:0] m185_102;
   assign m185_102 =10'b0;

   // m185_103 = W*in
   wire signed [9:0] m185_103;
   assign m185_103 =10'b0;

   // m185_104 = W*in
   wire signed [9:0] m185_104;
   assign m185_104 =10'b0;

   // m185_105 = W*in
   wire signed [9:0] m185_105;
   assign m185_105 =10'b0;

   // m185_106 = W*in
   wire signed [9:0] m185_106;
   assign m185_106 =10'b0;

   // m185_107 = W*in
   wire signed [9:0] m185_107;
   assign m185_107 =10'b0;

   // m185_108 = W*in
   wire signed [9:0] m185_108;
   assign m185_108 =10'b0;

   // m185_109 = W*in
   wire signed [9:0] m185_109;
   assign m185_109 =10'b0;

   // m185_110 = W*in
   wire signed [9:0] m185_110;
   assign m185_110 =10'b0;

   // m185_111 = W*in
   wire signed [9:0] m185_111;
   assign m185_111 =10'b0;

   // m185_112 = W*in
   wire signed [9:0] m185_112;
   assign m185_112 =10'b0;

   // m185_113 = W*in
   wire signed [9:0] m185_113;
   assign m185_113 =10'b0;

   // m185_114 = W*in
   wire signed [9:0] m185_114;
   assign m185_114 ={ {5{in185[5]}} , in185[5:1] };

   // m185_115 = W*in
   wire signed [9:0] m185_115;
   assign m185_115 =10'b0;

   // m185_116 = W*in
   wire signed [9:0] m185_116;
   assign m185_116 =10'b0;

   // m185_117 = W*in
   wire signed [9:0] m185_117;
   assign m185_117 =10'b0;

   // m186_1 = W*in
   wire signed [9:0] m186_1;
   assign m186_1 =10'b0;

   // m186_2 = W*in
   wire signed [9:0] m186_2;
   assign m186_2 =10'b0;

   // m186_3 = W*in
   wire signed [9:0] m186_3;
   assign m186_3 =10'b0;

   // m186_4 = W*in
   wire signed [9:0] m186_4;
   assign m186_4 =10'b0;

   // m186_5 = W*in
   wire signed [9:0] m186_5;
   assign m186_5 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_6 = W*in
   wire signed [9:0] m186_6;
   assign m186_6 =10'b0;

   // m186_7 = W*in
   wire signed [9:0] m186_7;
   assign m186_7 =10'b0;

   // m186_8 = W*in
   wire signed [9:0] m186_8;
   assign m186_8 =10'b0;

   // m186_9 = W*in
   wire signed [9:0] m186_9;
   assign m186_9 =10'b0;

   // m186_10 = W*in
   wire signed [9:0] m186_10;
   assign m186_10 =10'b0;

   // m186_11 = W*in
   wire signed [9:0] m186_11;
   assign m186_11 =10'b0;

   // m186_12 = W*in
   wire signed [9:0] m186_12;
   assign m186_12 ={ {4{in186[5]}} , in186[5:0] };

   // m186_13 = W*in
   wire signed [9:0] m186_13;
   assign m186_13 =10'b0;

   // m186_14 = W*in
   wire signed [9:0] m186_14;
   assign m186_14 =10'b0;

   // m186_15 = W*in
   wire signed [9:0] m186_15;
   assign m186_15 =10'b0;

   // m186_16 = W*in
   wire signed [9:0] m186_16;
   assign m186_16 =10'b0;

   // m186_17 = W*in
   wire signed [9:0] m186_17;
   assign m186_17 ={ {4{in186[5]}} , in186[5:0] };

   // m186_18 = W*in
   wire signed [9:0] m186_18;
   assign m186_18 ={ {4{in186[5]}} , in186[5:0] };

   // m186_19 = W*in
   wire signed [9:0] m186_19;
   assign m186_19 =10'b0;

   // m186_20 = W*in
   wire signed [9:0] m186_20;
   assign m186_20 ={ {5{neg186[5]}} , neg186[5:1] };

   // m186_21 = W*in
   wire signed [9:0] m186_21;
   assign m186_21 =10'b0;

   // m186_22 = W*in
   wire signed [9:0] m186_22;
   assign m186_22 =10'b0;

   // m186_23 = W*in
   wire signed [9:0] m186_23;
   assign m186_23 =10'b0;

   // m186_24 = W*in
   wire signed [9:0] m186_24;
   assign m186_24 =10'b0;

   // m186_25 = W*in
   wire signed [9:0] m186_25;
   assign m186_25 ={ {5{neg186[5]}} , neg186[5:1] };

   // m186_26 = W*in
   wire signed [9:0] m186_26;
   assign m186_26 ={ {4{in186[5]}} , in186[5:0] };

   // m186_27 = W*in
   wire signed [9:0] m186_27;
   assign m186_27 ={ {5{in186[5]}} , in186[5:1] };

   // m186_28 = W*in
   wire signed [9:0] m186_28;
   assign m186_28 =10'b0;

   // m186_29 = W*in
   wire signed [9:0] m186_29;
   assign m186_29 =10'b0;

   // m186_30 = W*in
   wire signed [9:0] m186_30;
   assign m186_30 =10'b0;

   // m186_31 = W*in
   wire signed [9:0] m186_31;
   assign m186_31 ={ {4{in186[5]}} , in186[5:0] };

   // m186_32 = W*in
   wire signed [9:0] m186_32;
   assign m186_32 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_33 = W*in
   wire signed [9:0] m186_33;
   assign m186_33 =10'b0;

   // m186_34 = W*in
   wire signed [9:0] m186_34;
   assign m186_34 =10'b0;

   // m186_35 = W*in
   wire signed [9:0] m186_35;
   assign m186_35 ={ {5{neg186[5]}} , neg186[5:1] };

   // m186_36 = W*in
   wire signed [9:0] m186_36;
   assign m186_36 =10'b0;

   // m186_37 = W*in
   wire signed [9:0] m186_37;
   assign m186_37 =10'b0;

   // m186_38 = W*in
   wire signed [9:0] m186_38;
   assign m186_38 =10'b0;

   // m186_39 = W*in
   wire signed [9:0] m186_39;
   assign m186_39 =10'b0;

   // m186_40 = W*in
   wire signed [9:0] m186_40;
   assign m186_40 =10'b0;

   // m186_41 = W*in
   wire signed [9:0] m186_41;
   assign m186_41 =10'b0;

   // m186_42 = W*in
   wire signed [9:0] m186_42;
   assign m186_42 ={ {3{in186[5]}} , in186 , {1{1'b0}} };

   // m186_43 = W*in
   wire signed [9:0] m186_43;
   assign m186_43 =10'b0;

   // m186_44 = W*in
   wire signed [9:0] m186_44;
   assign m186_44 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_45 = W*in
   wire signed [9:0] m186_45;
   assign m186_45 ={ {4{in186[5]}} , in186[5:0] };

   // m186_46 = W*in
   wire signed [9:0] m186_46;
   assign m186_46 =10'b0;

   // m186_47 = W*in
   wire signed [9:0] m186_47;
   assign m186_47 =10'b0;

   // m186_48 = W*in
   wire signed [9:0] m186_48;
   assign m186_48 =10'b0;

   // m186_49 = W*in
   wire signed [9:0] m186_49;
   assign m186_49 =10'b0;

   // m186_50 = W*in
   wire signed [9:0] m186_50;
   assign m186_50 =10'b0;

   // m186_51 = W*in
   wire signed [9:0] m186_51;
   assign m186_51 ={ {4{in186[5]}} , in186[5:0] };

   // m186_52 = W*in
   wire signed [9:0] m186_52;
   assign m186_52 ={ {4{in186[5]}} , in186[5:0] };

   // m186_53 = W*in
   wire signed [9:0] m186_53;
   assign m186_53 =10'b0;

   // m186_54 = W*in
   wire signed [9:0] m186_54;
   assign m186_54 =10'b0;

   // m186_55 = W*in
   wire signed [9:0] m186_55;
   assign m186_55 =10'b0;

   // m186_56 = W*in
   wire signed [9:0] m186_56;
   assign m186_56 =10'b0;

   // m186_57 = W*in
   wire signed [9:0] m186_57;
   assign m186_57 =10'b0;

   // m186_58 = W*in
   wire signed [9:0] m186_58;
   assign m186_58 =10'b0;

   // m186_59 = W*in
   wire signed [9:0] m186_59;
   assign m186_59 =10'b0;

   // m186_60 = W*in
   wire signed [9:0] m186_60;
   assign m186_60 =10'b0;

   // m186_61 = W*in
   wire signed [9:0] m186_61;
   assign m186_61 =10'b0;

   // m186_62 = W*in
   wire signed [9:0] m186_62;
   assign m186_62 =10'b0;

   // m186_63 = W*in
   wire signed [9:0] m186_63;
   assign m186_63 ={ {3{neg186[5]}} , neg186 , {1{1'b0}} };

   // m186_64 = W*in
   wire signed [9:0] m186_64;
   assign m186_64 ={ {3{in186[5]}} , in186 , {1{1'b0}} };

   // m186_65 = W*in
   wire signed [9:0] m186_65;
   assign m186_65 =10'b0;

   // m186_66 = W*in
   wire signed [9:0] m186_66;
   assign m186_66 =10'b0;

   // m186_67 = W*in
   wire signed [9:0] m186_67;
   assign m186_67 =10'b0;

   // m186_68 = W*in
   wire signed [9:0] m186_68;
   assign m186_68 =10'b0;

   // m186_69 = W*in
   wire signed [9:0] m186_69;
   assign m186_69 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_70 = W*in
   wire signed [9:0] m186_70;
   assign m186_70 =10'b0;

   // m186_71 = W*in
   wire signed [9:0] m186_71;
   assign m186_71 =10'b0;

   // m186_72 = W*in
   wire signed [9:0] m186_72;
   assign m186_72 =10'b0;

   // m186_73 = W*in
   wire signed [9:0] m186_73;
   assign m186_73 =10'b0;

   // m186_74 = W*in
   wire signed [9:0] m186_74;
   assign m186_74 =10'b0;

   // m186_75 = W*in
   wire signed [9:0] m186_75;
   assign m186_75 =10'b0;

   // m186_76 = W*in
   wire signed [9:0] m186_76;
   assign m186_76 =10'b0;

   // m186_77 = W*in
   wire signed [9:0] m186_77;
   assign m186_77 ={ {4{in186[5]}} , in186[5:0] };

   // m186_78 = W*in
   wire signed [9:0] m186_78;
   assign m186_78 =10'b0;

   // m186_79 = W*in
   wire signed [9:0] m186_79;
   assign m186_79 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_80 = W*in
   wire signed [9:0] m186_80;
   assign m186_80 =10'b0;

   // m186_81 = W*in
   wire signed [9:0] m186_81;
   assign m186_81 ={ {4{in186[5]}} , in186[5:0] };

   // m186_82 = W*in
   wire signed [9:0] m186_82;
   assign m186_82 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_83 = W*in
   wire signed [9:0] m186_83;
   assign m186_83 ={ {4{in186[5]}} , in186[5:0] };

   // m186_84 = W*in
   wire signed [9:0] m186_84;
   assign m186_84 =10'b0;

   // m186_85 = W*in
   wire signed [9:0] m186_85;
   assign m186_85 =10'b0;

   // m186_86 = W*in
   wire signed [9:0] m186_86;
   assign m186_86 =10'b0;

   // m186_87 = W*in
   wire signed [9:0] m186_87;
   assign m186_87 =10'b0;

   // m186_88 = W*in
   wire signed [9:0] m186_88;
   assign m186_88 =10'b0;

   // m186_89 = W*in
   wire signed [9:0] m186_89;
   assign m186_89 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_90 = W*in
   wire signed [9:0] m186_90;
   assign m186_90 =10'b0;

   // m186_91 = W*in
   wire signed [9:0] m186_91;
   assign m186_91 =10'b0;

   // m186_92 = W*in
   wire signed [9:0] m186_92;
   assign m186_92 =10'b0;

   // m186_93 = W*in
   wire signed [9:0] m186_93;
   assign m186_93 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_94 = W*in
   wire signed [9:0] m186_94;
   assign m186_94 ={ {4{in186[5]}} , in186[5:0] };

   // m186_95 = W*in
   wire signed [9:0] m186_95;
   assign m186_95 =10'b0;

   // m186_96 = W*in
   wire signed [9:0] m186_96;
   assign m186_96 =10'b0;

   // m186_97 = W*in
   wire signed [9:0] m186_97;
   assign m186_97 ={ {4{in186[5]}} , in186[5:0] };

   // m186_98 = W*in
   wire signed [9:0] m186_98;
   assign m186_98 =10'b0;

   // m186_99 = W*in
   wire signed [9:0] m186_99;
   assign m186_99 =10'b0;

   // m186_100 = W*in
   wire signed [9:0] m186_100;
   assign m186_100 ={ {4{in186[5]}} , in186[5:0] };

   // m186_101 = W*in
   wire signed [9:0] m186_101;
   assign m186_101 =10'b0;

   // m186_102 = W*in
   wire signed [9:0] m186_102;
   assign m186_102 =10'b0;

   // m186_103 = W*in
   wire signed [9:0] m186_103;
   assign m186_103 =10'b0;

   // m186_104 = W*in
   wire signed [9:0] m186_104;
   assign m186_104 =10'b0;

   // m186_105 = W*in
   wire signed [9:0] m186_105;
   assign m186_105 =10'b0;

   // m186_106 = W*in
   wire signed [9:0] m186_106;
   assign m186_106 =10'b0;

   // m186_107 = W*in
   wire signed [9:0] m186_107;
   assign m186_107 ={ {4{in186[5]}} , in186[5:0] };

   // m186_108 = W*in
   wire signed [9:0] m186_108;
   assign m186_108 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_109 = W*in
   wire signed [9:0] m186_109;
   assign m186_109 ={ {4{neg186[5]}} , neg186[5:0] };

   // m186_110 = W*in
   wire signed [9:0] m186_110;
   assign m186_110 =10'b0;

   // m186_111 = W*in
   wire signed [9:0] m186_111;
   assign m186_111 =10'b0;

   // m186_112 = W*in
   wire signed [9:0] m186_112;
   assign m186_112 ={ {4{in186[5]}} , in186[5:0] };

   // m186_113 = W*in
   wire signed [9:0] m186_113;
   assign m186_113 =10'b0;

   // m186_114 = W*in
   wire signed [9:0] m186_114;
   assign m186_114 =10'b0;

   // m186_115 = W*in
   wire signed [9:0] m186_115;
   assign m186_115 =10'b0;

   // m186_116 = W*in
   wire signed [9:0] m186_116;
   assign m186_116 =10'b0;

   // m186_117 = W*in
   wire signed [9:0] m186_117;
   assign m186_117 =10'b0;

   // m187_1 = W*in
   wire signed [9:0] m187_1;
   assign m187_1 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_2 = W*in
   wire signed [9:0] m187_2;
   assign m187_2 =10'b0;

   // m187_3 = W*in
   wire signed [9:0] m187_3;
   assign m187_3 =10'b0;

   // m187_4 = W*in
   wire signed [9:0] m187_4;
   assign m187_4 =10'b0;

   // m187_5 = W*in
   wire signed [9:0] m187_5;
   assign m187_5 =10'b0;

   // m187_6 = W*in
   wire signed [9:0] m187_6;
   assign m187_6 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_7 = W*in
   wire signed [9:0] m187_7;
   assign m187_7 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_8 = W*in
   wire signed [9:0] m187_8;
   assign m187_8 =10'b0;

   // m187_9 = W*in
   wire signed [9:0] m187_9;
   assign m187_9 =10'b0;

   // m187_10 = W*in
   wire signed [9:0] m187_10;
   assign m187_10 =10'b0;

   // m187_11 = W*in
   wire signed [9:0] m187_11;
   assign m187_11 =10'b0;

   // m187_12 = W*in
   wire signed [9:0] m187_12;
   assign m187_12 ={ {5{in187[5]}} , in187[5:1] };

   // m187_13 = W*in
   wire signed [9:0] m187_13;
   assign m187_13 =10'b0;

   // m187_14 = W*in
   wire signed [9:0] m187_14;
   assign m187_14 =10'b0;

   // m187_15 = W*in
   wire signed [9:0] m187_15;
   assign m187_15 ={ {4{in187[5]}} , in187[5:0] };

   // m187_16 = W*in
   wire signed [9:0] m187_16;
   assign m187_16 =10'b0;

   // m187_17 = W*in
   wire signed [9:0] m187_17;
   assign m187_17 =10'b0;

   // m187_18 = W*in
   wire signed [9:0] m187_18;
   assign m187_18 =10'b0;

   // m187_19 = W*in
   wire signed [9:0] m187_19;
   assign m187_19 =10'b0;

   // m187_20 = W*in
   wire signed [9:0] m187_20;
   assign m187_20 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_21 = W*in
   wire signed [9:0] m187_21;
   assign m187_21 =10'b0;

   // m187_22 = W*in
   wire signed [9:0] m187_22;
   assign m187_22 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_23 = W*in
   wire signed [9:0] m187_23;
   assign m187_23 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_24 = W*in
   wire signed [9:0] m187_24;
   assign m187_24 =10'b0;

   // m187_25 = W*in
   wire signed [9:0] m187_25;
   assign m187_25 =10'b0;

   // m187_26 = W*in
   wire signed [9:0] m187_26;
   assign m187_26 ={ {4{in187[5]}} , in187[5:0] };

   // m187_27 = W*in
   wire signed [9:0] m187_27;
   assign m187_27 =10'b0;

   // m187_28 = W*in
   wire signed [9:0] m187_28;
   assign m187_28 =10'b0;

   // m187_29 = W*in
   wire signed [9:0] m187_29;
   assign m187_29 =10'b0;

   // m187_30 = W*in
   wire signed [9:0] m187_30;
   assign m187_30 =10'b0;

   // m187_31 = W*in
   wire signed [9:0] m187_31;
   assign m187_31 =10'b0;

   // m187_32 = W*in
   wire signed [9:0] m187_32;
   assign m187_32 =10'b0;

   // m187_33 = W*in
   wire signed [9:0] m187_33;
   assign m187_33 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_34 = W*in
   wire signed [9:0] m187_34;
   assign m187_34 =10'b0;

   // m187_35 = W*in
   wire signed [9:0] m187_35;
   assign m187_35 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_36 = W*in
   wire signed [9:0] m187_36;
   assign m187_36 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_37 = W*in
   wire signed [9:0] m187_37;
   assign m187_37 =10'b0;

   // m187_38 = W*in
   wire signed [9:0] m187_38;
   assign m187_38 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_39 = W*in
   wire signed [9:0] m187_39;
   assign m187_39 =10'b0;

   // m187_40 = W*in
   wire signed [9:0] m187_40;
   assign m187_40 =10'b0;

   // m187_41 = W*in
   wire signed [9:0] m187_41;
   assign m187_41 =10'b0;

   // m187_42 = W*in
   wire signed [9:0] m187_42;
   assign m187_42 =10'b0;

   // m187_43 = W*in
   wire signed [9:0] m187_43;
   assign m187_43 =10'b0;

   // m187_44 = W*in
   wire signed [9:0] m187_44;
   assign m187_44 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_45 = W*in
   wire signed [9:0] m187_45;
   assign m187_45 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_46 = W*in
   wire signed [9:0] m187_46;
   assign m187_46 =10'b0;

   // m187_47 = W*in
   wire signed [9:0] m187_47;
   assign m187_47 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_48 = W*in
   wire signed [9:0] m187_48;
   assign m187_48 ={ {4{in187[5]}} , in187[5:0] };

   // m187_49 = W*in
   wire signed [9:0] m187_49;
   assign m187_49 =10'b0;

   // m187_50 = W*in
   wire signed [9:0] m187_50;
   assign m187_50 ={ {4{in187[5]}} , in187[5:0] };

   // m187_51 = W*in
   wire signed [9:0] m187_51;
   assign m187_51 =10'b0;

   // m187_52 = W*in
   wire signed [9:0] m187_52;
   assign m187_52 =10'b0;

   // m187_53 = W*in
   wire signed [9:0] m187_53;
   assign m187_53 =10'b0;

   // m187_54 = W*in
   wire signed [9:0] m187_54;
   assign m187_54 =10'b0;

   // m187_55 = W*in
   wire signed [9:0] m187_55;
   assign m187_55 =10'b0;

   // m187_56 = W*in
   wire signed [9:0] m187_56;
   assign m187_56 =10'b0;

   // m187_57 = W*in
   wire signed [9:0] m187_57;
   assign m187_57 =10'b0;

   // m187_58 = W*in
   wire signed [9:0] m187_58;
   assign m187_58 =10'b0;

   // m187_59 = W*in
   wire signed [9:0] m187_59;
   assign m187_59 =10'b0;

   // m187_60 = W*in
   wire signed [9:0] m187_60;
   assign m187_60 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_61 = W*in
   wire signed [9:0] m187_61;
   assign m187_61 =10'b0;

   // m187_62 = W*in
   wire signed [9:0] m187_62;
   assign m187_62 =10'b0;

   // m187_63 = W*in
   wire signed [9:0] m187_63;
   assign m187_63 =10'b0;

   // m187_64 = W*in
   wire signed [9:0] m187_64;
   assign m187_64 =10'b0;

   // m187_65 = W*in
   wire signed [9:0] m187_65;
   assign m187_65 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_66 = W*in
   wire signed [9:0] m187_66;
   assign m187_66 =10'b0;

   // m187_67 = W*in
   wire signed [9:0] m187_67;
   assign m187_67 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_68 = W*in
   wire signed [9:0] m187_68;
   assign m187_68 ={ {4{in187[5]}} , in187[5:0] };

   // m187_69 = W*in
   wire signed [9:0] m187_69;
   assign m187_69 =10'b0;

   // m187_70 = W*in
   wire signed [9:0] m187_70;
   assign m187_70 =10'b0;

   // m187_71 = W*in
   wire signed [9:0] m187_71;
   assign m187_71 =10'b0;

   // m187_72 = W*in
   wire signed [9:0] m187_72;
   assign m187_72 ={ {4{in187[5]}} , in187[5:0] };

   // m187_73 = W*in
   wire signed [9:0] m187_73;
   assign m187_73 =10'b0;

   // m187_74 = W*in
   wire signed [9:0] m187_74;
   assign m187_74 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_75 = W*in
   wire signed [9:0] m187_75;
   assign m187_75 =10'b0;

   // m187_76 = W*in
   wire signed [9:0] m187_76;
   assign m187_76 =10'b0;

   // m187_77 = W*in
   wire signed [9:0] m187_77;
   assign m187_77 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_78 = W*in
   wire signed [9:0] m187_78;
   assign m187_78 =10'b0;

   // m187_79 = W*in
   wire signed [9:0] m187_79;
   assign m187_79 =10'b0;

   // m187_80 = W*in
   wire signed [9:0] m187_80;
   assign m187_80 =10'b0;

   // m187_81 = W*in
   wire signed [9:0] m187_81;
   assign m187_81 =10'b0;

   // m187_82 = W*in
   wire signed [9:0] m187_82;
   assign m187_82 =10'b0;

   // m187_83 = W*in
   wire signed [9:0] m187_83;
   assign m187_83 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_84 = W*in
   wire signed [9:0] m187_84;
   assign m187_84 =10'b0;

   // m187_85 = W*in
   wire signed [9:0] m187_85;
   assign m187_85 =10'b0;

   // m187_86 = W*in
   wire signed [9:0] m187_86;
   assign m187_86 =10'b0;

   // m187_87 = W*in
   wire signed [9:0] m187_87;
   assign m187_87 =10'b0;

   // m187_88 = W*in
   wire signed [9:0] m187_88;
   assign m187_88 =10'b0;

   // m187_89 = W*in
   wire signed [9:0] m187_89;
   assign m187_89 =10'b0;

   // m187_90 = W*in
   wire signed [9:0] m187_90;
   assign m187_90 ={ {4{in187[5]}} , in187[5:0] };

   // m187_91 = W*in
   wire signed [9:0] m187_91;
   assign m187_91 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_92 = W*in
   wire signed [9:0] m187_92;
   assign m187_92 ={ {3{in187[5]}} , in187 , {1{1'b0}} };

   // m187_93 = W*in
   wire signed [9:0] m187_93;
   assign m187_93 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_94 = W*in
   wire signed [9:0] m187_94;
   assign m187_94 =10'b0;

   // m187_95 = W*in
   wire signed [9:0] m187_95;
   assign m187_95 =10'b0;

   // m187_96 = W*in
   wire signed [9:0] m187_96;
   assign m187_96 =10'b0;

   // m187_97 = W*in
   wire signed [9:0] m187_97;
   assign m187_97 =10'b0;

   // m187_98 = W*in
   wire signed [9:0] m187_98;
   assign m187_98 =10'b0;

   // m187_99 = W*in
   wire signed [9:0] m187_99;
   assign m187_99 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_100 = W*in
   wire signed [9:0] m187_100;
   assign m187_100 =10'b0;

   // m187_101 = W*in
   wire signed [9:0] m187_101;
   assign m187_101 =10'b0;

   // m187_102 = W*in
   wire signed [9:0] m187_102;
   assign m187_102 =10'b0;

   // m187_103 = W*in
   wire signed [9:0] m187_103;
   assign m187_103 =10'b0;

   // m187_104 = W*in
   wire signed [9:0] m187_104;
   assign m187_104 =10'b0;

   // m187_105 = W*in
   wire signed [9:0] m187_105;
   assign m187_105 =10'b0;

   // m187_106 = W*in
   wire signed [9:0] m187_106;
   assign m187_106 =10'b0;

   // m187_107 = W*in
   wire signed [9:0] m187_107;
   assign m187_107 =10'b0;

   // m187_108 = W*in
   wire signed [9:0] m187_108;
   assign m187_108 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_109 = W*in
   wire signed [9:0] m187_109;
   assign m187_109 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_110 = W*in
   wire signed [9:0] m187_110;
   assign m187_110 =10'b0;

   // m187_111 = W*in
   wire signed [9:0] m187_111;
   assign m187_111 =10'b0;

   // m187_112 = W*in
   wire signed [9:0] m187_112;
   assign m187_112 =10'b0;

   // m187_113 = W*in
   wire signed [9:0] m187_113;
   assign m187_113 ={ {4{in187[5]}} , in187[5:0] };

   // m187_114 = W*in
   wire signed [9:0] m187_114;
   assign m187_114 ={ {4{neg187[5]}} , neg187[5:0] };

   // m187_115 = W*in
   wire signed [9:0] m187_115;
   assign m187_115 ={ {5{neg187[5]}} , neg187[5:1] };

   // m187_116 = W*in
   wire signed [9:0] m187_116;
   assign m187_116 =10'b0;

   // m187_117 = W*in
   wire signed [9:0] m187_117;
   assign m187_117 ={ {4{neg187[5]}} , neg187[5:0] };

   // m188_1 = W*in
   wire signed [9:0] m188_1;
   assign m188_1 =10'b0;

   // m188_2 = W*in
   wire signed [9:0] m188_2;
   assign m188_2 =10'b0;

   // m188_3 = W*in
   wire signed [9:0] m188_3;
   assign m188_3 =10'b0;

   // m188_4 = W*in
   wire signed [9:0] m188_4;
   assign m188_4 =10'b0;

   // m188_5 = W*in
   wire signed [9:0] m188_5;
   assign m188_5 ={ {4{in188[5]}} , in188[5:0] };

   // m188_6 = W*in
   wire signed [9:0] m188_6;
   assign m188_6 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_7 = W*in
   wire signed [9:0] m188_7;
   assign m188_7 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_8 = W*in
   wire signed [9:0] m188_8;
   assign m188_8 =10'b0;

   // m188_9 = W*in
   wire signed [9:0] m188_9;
   assign m188_9 =10'b0;

   // m188_10 = W*in
   wire signed [9:0] m188_10;
   assign m188_10 =10'b0;

   // m188_11 = W*in
   wire signed [9:0] m188_11;
   assign m188_11 =10'b0;

   // m188_12 = W*in
   wire signed [9:0] m188_12;
   assign m188_12 =10'b0;

   // m188_13 = W*in
   wire signed [9:0] m188_13;
   assign m188_13 =10'b0;

   // m188_14 = W*in
   wire signed [9:0] m188_14;
   assign m188_14 =10'b0;

   // m188_15 = W*in
   wire signed [9:0] m188_15;
   assign m188_15 ={ {4{in188[5]}} , in188[5:0] };

   // m188_16 = W*in
   wire signed [9:0] m188_16;
   assign m188_16 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_17 = W*in
   wire signed [9:0] m188_17;
   assign m188_17 =10'b0;

   // m188_18 = W*in
   wire signed [9:0] m188_18;
   assign m188_18 =10'b0;

   // m188_19 = W*in
   wire signed [9:0] m188_19;
   assign m188_19 =10'b0;

   // m188_20 = W*in
   wire signed [9:0] m188_20;
   assign m188_20 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_21 = W*in
   wire signed [9:0] m188_21;
   assign m188_21 =10'b0;

   // m188_22 = W*in
   wire signed [9:0] m188_22;
   assign m188_22 =10'b0;

   // m188_23 = W*in
   wire signed [9:0] m188_23;
   assign m188_23 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_24 = W*in
   wire signed [9:0] m188_24;
   assign m188_24 =10'b0;

   // m188_25 = W*in
   wire signed [9:0] m188_25;
   assign m188_25 =10'b0;

   // m188_26 = W*in
   wire signed [9:0] m188_26;
   assign m188_26 ={ {4{in188[5]}} , in188[5:0] };

   // m188_27 = W*in
   wire signed [9:0] m188_27;
   assign m188_27 =10'b0;

   // m188_28 = W*in
   wire signed [9:0] m188_28;
   assign m188_28 =10'b0;

   // m188_29 = W*in
   wire signed [9:0] m188_29;
   assign m188_29 =10'b0;

   // m188_30 = W*in
   wire signed [9:0] m188_30;
   assign m188_30 =10'b0;

   // m188_31 = W*in
   wire signed [9:0] m188_31;
   assign m188_31 ={ {5{in188[5]}} , in188[5:1] };

   // m188_32 = W*in
   wire signed [9:0] m188_32;
   assign m188_32 =10'b0;

   // m188_33 = W*in
   wire signed [9:0] m188_33;
   assign m188_33 =10'b0;

   // m188_34 = W*in
   wire signed [9:0] m188_34;
   assign m188_34 =10'b0;

   // m188_35 = W*in
   wire signed [9:0] m188_35;
   assign m188_35 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_36 = W*in
   wire signed [9:0] m188_36;
   assign m188_36 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_37 = W*in
   wire signed [9:0] m188_37;
   assign m188_37 =10'b0;

   // m188_38 = W*in
   wire signed [9:0] m188_38;
   assign m188_38 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_39 = W*in
   wire signed [9:0] m188_39;
   assign m188_39 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_40 = W*in
   wire signed [9:0] m188_40;
   assign m188_40 =10'b0;

   // m188_41 = W*in
   wire signed [9:0] m188_41;
   assign m188_41 =10'b0;

   // m188_42 = W*in
   wire signed [9:0] m188_42;
   assign m188_42 =10'b0;

   // m188_43 = W*in
   wire signed [9:0] m188_43;
   assign m188_43 =10'b0;

   // m188_44 = W*in
   wire signed [9:0] m188_44;
   assign m188_44 =10'b0;

   // m188_45 = W*in
   wire signed [9:0] m188_45;
   assign m188_45 =10'b0;

   // m188_46 = W*in
   wire signed [9:0] m188_46;
   assign m188_46 =10'b0;

   // m188_47 = W*in
   wire signed [9:0] m188_47;
   assign m188_47 =10'b0;

   // m188_48 = W*in
   wire signed [9:0] m188_48;
   assign m188_48 =10'b0;

   // m188_49 = W*in
   wire signed [9:0] m188_49;
   assign m188_49 =10'b0;

   // m188_50 = W*in
   wire signed [9:0] m188_50;
   assign m188_50 =10'b0;

   // m188_51 = W*in
   wire signed [9:0] m188_51;
   assign m188_51 ={ {4{in188[5]}} , in188[5:0] };

   // m188_52 = W*in
   wire signed [9:0] m188_52;
   assign m188_52 ={ {4{in188[5]}} , in188[5:0] };

   // m188_53 = W*in
   wire signed [9:0] m188_53;
   assign m188_53 =10'b0;

   // m188_54 = W*in
   wire signed [9:0] m188_54;
   assign m188_54 =10'b0;

   // m188_55 = W*in
   wire signed [9:0] m188_55;
   assign m188_55 =10'b0;

   // m188_56 = W*in
   wire signed [9:0] m188_56;
   assign m188_56 =10'b0;

   // m188_57 = W*in
   wire signed [9:0] m188_57;
   assign m188_57 =10'b0;

   // m188_58 = W*in
   wire signed [9:0] m188_58;
   assign m188_58 =10'b0;

   // m188_59 = W*in
   wire signed [9:0] m188_59;
   assign m188_59 =10'b0;

   // m188_60 = W*in
   wire signed [9:0] m188_60;
   assign m188_60 =10'b0;

   // m188_61 = W*in
   wire signed [9:0] m188_61;
   assign m188_61 =10'b0;

   // m188_62 = W*in
   wire signed [9:0] m188_62;
   assign m188_62 =10'b0;

   // m188_63 = W*in
   wire signed [9:0] m188_63;
   assign m188_63 =10'b0;

   // m188_64 = W*in
   wire signed [9:0] m188_64;
   assign m188_64 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_65 = W*in
   wire signed [9:0] m188_65;
   assign m188_65 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_66 = W*in
   wire signed [9:0] m188_66;
   assign m188_66 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_67 = W*in
   wire signed [9:0] m188_67;
   assign m188_67 =10'b0;

   // m188_68 = W*in
   wire signed [9:0] m188_68;
   assign m188_68 ={ {4{in188[5]}} , in188[5:0] };

   // m188_69 = W*in
   wire signed [9:0] m188_69;
   assign m188_69 =10'b0;

   // m188_70 = W*in
   wire signed [9:0] m188_70;
   assign m188_70 =10'b0;

   // m188_71 = W*in
   wire signed [9:0] m188_71;
   assign m188_71 =10'b0;

   // m188_72 = W*in
   wire signed [9:0] m188_72;
   assign m188_72 =10'b0;

   // m188_73 = W*in
   wire signed [9:0] m188_73;
   assign m188_73 =10'b0;

   // m188_74 = W*in
   wire signed [9:0] m188_74;
   assign m188_74 =10'b0;

   // m188_75 = W*in
   wire signed [9:0] m188_75;
   assign m188_75 =10'b0;

   // m188_76 = W*in
   wire signed [9:0] m188_76;
   assign m188_76 =10'b0;

   // m188_77 = W*in
   wire signed [9:0] m188_77;
   assign m188_77 =10'b0;

   // m188_78 = W*in
   wire signed [9:0] m188_78;
   assign m188_78 ={ {5{in188[5]}} , in188[5:1] };

   // m188_79 = W*in
   wire signed [9:0] m188_79;
   assign m188_79 =10'b0;

   // m188_80 = W*in
   wire signed [9:0] m188_80;
   assign m188_80 =10'b0;

   // m188_81 = W*in
   wire signed [9:0] m188_81;
   assign m188_81 =10'b0;

   // m188_82 = W*in
   wire signed [9:0] m188_82;
   assign m188_82 ={ {5{in188[5]}} , in188[5:1] };

   // m188_83 = W*in
   wire signed [9:0] m188_83;
   assign m188_83 =10'b0;

   // m188_84 = W*in
   wire signed [9:0] m188_84;
   assign m188_84 =10'b0;

   // m188_85 = W*in
   wire signed [9:0] m188_85;
   assign m188_85 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_86 = W*in
   wire signed [9:0] m188_86;
   assign m188_86 =10'b0;

   // m188_87 = W*in
   wire signed [9:0] m188_87;
   assign m188_87 =10'b0;

   // m188_88 = W*in
   wire signed [9:0] m188_88;
   assign m188_88 =10'b0;

   // m188_89 = W*in
   wire signed [9:0] m188_89;
   assign m188_89 =10'b0;

   // m188_90 = W*in
   wire signed [9:0] m188_90;
   assign m188_90 =10'b0;

   // m188_91 = W*in
   wire signed [9:0] m188_91;
   assign m188_91 =10'b0;

   // m188_92 = W*in
   wire signed [9:0] m188_92;
   assign m188_92 =10'b0;

   // m188_93 = W*in
   wire signed [9:0] m188_93;
   assign m188_93 =10'b0;

   // m188_94 = W*in
   wire signed [9:0] m188_94;
   assign m188_94 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_95 = W*in
   wire signed [9:0] m188_95;
   assign m188_95 =10'b0;

   // m188_96 = W*in
   wire signed [9:0] m188_96;
   assign m188_96 =10'b0;

   // m188_97 = W*in
   wire signed [9:0] m188_97;
   assign m188_97 =10'b0;

   // m188_98 = W*in
   wire signed [9:0] m188_98;
   assign m188_98 =10'b0;

   // m188_99 = W*in
   wire signed [9:0] m188_99;
   assign m188_99 =10'b0;

   // m188_100 = W*in
   wire signed [9:0] m188_100;
   assign m188_100 =10'b0;

   // m188_101 = W*in
   wire signed [9:0] m188_101;
   assign m188_101 =10'b0;

   // m188_102 = W*in
   wire signed [9:0] m188_102;
   assign m188_102 =10'b0;

   // m188_103 = W*in
   wire signed [9:0] m188_103;
   assign m188_103 =10'b0;

   // m188_104 = W*in
   wire signed [9:0] m188_104;
   assign m188_104 =10'b0;

   // m188_105 = W*in
   wire signed [9:0] m188_105;
   assign m188_105 =10'b0;

   // m188_106 = W*in
   wire signed [9:0] m188_106;
   assign m188_106 =10'b0;

   // m188_107 = W*in
   wire signed [9:0] m188_107;
   assign m188_107 =10'b0;

   // m188_108 = W*in
   wire signed [9:0] m188_108;
   assign m188_108 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_109 = W*in
   wire signed [9:0] m188_109;
   assign m188_109 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_110 = W*in
   wire signed [9:0] m188_110;
   assign m188_110 ={ {4{neg188[5]}} , neg188[5:0] };

   // m188_111 = W*in
   wire signed [9:0] m188_111;
   assign m188_111 =10'b0;

   // m188_112 = W*in
   wire signed [9:0] m188_112;
   assign m188_112 =10'b0;

   // m188_113 = W*in
   wire signed [9:0] m188_113;
   assign m188_113 =10'b0;

   // m188_114 = W*in
   wire signed [9:0] m188_114;
   assign m188_114 ={ {5{neg188[5]}} , neg188[5:1] };

   // m188_115 = W*in
   wire signed [9:0] m188_115;
   assign m188_115 =10'b0;

   // m188_116 = W*in
   wire signed [9:0] m188_116;
   assign m188_116 =10'b0;

   // m188_117 = W*in
   wire signed [9:0] m188_117;
   assign m188_117 =10'b0;

   // m189_1 = W*in
   wire signed [9:0] m189_1;
   assign m189_1 =10'b0;

   // m189_2 = W*in
   wire signed [9:0] m189_2;
   assign m189_2 =10'b0;

   // m189_3 = W*in
   wire signed [9:0] m189_3;
   assign m189_3 =10'b0;

   // m189_4 = W*in
   wire signed [9:0] m189_4;
   assign m189_4 =10'b0;

   // m189_5 = W*in
   wire signed [9:0] m189_5;
   assign m189_5 =10'b0;

   // m189_6 = W*in
   wire signed [9:0] m189_6;
   assign m189_6 =10'b0;

   // m189_7 = W*in
   wire signed [9:0] m189_7;
   assign m189_7 =10'b0;

   // m189_8 = W*in
   wire signed [9:0] m189_8;
   assign m189_8 =10'b0;

   // m189_9 = W*in
   wire signed [9:0] m189_9;
   assign m189_9 =10'b0;

   // m189_10 = W*in
   wire signed [9:0] m189_10;
   assign m189_10 =10'b0;

   // m189_11 = W*in
   wire signed [9:0] m189_11;
   assign m189_11 =10'b0;

   // m189_12 = W*in
   wire signed [9:0] m189_12;
   assign m189_12 =10'b0;

   // m189_13 = W*in
   wire signed [9:0] m189_13;
   assign m189_13 =10'b0;

   // m189_14 = W*in
   wire signed [9:0] m189_14;
   assign m189_14 =10'b0;

   // m189_15 = W*in
   wire signed [9:0] m189_15;
   assign m189_15 =10'b0;

   // m189_16 = W*in
   wire signed [9:0] m189_16;
   assign m189_16 =10'b0;

   // m189_17 = W*in
   wire signed [9:0] m189_17;
   assign m189_17 =10'b0;

   // m189_18 = W*in
   wire signed [9:0] m189_18;
   assign m189_18 =10'b0;

   // m189_19 = W*in
   wire signed [9:0] m189_19;
   assign m189_19 =10'b0;

   // m189_20 = W*in
   wire signed [9:0] m189_20;
   assign m189_20 =10'b0;

   // m189_21 = W*in
   wire signed [9:0] m189_21;
   assign m189_21 =10'b0;

   // m189_22 = W*in
   wire signed [9:0] m189_22;
   assign m189_22 =10'b0;

   // m189_23 = W*in
   wire signed [9:0] m189_23;
   assign m189_23 =10'b0;

   // m189_24 = W*in
   wire signed [9:0] m189_24;
   assign m189_24 =10'b0;

   // m189_25 = W*in
   wire signed [9:0] m189_25;
   assign m189_25 =10'b0;

   // m189_26 = W*in
   wire signed [9:0] m189_26;
   assign m189_26 =10'b0;

   // m189_27 = W*in
   wire signed [9:0] m189_27;
   assign m189_27 =10'b0;

   // m189_28 = W*in
   wire signed [9:0] m189_28;
   assign m189_28 =10'b0;

   // m189_29 = W*in
   wire signed [9:0] m189_29;
   assign m189_29 =10'b0;

   // m189_30 = W*in
   wire signed [9:0] m189_30;
   assign m189_30 =10'b0;

   // m189_31 = W*in
   wire signed [9:0] m189_31;
   assign m189_31 =10'b0;

   // m189_32 = W*in
   wire signed [9:0] m189_32;
   assign m189_32 =10'b0;

   // m189_33 = W*in
   wire signed [9:0] m189_33;
   assign m189_33 =10'b0;

   // m189_34 = W*in
   wire signed [9:0] m189_34;
   assign m189_34 =10'b0;

   // m189_35 = W*in
   wire signed [9:0] m189_35;
   assign m189_35 =10'b0;

   // m189_36 = W*in
   wire signed [9:0] m189_36;
   assign m189_36 =10'b0;

   // m189_37 = W*in
   wire signed [9:0] m189_37;
   assign m189_37 =10'b0;

   // m189_38 = W*in
   wire signed [9:0] m189_38;
   assign m189_38 =10'b0;

   // m189_39 = W*in
   wire signed [9:0] m189_39;
   assign m189_39 =10'b0;

   // m189_40 = W*in
   wire signed [9:0] m189_40;
   assign m189_40 =10'b0;

   // m189_41 = W*in
   wire signed [9:0] m189_41;
   assign m189_41 =10'b0;

   // m189_42 = W*in
   wire signed [9:0] m189_42;
   assign m189_42 =10'b0;

   // m189_43 = W*in
   wire signed [9:0] m189_43;
   assign m189_43 =10'b0;

   // m189_44 = W*in
   wire signed [9:0] m189_44;
   assign m189_44 =10'b0;

   // m189_45 = W*in
   wire signed [9:0] m189_45;
   assign m189_45 =10'b0;

   // m189_46 = W*in
   wire signed [9:0] m189_46;
   assign m189_46 =10'b0;

   // m189_47 = W*in
   wire signed [9:0] m189_47;
   assign m189_47 =10'b0;

   // m189_48 = W*in
   wire signed [9:0] m189_48;
   assign m189_48 =10'b0;

   // m189_49 = W*in
   wire signed [9:0] m189_49;
   assign m189_49 =10'b0;

   // m189_50 = W*in
   wire signed [9:0] m189_50;
   assign m189_50 =10'b0;

   // m189_51 = W*in
   wire signed [9:0] m189_51;
   assign m189_51 =10'b0;

   // m189_52 = W*in
   wire signed [9:0] m189_52;
   assign m189_52 =10'b0;

   // m189_53 = W*in
   wire signed [9:0] m189_53;
   assign m189_53 =10'b0;

   // m189_54 = W*in
   wire signed [9:0] m189_54;
   assign m189_54 =10'b0;

   // m189_55 = W*in
   wire signed [9:0] m189_55;
   assign m189_55 =10'b0;

   // m189_56 = W*in
   wire signed [9:0] m189_56;
   assign m189_56 =10'b0;

   // m189_57 = W*in
   wire signed [9:0] m189_57;
   assign m189_57 =10'b0;

   // m189_58 = W*in
   wire signed [9:0] m189_58;
   assign m189_58 =10'b0;

   // m189_59 = W*in
   wire signed [9:0] m189_59;
   assign m189_59 =10'b0;

   // m189_60 = W*in
   wire signed [9:0] m189_60;
   assign m189_60 =10'b0;

   // m189_61 = W*in
   wire signed [9:0] m189_61;
   assign m189_61 =10'b0;

   // m189_62 = W*in
   wire signed [9:0] m189_62;
   assign m189_62 =10'b0;

   // m189_63 = W*in
   wire signed [9:0] m189_63;
   assign m189_63 =10'b0;

   // m189_64 = W*in
   wire signed [9:0] m189_64;
   assign m189_64 =10'b0;

   // m189_65 = W*in
   wire signed [9:0] m189_65;
   assign m189_65 =10'b0;

   // m189_66 = W*in
   wire signed [9:0] m189_66;
   assign m189_66 =10'b0;

   // m189_67 = W*in
   wire signed [9:0] m189_67;
   assign m189_67 =10'b0;

   // m189_68 = W*in
   wire signed [9:0] m189_68;
   assign m189_68 =10'b0;

   // m189_69 = W*in
   wire signed [9:0] m189_69;
   assign m189_69 =10'b0;

   // m189_70 = W*in
   wire signed [9:0] m189_70;
   assign m189_70 =10'b0;

   // m189_71 = W*in
   wire signed [9:0] m189_71;
   assign m189_71 =10'b0;

   // m189_72 = W*in
   wire signed [9:0] m189_72;
   assign m189_72 =10'b0;

   // m189_73 = W*in
   wire signed [9:0] m189_73;
   assign m189_73 =10'b0;

   // m189_74 = W*in
   wire signed [9:0] m189_74;
   assign m189_74 =10'b0;

   // m189_75 = W*in
   wire signed [9:0] m189_75;
   assign m189_75 =10'b0;

   // m189_76 = W*in
   wire signed [9:0] m189_76;
   assign m189_76 =10'b0;

   // m189_77 = W*in
   wire signed [9:0] m189_77;
   assign m189_77 =10'b0;

   // m189_78 = W*in
   wire signed [9:0] m189_78;
   assign m189_78 =10'b0;

   // m189_79 = W*in
   wire signed [9:0] m189_79;
   assign m189_79 =10'b0;

   // m189_80 = W*in
   wire signed [9:0] m189_80;
   assign m189_80 =10'b0;

   // m189_81 = W*in
   wire signed [9:0] m189_81;
   assign m189_81 =10'b0;

   // m189_82 = W*in
   wire signed [9:0] m189_82;
   assign m189_82 =10'b0;

   // m189_83 = W*in
   wire signed [9:0] m189_83;
   assign m189_83 =10'b0;

   // m189_84 = W*in
   wire signed [9:0] m189_84;
   assign m189_84 =10'b0;

   // m189_85 = W*in
   wire signed [9:0] m189_85;
   assign m189_85 =10'b0;

   // m189_86 = W*in
   wire signed [9:0] m189_86;
   assign m189_86 =10'b0;

   // m189_87 = W*in
   wire signed [9:0] m189_87;
   assign m189_87 =10'b0;

   // m189_88 = W*in
   wire signed [9:0] m189_88;
   assign m189_88 =10'b0;

   // m189_89 = W*in
   wire signed [9:0] m189_89;
   assign m189_89 =10'b0;

   // m189_90 = W*in
   wire signed [9:0] m189_90;
   assign m189_90 =10'b0;

   // m189_91 = W*in
   wire signed [9:0] m189_91;
   assign m189_91 =10'b0;

   // m189_92 = W*in
   wire signed [9:0] m189_92;
   assign m189_92 =10'b0;

   // m189_93 = W*in
   wire signed [9:0] m189_93;
   assign m189_93 =10'b0;

   // m189_94 = W*in
   wire signed [9:0] m189_94;
   assign m189_94 =10'b0;

   // m189_95 = W*in
   wire signed [9:0] m189_95;
   assign m189_95 =10'b0;

   // m189_96 = W*in
   wire signed [9:0] m189_96;
   assign m189_96 =10'b0;

   // m189_97 = W*in
   wire signed [9:0] m189_97;
   assign m189_97 =10'b0;

   // m189_98 = W*in
   wire signed [9:0] m189_98;
   assign m189_98 =10'b0;

   // m189_99 = W*in
   wire signed [9:0] m189_99;
   assign m189_99 =10'b0;

   // m189_100 = W*in
   wire signed [9:0] m189_100;
   assign m189_100 =10'b0;

   // m189_101 = W*in
   wire signed [9:0] m189_101;
   assign m189_101 =10'b0;

   // m189_102 = W*in
   wire signed [9:0] m189_102;
   assign m189_102 =10'b0;

   // m189_103 = W*in
   wire signed [9:0] m189_103;
   assign m189_103 =10'b0;

   // m189_104 = W*in
   wire signed [9:0] m189_104;
   assign m189_104 =10'b0;

   // m189_105 = W*in
   wire signed [9:0] m189_105;
   assign m189_105 =10'b0;

   // m189_106 = W*in
   wire signed [9:0] m189_106;
   assign m189_106 =10'b0;

   // m189_107 = W*in
   wire signed [9:0] m189_107;
   assign m189_107 =10'b0;

   // m189_108 = W*in
   wire signed [9:0] m189_108;
   assign m189_108 =10'b0;

   // m189_109 = W*in
   wire signed [9:0] m189_109;
   assign m189_109 ={ {5{neg189[5]}} , neg189[5:1] };

   // m189_110 = W*in
   wire signed [9:0] m189_110;
   assign m189_110 =10'b0;

   // m189_111 = W*in
   wire signed [9:0] m189_111;
   assign m189_111 =10'b0;

   // m189_112 = W*in
   wire signed [9:0] m189_112;
   assign m189_112 =10'b0;

   // m189_113 = W*in
   wire signed [9:0] m189_113;
   assign m189_113 =10'b0;

   // m189_114 = W*in
   wire signed [9:0] m189_114;
   assign m189_114 =10'b0;

   // m189_115 = W*in
   wire signed [9:0] m189_115;
   assign m189_115 =10'b0;

   // m189_116 = W*in
   wire signed [9:0] m189_116;
   assign m189_116 =10'b0;

   // m189_117 = W*in
   wire signed [9:0] m189_117;
   assign m189_117 =10'b0;

   // m190_1 = W*in
   wire signed [9:0] m190_1;
   assign m190_1 =10'b0;

   // m190_2 = W*in
   wire signed [9:0] m190_2;
   assign m190_2 =10'b0;

   // m190_3 = W*in
   wire signed [9:0] m190_3;
   assign m190_3 =10'b0;

   // m190_4 = W*in
   wire signed [9:0] m190_4;
   assign m190_4 =10'b0;

   // m190_5 = W*in
   wire signed [9:0] m190_5;
   assign m190_5 =10'b0;

   // m190_6 = W*in
   wire signed [9:0] m190_6;
   assign m190_6 =10'b0;

   // m190_7 = W*in
   wire signed [9:0] m190_7;
   assign m190_7 =10'b0;

   // m190_8 = W*in
   wire signed [9:0] m190_8;
   assign m190_8 =10'b0;

   // m190_9 = W*in
   wire signed [9:0] m190_9;
   assign m190_9 =10'b0;

   // m190_10 = W*in
   wire signed [9:0] m190_10;
   assign m190_10 =10'b0;

   // m190_11 = W*in
   wire signed [9:0] m190_11;
   assign m190_11 =10'b0;

   // m190_12 = W*in
   wire signed [9:0] m190_12;
   assign m190_12 =10'b0;

   // m190_13 = W*in
   wire signed [9:0] m190_13;
   assign m190_13 =10'b0;

   // m190_14 = W*in
   wire signed [9:0] m190_14;
   assign m190_14 =10'b0;

   // m190_15 = W*in
   wire signed [9:0] m190_15;
   assign m190_15 =10'b0;

   // m190_16 = W*in
   wire signed [9:0] m190_16;
   assign m190_16 =10'b0;

   // m190_17 = W*in
   wire signed [9:0] m190_17;
   assign m190_17 =10'b0;

   // m190_18 = W*in
   wire signed [9:0] m190_18;
   assign m190_18 =10'b0;

   // m190_19 = W*in
   wire signed [9:0] m190_19;
   assign m190_19 =10'b0;

   // m190_20 = W*in
   wire signed [9:0] m190_20;
   assign m190_20 =10'b0;

   // m190_21 = W*in
   wire signed [9:0] m190_21;
   assign m190_21 =10'b0;

   // m190_22 = W*in
   wire signed [9:0] m190_22;
   assign m190_22 ={ {5{in190[5]}} , in190[5:1] };

   // m190_23 = W*in
   wire signed [9:0] m190_23;
   assign m190_23 ={ {5{in190[5]}} , in190[5:1] };

   // m190_24 = W*in
   wire signed [9:0] m190_24;
   assign m190_24 =10'b0;

   // m190_25 = W*in
   wire signed [9:0] m190_25;
   assign m190_25 =10'b0;

   // m190_26 = W*in
   wire signed [9:0] m190_26;
   assign m190_26 =10'b0;

   // m190_27 = W*in
   wire signed [9:0] m190_27;
   assign m190_27 ={ {5{in190[5]}} , in190[5:1] };

   // m190_28 = W*in
   wire signed [9:0] m190_28;
   assign m190_28 =10'b0;

   // m190_29 = W*in
   wire signed [9:0] m190_29;
   assign m190_29 =10'b0;

   // m190_30 = W*in
   wire signed [9:0] m190_30;
   assign m190_30 =10'b0;

   // m190_31 = W*in
   wire signed [9:0] m190_31;
   assign m190_31 =10'b0;

   // m190_32 = W*in
   wire signed [9:0] m190_32;
   assign m190_32 =10'b0;

   // m190_33 = W*in
   wire signed [9:0] m190_33;
   assign m190_33 =10'b0;

   // m190_34 = W*in
   wire signed [9:0] m190_34;
   assign m190_34 =10'b0;

   // m190_35 = W*in
   wire signed [9:0] m190_35;
   assign m190_35 =10'b0;

   // m190_36 = W*in
   wire signed [9:0] m190_36;
   assign m190_36 =10'b0;

   // m190_37 = W*in
   wire signed [9:0] m190_37;
   assign m190_37 =10'b0;

   // m190_38 = W*in
   wire signed [9:0] m190_38;
   assign m190_38 =10'b0;

   // m190_39 = W*in
   wire signed [9:0] m190_39;
   assign m190_39 =10'b0;

   // m190_40 = W*in
   wire signed [9:0] m190_40;
   assign m190_40 =10'b0;

   // m190_41 = W*in
   wire signed [9:0] m190_41;
   assign m190_41 =10'b0;

   // m190_42 = W*in
   wire signed [9:0] m190_42;
   assign m190_42 =10'b0;

   // m190_43 = W*in
   wire signed [9:0] m190_43;
   assign m190_43 =10'b0;

   // m190_44 = W*in
   wire signed [9:0] m190_44;
   assign m190_44 =10'b0;

   // m190_45 = W*in
   wire signed [9:0] m190_45;
   assign m190_45 =10'b0;

   // m190_46 = W*in
   wire signed [9:0] m190_46;
   assign m190_46 =10'b0;

   // m190_47 = W*in
   wire signed [9:0] m190_47;
   assign m190_47 =10'b0;

   // m190_48 = W*in
   wire signed [9:0] m190_48;
   assign m190_48 =10'b0;

   // m190_49 = W*in
   wire signed [9:0] m190_49;
   assign m190_49 =10'b0;

   // m190_50 = W*in
   wire signed [9:0] m190_50;
   assign m190_50 =10'b0;

   // m190_51 = W*in
   wire signed [9:0] m190_51;
   assign m190_51 =10'b0;

   // m190_52 = W*in
   wire signed [9:0] m190_52;
   assign m190_52 =10'b0;

   // m190_53 = W*in
   wire signed [9:0] m190_53;
   assign m190_53 =10'b0;

   // m190_54 = W*in
   wire signed [9:0] m190_54;
   assign m190_54 =10'b0;

   // m190_55 = W*in
   wire signed [9:0] m190_55;
   assign m190_55 =10'b0;

   // m190_56 = W*in
   wire signed [9:0] m190_56;
   assign m190_56 =10'b0;

   // m190_57 = W*in
   wire signed [9:0] m190_57;
   assign m190_57 =10'b0;

   // m190_58 = W*in
   wire signed [9:0] m190_58;
   assign m190_58 =10'b0;

   // m190_59 = W*in
   wire signed [9:0] m190_59;
   assign m190_59 =10'b0;

   // m190_60 = W*in
   wire signed [9:0] m190_60;
   assign m190_60 =10'b0;

   // m190_61 = W*in
   wire signed [9:0] m190_61;
   assign m190_61 =10'b0;

   // m190_62 = W*in
   wire signed [9:0] m190_62;
   assign m190_62 =10'b0;

   // m190_63 = W*in
   wire signed [9:0] m190_63;
   assign m190_63 =10'b0;

   // m190_64 = W*in
   wire signed [9:0] m190_64;
   assign m190_64 =10'b0;

   // m190_65 = W*in
   wire signed [9:0] m190_65;
   assign m190_65 =10'b0;

   // m190_66 = W*in
   wire signed [9:0] m190_66;
   assign m190_66 ={ {5{neg190[5]}} , neg190[5:1] };

   // m190_67 = W*in
   wire signed [9:0] m190_67;
   assign m190_67 =10'b0;

   // m190_68 = W*in
   wire signed [9:0] m190_68;
   assign m190_68 =10'b0;

   // m190_69 = W*in
   wire signed [9:0] m190_69;
   assign m190_69 =10'b0;

   // m190_70 = W*in
   wire signed [9:0] m190_70;
   assign m190_70 ={ {5{neg190[5]}} , neg190[5:1] };

   // m190_71 = W*in
   wire signed [9:0] m190_71;
   assign m190_71 =10'b0;

   // m190_72 = W*in
   wire signed [9:0] m190_72;
   assign m190_72 =10'b0;

   // m190_73 = W*in
   wire signed [9:0] m190_73;
   assign m190_73 =10'b0;

   // m190_74 = W*in
   wire signed [9:0] m190_74;
   assign m190_74 =10'b0;

   // m190_75 = W*in
   wire signed [9:0] m190_75;
   assign m190_75 =10'b0;

   // m190_76 = W*in
   wire signed [9:0] m190_76;
   assign m190_76 =10'b0;

   // m190_77 = W*in
   wire signed [9:0] m190_77;
   assign m190_77 =10'b0;

   // m190_78 = W*in
   wire signed [9:0] m190_78;
   assign m190_78 =10'b0;

   // m190_79 = W*in
   wire signed [9:0] m190_79;
   assign m190_79 =10'b0;

   // m190_80 = W*in
   wire signed [9:0] m190_80;
   assign m190_80 =10'b0;

   // m190_81 = W*in
   wire signed [9:0] m190_81;
   assign m190_81 =10'b0;

   // m190_82 = W*in
   wire signed [9:0] m190_82;
   assign m190_82 =10'b0;

   // m190_83 = W*in
   wire signed [9:0] m190_83;
   assign m190_83 =10'b0;

   // m190_84 = W*in
   wire signed [9:0] m190_84;
   assign m190_84 =10'b0;

   // m190_85 = W*in
   wire signed [9:0] m190_85;
   assign m190_85 =10'b0;

   // m190_86 = W*in
   wire signed [9:0] m190_86;
   assign m190_86 =10'b0;

   // m190_87 = W*in
   wire signed [9:0] m190_87;
   assign m190_87 =10'b0;

   // m190_88 = W*in
   wire signed [9:0] m190_88;
   assign m190_88 =10'b0;

   // m190_89 = W*in
   wire signed [9:0] m190_89;
   assign m190_89 =10'b0;

   // m190_90 = W*in
   wire signed [9:0] m190_90;
   assign m190_90 =10'b0;

   // m190_91 = W*in
   wire signed [9:0] m190_91;
   assign m190_91 =10'b0;

   // m190_92 = W*in
   wire signed [9:0] m190_92;
   assign m190_92 ={ {4{neg190[5]}} , neg190[5:0] };

   // m190_93 = W*in
   wire signed [9:0] m190_93;
   assign m190_93 =10'b0;

   // m190_94 = W*in
   wire signed [9:0] m190_94;
   assign m190_94 =10'b0;

   // m190_95 = W*in
   wire signed [9:0] m190_95;
   assign m190_95 =10'b0;

   // m190_96 = W*in
   wire signed [9:0] m190_96;
   assign m190_96 =10'b0;

   // m190_97 = W*in
   wire signed [9:0] m190_97;
   assign m190_97 =10'b0;

   // m190_98 = W*in
   wire signed [9:0] m190_98;
   assign m190_98 =10'b0;

   // m190_99 = W*in
   wire signed [9:0] m190_99;
   assign m190_99 =10'b0;

   // m190_100 = W*in
   wire signed [9:0] m190_100;
   assign m190_100 =10'b0;

   // m190_101 = W*in
   wire signed [9:0] m190_101;
   assign m190_101 =10'b0;

   // m190_102 = W*in
   wire signed [9:0] m190_102;
   assign m190_102 =10'b0;

   // m190_103 = W*in
   wire signed [9:0] m190_103;
   assign m190_103 =10'b0;

   // m190_104 = W*in
   wire signed [9:0] m190_104;
   assign m190_104 =10'b0;

   // m190_105 = W*in
   wire signed [9:0] m190_105;
   assign m190_105 =10'b0;

   // m190_106 = W*in
   wire signed [9:0] m190_106;
   assign m190_106 =10'b0;

   // m190_107 = W*in
   wire signed [9:0] m190_107;
   assign m190_107 =10'b0;

   // m190_108 = W*in
   wire signed [9:0] m190_108;
   assign m190_108 ={ {5{neg190[5]}} , neg190[5:1] };

   // m190_109 = W*in
   wire signed [9:0] m190_109;
   assign m190_109 =10'b0;

   // m190_110 = W*in
   wire signed [9:0] m190_110;
   assign m190_110 =10'b0;

   // m190_111 = W*in
   wire signed [9:0] m190_111;
   assign m190_111 =10'b0;

   // m190_112 = W*in
   wire signed [9:0] m190_112;
   assign m190_112 =10'b0;

   // m190_113 = W*in
   wire signed [9:0] m190_113;
   assign m190_113 =10'b0;

   // m190_114 = W*in
   wire signed [9:0] m190_114;
   assign m190_114 =10'b0;

   // m190_115 = W*in
   wire signed [9:0] m190_115;
   assign m190_115 ={ {5{neg190[5]}} , neg190[5:1] };

   // m190_116 = W*in
   wire signed [9:0] m190_116;
   assign m190_116 =10'b0;

   // m190_117 = W*in
   wire signed [9:0] m190_117;
   assign m190_117 =10'b0;

   // m191_1 = W*in
   wire signed [9:0] m191_1;
   assign m191_1 =10'b0;

   // m191_2 = W*in
   wire signed [9:0] m191_2;
   assign m191_2 =10'b0;

   // m191_3 = W*in
   wire signed [9:0] m191_3;
   assign m191_3 =10'b0;

   // m191_4 = W*in
   wire signed [9:0] m191_4;
   assign m191_4 =10'b0;

   // m191_5 = W*in
   wire signed [9:0] m191_5;
   assign m191_5 =10'b0;

   // m191_6 = W*in
   wire signed [9:0] m191_6;
   assign m191_6 =10'b0;

   // m191_7 = W*in
   wire signed [9:0] m191_7;
   assign m191_7 =10'b0;

   // m191_8 = W*in
   wire signed [9:0] m191_8;
   assign m191_8 =10'b0;

   // m191_9 = W*in
   wire signed [9:0] m191_9;
   assign m191_9 =10'b0;

   // m191_10 = W*in
   wire signed [9:0] m191_10;
   assign m191_10 =10'b0;

   // m191_11 = W*in
   wire signed [9:0] m191_11;
   assign m191_11 =10'b0;

   // m191_12 = W*in
   wire signed [9:0] m191_12;
   assign m191_12 =10'b0;

   // m191_13 = W*in
   wire signed [9:0] m191_13;
   assign m191_13 =10'b0;

   // m191_14 = W*in
   wire signed [9:0] m191_14;
   assign m191_14 =10'b0;

   // m191_15 = W*in
   wire signed [9:0] m191_15;
   assign m191_15 =10'b0;

   // m191_16 = W*in
   wire signed [9:0] m191_16;
   assign m191_16 =10'b0;

   // m191_17 = W*in
   wire signed [9:0] m191_17;
   assign m191_17 =10'b0;

   // m191_18 = W*in
   wire signed [9:0] m191_18;
   assign m191_18 ={ {5{neg191[5]}} , neg191[5:1] };

   // m191_19 = W*in
   wire signed [9:0] m191_19;
   assign m191_19 =10'b0;

   // m191_20 = W*in
   wire signed [9:0] m191_20;
   assign m191_20 =10'b0;

   // m191_21 = W*in
   wire signed [9:0] m191_21;
   assign m191_21 =10'b0;

   // m191_22 = W*in
   wire signed [9:0] m191_22;
   assign m191_22 ={ {5{in191[5]}} , in191[5:1] };

   // m191_23 = W*in
   wire signed [9:0] m191_23;
   assign m191_23 ={ {5{in191[5]}} , in191[5:1] };

   // m191_24 = W*in
   wire signed [9:0] m191_24;
   assign m191_24 =10'b0;

   // m191_25 = W*in
   wire signed [9:0] m191_25;
   assign m191_25 =10'b0;

   // m191_26 = W*in
   wire signed [9:0] m191_26;
   assign m191_26 ={ {5{neg191[5]}} , neg191[5:1] };

   // m191_27 = W*in
   wire signed [9:0] m191_27;
   assign m191_27 =10'b0;

   // m191_28 = W*in
   wire signed [9:0] m191_28;
   assign m191_28 =10'b0;

   // m191_29 = W*in
   wire signed [9:0] m191_29;
   assign m191_29 =10'b0;

   // m191_30 = W*in
   wire signed [9:0] m191_30;
   assign m191_30 =10'b0;

   // m191_31 = W*in
   wire signed [9:0] m191_31;
   assign m191_31 =10'b0;

   // m191_32 = W*in
   wire signed [9:0] m191_32;
   assign m191_32 =10'b0;

   // m191_33 = W*in
   wire signed [9:0] m191_33;
   assign m191_33 =10'b0;

   // m191_34 = W*in
   wire signed [9:0] m191_34;
   assign m191_34 =10'b0;

   // m191_35 = W*in
   wire signed [9:0] m191_35;
   assign m191_35 =10'b0;

   // m191_36 = W*in
   wire signed [9:0] m191_36;
   assign m191_36 =10'b0;

   // m191_37 = W*in
   wire signed [9:0] m191_37;
   assign m191_37 =10'b0;

   // m191_38 = W*in
   wire signed [9:0] m191_38;
   assign m191_38 =10'b0;

   // m191_39 = W*in
   wire signed [9:0] m191_39;
   assign m191_39 =10'b0;

   // m191_40 = W*in
   wire signed [9:0] m191_40;
   assign m191_40 =10'b0;

   // m191_41 = W*in
   wire signed [9:0] m191_41;
   assign m191_41 =10'b0;

   // m191_42 = W*in
   wire signed [9:0] m191_42;
   assign m191_42 =10'b0;

   // m191_43 = W*in
   wire signed [9:0] m191_43;
   assign m191_43 =10'b0;

   // m191_44 = W*in
   wire signed [9:0] m191_44;
   assign m191_44 =10'b0;

   // m191_45 = W*in
   wire signed [9:0] m191_45;
   assign m191_45 =10'b0;

   // m191_46 = W*in
   wire signed [9:0] m191_46;
   assign m191_46 =10'b0;

   // m191_47 = W*in
   wire signed [9:0] m191_47;
   assign m191_47 =10'b0;

   // m191_48 = W*in
   wire signed [9:0] m191_48;
   assign m191_48 =10'b0;

   // m191_49 = W*in
   wire signed [9:0] m191_49;
   assign m191_49 =10'b0;

   // m191_50 = W*in
   wire signed [9:0] m191_50;
   assign m191_50 =10'b0;

   // m191_51 = W*in
   wire signed [9:0] m191_51;
   assign m191_51 =10'b0;

   // m191_52 = W*in
   wire signed [9:0] m191_52;
   assign m191_52 =10'b0;

   // m191_53 = W*in
   wire signed [9:0] m191_53;
   assign m191_53 =10'b0;

   // m191_54 = W*in
   wire signed [9:0] m191_54;
   assign m191_54 =10'b0;

   // m191_55 = W*in
   wire signed [9:0] m191_55;
   assign m191_55 =10'b0;

   // m191_56 = W*in
   wire signed [9:0] m191_56;
   assign m191_56 =10'b0;

   // m191_57 = W*in
   wire signed [9:0] m191_57;
   assign m191_57 =10'b0;

   // m191_58 = W*in
   wire signed [9:0] m191_58;
   assign m191_58 =10'b0;

   // m191_59 = W*in
   wire signed [9:0] m191_59;
   assign m191_59 =10'b0;

   // m191_60 = W*in
   wire signed [9:0] m191_60;
   assign m191_60 =10'b0;

   // m191_61 = W*in
   wire signed [9:0] m191_61;
   assign m191_61 =10'b0;

   // m191_62 = W*in
   wire signed [9:0] m191_62;
   assign m191_62 =10'b0;

   // m191_63 = W*in
   wire signed [9:0] m191_63;
   assign m191_63 =10'b0;

   // m191_64 = W*in
   wire signed [9:0] m191_64;
   assign m191_64 ={ {5{neg191[5]}} , neg191[5:1] };

   // m191_65 = W*in
   wire signed [9:0] m191_65;
   assign m191_65 =10'b0;

   // m191_66 = W*in
   wire signed [9:0] m191_66;
   assign m191_66 ={ {5{neg191[5]}} , neg191[5:1] };

   // m191_67 = W*in
   wire signed [9:0] m191_67;
   assign m191_67 =10'b0;

   // m191_68 = W*in
   wire signed [9:0] m191_68;
   assign m191_68 =10'b0;

   // m191_69 = W*in
   wire signed [9:0] m191_69;
   assign m191_69 =10'b0;

   // m191_70 = W*in
   wire signed [9:0] m191_70;
   assign m191_70 =10'b0;

   // m191_71 = W*in
   wire signed [9:0] m191_71;
   assign m191_71 =10'b0;

   // m191_72 = W*in
   wire signed [9:0] m191_72;
   assign m191_72 =10'b0;

   // m191_73 = W*in
   wire signed [9:0] m191_73;
   assign m191_73 =10'b0;

   // m191_74 = W*in
   wire signed [9:0] m191_74;
   assign m191_74 =10'b0;

   // m191_75 = W*in
   wire signed [9:0] m191_75;
   assign m191_75 =10'b0;

   // m191_76 = W*in
   wire signed [9:0] m191_76;
   assign m191_76 =10'b0;

   // m191_77 = W*in
   wire signed [9:0] m191_77;
   assign m191_77 =10'b0;

   // m191_78 = W*in
   wire signed [9:0] m191_78;
   assign m191_78 =10'b0;

   // m191_79 = W*in
   wire signed [9:0] m191_79;
   assign m191_79 =10'b0;

   // m191_80 = W*in
   wire signed [9:0] m191_80;
   assign m191_80 =10'b0;

   // m191_81 = W*in
   wire signed [9:0] m191_81;
   assign m191_81 =10'b0;

   // m191_82 = W*in
   wire signed [9:0] m191_82;
   assign m191_82 =10'b0;

   // m191_83 = W*in
   wire signed [9:0] m191_83;
   assign m191_83 =10'b0;

   // m191_84 = W*in
   wire signed [9:0] m191_84;
   assign m191_84 =10'b0;

   // m191_85 = W*in
   wire signed [9:0] m191_85;
   assign m191_85 =10'b0;

   // m191_86 = W*in
   wire signed [9:0] m191_86;
   assign m191_86 =10'b0;

   // m191_87 = W*in
   wire signed [9:0] m191_87;
   assign m191_87 =10'b0;

   // m191_88 = W*in
   wire signed [9:0] m191_88;
   assign m191_88 =10'b0;

   // m191_89 = W*in
   wire signed [9:0] m191_89;
   assign m191_89 =10'b0;

   // m191_90 = W*in
   wire signed [9:0] m191_90;
   assign m191_90 =10'b0;

   // m191_91 = W*in
   wire signed [9:0] m191_91;
   assign m191_91 =10'b0;

   // m191_92 = W*in
   wire signed [9:0] m191_92;
   assign m191_92 =10'b0;

   // m191_93 = W*in
   wire signed [9:0] m191_93;
   assign m191_93 =10'b0;

   // m191_94 = W*in
   wire signed [9:0] m191_94;
   assign m191_94 =10'b0;

   // m191_95 = W*in
   wire signed [9:0] m191_95;
   assign m191_95 =10'b0;

   // m191_96 = W*in
   wire signed [9:0] m191_96;
   assign m191_96 =10'b0;

   // m191_97 = W*in
   wire signed [9:0] m191_97;
   assign m191_97 =10'b0;

   // m191_98 = W*in
   wire signed [9:0] m191_98;
   assign m191_98 =10'b0;

   // m191_99 = W*in
   wire signed [9:0] m191_99;
   assign m191_99 =10'b0;

   // m191_100 = W*in
   wire signed [9:0] m191_100;
   assign m191_100 =10'b0;

   // m191_101 = W*in
   wire signed [9:0] m191_101;
   assign m191_101 =10'b0;

   // m191_102 = W*in
   wire signed [9:0] m191_102;
   assign m191_102 =10'b0;

   // m191_103 = W*in
   wire signed [9:0] m191_103;
   assign m191_103 =10'b0;

   // m191_104 = W*in
   wire signed [9:0] m191_104;
   assign m191_104 =10'b0;

   // m191_105 = W*in
   wire signed [9:0] m191_105;
   assign m191_105 =10'b0;

   // m191_106 = W*in
   wire signed [9:0] m191_106;
   assign m191_106 =10'b0;

   // m191_107 = W*in
   wire signed [9:0] m191_107;
   assign m191_107 =10'b0;

   // m191_108 = W*in
   wire signed [9:0] m191_108;
   assign m191_108 =10'b0;

   // m191_109 = W*in
   wire signed [9:0] m191_109;
   assign m191_109 ={ {5{in191[5]}} , in191[5:1] };

   // m191_110 = W*in
   wire signed [9:0] m191_110;
   assign m191_110 =10'b0;

   // m191_111 = W*in
   wire signed [9:0] m191_111;
   assign m191_111 =10'b0;

   // m191_112 = W*in
   wire signed [9:0] m191_112;
   assign m191_112 =10'b0;

   // m191_113 = W*in
   wire signed [9:0] m191_113;
   assign m191_113 =10'b0;

   // m191_114 = W*in
   wire signed [9:0] m191_114;
   assign m191_114 =10'b0;

   // m191_115 = W*in
   wire signed [9:0] m191_115;
   assign m191_115 =10'b0;

   // m191_116 = W*in
   wire signed [9:0] m191_116;
   assign m191_116 =10'b0;

   // m191_117 = W*in
   wire signed [9:0] m191_117;
   assign m191_117 =10'b0;

   // m192_1 = W*in
   wire signed [9:0] m192_1;
   assign m192_1 =10'b0;

   // m192_2 = W*in
   wire signed [9:0] m192_2;
   assign m192_2 =10'b0;

   // m192_3 = W*in
   wire signed [9:0] m192_3;
   assign m192_3 =10'b0;

   // m192_4 = W*in
   wire signed [9:0] m192_4;
   assign m192_4 =10'b0;

   // m192_5 = W*in
   wire signed [9:0] m192_5;
   assign m192_5 =10'b0;

   // m192_6 = W*in
   wire signed [9:0] m192_6;
   assign m192_6 =10'b0;

   // m192_7 = W*in
   wire signed [9:0] m192_7;
   assign m192_7 =10'b0;

   // m192_8 = W*in
   wire signed [9:0] m192_8;
   assign m192_8 =10'b0;

   // m192_9 = W*in
   wire signed [9:0] m192_9;
   assign m192_9 =10'b0;

   // m192_10 = W*in
   wire signed [9:0] m192_10;
   assign m192_10 =10'b0;

   // m192_11 = W*in
   wire signed [9:0] m192_11;
   assign m192_11 =10'b0;

   // m192_12 = W*in
   wire signed [9:0] m192_12;
   assign m192_12 =10'b0;

   // m192_13 = W*in
   wire signed [9:0] m192_13;
   assign m192_13 =10'b0;

   // m192_14 = W*in
   wire signed [9:0] m192_14;
   assign m192_14 =10'b0;

   // m192_15 = W*in
   wire signed [9:0] m192_15;
   assign m192_15 =10'b0;

   // m192_16 = W*in
   wire signed [9:0] m192_16;
   assign m192_16 =10'b0;

   // m192_17 = W*in
   wire signed [9:0] m192_17;
   assign m192_17 =10'b0;

   // m192_18 = W*in
   wire signed [9:0] m192_18;
   assign m192_18 ={ {5{in192[5]}} , in192[5:1] };

   // m192_19 = W*in
   wire signed [9:0] m192_19;
   assign m192_19 ={ {5{neg192[5]}} , neg192[5:1] };

   // m192_20 = W*in
   wire signed [9:0] m192_20;
   assign m192_20 =10'b0;

   // m192_21 = W*in
   wire signed [9:0] m192_21;
   assign m192_21 =10'b0;

   // m192_22 = W*in
   wire signed [9:0] m192_22;
   assign m192_22 =10'b0;

   // m192_23 = W*in
   wire signed [9:0] m192_23;
   assign m192_23 =10'b0;

   // m192_24 = W*in
   wire signed [9:0] m192_24;
   assign m192_24 =10'b0;

   // m192_25 = W*in
   wire signed [9:0] m192_25;
   assign m192_25 =10'b0;

   // m192_26 = W*in
   wire signed [9:0] m192_26;
   assign m192_26 ={ {5{in192[5]}} , in192[5:1] };

   // m192_27 = W*in
   wire signed [9:0] m192_27;
   assign m192_27 =10'b0;

   // m192_28 = W*in
   wire signed [9:0] m192_28;
   assign m192_28 =10'b0;

   // m192_29 = W*in
   wire signed [9:0] m192_29;
   assign m192_29 =10'b0;

   // m192_30 = W*in
   wire signed [9:0] m192_30;
   assign m192_30 =10'b0;

   // m192_31 = W*in
   wire signed [9:0] m192_31;
   assign m192_31 =10'b0;

   // m192_32 = W*in
   wire signed [9:0] m192_32;
   assign m192_32 =10'b0;

   // m192_33 = W*in
   wire signed [9:0] m192_33;
   assign m192_33 =10'b0;

   // m192_34 = W*in
   wire signed [9:0] m192_34;
   assign m192_34 =10'b0;

   // m192_35 = W*in
   wire signed [9:0] m192_35;
   assign m192_35 =10'b0;

   // m192_36 = W*in
   wire signed [9:0] m192_36;
   assign m192_36 =10'b0;

   // m192_37 = W*in
   wire signed [9:0] m192_37;
   assign m192_37 =10'b0;

   // m192_38 = W*in
   wire signed [9:0] m192_38;
   assign m192_38 =10'b0;

   // m192_39 = W*in
   wire signed [9:0] m192_39;
   assign m192_39 =10'b0;

   // m192_40 = W*in
   wire signed [9:0] m192_40;
   assign m192_40 =10'b0;

   // m192_41 = W*in
   wire signed [9:0] m192_41;
   assign m192_41 =10'b0;

   // m192_42 = W*in
   wire signed [9:0] m192_42;
   assign m192_42 =10'b0;

   // m192_43 = W*in
   wire signed [9:0] m192_43;
   assign m192_43 =10'b0;

   // m192_44 = W*in
   wire signed [9:0] m192_44;
   assign m192_44 =10'b0;

   // m192_45 = W*in
   wire signed [9:0] m192_45;
   assign m192_45 =10'b0;

   // m192_46 = W*in
   wire signed [9:0] m192_46;
   assign m192_46 =10'b0;

   // m192_47 = W*in
   wire signed [9:0] m192_47;
   assign m192_47 =10'b0;

   // m192_48 = W*in
   wire signed [9:0] m192_48;
   assign m192_48 =10'b0;

   // m192_49 = W*in
   wire signed [9:0] m192_49;
   assign m192_49 =10'b0;

   // m192_50 = W*in
   wire signed [9:0] m192_50;
   assign m192_50 =10'b0;

   // m192_51 = W*in
   wire signed [9:0] m192_51;
   assign m192_51 =10'b0;

   // m192_52 = W*in
   wire signed [9:0] m192_52;
   assign m192_52 =10'b0;

   // m192_53 = W*in
   wire signed [9:0] m192_53;
   assign m192_53 =10'b0;

   // m192_54 = W*in
   wire signed [9:0] m192_54;
   assign m192_54 =10'b0;

   // m192_55 = W*in
   wire signed [9:0] m192_55;
   assign m192_55 =10'b0;

   // m192_56 = W*in
   wire signed [9:0] m192_56;
   assign m192_56 =10'b0;

   // m192_57 = W*in
   wire signed [9:0] m192_57;
   assign m192_57 =10'b0;

   // m192_58 = W*in
   wire signed [9:0] m192_58;
   assign m192_58 =10'b0;

   // m192_59 = W*in
   wire signed [9:0] m192_59;
   assign m192_59 =10'b0;

   // m192_60 = W*in
   wire signed [9:0] m192_60;
   assign m192_60 =10'b0;

   // m192_61 = W*in
   wire signed [9:0] m192_61;
   assign m192_61 =10'b0;

   // m192_62 = W*in
   wire signed [9:0] m192_62;
   assign m192_62 =10'b0;

   // m192_63 = W*in
   wire signed [9:0] m192_63;
   assign m192_63 =10'b0;

   // m192_64 = W*in
   wire signed [9:0] m192_64;
   assign m192_64 =10'b0;

   // m192_65 = W*in
   wire signed [9:0] m192_65;
   assign m192_65 =10'b0;

   // m192_66 = W*in
   wire signed [9:0] m192_66;
   assign m192_66 =10'b0;

   // m192_67 = W*in
   wire signed [9:0] m192_67;
   assign m192_67 =10'b0;

   // m192_68 = W*in
   wire signed [9:0] m192_68;
   assign m192_68 =10'b0;

   // m192_69 = W*in
   wire signed [9:0] m192_69;
   assign m192_69 =10'b0;

   // m192_70 = W*in
   wire signed [9:0] m192_70;
   assign m192_70 =10'b0;

   // m192_71 = W*in
   wire signed [9:0] m192_71;
   assign m192_71 =10'b0;

   // m192_72 = W*in
   wire signed [9:0] m192_72;
   assign m192_72 ={ {5{in192[5]}} , in192[5:1] };

   // m192_73 = W*in
   wire signed [9:0] m192_73;
   assign m192_73 =10'b0;

   // m192_74 = W*in
   wire signed [9:0] m192_74;
   assign m192_74 =10'b0;

   // m192_75 = W*in
   wire signed [9:0] m192_75;
   assign m192_75 =10'b0;

   // m192_76 = W*in
   wire signed [9:0] m192_76;
   assign m192_76 =10'b0;

   // m192_77 = W*in
   wire signed [9:0] m192_77;
   assign m192_77 =10'b0;

   // m192_78 = W*in
   wire signed [9:0] m192_78;
   assign m192_78 ={ {5{in192[5]}} , in192[5:1] };

   // m192_79 = W*in
   wire signed [9:0] m192_79;
   assign m192_79 =10'b0;

   // m192_80 = W*in
   wire signed [9:0] m192_80;
   assign m192_80 =10'b0;

   // m192_81 = W*in
   wire signed [9:0] m192_81;
   assign m192_81 =10'b0;

   // m192_82 = W*in
   wire signed [9:0] m192_82;
   assign m192_82 =10'b0;

   // m192_83 = W*in
   wire signed [9:0] m192_83;
   assign m192_83 =10'b0;

   // m192_84 = W*in
   wire signed [9:0] m192_84;
   assign m192_84 =10'b0;

   // m192_85 = W*in
   wire signed [9:0] m192_85;
   assign m192_85 =10'b0;

   // m192_86 = W*in
   wire signed [9:0] m192_86;
   assign m192_86 =10'b0;

   // m192_87 = W*in
   wire signed [9:0] m192_87;
   assign m192_87 =10'b0;

   // m192_88 = W*in
   wire signed [9:0] m192_88;
   assign m192_88 =10'b0;

   // m192_89 = W*in
   wire signed [9:0] m192_89;
   assign m192_89 =10'b0;

   // m192_90 = W*in
   wire signed [9:0] m192_90;
   assign m192_90 =10'b0;

   // m192_91 = W*in
   wire signed [9:0] m192_91;
   assign m192_91 =10'b0;

   // m192_92 = W*in
   wire signed [9:0] m192_92;
   assign m192_92 =10'b0;

   // m192_93 = W*in
   wire signed [9:0] m192_93;
   assign m192_93 =10'b0;

   // m192_94 = W*in
   wire signed [9:0] m192_94;
   assign m192_94 =10'b0;

   // m192_95 = W*in
   wire signed [9:0] m192_95;
   assign m192_95 =10'b0;

   // m192_96 = W*in
   wire signed [9:0] m192_96;
   assign m192_96 =10'b0;

   // m192_97 = W*in
   wire signed [9:0] m192_97;
   assign m192_97 =10'b0;

   // m192_98 = W*in
   wire signed [9:0] m192_98;
   assign m192_98 =10'b0;

   // m192_99 = W*in
   wire signed [9:0] m192_99;
   assign m192_99 =10'b0;

   // m192_100 = W*in
   wire signed [9:0] m192_100;
   assign m192_100 =10'b0;

   // m192_101 = W*in
   wire signed [9:0] m192_101;
   assign m192_101 =10'b0;

   // m192_102 = W*in
   wire signed [9:0] m192_102;
   assign m192_102 =10'b0;

   // m192_103 = W*in
   wire signed [9:0] m192_103;
   assign m192_103 =10'b0;

   // m192_104 = W*in
   wire signed [9:0] m192_104;
   assign m192_104 =10'b0;

   // m192_105 = W*in
   wire signed [9:0] m192_105;
   assign m192_105 =10'b0;

   // m192_106 = W*in
   wire signed [9:0] m192_106;
   assign m192_106 =10'b0;

   // m192_107 = W*in
   wire signed [9:0] m192_107;
   assign m192_107 =10'b0;

   // m192_108 = W*in
   wire signed [9:0] m192_108;
   assign m192_108 =10'b0;

   // m192_109 = W*in
   wire signed [9:0] m192_109;
   assign m192_109 =10'b0;

   // m192_110 = W*in
   wire signed [9:0] m192_110;
   assign m192_110 =10'b0;

   // m192_111 = W*in
   wire signed [9:0] m192_111;
   assign m192_111 =10'b0;

   // m192_112 = W*in
   wire signed [9:0] m192_112;
   assign m192_112 =10'b0;

   // m192_113 = W*in
   wire signed [9:0] m192_113;
   assign m192_113 =10'b0;

   // m192_114 = W*in
   wire signed [9:0] m192_114;
   assign m192_114 =10'b0;

   // m192_115 = W*in
   wire signed [9:0] m192_115;
   assign m192_115 =10'b0;

   // m192_116 = W*in
   wire signed [9:0] m192_116;
   assign m192_116 =10'b0;

   // m192_117 = W*in
   wire signed [9:0] m192_117;
   assign m192_117 =10'b0;

   // m193_1 = W*in
   wire signed [9:0] m193_1;
   assign m193_1 =10'b0;

   // m193_2 = W*in
   wire signed [9:0] m193_2;
   assign m193_2 =10'b0;

   // m193_3 = W*in
   wire signed [9:0] m193_3;
   assign m193_3 =10'b0;

   // m193_4 = W*in
   wire signed [9:0] m193_4;
   assign m193_4 =10'b0;

   // m193_5 = W*in
   wire signed [9:0] m193_5;
   assign m193_5 =10'b0;

   // m193_6 = W*in
   wire signed [9:0] m193_6;
   assign m193_6 =10'b0;

   // m193_7 = W*in
   wire signed [9:0] m193_7;
   assign m193_7 =10'b0;

   // m193_8 = W*in
   wire signed [9:0] m193_8;
   assign m193_8 =10'b0;

   // m193_9 = W*in
   wire signed [9:0] m193_9;
   assign m193_9 =10'b0;

   // m193_10 = W*in
   wire signed [9:0] m193_10;
   assign m193_10 =10'b0;

   // m193_11 = W*in
   wire signed [9:0] m193_11;
   assign m193_11 =10'b0;

   // m193_12 = W*in
   wire signed [9:0] m193_12;
   assign m193_12 =10'b0;

   // m193_13 = W*in
   wire signed [9:0] m193_13;
   assign m193_13 =10'b0;

   // m193_14 = W*in
   wire signed [9:0] m193_14;
   assign m193_14 =10'b0;

   // m193_15 = W*in
   wire signed [9:0] m193_15;
   assign m193_15 =10'b0;

   // m193_16 = W*in
   wire signed [9:0] m193_16;
   assign m193_16 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_17 = W*in
   wire signed [9:0] m193_17;
   assign m193_17 =10'b0;

   // m193_18 = W*in
   wire signed [9:0] m193_18;
   assign m193_18 ={ {4{in193[5]}} , in193[5:0] };

   // m193_19 = W*in
   wire signed [9:0] m193_19;
   assign m193_19 =10'b0;

   // m193_20 = W*in
   wire signed [9:0] m193_20;
   assign m193_20 =10'b0;

   // m193_21 = W*in
   wire signed [9:0] m193_21;
   assign m193_21 =10'b0;

   // m193_22 = W*in
   wire signed [9:0] m193_22;
   assign m193_22 =10'b0;

   // m193_23 = W*in
   wire signed [9:0] m193_23;
   assign m193_23 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_24 = W*in
   wire signed [9:0] m193_24;
   assign m193_24 =10'b0;

   // m193_25 = W*in
   wire signed [9:0] m193_25;
   assign m193_25 =10'b0;

   // m193_26 = W*in
   wire signed [9:0] m193_26;
   assign m193_26 ={ {4{in193[5]}} , in193[5:0] };

   // m193_27 = W*in
   wire signed [9:0] m193_27;
   assign m193_27 =10'b0;

   // m193_28 = W*in
   wire signed [9:0] m193_28;
   assign m193_28 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_29 = W*in
   wire signed [9:0] m193_29;
   assign m193_29 =10'b0;

   // m193_30 = W*in
   wire signed [9:0] m193_30;
   assign m193_30 =10'b0;

   // m193_31 = W*in
   wire signed [9:0] m193_31;
   assign m193_31 =10'b0;

   // m193_32 = W*in
   wire signed [9:0] m193_32;
   assign m193_32 =10'b0;

   // m193_33 = W*in
   wire signed [9:0] m193_33;
   assign m193_33 =10'b0;

   // m193_34 = W*in
   wire signed [9:0] m193_34;
   assign m193_34 =10'b0;

   // m193_35 = W*in
   wire signed [9:0] m193_35;
   assign m193_35 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_36 = W*in
   wire signed [9:0] m193_36;
   assign m193_36 =10'b0;

   // m193_37 = W*in
   wire signed [9:0] m193_37;
   assign m193_37 =10'b0;

   // m193_38 = W*in
   wire signed [9:0] m193_38;
   assign m193_38 =10'b0;

   // m193_39 = W*in
   wire signed [9:0] m193_39;
   assign m193_39 =10'b0;

   // m193_40 = W*in
   wire signed [9:0] m193_40;
   assign m193_40 =10'b0;

   // m193_41 = W*in
   wire signed [9:0] m193_41;
   assign m193_41 =10'b0;

   // m193_42 = W*in
   wire signed [9:0] m193_42;
   assign m193_42 =10'b0;

   // m193_43 = W*in
   wire signed [9:0] m193_43;
   assign m193_43 =10'b0;

   // m193_44 = W*in
   wire signed [9:0] m193_44;
   assign m193_44 =10'b0;

   // m193_45 = W*in
   wire signed [9:0] m193_45;
   assign m193_45 =10'b0;

   // m193_46 = W*in
   wire signed [9:0] m193_46;
   assign m193_46 =10'b0;

   // m193_47 = W*in
   wire signed [9:0] m193_47;
   assign m193_47 =10'b0;

   // m193_48 = W*in
   wire signed [9:0] m193_48;
   assign m193_48 =10'b0;

   // m193_49 = W*in
   wire signed [9:0] m193_49;
   assign m193_49 =10'b0;

   // m193_50 = W*in
   wire signed [9:0] m193_50;
   assign m193_50 =10'b0;

   // m193_51 = W*in
   wire signed [9:0] m193_51;
   assign m193_51 =10'b0;

   // m193_52 = W*in
   wire signed [9:0] m193_52;
   assign m193_52 =10'b0;

   // m193_53 = W*in
   wire signed [9:0] m193_53;
   assign m193_53 =10'b0;

   // m193_54 = W*in
   wire signed [9:0] m193_54;
   assign m193_54 =10'b0;

   // m193_55 = W*in
   wire signed [9:0] m193_55;
   assign m193_55 =10'b0;

   // m193_56 = W*in
   wire signed [9:0] m193_56;
   assign m193_56 =10'b0;

   // m193_57 = W*in
   wire signed [9:0] m193_57;
   assign m193_57 =10'b0;

   // m193_58 = W*in
   wire signed [9:0] m193_58;
   assign m193_58 =10'b0;

   // m193_59 = W*in
   wire signed [9:0] m193_59;
   assign m193_59 =10'b0;

   // m193_60 = W*in
   wire signed [9:0] m193_60;
   assign m193_60 =10'b0;

   // m193_61 = W*in
   wire signed [9:0] m193_61;
   assign m193_61 =10'b0;

   // m193_62 = W*in
   wire signed [9:0] m193_62;
   assign m193_62 =10'b0;

   // m193_63 = W*in
   wire signed [9:0] m193_63;
   assign m193_63 =10'b0;

   // m193_64 = W*in
   wire signed [9:0] m193_64;
   assign m193_64 =10'b0;

   // m193_65 = W*in
   wire signed [9:0] m193_65;
   assign m193_65 =10'b0;

   // m193_66 = W*in
   wire signed [9:0] m193_66;
   assign m193_66 =10'b0;

   // m193_67 = W*in
   wire signed [9:0] m193_67;
   assign m193_67 =10'b0;

   // m193_68 = W*in
   wire signed [9:0] m193_68;
   assign m193_68 =10'b0;

   // m193_69 = W*in
   wire signed [9:0] m193_69;
   assign m193_69 =10'b0;

   // m193_70 = W*in
   wire signed [9:0] m193_70;
   assign m193_70 =10'b0;

   // m193_71 = W*in
   wire signed [9:0] m193_71;
   assign m193_71 ={ {5{in193[5]}} , in193[5:1] };

   // m193_72 = W*in
   wire signed [9:0] m193_72;
   assign m193_72 =10'b0;

   // m193_73 = W*in
   wire signed [9:0] m193_73;
   assign m193_73 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_74 = W*in
   wire signed [9:0] m193_74;
   assign m193_74 =10'b0;

   // m193_75 = W*in
   wire signed [9:0] m193_75;
   assign m193_75 =10'b0;

   // m193_76 = W*in
   wire signed [9:0] m193_76;
   assign m193_76 =10'b0;

   // m193_77 = W*in
   wire signed [9:0] m193_77;
   assign m193_77 =10'b0;

   // m193_78 = W*in
   wire signed [9:0] m193_78;
   assign m193_78 ={ {5{in193[5]}} , in193[5:1] };

   // m193_79 = W*in
   wire signed [9:0] m193_79;
   assign m193_79 =10'b0;

   // m193_80 = W*in
   wire signed [9:0] m193_80;
   assign m193_80 =10'b0;

   // m193_81 = W*in
   wire signed [9:0] m193_81;
   assign m193_81 =10'b0;

   // m193_82 = W*in
   wire signed [9:0] m193_82;
   assign m193_82 =10'b0;

   // m193_83 = W*in
   wire signed [9:0] m193_83;
   assign m193_83 =10'b0;

   // m193_84 = W*in
   wire signed [9:0] m193_84;
   assign m193_84 =10'b0;

   // m193_85 = W*in
   wire signed [9:0] m193_85;
   assign m193_85 =10'b0;

   // m193_86 = W*in
   wire signed [9:0] m193_86;
   assign m193_86 =10'b0;

   // m193_87 = W*in
   wire signed [9:0] m193_87;
   assign m193_87 =10'b0;

   // m193_88 = W*in
   wire signed [9:0] m193_88;
   assign m193_88 =10'b0;

   // m193_89 = W*in
   wire signed [9:0] m193_89;
   assign m193_89 =10'b0;

   // m193_90 = W*in
   wire signed [9:0] m193_90;
   assign m193_90 =10'b0;

   // m193_91 = W*in
   wire signed [9:0] m193_91;
   assign m193_91 =10'b0;

   // m193_92 = W*in
   wire signed [9:0] m193_92;
   assign m193_92 ={ {4{in193[5]}} , in193[5:0] };

   // m193_93 = W*in
   wire signed [9:0] m193_93;
   assign m193_93 =10'b0;

   // m193_94 = W*in
   wire signed [9:0] m193_94;
   assign m193_94 =10'b0;

   // m193_95 = W*in
   wire signed [9:0] m193_95;
   assign m193_95 =10'b0;

   // m193_96 = W*in
   wire signed [9:0] m193_96;
   assign m193_96 =10'b0;

   // m193_97 = W*in
   wire signed [9:0] m193_97;
   assign m193_97 =10'b0;

   // m193_98 = W*in
   wire signed [9:0] m193_98;
   assign m193_98 =10'b0;

   // m193_99 = W*in
   wire signed [9:0] m193_99;
   assign m193_99 =10'b0;

   // m193_100 = W*in
   wire signed [9:0] m193_100;
   assign m193_100 =10'b0;

   // m193_101 = W*in
   wire signed [9:0] m193_101;
   assign m193_101 =10'b0;

   // m193_102 = W*in
   wire signed [9:0] m193_102;
   assign m193_102 =10'b0;

   // m193_103 = W*in
   wire signed [9:0] m193_103;
   assign m193_103 =10'b0;

   // m193_104 = W*in
   wire signed [9:0] m193_104;
   assign m193_104 =10'b0;

   // m193_105 = W*in
   wire signed [9:0] m193_105;
   assign m193_105 =10'b0;

   // m193_106 = W*in
   wire signed [9:0] m193_106;
   assign m193_106 =10'b0;

   // m193_107 = W*in
   wire signed [9:0] m193_107;
   assign m193_107 =10'b0;

   // m193_108 = W*in
   wire signed [9:0] m193_108;
   assign m193_108 =10'b0;

   // m193_109 = W*in
   wire signed [9:0] m193_109;
   assign m193_109 =10'b0;

   // m193_110 = W*in
   wire signed [9:0] m193_110;
   assign m193_110 =10'b0;

   // m193_111 = W*in
   wire signed [9:0] m193_111;
   assign m193_111 =10'b0;

   // m193_112 = W*in
   wire signed [9:0] m193_112;
   assign m193_112 =10'b0;

   // m193_113 = W*in
   wire signed [9:0] m193_113;
   assign m193_113 =10'b0;

   // m193_114 = W*in
   wire signed [9:0] m193_114;
   assign m193_114 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_115 = W*in
   wire signed [9:0] m193_115;
   assign m193_115 ={ {5{neg193[5]}} , neg193[5:1] };

   // m193_116 = W*in
   wire signed [9:0] m193_116;
   assign m193_116 =10'b0;

   // m193_117 = W*in
   wire signed [9:0] m193_117;
   assign m193_117 =10'b0;

   // m194_1 = W*in
   wire signed [9:0] m194_1;
   assign m194_1 =10'b0;

   // m194_2 = W*in
   wire signed [9:0] m194_2;
   assign m194_2 =10'b0;

   // m194_3 = W*in
   wire signed [9:0] m194_3;
   assign m194_3 =10'b0;

   // m194_4 = W*in
   wire signed [9:0] m194_4;
   assign m194_4 =10'b0;

   // m194_5 = W*in
   wire signed [9:0] m194_5;
   assign m194_5 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_6 = W*in
   wire signed [9:0] m194_6;
   assign m194_6 =10'b0;

   // m194_7 = W*in
   wire signed [9:0] m194_7;
   assign m194_7 =10'b0;

   // m194_8 = W*in
   wire signed [9:0] m194_8;
   assign m194_8 =10'b0;

   // m194_9 = W*in
   wire signed [9:0] m194_9;
   assign m194_9 =10'b0;

   // m194_10 = W*in
   wire signed [9:0] m194_10;
   assign m194_10 =10'b0;

   // m194_11 = W*in
   wire signed [9:0] m194_11;
   assign m194_11 =10'b0;

   // m194_12 = W*in
   wire signed [9:0] m194_12;
   assign m194_12 =10'b0;

   // m194_13 = W*in
   wire signed [9:0] m194_13;
   assign m194_13 =10'b0;

   // m194_14 = W*in
   wire signed [9:0] m194_14;
   assign m194_14 =10'b0;

   // m194_15 = W*in
   wire signed [9:0] m194_15;
   assign m194_15 =10'b0;

   // m194_16 = W*in
   wire signed [9:0] m194_16;
   assign m194_16 ={ {5{neg194[5]}} , neg194[5:1] };

   // m194_17 = W*in
   wire signed [9:0] m194_17;
   assign m194_17 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_18 = W*in
   wire signed [9:0] m194_18;
   assign m194_18 =10'b0;

   // m194_19 = W*in
   wire signed [9:0] m194_19;
   assign m194_19 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_20 = W*in
   wire signed [9:0] m194_20;
   assign m194_20 ={ {5{in194[5]}} , in194[5:1] };

   // m194_21 = W*in
   wire signed [9:0] m194_21;
   assign m194_21 =10'b0;

   // m194_22 = W*in
   wire signed [9:0] m194_22;
   assign m194_22 =10'b0;

   // m194_23 = W*in
   wire signed [9:0] m194_23;
   assign m194_23 ={ {5{in194[5]}} , in194[5:1] };

   // m194_24 = W*in
   wire signed [9:0] m194_24;
   assign m194_24 =10'b0;

   // m194_25 = W*in
   wire signed [9:0] m194_25;
   assign m194_25 =10'b0;

   // m194_26 = W*in
   wire signed [9:0] m194_26;
   assign m194_26 ={ {4{in194[5]}} , in194[5:0] };

   // m194_27 = W*in
   wire signed [9:0] m194_27;
   assign m194_27 =10'b0;

   // m194_28 = W*in
   wire signed [9:0] m194_28;
   assign m194_28 =10'b0;

   // m194_29 = W*in
   wire signed [9:0] m194_29;
   assign m194_29 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_30 = W*in
   wire signed [9:0] m194_30;
   assign m194_30 =10'b0;

   // m194_31 = W*in
   wire signed [9:0] m194_31;
   assign m194_31 ={ {5{neg194[5]}} , neg194[5:1] };

   // m194_32 = W*in
   wire signed [9:0] m194_32;
   assign m194_32 =10'b0;

   // m194_33 = W*in
   wire signed [9:0] m194_33;
   assign m194_33 =10'b0;

   // m194_34 = W*in
   wire signed [9:0] m194_34;
   assign m194_34 =10'b0;

   // m194_35 = W*in
   wire signed [9:0] m194_35;
   assign m194_35 ={ {5{in194[5]}} , in194[5:1] };

   // m194_36 = W*in
   wire signed [9:0] m194_36;
   assign m194_36 ={ {5{neg194[5]}} , neg194[5:1] };

   // m194_37 = W*in
   wire signed [9:0] m194_37;
   assign m194_37 =10'b0;

   // m194_38 = W*in
   wire signed [9:0] m194_38;
   assign m194_38 =10'b0;

   // m194_39 = W*in
   wire signed [9:0] m194_39;
   assign m194_39 =10'b0;

   // m194_40 = W*in
   wire signed [9:0] m194_40;
   assign m194_40 =10'b0;

   // m194_41 = W*in
   wire signed [9:0] m194_41;
   assign m194_41 =10'b0;

   // m194_42 = W*in
   wire signed [9:0] m194_42;
   assign m194_42 =10'b0;

   // m194_43 = W*in
   wire signed [9:0] m194_43;
   assign m194_43 =10'b0;

   // m194_44 = W*in
   wire signed [9:0] m194_44;
   assign m194_44 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_45 = W*in
   wire signed [9:0] m194_45;
   assign m194_45 =10'b0;

   // m194_46 = W*in
   wire signed [9:0] m194_46;
   assign m194_46 =10'b0;

   // m194_47 = W*in
   wire signed [9:0] m194_47;
   assign m194_47 =10'b0;

   // m194_48 = W*in
   wire signed [9:0] m194_48;
   assign m194_48 ={ {4{in194[5]}} , in194[5:0] };

   // m194_49 = W*in
   wire signed [9:0] m194_49;
   assign m194_49 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_50 = W*in
   wire signed [9:0] m194_50;
   assign m194_50 =10'b0;

   // m194_51 = W*in
   wire signed [9:0] m194_51;
   assign m194_51 =10'b0;

   // m194_52 = W*in
   wire signed [9:0] m194_52;
   assign m194_52 =10'b0;

   // m194_53 = W*in
   wire signed [9:0] m194_53;
   assign m194_53 ={ {3{neg194[5]}} , neg194 , {1{1'b0}} };

   // m194_54 = W*in
   wire signed [9:0] m194_54;
   assign m194_54 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_55 = W*in
   wire signed [9:0] m194_55;
   assign m194_55 =10'b0;

   // m194_56 = W*in
   wire signed [9:0] m194_56;
   assign m194_56 =10'b0;

   // m194_57 = W*in
   wire signed [9:0] m194_57;
   assign m194_57 =10'b0;

   // m194_58 = W*in
   wire signed [9:0] m194_58;
   assign m194_58 =10'b0;

   // m194_59 = W*in
   wire signed [9:0] m194_59;
   assign m194_59 =10'b0;

   // m194_60 = W*in
   wire signed [9:0] m194_60;
   assign m194_60 =10'b0;

   // m194_61 = W*in
   wire signed [9:0] m194_61;
   assign m194_61 =10'b0;

   // m194_62 = W*in
   wire signed [9:0] m194_62;
   assign m194_62 =10'b0;

   // m194_63 = W*in
   wire signed [9:0] m194_63;
   assign m194_63 =10'b0;

   // m194_64 = W*in
   wire signed [9:0] m194_64;
   assign m194_64 =10'b0;

   // m194_65 = W*in
   wire signed [9:0] m194_65;
   assign m194_65 =10'b0;

   // m194_66 = W*in
   wire signed [9:0] m194_66;
   assign m194_66 =10'b0;

   // m194_67 = W*in
   wire signed [9:0] m194_67;
   assign m194_67 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_68 = W*in
   wire signed [9:0] m194_68;
   assign m194_68 =10'b0;

   // m194_69 = W*in
   wire signed [9:0] m194_69;
   assign m194_69 =10'b0;

   // m194_70 = W*in
   wire signed [9:0] m194_70;
   assign m194_70 =10'b0;

   // m194_71 = W*in
   wire signed [9:0] m194_71;
   assign m194_71 ={ {5{in194[5]}} , in194[5:1] };

   // m194_72 = W*in
   wire signed [9:0] m194_72;
   assign m194_72 ={ {5{in194[5]}} , in194[5:1] };

   // m194_73 = W*in
   wire signed [9:0] m194_73;
   assign m194_73 ={ {5{neg194[5]}} , neg194[5:1] };

   // m194_74 = W*in
   wire signed [9:0] m194_74;
   assign m194_74 =10'b0;

   // m194_75 = W*in
   wire signed [9:0] m194_75;
   assign m194_75 ={ {4{in194[5]}} , in194[5:0] };

   // m194_76 = W*in
   wire signed [9:0] m194_76;
   assign m194_76 =10'b0;

   // m194_77 = W*in
   wire signed [9:0] m194_77;
   assign m194_77 =10'b0;

   // m194_78 = W*in
   wire signed [9:0] m194_78;
   assign m194_78 ={ {5{in194[5]}} , in194[5:1] };

   // m194_79 = W*in
   wire signed [9:0] m194_79;
   assign m194_79 =10'b0;

   // m194_80 = W*in
   wire signed [9:0] m194_80;
   assign m194_80 =10'b0;

   // m194_81 = W*in
   wire signed [9:0] m194_81;
   assign m194_81 =10'b0;

   // m194_82 = W*in
   wire signed [9:0] m194_82;
   assign m194_82 =10'b0;

   // m194_83 = W*in
   wire signed [9:0] m194_83;
   assign m194_83 =10'b0;

   // m194_84 = W*in
   wire signed [9:0] m194_84;
   assign m194_84 =10'b0;

   // m194_85 = W*in
   wire signed [9:0] m194_85;
   assign m194_85 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_86 = W*in
   wire signed [9:0] m194_86;
   assign m194_86 =10'b0;

   // m194_87 = W*in
   wire signed [9:0] m194_87;
   assign m194_87 ={ {4{in194[5]}} , in194[5:0] };

   // m194_88 = W*in
   wire signed [9:0] m194_88;
   assign m194_88 ={ {4{in194[5]}} , in194[5:0] };

   // m194_89 = W*in
   wire signed [9:0] m194_89;
   assign m194_89 =10'b0;

   // m194_90 = W*in
   wire signed [9:0] m194_90;
   assign m194_90 =10'b0;

   // m194_91 = W*in
   wire signed [9:0] m194_91;
   assign m194_91 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_92 = W*in
   wire signed [9:0] m194_92;
   assign m194_92 =10'b0;

   // m194_93 = W*in
   wire signed [9:0] m194_93;
   assign m194_93 =10'b0;

   // m194_94 = W*in
   wire signed [9:0] m194_94;
   assign m194_94 =10'b0;

   // m194_95 = W*in
   wire signed [9:0] m194_95;
   assign m194_95 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_96 = W*in
   wire signed [9:0] m194_96;
   assign m194_96 =10'b0;

   // m194_97 = W*in
   wire signed [9:0] m194_97;
   assign m194_97 =10'b0;

   // m194_98 = W*in
   wire signed [9:0] m194_98;
   assign m194_98 =10'b0;

   // m194_99 = W*in
   wire signed [9:0] m194_99;
   assign m194_99 =10'b0;

   // m194_100 = W*in
   wire signed [9:0] m194_100;
   assign m194_100 =10'b0;

   // m194_101 = W*in
   wire signed [9:0] m194_101;
   assign m194_101 =10'b0;

   // m194_102 = W*in
   wire signed [9:0] m194_102;
   assign m194_102 =10'b0;

   // m194_103 = W*in
   wire signed [9:0] m194_103;
   assign m194_103 =10'b0;

   // m194_104 = W*in
   wire signed [9:0] m194_104;
   assign m194_104 =10'b0;

   // m194_105 = W*in
   wire signed [9:0] m194_105;
   assign m194_105 =10'b0;

   // m194_106 = W*in
   wire signed [9:0] m194_106;
   assign m194_106 =10'b0;

   // m194_107 = W*in
   wire signed [9:0] m194_107;
   assign m194_107 =10'b0;

   // m194_108 = W*in
   wire signed [9:0] m194_108;
   assign m194_108 ={ {4{in194[5]}} , in194[5:0] };

   // m194_109 = W*in
   wire signed [9:0] m194_109;
   assign m194_109 ={ {4{in194[5]}} , in194[5:0] };

   // m194_110 = W*in
   wire signed [9:0] m194_110;
   assign m194_110 ={ {4{neg194[5]}} , neg194[5:0] };

   // m194_111 = W*in
   wire signed [9:0] m194_111;
   assign m194_111 =10'b0;

   // m194_112 = W*in
   wire signed [9:0] m194_112;
   assign m194_112 =10'b0;

   // m194_113 = W*in
   wire signed [9:0] m194_113;
   assign m194_113 =10'b0;

   // m194_114 = W*in
   wire signed [9:0] m194_114;
   assign m194_114 =10'b0;

   // m194_115 = W*in
   wire signed [9:0] m194_115;
   assign m194_115 ={ {5{in194[5]}} , in194[5:1] };

   // m194_116 = W*in
   wire signed [9:0] m194_116;
   assign m194_116 ={ {4{in194[5]}} , in194[5:0] };

   // m194_117 = W*in
   wire signed [9:0] m194_117;
   assign m194_117 ={ {4{in194[5]}} , in194[5:0] };

   // m195_1 = W*in
   wire signed [9:0] m195_1;
   assign m195_1 =10'b0;

   // m195_2 = W*in
   wire signed [9:0] m195_2;
   assign m195_2 =10'b0;

   // m195_3 = W*in
   wire signed [9:0] m195_3;
   assign m195_3 =10'b0;

   // m195_4 = W*in
   wire signed [9:0] m195_4;
   assign m195_4 =10'b0;

   // m195_5 = W*in
   wire signed [9:0] m195_5;
   assign m195_5 =10'b0;

   // m195_6 = W*in
   wire signed [9:0] m195_6;
   assign m195_6 =10'b0;

   // m195_7 = W*in
   wire signed [9:0] m195_7;
   assign m195_7 =10'b0;

   // m195_8 = W*in
   wire signed [9:0] m195_8;
   assign m195_8 =10'b0;

   // m195_9 = W*in
   wire signed [9:0] m195_9;
   assign m195_9 =10'b0;

   // m195_10 = W*in
   wire signed [9:0] m195_10;
   assign m195_10 =10'b0;

   // m195_11 = W*in
   wire signed [9:0] m195_11;
   assign m195_11 =10'b0;

   // m195_12 = W*in
   wire signed [9:0] m195_12;
   assign m195_12 =10'b0;

   // m195_13 = W*in
   wire signed [9:0] m195_13;
   assign m195_13 =10'b0;

   // m195_14 = W*in
   wire signed [9:0] m195_14;
   assign m195_14 =10'b0;

   // m195_15 = W*in
   wire signed [9:0] m195_15;
   assign m195_15 =10'b0;

   // m195_16 = W*in
   wire signed [9:0] m195_16;
   assign m195_16 =10'b0;

   // m195_17 = W*in
   wire signed [9:0] m195_17;
   assign m195_17 =10'b0;

   // m195_18 = W*in
   wire signed [9:0] m195_18;
   assign m195_18 =10'b0;

   // m195_19 = W*in
   wire signed [9:0] m195_19;
   assign m195_19 =10'b0;

   // m195_20 = W*in
   wire signed [9:0] m195_20;
   assign m195_20 ={ {5{in195[5]}} , in195[5:1] };

   // m195_21 = W*in
   wire signed [9:0] m195_21;
   assign m195_21 =10'b0;

   // m195_22 = W*in
   wire signed [9:0] m195_22;
   assign m195_22 ={ {5{in195[5]}} , in195[5:1] };

   // m195_23 = W*in
   wire signed [9:0] m195_23;
   assign m195_23 =10'b0;

   // m195_24 = W*in
   wire signed [9:0] m195_24;
   assign m195_24 =10'b0;

   // m195_25 = W*in
   wire signed [9:0] m195_25;
   assign m195_25 =10'b0;

   // m195_26 = W*in
   wire signed [9:0] m195_26;
   assign m195_26 =10'b0;

   // m195_27 = W*in
   wire signed [9:0] m195_27;
   assign m195_27 =10'b0;

   // m195_28 = W*in
   wire signed [9:0] m195_28;
   assign m195_28 =10'b0;

   // m195_29 = W*in
   wire signed [9:0] m195_29;
   assign m195_29 =10'b0;

   // m195_30 = W*in
   wire signed [9:0] m195_30;
   assign m195_30 =10'b0;

   // m195_31 = W*in
   wire signed [9:0] m195_31;
   assign m195_31 ={ {5{neg195[5]}} , neg195[5:1] };

   // m195_32 = W*in
   wire signed [9:0] m195_32;
   assign m195_32 =10'b0;

   // m195_33 = W*in
   wire signed [9:0] m195_33;
   assign m195_33 =10'b0;

   // m195_34 = W*in
   wire signed [9:0] m195_34;
   assign m195_34 =10'b0;

   // m195_35 = W*in
   wire signed [9:0] m195_35;
   assign m195_35 =10'b0;

   // m195_36 = W*in
   wire signed [9:0] m195_36;
   assign m195_36 =10'b0;

   // m195_37 = W*in
   wire signed [9:0] m195_37;
   assign m195_37 =10'b0;

   // m195_38 = W*in
   wire signed [9:0] m195_38;
   assign m195_38 =10'b0;

   // m195_39 = W*in
   wire signed [9:0] m195_39;
   assign m195_39 =10'b0;

   // m195_40 = W*in
   wire signed [9:0] m195_40;
   assign m195_40 =10'b0;

   // m195_41 = W*in
   wire signed [9:0] m195_41;
   assign m195_41 =10'b0;

   // m195_42 = W*in
   wire signed [9:0] m195_42;
   assign m195_42 =10'b0;

   // m195_43 = W*in
   wire signed [9:0] m195_43;
   assign m195_43 =10'b0;

   // m195_44 = W*in
   wire signed [9:0] m195_44;
   assign m195_44 =10'b0;

   // m195_45 = W*in
   wire signed [9:0] m195_45;
   assign m195_45 =10'b0;

   // m195_46 = W*in
   wire signed [9:0] m195_46;
   assign m195_46 =10'b0;

   // m195_47 = W*in
   wire signed [9:0] m195_47;
   assign m195_47 =10'b0;

   // m195_48 = W*in
   wire signed [9:0] m195_48;
   assign m195_48 =10'b0;

   // m195_49 = W*in
   wire signed [9:0] m195_49;
   assign m195_49 =10'b0;

   // m195_50 = W*in
   wire signed [9:0] m195_50;
   assign m195_50 =10'b0;

   // m195_51 = W*in
   wire signed [9:0] m195_51;
   assign m195_51 =10'b0;

   // m195_52 = W*in
   wire signed [9:0] m195_52;
   assign m195_52 =10'b0;

   // m195_53 = W*in
   wire signed [9:0] m195_53;
   assign m195_53 =10'b0;

   // m195_54 = W*in
   wire signed [9:0] m195_54;
   assign m195_54 =10'b0;

   // m195_55 = W*in
   wire signed [9:0] m195_55;
   assign m195_55 =10'b0;

   // m195_56 = W*in
   wire signed [9:0] m195_56;
   assign m195_56 =10'b0;

   // m195_57 = W*in
   wire signed [9:0] m195_57;
   assign m195_57 =10'b0;

   // m195_58 = W*in
   wire signed [9:0] m195_58;
   assign m195_58 =10'b0;

   // m195_59 = W*in
   wire signed [9:0] m195_59;
   assign m195_59 =10'b0;

   // m195_60 = W*in
   wire signed [9:0] m195_60;
   assign m195_60 =10'b0;

   // m195_61 = W*in
   wire signed [9:0] m195_61;
   assign m195_61 =10'b0;

   // m195_62 = W*in
   wire signed [9:0] m195_62;
   assign m195_62 =10'b0;

   // m195_63 = W*in
   wire signed [9:0] m195_63;
   assign m195_63 =10'b0;

   // m195_64 = W*in
   wire signed [9:0] m195_64;
   assign m195_64 ={ {5{neg195[5]}} , neg195[5:1] };

   // m195_65 = W*in
   wire signed [9:0] m195_65;
   assign m195_65 =10'b0;

   // m195_66 = W*in
   wire signed [9:0] m195_66;
   assign m195_66 ={ {5{neg195[5]}} , neg195[5:1] };

   // m195_67 = W*in
   wire signed [9:0] m195_67;
   assign m195_67 =10'b0;

   // m195_68 = W*in
   wire signed [9:0] m195_68;
   assign m195_68 =10'b0;

   // m195_69 = W*in
   wire signed [9:0] m195_69;
   assign m195_69 =10'b0;

   // m195_70 = W*in
   wire signed [9:0] m195_70;
   assign m195_70 =10'b0;

   // m195_71 = W*in
   wire signed [9:0] m195_71;
   assign m195_71 =10'b0;

   // m195_72 = W*in
   wire signed [9:0] m195_72;
   assign m195_72 =10'b0;

   // m195_73 = W*in
   wire signed [9:0] m195_73;
   assign m195_73 ={ {5{neg195[5]}} , neg195[5:1] };

   // m195_74 = W*in
   wire signed [9:0] m195_74;
   assign m195_74 =10'b0;

   // m195_75 = W*in
   wire signed [9:0] m195_75;
   assign m195_75 =10'b0;

   // m195_76 = W*in
   wire signed [9:0] m195_76;
   assign m195_76 =10'b0;

   // m195_77 = W*in
   wire signed [9:0] m195_77;
   assign m195_77 =10'b0;

   // m195_78 = W*in
   wire signed [9:0] m195_78;
   assign m195_78 =10'b0;

   // m195_79 = W*in
   wire signed [9:0] m195_79;
   assign m195_79 =10'b0;

   // m195_80 = W*in
   wire signed [9:0] m195_80;
   assign m195_80 =10'b0;

   // m195_81 = W*in
   wire signed [9:0] m195_81;
   assign m195_81 =10'b0;

   // m195_82 = W*in
   wire signed [9:0] m195_82;
   assign m195_82 =10'b0;

   // m195_83 = W*in
   wire signed [9:0] m195_83;
   assign m195_83 =10'b0;

   // m195_84 = W*in
   wire signed [9:0] m195_84;
   assign m195_84 =10'b0;

   // m195_85 = W*in
   wire signed [9:0] m195_85;
   assign m195_85 ={ {5{neg195[5]}} , neg195[5:1] };

   // m195_86 = W*in
   wire signed [9:0] m195_86;
   assign m195_86 =10'b0;

   // m195_87 = W*in
   wire signed [9:0] m195_87;
   assign m195_87 =10'b0;

   // m195_88 = W*in
   wire signed [9:0] m195_88;
   assign m195_88 =10'b0;

   // m195_89 = W*in
   wire signed [9:0] m195_89;
   assign m195_89 =10'b0;

   // m195_90 = W*in
   wire signed [9:0] m195_90;
   assign m195_90 =10'b0;

   // m195_91 = W*in
   wire signed [9:0] m195_91;
   assign m195_91 =10'b0;

   // m195_92 = W*in
   wire signed [9:0] m195_92;
   assign m195_92 =10'b0;

   // m195_93 = W*in
   wire signed [9:0] m195_93;
   assign m195_93 =10'b0;

   // m195_94 = W*in
   wire signed [9:0] m195_94;
   assign m195_94 =10'b0;

   // m195_95 = W*in
   wire signed [9:0] m195_95;
   assign m195_95 =10'b0;

   // m195_96 = W*in
   wire signed [9:0] m195_96;
   assign m195_96 =10'b0;

   // m195_97 = W*in
   wire signed [9:0] m195_97;
   assign m195_97 =10'b0;

   // m195_98 = W*in
   wire signed [9:0] m195_98;
   assign m195_98 =10'b0;

   // m195_99 = W*in
   wire signed [9:0] m195_99;
   assign m195_99 =10'b0;

   // m195_100 = W*in
   wire signed [9:0] m195_100;
   assign m195_100 =10'b0;

   // m195_101 = W*in
   wire signed [9:0] m195_101;
   assign m195_101 =10'b0;

   // m195_102 = W*in
   wire signed [9:0] m195_102;
   assign m195_102 =10'b0;

   // m195_103 = W*in
   wire signed [9:0] m195_103;
   assign m195_103 =10'b0;

   // m195_104 = W*in
   wire signed [9:0] m195_104;
   assign m195_104 =10'b0;

   // m195_105 = W*in
   wire signed [9:0] m195_105;
   assign m195_105 =10'b0;

   // m195_106 = W*in
   wire signed [9:0] m195_106;
   assign m195_106 =10'b0;

   // m195_107 = W*in
   wire signed [9:0] m195_107;
   assign m195_107 =10'b0;

   // m195_108 = W*in
   wire signed [9:0] m195_108;
   assign m195_108 =10'b0;

   // m195_109 = W*in
   wire signed [9:0] m195_109;
   assign m195_109 ={ {5{in195[5]}} , in195[5:1] };

   // m195_110 = W*in
   wire signed [9:0] m195_110;
   assign m195_110 =10'b0;

   // m195_111 = W*in
   wire signed [9:0] m195_111;
   assign m195_111 =10'b0;

   // m195_112 = W*in
   wire signed [9:0] m195_112;
   assign m195_112 =10'b0;

   // m195_113 = W*in
   wire signed [9:0] m195_113;
   assign m195_113 =10'b0;

   // m195_114 = W*in
   wire signed [9:0] m195_114;
   assign m195_114 =10'b0;

   // m195_115 = W*in
   wire signed [9:0] m195_115;
   assign m195_115 =10'b0;

   // m195_116 = W*in
   wire signed [9:0] m195_116;
   assign m195_116 =10'b0;

   // m195_117 = W*in
   wire signed [9:0] m195_117;
   assign m195_117 =10'b0;

   // m196_1 = W*in
   wire signed [9:0] m196_1;
   assign m196_1 =10'b0;

   // m196_2 = W*in
   wire signed [9:0] m196_2;
   assign m196_2 =10'b0;

   // m196_3 = W*in
   wire signed [9:0] m196_3;
   assign m196_3 =10'b0;

   // m196_4 = W*in
   wire signed [9:0] m196_4;
   assign m196_4 =10'b0;

   // m196_5 = W*in
   wire signed [9:0] m196_5;
   assign m196_5 =10'b0;

   // m196_6 = W*in
   wire signed [9:0] m196_6;
   assign m196_6 =10'b0;

   // m196_7 = W*in
   wire signed [9:0] m196_7;
   assign m196_7 ={ {4{in196[5]}} , in196[5:0] };

   // m196_8 = W*in
   wire signed [9:0] m196_8;
   assign m196_8 =10'b0;

   // m196_9 = W*in
   wire signed [9:0] m196_9;
   assign m196_9 =10'b0;

   // m196_10 = W*in
   wire signed [9:0] m196_10;
   assign m196_10 =10'b0;

   // m196_11 = W*in
   wire signed [9:0] m196_11;
   assign m196_11 =10'b0;

   // m196_12 = W*in
   wire signed [9:0] m196_12;
   assign m196_12 =10'b0;

   // m196_13 = W*in
   wire signed [9:0] m196_13;
   assign m196_13 =10'b0;

   // m196_14 = W*in
   wire signed [9:0] m196_14;
   assign m196_14 =10'b0;

   // m196_15 = W*in
   wire signed [9:0] m196_15;
   assign m196_15 =10'b0;

   // m196_16 = W*in
   wire signed [9:0] m196_16;
   assign m196_16 ={ {5{in196[5]}} , in196[5:1] };

   // m196_17 = W*in
   wire signed [9:0] m196_17;
   assign m196_17 =10'b0;

   // m196_18 = W*in
   wire signed [9:0] m196_18;
   assign m196_18 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_19 = W*in
   wire signed [9:0] m196_19;
   assign m196_19 =10'b0;

   // m196_20 = W*in
   wire signed [9:0] m196_20;
   assign m196_20 =10'b0;

   // m196_21 = W*in
   wire signed [9:0] m196_21;
   assign m196_21 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_22 = W*in
   wire signed [9:0] m196_22;
   assign m196_22 ={ {5{in196[5]}} , in196[5:1] };

   // m196_23 = W*in
   wire signed [9:0] m196_23;
   assign m196_23 =10'b0;

   // m196_24 = W*in
   wire signed [9:0] m196_24;
   assign m196_24 =10'b0;

   // m196_25 = W*in
   wire signed [9:0] m196_25;
   assign m196_25 =10'b0;

   // m196_26 = W*in
   wire signed [9:0] m196_26;
   assign m196_26 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_27 = W*in
   wire signed [9:0] m196_27;
   assign m196_27 =10'b0;

   // m196_28 = W*in
   wire signed [9:0] m196_28;
   assign m196_28 =10'b0;

   // m196_29 = W*in
   wire signed [9:0] m196_29;
   assign m196_29 =10'b0;

   // m196_30 = W*in
   wire signed [9:0] m196_30;
   assign m196_30 =10'b0;

   // m196_31 = W*in
   wire signed [9:0] m196_31;
   assign m196_31 =10'b0;

   // m196_32 = W*in
   wire signed [9:0] m196_32;
   assign m196_32 =10'b0;

   // m196_33 = W*in
   wire signed [9:0] m196_33;
   assign m196_33 =10'b0;

   // m196_34 = W*in
   wire signed [9:0] m196_34;
   assign m196_34 =10'b0;

   // m196_35 = W*in
   wire signed [9:0] m196_35;
   assign m196_35 =10'b0;

   // m196_36 = W*in
   wire signed [9:0] m196_36;
   assign m196_36 ={ {5{in196[5]}} , in196[5:1] };

   // m196_37 = W*in
   wire signed [9:0] m196_37;
   assign m196_37 =10'b0;

   // m196_38 = W*in
   wire signed [9:0] m196_38;
   assign m196_38 =10'b0;

   // m196_39 = W*in
   wire signed [9:0] m196_39;
   assign m196_39 =10'b0;

   // m196_40 = W*in
   wire signed [9:0] m196_40;
   assign m196_40 =10'b0;

   // m196_41 = W*in
   wire signed [9:0] m196_41;
   assign m196_41 =10'b0;

   // m196_42 = W*in
   wire signed [9:0] m196_42;
   assign m196_42 =10'b0;

   // m196_43 = W*in
   wire signed [9:0] m196_43;
   assign m196_43 =10'b0;

   // m196_44 = W*in
   wire signed [9:0] m196_44;
   assign m196_44 =10'b0;

   // m196_45 = W*in
   wire signed [9:0] m196_45;
   assign m196_45 =10'b0;

   // m196_46 = W*in
   wire signed [9:0] m196_46;
   assign m196_46 =10'b0;

   // m196_47 = W*in
   wire signed [9:0] m196_47;
   assign m196_47 =10'b0;

   // m196_48 = W*in
   wire signed [9:0] m196_48;
   assign m196_48 =10'b0;

   // m196_49 = W*in
   wire signed [9:0] m196_49;
   assign m196_49 =10'b0;

   // m196_50 = W*in
   wire signed [9:0] m196_50;
   assign m196_50 =10'b0;

   // m196_51 = W*in
   wire signed [9:0] m196_51;
   assign m196_51 =10'b0;

   // m196_52 = W*in
   wire signed [9:0] m196_52;
   assign m196_52 =10'b0;

   // m196_53 = W*in
   wire signed [9:0] m196_53;
   assign m196_53 =10'b0;

   // m196_54 = W*in
   wire signed [9:0] m196_54;
   assign m196_54 =10'b0;

   // m196_55 = W*in
   wire signed [9:0] m196_55;
   assign m196_55 =10'b0;

   // m196_56 = W*in
   wire signed [9:0] m196_56;
   assign m196_56 ={ {4{in196[5]}} , in196[5:0] };

   // m196_57 = W*in
   wire signed [9:0] m196_57;
   assign m196_57 =10'b0;

   // m196_58 = W*in
   wire signed [9:0] m196_58;
   assign m196_58 =10'b0;

   // m196_59 = W*in
   wire signed [9:0] m196_59;
   assign m196_59 =10'b0;

   // m196_60 = W*in
   wire signed [9:0] m196_60;
   assign m196_60 =10'b0;

   // m196_61 = W*in
   wire signed [9:0] m196_61;
   assign m196_61 =10'b0;

   // m196_62 = W*in
   wire signed [9:0] m196_62;
   assign m196_62 =10'b0;

   // m196_63 = W*in
   wire signed [9:0] m196_63;
   assign m196_63 =10'b0;

   // m196_64 = W*in
   wire signed [9:0] m196_64;
   assign m196_64 =10'b0;

   // m196_65 = W*in
   wire signed [9:0] m196_65;
   assign m196_65 =10'b0;

   // m196_66 = W*in
   wire signed [9:0] m196_66;
   assign m196_66 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_67 = W*in
   wire signed [9:0] m196_67;
   assign m196_67 =10'b0;

   // m196_68 = W*in
   wire signed [9:0] m196_68;
   assign m196_68 =10'b0;

   // m196_69 = W*in
   wire signed [9:0] m196_69;
   assign m196_69 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_70 = W*in
   wire signed [9:0] m196_70;
   assign m196_70 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_71 = W*in
   wire signed [9:0] m196_71;
   assign m196_71 =10'b0;

   // m196_72 = W*in
   wire signed [9:0] m196_72;
   assign m196_72 =10'b0;

   // m196_73 = W*in
   wire signed [9:0] m196_73;
   assign m196_73 ={ {5{in196[5]}} , in196[5:1] };

   // m196_74 = W*in
   wire signed [9:0] m196_74;
   assign m196_74 ={ {5{neg196[5]}} , neg196[5:1] };

   // m196_75 = W*in
   wire signed [9:0] m196_75;
   assign m196_75 =10'b0;

   // m196_76 = W*in
   wire signed [9:0] m196_76;
   assign m196_76 =10'b0;

   // m196_77 = W*in
   wire signed [9:0] m196_77;
   assign m196_77 =10'b0;

   // m196_78 = W*in
   wire signed [9:0] m196_78;
   assign m196_78 =10'b0;

   // m196_79 = W*in
   wire signed [9:0] m196_79;
   assign m196_79 =10'b0;

   // m196_80 = W*in
   wire signed [9:0] m196_80;
   assign m196_80 =10'b0;

   // m196_81 = W*in
   wire signed [9:0] m196_81;
   assign m196_81 =10'b0;

   // m196_82 = W*in
   wire signed [9:0] m196_82;
   assign m196_82 =10'b0;

   // m196_83 = W*in
   wire signed [9:0] m196_83;
   assign m196_83 =10'b0;

   // m196_84 = W*in
   wire signed [9:0] m196_84;
   assign m196_84 =10'b0;

   // m196_85 = W*in
   wire signed [9:0] m196_85;
   assign m196_85 =10'b0;

   // m196_86 = W*in
   wire signed [9:0] m196_86;
   assign m196_86 =10'b0;

   // m196_87 = W*in
   wire signed [9:0] m196_87;
   assign m196_87 =10'b0;

   // m196_88 = W*in
   wire signed [9:0] m196_88;
   assign m196_88 =10'b0;

   // m196_89 = W*in
   wire signed [9:0] m196_89;
   assign m196_89 =10'b0;

   // m196_90 = W*in
   wire signed [9:0] m196_90;
   assign m196_90 =10'b0;

   // m196_91 = W*in
   wire signed [9:0] m196_91;
   assign m196_91 =10'b0;

   // m196_92 = W*in
   wire signed [9:0] m196_92;
   assign m196_92 =10'b0;

   // m196_93 = W*in
   wire signed [9:0] m196_93;
   assign m196_93 =10'b0;

   // m196_94 = W*in
   wire signed [9:0] m196_94;
   assign m196_94 =10'b0;

   // m196_95 = W*in
   wire signed [9:0] m196_95;
   assign m196_95 =10'b0;

   // m196_96 = W*in
   wire signed [9:0] m196_96;
   assign m196_96 =10'b0;

   // m196_97 = W*in
   wire signed [9:0] m196_97;
   assign m196_97 =10'b0;

   // m196_98 = W*in
   wire signed [9:0] m196_98;
   assign m196_98 =10'b0;

   // m196_99 = W*in
   wire signed [9:0] m196_99;
   assign m196_99 =10'b0;

   // m196_100 = W*in
   wire signed [9:0] m196_100;
   assign m196_100 =10'b0;

   // m196_101 = W*in
   wire signed [9:0] m196_101;
   assign m196_101 =10'b0;

   // m196_102 = W*in
   wire signed [9:0] m196_102;
   assign m196_102 =10'b0;

   // m196_103 = W*in
   wire signed [9:0] m196_103;
   assign m196_103 =10'b0;

   // m196_104 = W*in
   wire signed [9:0] m196_104;
   assign m196_104 =10'b0;

   // m196_105 = W*in
   wire signed [9:0] m196_105;
   assign m196_105 =10'b0;

   // m196_106 = W*in
   wire signed [9:0] m196_106;
   assign m196_106 =10'b0;

   // m196_107 = W*in
   wire signed [9:0] m196_107;
   assign m196_107 =10'b0;

   // m196_108 = W*in
   wire signed [9:0] m196_108;
   assign m196_108 =10'b0;

   // m196_109 = W*in
   wire signed [9:0] m196_109;
   assign m196_109 =10'b0;

   // m196_110 = W*in
   wire signed [9:0] m196_110;
   assign m196_110 =10'b0;

   // m196_111 = W*in
   wire signed [9:0] m196_111;
   assign m196_111 =10'b0;

   // m196_112 = W*in
   wire signed [9:0] m196_112;
   assign m196_112 =10'b0;

   // m196_113 = W*in
   wire signed [9:0] m196_113;
   assign m196_113 =10'b0;

   // m196_114 = W*in
   wire signed [9:0] m196_114;
   assign m196_114 =10'b0;

   // m196_115 = W*in
   wire signed [9:0] m196_115;
   assign m196_115 ={ {5{in196[5]}} , in196[5:1] };

   // m196_116 = W*in
   wire signed [9:0] m196_116;
   assign m196_116 =10'b0;

   // m196_117 = W*in
   wire signed [9:0] m196_117;
   assign m196_117 =10'b0;

   // m197_1 = W*in
   wire signed [9:0] m197_1;
   assign m197_1 =10'b0;

   // m197_2 = W*in
   wire signed [9:0] m197_2;
   assign m197_2 =10'b0;

   // m197_3 = W*in
   wire signed [9:0] m197_3;
   assign m197_3 =10'b0;

   // m197_4 = W*in
   wire signed [9:0] m197_4;
   assign m197_4 =10'b0;

   // m197_5 = W*in
   wire signed [9:0] m197_5;
   assign m197_5 =10'b0;

   // m197_6 = W*in
   wire signed [9:0] m197_6;
   assign m197_6 =10'b0;

   // m197_7 = W*in
   wire signed [9:0] m197_7;
   assign m197_7 =10'b0;

   // m197_8 = W*in
   wire signed [9:0] m197_8;
   assign m197_8 =10'b0;

   // m197_9 = W*in
   wire signed [9:0] m197_9;
   assign m197_9 =10'b0;

   // m197_10 = W*in
   wire signed [9:0] m197_10;
   assign m197_10 =10'b0;

   // m197_11 = W*in
   wire signed [9:0] m197_11;
   assign m197_11 =10'b0;

   // m197_12 = W*in
   wire signed [9:0] m197_12;
   assign m197_12 =10'b0;

   // m197_13 = W*in
   wire signed [9:0] m197_13;
   assign m197_13 =10'b0;

   // m197_14 = W*in
   wire signed [9:0] m197_14;
   assign m197_14 =10'b0;

   // m197_15 = W*in
   wire signed [9:0] m197_15;
   assign m197_15 =10'b0;

   // m197_16 = W*in
   wire signed [9:0] m197_16;
   assign m197_16 =10'b0;

   // m197_17 = W*in
   wire signed [9:0] m197_17;
   assign m197_17 =10'b0;

   // m197_18 = W*in
   wire signed [9:0] m197_18;
   assign m197_18 =10'b0;

   // m197_19 = W*in
   wire signed [9:0] m197_19;
   assign m197_19 =10'b0;

   // m197_20 = W*in
   wire signed [9:0] m197_20;
   assign m197_20 ={ {5{in197[5]}} , in197[5:1] };

   // m197_21 = W*in
   wire signed [9:0] m197_21;
   assign m197_21 =10'b0;

   // m197_22 = W*in
   wire signed [9:0] m197_22;
   assign m197_22 =10'b0;

   // m197_23 = W*in
   wire signed [9:0] m197_23;
   assign m197_23 =10'b0;

   // m197_24 = W*in
   wire signed [9:0] m197_24;
   assign m197_24 =10'b0;

   // m197_25 = W*in
   wire signed [9:0] m197_25;
   assign m197_25 =10'b0;

   // m197_26 = W*in
   wire signed [9:0] m197_26;
   assign m197_26 =10'b0;

   // m197_27 = W*in
   wire signed [9:0] m197_27;
   assign m197_27 =10'b0;

   // m197_28 = W*in
   wire signed [9:0] m197_28;
   assign m197_28 =10'b0;

   // m197_29 = W*in
   wire signed [9:0] m197_29;
   assign m197_29 =10'b0;

   // m197_30 = W*in
   wire signed [9:0] m197_30;
   assign m197_30 =10'b0;

   // m197_31 = W*in
   wire signed [9:0] m197_31;
   assign m197_31 =10'b0;

   // m197_32 = W*in
   wire signed [9:0] m197_32;
   assign m197_32 =10'b0;

   // m197_33 = W*in
   wire signed [9:0] m197_33;
   assign m197_33 =10'b0;

   // m197_34 = W*in
   wire signed [9:0] m197_34;
   assign m197_34 =10'b0;

   // m197_35 = W*in
   wire signed [9:0] m197_35;
   assign m197_35 =10'b0;

   // m197_36 = W*in
   wire signed [9:0] m197_36;
   assign m197_36 =10'b0;

   // m197_37 = W*in
   wire signed [9:0] m197_37;
   assign m197_37 =10'b0;

   // m197_38 = W*in
   wire signed [9:0] m197_38;
   assign m197_38 =10'b0;

   // m197_39 = W*in
   wire signed [9:0] m197_39;
   assign m197_39 =10'b0;

   // m197_40 = W*in
   wire signed [9:0] m197_40;
   assign m197_40 =10'b0;

   // m197_41 = W*in
   wire signed [9:0] m197_41;
   assign m197_41 =10'b0;

   // m197_42 = W*in
   wire signed [9:0] m197_42;
   assign m197_42 =10'b0;

   // m197_43 = W*in
   wire signed [9:0] m197_43;
   assign m197_43 =10'b0;

   // m197_44 = W*in
   wire signed [9:0] m197_44;
   assign m197_44 =10'b0;

   // m197_45 = W*in
   wire signed [9:0] m197_45;
   assign m197_45 =10'b0;

   // m197_46 = W*in
   wire signed [9:0] m197_46;
   assign m197_46 =10'b0;

   // m197_47 = W*in
   wire signed [9:0] m197_47;
   assign m197_47 =10'b0;

   // m197_48 = W*in
   wire signed [9:0] m197_48;
   assign m197_48 =10'b0;

   // m197_49 = W*in
   wire signed [9:0] m197_49;
   assign m197_49 =10'b0;

   // m197_50 = W*in
   wire signed [9:0] m197_50;
   assign m197_50 =10'b0;

   // m197_51 = W*in
   wire signed [9:0] m197_51;
   assign m197_51 =10'b0;

   // m197_52 = W*in
   wire signed [9:0] m197_52;
   assign m197_52 =10'b0;

   // m197_53 = W*in
   wire signed [9:0] m197_53;
   assign m197_53 =10'b0;

   // m197_54 = W*in
   wire signed [9:0] m197_54;
   assign m197_54 =10'b0;

   // m197_55 = W*in
   wire signed [9:0] m197_55;
   assign m197_55 =10'b0;

   // m197_56 = W*in
   wire signed [9:0] m197_56;
   assign m197_56 =10'b0;

   // m197_57 = W*in
   wire signed [9:0] m197_57;
   assign m197_57 =10'b0;

   // m197_58 = W*in
   wire signed [9:0] m197_58;
   assign m197_58 =10'b0;

   // m197_59 = W*in
   wire signed [9:0] m197_59;
   assign m197_59 =10'b0;

   // m197_60 = W*in
   wire signed [9:0] m197_60;
   assign m197_60 =10'b0;

   // m197_61 = W*in
   wire signed [9:0] m197_61;
   assign m197_61 =10'b0;

   // m197_62 = W*in
   wire signed [9:0] m197_62;
   assign m197_62 =10'b0;

   // m197_63 = W*in
   wire signed [9:0] m197_63;
   assign m197_63 =10'b0;

   // m197_64 = W*in
   wire signed [9:0] m197_64;
   assign m197_64 =10'b0;

   // m197_65 = W*in
   wire signed [9:0] m197_65;
   assign m197_65 =10'b0;

   // m197_66 = W*in
   wire signed [9:0] m197_66;
   assign m197_66 ={ {5{neg197[5]}} , neg197[5:1] };

   // m197_67 = W*in
   wire signed [9:0] m197_67;
   assign m197_67 =10'b0;

   // m197_68 = W*in
   wire signed [9:0] m197_68;
   assign m197_68 =10'b0;

   // m197_69 = W*in
   wire signed [9:0] m197_69;
   assign m197_69 =10'b0;

   // m197_70 = W*in
   wire signed [9:0] m197_70;
   assign m197_70 =10'b0;

   // m197_71 = W*in
   wire signed [9:0] m197_71;
   assign m197_71 =10'b0;

   // m197_72 = W*in
   wire signed [9:0] m197_72;
   assign m197_72 ={ {5{in197[5]}} , in197[5:1] };

   // m197_73 = W*in
   wire signed [9:0] m197_73;
   assign m197_73 =10'b0;

   // m197_74 = W*in
   wire signed [9:0] m197_74;
   assign m197_74 =10'b0;

   // m197_75 = W*in
   wire signed [9:0] m197_75;
   assign m197_75 =10'b0;

   // m197_76 = W*in
   wire signed [9:0] m197_76;
   assign m197_76 =10'b0;

   // m197_77 = W*in
   wire signed [9:0] m197_77;
   assign m197_77 =10'b0;

   // m197_78 = W*in
   wire signed [9:0] m197_78;
   assign m197_78 =10'b0;

   // m197_79 = W*in
   wire signed [9:0] m197_79;
   assign m197_79 =10'b0;

   // m197_80 = W*in
   wire signed [9:0] m197_80;
   assign m197_80 =10'b0;

   // m197_81 = W*in
   wire signed [9:0] m197_81;
   assign m197_81 =10'b0;

   // m197_82 = W*in
   wire signed [9:0] m197_82;
   assign m197_82 =10'b0;

   // m197_83 = W*in
   wire signed [9:0] m197_83;
   assign m197_83 =10'b0;

   // m197_84 = W*in
   wire signed [9:0] m197_84;
   assign m197_84 =10'b0;

   // m197_85 = W*in
   wire signed [9:0] m197_85;
   assign m197_85 ={ {5{neg197[5]}} , neg197[5:1] };

   // m197_86 = W*in
   wire signed [9:0] m197_86;
   assign m197_86 =10'b0;

   // m197_87 = W*in
   wire signed [9:0] m197_87;
   assign m197_87 =10'b0;

   // m197_88 = W*in
   wire signed [9:0] m197_88;
   assign m197_88 =10'b0;

   // m197_89 = W*in
   wire signed [9:0] m197_89;
   assign m197_89 =10'b0;

   // m197_90 = W*in
   wire signed [9:0] m197_90;
   assign m197_90 =10'b0;

   // m197_91 = W*in
   wire signed [9:0] m197_91;
   assign m197_91 =10'b0;

   // m197_92 = W*in
   wire signed [9:0] m197_92;
   assign m197_92 =10'b0;

   // m197_93 = W*in
   wire signed [9:0] m197_93;
   assign m197_93 =10'b0;

   // m197_94 = W*in
   wire signed [9:0] m197_94;
   assign m197_94 =10'b0;

   // m197_95 = W*in
   wire signed [9:0] m197_95;
   assign m197_95 =10'b0;

   // m197_96 = W*in
   wire signed [9:0] m197_96;
   assign m197_96 =10'b0;

   // m197_97 = W*in
   wire signed [9:0] m197_97;
   assign m197_97 =10'b0;

   // m197_98 = W*in
   wire signed [9:0] m197_98;
   assign m197_98 =10'b0;

   // m197_99 = W*in
   wire signed [9:0] m197_99;
   assign m197_99 =10'b0;

   // m197_100 = W*in
   wire signed [9:0] m197_100;
   assign m197_100 =10'b0;

   // m197_101 = W*in
   wire signed [9:0] m197_101;
   assign m197_101 =10'b0;

   // m197_102 = W*in
   wire signed [9:0] m197_102;
   assign m197_102 =10'b0;

   // m197_103 = W*in
   wire signed [9:0] m197_103;
   assign m197_103 =10'b0;

   // m197_104 = W*in
   wire signed [9:0] m197_104;
   assign m197_104 =10'b0;

   // m197_105 = W*in
   wire signed [9:0] m197_105;
   assign m197_105 =10'b0;

   // m197_106 = W*in
   wire signed [9:0] m197_106;
   assign m197_106 =10'b0;

   // m197_107 = W*in
   wire signed [9:0] m197_107;
   assign m197_107 =10'b0;

   // m197_108 = W*in
   wire signed [9:0] m197_108;
   assign m197_108 =10'b0;

   // m197_109 = W*in
   wire signed [9:0] m197_109;
   assign m197_109 =10'b0;

   // m197_110 = W*in
   wire signed [9:0] m197_110;
   assign m197_110 =10'b0;

   // m197_111 = W*in
   wire signed [9:0] m197_111;
   assign m197_111 =10'b0;

   // m197_112 = W*in
   wire signed [9:0] m197_112;
   assign m197_112 =10'b0;

   // m197_113 = W*in
   wire signed [9:0] m197_113;
   assign m197_113 =10'b0;

   // m197_114 = W*in
   wire signed [9:0] m197_114;
   assign m197_114 =10'b0;

   // m197_115 = W*in
   wire signed [9:0] m197_115;
   assign m197_115 ={ {5{in197[5]}} , in197[5:1] };

   // m197_116 = W*in
   wire signed [9:0] m197_116;
   assign m197_116 =10'b0;

   // m197_117 = W*in
   wire signed [9:0] m197_117;
   assign m197_117 =10'b0;

   // m198_1 = W*in
   wire signed [9:0] m198_1;
   assign m198_1 =10'b0;

   // m198_2 = W*in
   wire signed [9:0] m198_2;
   assign m198_2 =10'b0;

   // m198_3 = W*in
   wire signed [9:0] m198_3;
   assign m198_3 =10'b0;

   // m198_4 = W*in
   wire signed [9:0] m198_4;
   assign m198_4 =10'b0;

   // m198_5 = W*in
   wire signed [9:0] m198_5;
   assign m198_5 =10'b0;

   // m198_6 = W*in
   wire signed [9:0] m198_6;
   assign m198_6 =10'b0;

   // m198_7 = W*in
   wire signed [9:0] m198_7;
   assign m198_7 =10'b0;

   // m198_8 = W*in
   wire signed [9:0] m198_8;
   assign m198_8 =10'b0;

   // m198_9 = W*in
   wire signed [9:0] m198_9;
   assign m198_9 =10'b0;

   // m198_10 = W*in
   wire signed [9:0] m198_10;
   assign m198_10 =10'b0;

   // m198_11 = W*in
   wire signed [9:0] m198_11;
   assign m198_11 =10'b0;

   // m198_12 = W*in
   wire signed [9:0] m198_12;
   assign m198_12 =10'b0;

   // m198_13 = W*in
   wire signed [9:0] m198_13;
   assign m198_13 =10'b0;

   // m198_14 = W*in
   wire signed [9:0] m198_14;
   assign m198_14 =10'b0;

   // m198_15 = W*in
   wire signed [9:0] m198_15;
   assign m198_15 =10'b0;

   // m198_16 = W*in
   wire signed [9:0] m198_16;
   assign m198_16 =10'b0;

   // m198_17 = W*in
   wire signed [9:0] m198_17;
   assign m198_17 =10'b0;

   // m198_18 = W*in
   wire signed [9:0] m198_18;
   assign m198_18 =10'b0;

   // m198_19 = W*in
   wire signed [9:0] m198_19;
   assign m198_19 ={ {5{neg198[5]}} , neg198[5:1] };

   // m198_20 = W*in
   wire signed [9:0] m198_20;
   assign m198_20 =10'b0;

   // m198_21 = W*in
   wire signed [9:0] m198_21;
   assign m198_21 =10'b0;

   // m198_22 = W*in
   wire signed [9:0] m198_22;
   assign m198_22 =10'b0;

   // m198_23 = W*in
   wire signed [9:0] m198_23;
   assign m198_23 =10'b0;

   // m198_24 = W*in
   wire signed [9:0] m198_24;
   assign m198_24 =10'b0;

   // m198_25 = W*in
   wire signed [9:0] m198_25;
   assign m198_25 =10'b0;

   // m198_26 = W*in
   wire signed [9:0] m198_26;
   assign m198_26 ={ {5{in198[5]}} , in198[5:1] };

   // m198_27 = W*in
   wire signed [9:0] m198_27;
   assign m198_27 ={ {5{in198[5]}} , in198[5:1] };

   // m198_28 = W*in
   wire signed [9:0] m198_28;
   assign m198_28 =10'b0;

   // m198_29 = W*in
   wire signed [9:0] m198_29;
   assign m198_29 =10'b0;

   // m198_30 = W*in
   wire signed [9:0] m198_30;
   assign m198_30 =10'b0;

   // m198_31 = W*in
   wire signed [9:0] m198_31;
   assign m198_31 =10'b0;

   // m198_32 = W*in
   wire signed [9:0] m198_32;
   assign m198_32 =10'b0;

   // m198_33 = W*in
   wire signed [9:0] m198_33;
   assign m198_33 =10'b0;

   // m198_34 = W*in
   wire signed [9:0] m198_34;
   assign m198_34 =10'b0;

   // m198_35 = W*in
   wire signed [9:0] m198_35;
   assign m198_35 =10'b0;

   // m198_36 = W*in
   wire signed [9:0] m198_36;
   assign m198_36 =10'b0;

   // m198_37 = W*in
   wire signed [9:0] m198_37;
   assign m198_37 =10'b0;

   // m198_38 = W*in
   wire signed [9:0] m198_38;
   assign m198_38 =10'b0;

   // m198_39 = W*in
   wire signed [9:0] m198_39;
   assign m198_39 =10'b0;

   // m198_40 = W*in
   wire signed [9:0] m198_40;
   assign m198_40 =10'b0;

   // m198_41 = W*in
   wire signed [9:0] m198_41;
   assign m198_41 =10'b0;

   // m198_42 = W*in
   wire signed [9:0] m198_42;
   assign m198_42 =10'b0;

   // m198_43 = W*in
   wire signed [9:0] m198_43;
   assign m198_43 =10'b0;

   // m198_44 = W*in
   wire signed [9:0] m198_44;
   assign m198_44 =10'b0;

   // m198_45 = W*in
   wire signed [9:0] m198_45;
   assign m198_45 =10'b0;

   // m198_46 = W*in
   wire signed [9:0] m198_46;
   assign m198_46 =10'b0;

   // m198_47 = W*in
   wire signed [9:0] m198_47;
   assign m198_47 =10'b0;

   // m198_48 = W*in
   wire signed [9:0] m198_48;
   assign m198_48 =10'b0;

   // m198_49 = W*in
   wire signed [9:0] m198_49;
   assign m198_49 =10'b0;

   // m198_50 = W*in
   wire signed [9:0] m198_50;
   assign m198_50 =10'b0;

   // m198_51 = W*in
   wire signed [9:0] m198_51;
   assign m198_51 =10'b0;

   // m198_52 = W*in
   wire signed [9:0] m198_52;
   assign m198_52 =10'b0;

   // m198_53 = W*in
   wire signed [9:0] m198_53;
   assign m198_53 =10'b0;

   // m198_54 = W*in
   wire signed [9:0] m198_54;
   assign m198_54 =10'b0;

   // m198_55 = W*in
   wire signed [9:0] m198_55;
   assign m198_55 =10'b0;

   // m198_56 = W*in
   wire signed [9:0] m198_56;
   assign m198_56 =10'b0;

   // m198_57 = W*in
   wire signed [9:0] m198_57;
   assign m198_57 =10'b0;

   // m198_58 = W*in
   wire signed [9:0] m198_58;
   assign m198_58 =10'b0;

   // m198_59 = W*in
   wire signed [9:0] m198_59;
   assign m198_59 =10'b0;

   // m198_60 = W*in
   wire signed [9:0] m198_60;
   assign m198_60 ={ {4{in198[5]}} , in198[5:0] };

   // m198_61 = W*in
   wire signed [9:0] m198_61;
   assign m198_61 =10'b0;

   // m198_62 = W*in
   wire signed [9:0] m198_62;
   assign m198_62 =10'b0;

   // m198_63 = W*in
   wire signed [9:0] m198_63;
   assign m198_63 =10'b0;

   // m198_64 = W*in
   wire signed [9:0] m198_64;
   assign m198_64 =10'b0;

   // m198_65 = W*in
   wire signed [9:0] m198_65;
   assign m198_65 =10'b0;

   // m198_66 = W*in
   wire signed [9:0] m198_66;
   assign m198_66 =10'b0;

   // m198_67 = W*in
   wire signed [9:0] m198_67;
   assign m198_67 ={ {5{neg198[5]}} , neg198[5:1] };

   // m198_68 = W*in
   wire signed [9:0] m198_68;
   assign m198_68 =10'b0;

   // m198_69 = W*in
   wire signed [9:0] m198_69;
   assign m198_69 =10'b0;

   // m198_70 = W*in
   wire signed [9:0] m198_70;
   assign m198_70 =10'b0;

   // m198_71 = W*in
   wire signed [9:0] m198_71;
   assign m198_71 =10'b0;

   // m198_72 = W*in
   wire signed [9:0] m198_72;
   assign m198_72 ={ {5{in198[5]}} , in198[5:1] };

   // m198_73 = W*in
   wire signed [9:0] m198_73;
   assign m198_73 =10'b0;

   // m198_74 = W*in
   wire signed [9:0] m198_74;
   assign m198_74 =10'b0;

   // m198_75 = W*in
   wire signed [9:0] m198_75;
   assign m198_75 =10'b0;

   // m198_76 = W*in
   wire signed [9:0] m198_76;
   assign m198_76 =10'b0;

   // m198_77 = W*in
   wire signed [9:0] m198_77;
   assign m198_77 =10'b0;

   // m198_78 = W*in
   wire signed [9:0] m198_78;
   assign m198_78 =10'b0;

   // m198_79 = W*in
   wire signed [9:0] m198_79;
   assign m198_79 =10'b0;

   // m198_80 = W*in
   wire signed [9:0] m198_80;
   assign m198_80 =10'b0;

   // m198_81 = W*in
   wire signed [9:0] m198_81;
   assign m198_81 =10'b0;

   // m198_82 = W*in
   wire signed [9:0] m198_82;
   assign m198_82 =10'b0;

   // m198_83 = W*in
   wire signed [9:0] m198_83;
   assign m198_83 =10'b0;

   // m198_84 = W*in
   wire signed [9:0] m198_84;
   assign m198_84 =10'b0;

   // m198_85 = W*in
   wire signed [9:0] m198_85;
   assign m198_85 =10'b0;

   // m198_86 = W*in
   wire signed [9:0] m198_86;
   assign m198_86 =10'b0;

   // m198_87 = W*in
   wire signed [9:0] m198_87;
   assign m198_87 =10'b0;

   // m198_88 = W*in
   wire signed [9:0] m198_88;
   assign m198_88 =10'b0;

   // m198_89 = W*in
   wire signed [9:0] m198_89;
   assign m198_89 =10'b0;

   // m198_90 = W*in
   wire signed [9:0] m198_90;
   assign m198_90 =10'b0;

   // m198_91 = W*in
   wire signed [9:0] m198_91;
   assign m198_91 =10'b0;

   // m198_92 = W*in
   wire signed [9:0] m198_92;
   assign m198_92 =10'b0;

   // m198_93 = W*in
   wire signed [9:0] m198_93;
   assign m198_93 =10'b0;

   // m198_94 = W*in
   wire signed [9:0] m198_94;
   assign m198_94 =10'b0;

   // m198_95 = W*in
   wire signed [9:0] m198_95;
   assign m198_95 =10'b0;

   // m198_96 = W*in
   wire signed [9:0] m198_96;
   assign m198_96 =10'b0;

   // m198_97 = W*in
   wire signed [9:0] m198_97;
   assign m198_97 ={ {4{neg198[5]}} , neg198[5:0] };

   // m198_98 = W*in
   wire signed [9:0] m198_98;
   assign m198_98 =10'b0;

   // m198_99 = W*in
   wire signed [9:0] m198_99;
   assign m198_99 =10'b0;

   // m198_100 = W*in
   wire signed [9:0] m198_100;
   assign m198_100 =10'b0;

   // m198_101 = W*in
   wire signed [9:0] m198_101;
   assign m198_101 =10'b0;

   // m198_102 = W*in
   wire signed [9:0] m198_102;
   assign m198_102 =10'b0;

   // m198_103 = W*in
   wire signed [9:0] m198_103;
   assign m198_103 =10'b0;

   // m198_104 = W*in
   wire signed [9:0] m198_104;
   assign m198_104 =10'b0;

   // m198_105 = W*in
   wire signed [9:0] m198_105;
   assign m198_105 =10'b0;

   // m198_106 = W*in
   wire signed [9:0] m198_106;
   assign m198_106 =10'b0;

   // m198_107 = W*in
   wire signed [9:0] m198_107;
   assign m198_107 =10'b0;

   // m198_108 = W*in
   wire signed [9:0] m198_108;
   assign m198_108 =10'b0;

   // m198_109 = W*in
   wire signed [9:0] m198_109;
   assign m198_109 =10'b0;

   // m198_110 = W*in
   wire signed [9:0] m198_110;
   assign m198_110 =10'b0;

   // m198_111 = W*in
   wire signed [9:0] m198_111;
   assign m198_111 =10'b0;

   // m198_112 = W*in
   wire signed [9:0] m198_112;
   assign m198_112 =10'b0;

   // m198_113 = W*in
   wire signed [9:0] m198_113;
   assign m198_113 =10'b0;

   // m198_114 = W*in
   wire signed [9:0] m198_114;
   assign m198_114 =10'b0;

   // m198_115 = W*in
   wire signed [9:0] m198_115;
   assign m198_115 =10'b0;

   // m198_116 = W*in
   wire signed [9:0] m198_116;
   assign m198_116 =10'b0;

   // m198_117 = W*in
   wire signed [9:0] m198_117;
   assign m198_117 =10'b0;

   // m199_1 = W*in
   wire signed [9:0] m199_1;
   assign m199_1 =10'b0;

   // m199_2 = W*in
   wire signed [9:0] m199_2;
   assign m199_2 =10'b0;

   // m199_3 = W*in
   wire signed [9:0] m199_3;
   assign m199_3 =10'b0;

   // m199_4 = W*in
   wire signed [9:0] m199_4;
   assign m199_4 =10'b0;

   // m199_5 = W*in
   wire signed [9:0] m199_5;
   assign m199_5 =10'b0;

   // m199_6 = W*in
   wire signed [9:0] m199_6;
   assign m199_6 =10'b0;

   // m199_7 = W*in
   wire signed [9:0] m199_7;
   assign m199_7 =10'b0;

   // m199_8 = W*in
   wire signed [9:0] m199_8;
   assign m199_8 =10'b0;

   // m199_9 = W*in
   wire signed [9:0] m199_9;
   assign m199_9 =10'b0;

   // m199_10 = W*in
   wire signed [9:0] m199_10;
   assign m199_10 =10'b0;

   // m199_11 = W*in
   wire signed [9:0] m199_11;
   assign m199_11 =10'b0;

   // m199_12 = W*in
   wire signed [9:0] m199_12;
   assign m199_12 =10'b0;

   // m199_13 = W*in
   wire signed [9:0] m199_13;
   assign m199_13 =10'b0;

   // m199_14 = W*in
   wire signed [9:0] m199_14;
   assign m199_14 =10'b0;

   // m199_15 = W*in
   wire signed [9:0] m199_15;
   assign m199_15 =10'b0;

   // m199_16 = W*in
   wire signed [9:0] m199_16;
   assign m199_16 =10'b0;

   // m199_17 = W*in
   wire signed [9:0] m199_17;
   assign m199_17 =10'b0;

   // m199_18 = W*in
   wire signed [9:0] m199_18;
   assign m199_18 ={ {5{neg199[5]}} , neg199[5:1] };

   // m199_19 = W*in
   wire signed [9:0] m199_19;
   assign m199_19 =10'b0;

   // m199_20 = W*in
   wire signed [9:0] m199_20;
   assign m199_20 ={ {5{in199[5]}} , in199[5:1] };

   // m199_21 = W*in
   wire signed [9:0] m199_21;
   assign m199_21 =10'b0;

   // m199_22 = W*in
   wire signed [9:0] m199_22;
   assign m199_22 =10'b0;

   // m199_23 = W*in
   wire signed [9:0] m199_23;
   assign m199_23 =10'b0;

   // m199_24 = W*in
   wire signed [9:0] m199_24;
   assign m199_24 =10'b0;

   // m199_25 = W*in
   wire signed [9:0] m199_25;
   assign m199_25 =10'b0;

   // m199_26 = W*in
   wire signed [9:0] m199_26;
   assign m199_26 =10'b0;

   // m199_27 = W*in
   wire signed [9:0] m199_27;
   assign m199_27 ={ {5{in199[5]}} , in199[5:1] };

   // m199_28 = W*in
   wire signed [9:0] m199_28;
   assign m199_28 ={ {5{in199[5]}} , in199[5:1] };

   // m199_29 = W*in
   wire signed [9:0] m199_29;
   assign m199_29 =10'b0;

   // m199_30 = W*in
   wire signed [9:0] m199_30;
   assign m199_30 =10'b0;

   // m199_31 = W*in
   wire signed [9:0] m199_31;
   assign m199_31 =10'b0;

   // m199_32 = W*in
   wire signed [9:0] m199_32;
   assign m199_32 =10'b0;

   // m199_33 = W*in
   wire signed [9:0] m199_33;
   assign m199_33 =10'b0;

   // m199_34 = W*in
   wire signed [9:0] m199_34;
   assign m199_34 ={ {5{in199[5]}} , in199[5:1] };

   // m199_35 = W*in
   wire signed [9:0] m199_35;
   assign m199_35 ={ {5{in199[5]}} , in199[5:1] };

   // m199_36 = W*in
   wire signed [9:0] m199_36;
   assign m199_36 =10'b0;

   // m199_37 = W*in
   wire signed [9:0] m199_37;
   assign m199_37 =10'b0;

   // m199_38 = W*in
   wire signed [9:0] m199_38;
   assign m199_38 =10'b0;

   // m199_39 = W*in
   wire signed [9:0] m199_39;
   assign m199_39 =10'b0;

   // m199_40 = W*in
   wire signed [9:0] m199_40;
   assign m199_40 =10'b0;

   // m199_41 = W*in
   wire signed [9:0] m199_41;
   assign m199_41 ={ {4{in199[5]}} , in199[5:0] };

   // m199_42 = W*in
   wire signed [9:0] m199_42;
   assign m199_42 ={ {4{neg199[5]}} , neg199[5:0] };

   // m199_43 = W*in
   wire signed [9:0] m199_43;
   assign m199_43 =10'b0;

   // m199_44 = W*in
   wire signed [9:0] m199_44;
   assign m199_44 =10'b0;

   // m199_45 = W*in
   wire signed [9:0] m199_45;
   assign m199_45 =10'b0;

   // m199_46 = W*in
   wire signed [9:0] m199_46;
   assign m199_46 =10'b0;

   // m199_47 = W*in
   wire signed [9:0] m199_47;
   assign m199_47 =10'b0;

   // m199_48 = W*in
   wire signed [9:0] m199_48;
   assign m199_48 =10'b0;

   // m199_49 = W*in
   wire signed [9:0] m199_49;
   assign m199_49 =10'b0;

   // m199_50 = W*in
   wire signed [9:0] m199_50;
   assign m199_50 =10'b0;

   // m199_51 = W*in
   wire signed [9:0] m199_51;
   assign m199_51 =10'b0;

   // m199_52 = W*in
   wire signed [9:0] m199_52;
   assign m199_52 =10'b0;

   // m199_53 = W*in
   wire signed [9:0] m199_53;
   assign m199_53 =10'b0;

   // m199_54 = W*in
   wire signed [9:0] m199_54;
   assign m199_54 =10'b0;

   // m199_55 = W*in
   wire signed [9:0] m199_55;
   assign m199_55 =10'b0;

   // m199_56 = W*in
   wire signed [9:0] m199_56;
   assign m199_56 =10'b0;

   // m199_57 = W*in
   wire signed [9:0] m199_57;
   assign m199_57 =10'b0;

   // m199_58 = W*in
   wire signed [9:0] m199_58;
   assign m199_58 =10'b0;

   // m199_59 = W*in
   wire signed [9:0] m199_59;
   assign m199_59 =10'b0;

   // m199_60 = W*in
   wire signed [9:0] m199_60;
   assign m199_60 =10'b0;

   // m199_61 = W*in
   wire signed [9:0] m199_61;
   assign m199_61 =10'b0;

   // m199_62 = W*in
   wire signed [9:0] m199_62;
   assign m199_62 =10'b0;

   // m199_63 = W*in
   wire signed [9:0] m199_63;
   assign m199_63 =10'b0;

   // m199_64 = W*in
   wire signed [9:0] m199_64;
   assign m199_64 =10'b0;

   // m199_65 = W*in
   wire signed [9:0] m199_65;
   assign m199_65 =10'b0;

   // m199_66 = W*in
   wire signed [9:0] m199_66;
   assign m199_66 =10'b0;

   // m199_67 = W*in
   wire signed [9:0] m199_67;
   assign m199_67 =10'b0;

   // m199_68 = W*in
   wire signed [9:0] m199_68;
   assign m199_68 =10'b0;

   // m199_69 = W*in
   wire signed [9:0] m199_69;
   assign m199_69 =10'b0;

   // m199_70 = W*in
   wire signed [9:0] m199_70;
   assign m199_70 =10'b0;

   // m199_71 = W*in
   wire signed [9:0] m199_71;
   assign m199_71 =10'b0;

   // m199_72 = W*in
   wire signed [9:0] m199_72;
   assign m199_72 =10'b0;

   // m199_73 = W*in
   wire signed [9:0] m199_73;
   assign m199_73 ={ {5{neg199[5]}} , neg199[5:1] };

   // m199_74 = W*in
   wire signed [9:0] m199_74;
   assign m199_74 =10'b0;

   // m199_75 = W*in
   wire signed [9:0] m199_75;
   assign m199_75 =10'b0;

   // m199_76 = W*in
   wire signed [9:0] m199_76;
   assign m199_76 =10'b0;

   // m199_77 = W*in
   wire signed [9:0] m199_77;
   assign m199_77 ={ {4{neg199[5]}} , neg199[5:0] };

   // m199_78 = W*in
   wire signed [9:0] m199_78;
   assign m199_78 =10'b0;

   // m199_79 = W*in
   wire signed [9:0] m199_79;
   assign m199_79 =10'b0;

   // m199_80 = W*in
   wire signed [9:0] m199_80;
   assign m199_80 =10'b0;

   // m199_81 = W*in
   wire signed [9:0] m199_81;
   assign m199_81 =10'b0;

   // m199_82 = W*in
   wire signed [9:0] m199_82;
   assign m199_82 =10'b0;

   // m199_83 = W*in
   wire signed [9:0] m199_83;
   assign m199_83 =10'b0;

   // m199_84 = W*in
   wire signed [9:0] m199_84;
   assign m199_84 =10'b0;

   // m199_85 = W*in
   wire signed [9:0] m199_85;
   assign m199_85 =10'b0;

   // m199_86 = W*in
   wire signed [9:0] m199_86;
   assign m199_86 =10'b0;

   // m199_87 = W*in
   wire signed [9:0] m199_87;
   assign m199_87 =10'b0;

   // m199_88 = W*in
   wire signed [9:0] m199_88;
   assign m199_88 =10'b0;

   // m199_89 = W*in
   wire signed [9:0] m199_89;
   assign m199_89 =10'b0;

   // m199_90 = W*in
   wire signed [9:0] m199_90;
   assign m199_90 =10'b0;

   // m199_91 = W*in
   wire signed [9:0] m199_91;
   assign m199_91 =10'b0;

   // m199_92 = W*in
   wire signed [9:0] m199_92;
   assign m199_92 =10'b0;

   // m199_93 = W*in
   wire signed [9:0] m199_93;
   assign m199_93 =10'b0;

   // m199_94 = W*in
   wire signed [9:0] m199_94;
   assign m199_94 =10'b0;

   // m199_95 = W*in
   wire signed [9:0] m199_95;
   assign m199_95 =10'b0;

   // m199_96 = W*in
   wire signed [9:0] m199_96;
   assign m199_96 =10'b0;

   // m199_97 = W*in
   wire signed [9:0] m199_97;
   assign m199_97 =10'b0;

   // m199_98 = W*in
   wire signed [9:0] m199_98;
   assign m199_98 =10'b0;

   // m199_99 = W*in
   wire signed [9:0] m199_99;
   assign m199_99 =10'b0;

   // m199_100 = W*in
   wire signed [9:0] m199_100;
   assign m199_100 =10'b0;

   // m199_101 = W*in
   wire signed [9:0] m199_101;
   assign m199_101 =10'b0;

   // m199_102 = W*in
   wire signed [9:0] m199_102;
   assign m199_102 =10'b0;

   // m199_103 = W*in
   wire signed [9:0] m199_103;
   assign m199_103 =10'b0;

   // m199_104 = W*in
   wire signed [9:0] m199_104;
   assign m199_104 =10'b0;

   // m199_105 = W*in
   wire signed [9:0] m199_105;
   assign m199_105 =10'b0;

   // m199_106 = W*in
   wire signed [9:0] m199_106;
   assign m199_106 =10'b0;

   // m199_107 = W*in
   wire signed [9:0] m199_107;
   assign m199_107 =10'b0;

   // m199_108 = W*in
   wire signed [9:0] m199_108;
   assign m199_108 ={ {5{in199[5]}} , in199[5:1] };

   // m199_109 = W*in
   wire signed [9:0] m199_109;
   assign m199_109 =10'b0;

   // m199_110 = W*in
   wire signed [9:0] m199_110;
   assign m199_110 =10'b0;

   // m199_111 = W*in
   wire signed [9:0] m199_111;
   assign m199_111 =10'b0;

   // m199_112 = W*in
   wire signed [9:0] m199_112;
   assign m199_112 =10'b0;

   // m199_113 = W*in
   wire signed [9:0] m199_113;
   assign m199_113 =10'b0;

   // m199_114 = W*in
   wire signed [9:0] m199_114;
   assign m199_114 =10'b0;

   // m199_115 = W*in
   wire signed [9:0] m199_115;
   assign m199_115 =10'b0;

   // m199_116 = W*in
   wire signed [9:0] m199_116;
   assign m199_116 ={ {4{in199[5]}} , in199[5:0] };

   // m199_117 = W*in
   wire signed [9:0] m199_117;
   assign m199_117 =10'b0;

   // m200_1 = W*in
   wire signed [9:0] m200_1;
   assign m200_1 =10'b0;

   // m200_2 = W*in
   wire signed [9:0] m200_2;
   assign m200_2 =10'b0;

   // m200_3 = W*in
   wire signed [9:0] m200_3;
   assign m200_3 =10'b0;

   // m200_4 = W*in
   wire signed [9:0] m200_4;
   assign m200_4 =10'b0;

   // m200_5 = W*in
   wire signed [9:0] m200_5;
   assign m200_5 =10'b0;

   // m200_6 = W*in
   wire signed [9:0] m200_6;
   assign m200_6 =10'b0;

   // m200_7 = W*in
   wire signed [9:0] m200_7;
   assign m200_7 =10'b0;

   // m200_8 = W*in
   wire signed [9:0] m200_8;
   assign m200_8 =10'b0;

   // m200_9 = W*in
   wire signed [9:0] m200_9;
   assign m200_9 =10'b0;

   // m200_10 = W*in
   wire signed [9:0] m200_10;
   assign m200_10 =10'b0;

   // m200_11 = W*in
   wire signed [9:0] m200_11;
   assign m200_11 =10'b0;

   // m200_12 = W*in
   wire signed [9:0] m200_12;
   assign m200_12 =10'b0;

   // m200_13 = W*in
   wire signed [9:0] m200_13;
   assign m200_13 =10'b0;

   // m200_14 = W*in
   wire signed [9:0] m200_14;
   assign m200_14 =10'b0;

   // m200_15 = W*in
   wire signed [9:0] m200_15;
   assign m200_15 =10'b0;

   // m200_16 = W*in
   wire signed [9:0] m200_16;
   assign m200_16 ={ {4{in200[5]}} , in200[5:0] };

   // m200_17 = W*in
   wire signed [9:0] m200_17;
   assign m200_17 =10'b0;

   // m200_18 = W*in
   wire signed [9:0] m200_18;
   assign m200_18 =10'b0;

   // m200_19 = W*in
   wire signed [9:0] m200_19;
   assign m200_19 =10'b0;

   // m200_20 = W*in
   wire signed [9:0] m200_20;
   assign m200_20 =10'b0;

   // m200_21 = W*in
   wire signed [9:0] m200_21;
   assign m200_21 =10'b0;

   // m200_22 = W*in
   wire signed [9:0] m200_22;
   assign m200_22 =10'b0;

   // m200_23 = W*in
   wire signed [9:0] m200_23;
   assign m200_23 ={ {5{neg200[5]}} , neg200[5:1] };

   // m200_24 = W*in
   wire signed [9:0] m200_24;
   assign m200_24 =10'b0;

   // m200_25 = W*in
   wire signed [9:0] m200_25;
   assign m200_25 =10'b0;

   // m200_26 = W*in
   wire signed [9:0] m200_26;
   assign m200_26 ={ {5{neg200[5]}} , neg200[5:1] };

   // m200_27 = W*in
   wire signed [9:0] m200_27;
   assign m200_27 =10'b0;

   // m200_28 = W*in
   wire signed [9:0] m200_28;
   assign m200_28 ={ {5{in200[5]}} , in200[5:1] };

   // m200_29 = W*in
   wire signed [9:0] m200_29;
   assign m200_29 =10'b0;

   // m200_30 = W*in
   wire signed [9:0] m200_30;
   assign m200_30 =10'b0;

   // m200_31 = W*in
   wire signed [9:0] m200_31;
   assign m200_31 =10'b0;

   // m200_32 = W*in
   wire signed [9:0] m200_32;
   assign m200_32 =10'b0;

   // m200_33 = W*in
   wire signed [9:0] m200_33;
   assign m200_33 =10'b0;

   // m200_34 = W*in
   wire signed [9:0] m200_34;
   assign m200_34 ={ {4{neg200[5]}} , neg200[5:0] };

   // m200_35 = W*in
   wire signed [9:0] m200_35;
   assign m200_35 ={ {5{in200[5]}} , in200[5:1] };

   // m200_36 = W*in
   wire signed [9:0] m200_36;
   assign m200_36 =10'b0;

   // m200_37 = W*in
   wire signed [9:0] m200_37;
   assign m200_37 =10'b0;

   // m200_38 = W*in
   wire signed [9:0] m200_38;
   assign m200_38 =10'b0;

   // m200_39 = W*in
   wire signed [9:0] m200_39;
   assign m200_39 =10'b0;

   // m200_40 = W*in
   wire signed [9:0] m200_40;
   assign m200_40 =10'b0;

   // m200_41 = W*in
   wire signed [9:0] m200_41;
   assign m200_41 =10'b0;

   // m200_42 = W*in
   wire signed [9:0] m200_42;
   assign m200_42 =10'b0;

   // m200_43 = W*in
   wire signed [9:0] m200_43;
   assign m200_43 =10'b0;

   // m200_44 = W*in
   wire signed [9:0] m200_44;
   assign m200_44 =10'b0;

   // m200_45 = W*in
   wire signed [9:0] m200_45;
   assign m200_45 =10'b0;

   // m200_46 = W*in
   wire signed [9:0] m200_46;
   assign m200_46 =10'b0;

   // m200_47 = W*in
   wire signed [9:0] m200_47;
   assign m200_47 =10'b0;

   // m200_48 = W*in
   wire signed [9:0] m200_48;
   assign m200_48 =10'b0;

   // m200_49 = W*in
   wire signed [9:0] m200_49;
   assign m200_49 =10'b0;

   // m200_50 = W*in
   wire signed [9:0] m200_50;
   assign m200_50 =10'b0;

   // m200_51 = W*in
   wire signed [9:0] m200_51;
   assign m200_51 =10'b0;

   // m200_52 = W*in
   wire signed [9:0] m200_52;
   assign m200_52 =10'b0;

   // m200_53 = W*in
   wire signed [9:0] m200_53;
   assign m200_53 =10'b0;

   // m200_54 = W*in
   wire signed [9:0] m200_54;
   assign m200_54 =10'b0;

   // m200_55 = W*in
   wire signed [9:0] m200_55;
   assign m200_55 =10'b0;

   // m200_56 = W*in
   wire signed [9:0] m200_56;
   assign m200_56 ={ {4{in200[5]}} , in200[5:0] };

   // m200_57 = W*in
   wire signed [9:0] m200_57;
   assign m200_57 =10'b0;

   // m200_58 = W*in
   wire signed [9:0] m200_58;
   assign m200_58 =10'b0;

   // m200_59 = W*in
   wire signed [9:0] m200_59;
   assign m200_59 =10'b0;

   // m200_60 = W*in
   wire signed [9:0] m200_60;
   assign m200_60 =10'b0;

   // m200_61 = W*in
   wire signed [9:0] m200_61;
   assign m200_61 =10'b0;

   // m200_62 = W*in
   wire signed [9:0] m200_62;
   assign m200_62 =10'b0;

   // m200_63 = W*in
   wire signed [9:0] m200_63;
   assign m200_63 =10'b0;

   // m200_64 = W*in
   wire signed [9:0] m200_64;
   assign m200_64 =10'b0;

   // m200_65 = W*in
   wire signed [9:0] m200_65;
   assign m200_65 =10'b0;

   // m200_66 = W*in
   wire signed [9:0] m200_66;
   assign m200_66 ={ {5{in200[5]}} , in200[5:1] };

   // m200_67 = W*in
   wire signed [9:0] m200_67;
   assign m200_67 =10'b0;

   // m200_68 = W*in
   wire signed [9:0] m200_68;
   assign m200_68 =10'b0;

   // m200_69 = W*in
   wire signed [9:0] m200_69;
   assign m200_69 =10'b0;

   // m200_70 = W*in
   wire signed [9:0] m200_70;
   assign m200_70 ={ {5{neg200[5]}} , neg200[5:1] };

   // m200_71 = W*in
   wire signed [9:0] m200_71;
   assign m200_71 ={ {5{neg200[5]}} , neg200[5:1] };

   // m200_72 = W*in
   wire signed [9:0] m200_72;
   assign m200_72 ={ {5{neg200[5]}} , neg200[5:1] };

   // m200_73 = W*in
   wire signed [9:0] m200_73;
   assign m200_73 =10'b0;

   // m200_74 = W*in
   wire signed [9:0] m200_74;
   assign m200_74 =10'b0;

   // m200_75 = W*in
   wire signed [9:0] m200_75;
   assign m200_75 =10'b0;

   // m200_76 = W*in
   wire signed [9:0] m200_76;
   assign m200_76 =10'b0;

   // m200_77 = W*in
   wire signed [9:0] m200_77;
   assign m200_77 =10'b0;

   // m200_78 = W*in
   wire signed [9:0] m200_78;
   assign m200_78 =10'b0;

   // m200_79 = W*in
   wire signed [9:0] m200_79;
   assign m200_79 =10'b0;

   // m200_80 = W*in
   wire signed [9:0] m200_80;
   assign m200_80 =10'b0;

   // m200_81 = W*in
   wire signed [9:0] m200_81;
   assign m200_81 =10'b0;

   // m200_82 = W*in
   wire signed [9:0] m200_82;
   assign m200_82 =10'b0;

   // m200_83 = W*in
   wire signed [9:0] m200_83;
   assign m200_83 =10'b0;

   // m200_84 = W*in
   wire signed [9:0] m200_84;
   assign m200_84 =10'b0;

   // m200_85 = W*in
   wire signed [9:0] m200_85;
   assign m200_85 =10'b0;

   // m200_86 = W*in
   wire signed [9:0] m200_86;
   assign m200_86 =10'b0;

   // m200_87 = W*in
   wire signed [9:0] m200_87;
   assign m200_87 =10'b0;

   // m200_88 = W*in
   wire signed [9:0] m200_88;
   assign m200_88 =10'b0;

   // m200_89 = W*in
   wire signed [9:0] m200_89;
   assign m200_89 =10'b0;

   // m200_90 = W*in
   wire signed [9:0] m200_90;
   assign m200_90 =10'b0;

   // m200_91 = W*in
   wire signed [9:0] m200_91;
   assign m200_91 ={ {4{in200[5]}} , in200[5:0] };

   // m200_92 = W*in
   wire signed [9:0] m200_92;
   assign m200_92 =10'b0;

   // m200_93 = W*in
   wire signed [9:0] m200_93;
   assign m200_93 =10'b0;

   // m200_94 = W*in
   wire signed [9:0] m200_94;
   assign m200_94 =10'b0;

   // m200_95 = W*in
   wire signed [9:0] m200_95;
   assign m200_95 =10'b0;

   // m200_96 = W*in
   wire signed [9:0] m200_96;
   assign m200_96 =10'b0;

   // m200_97 = W*in
   wire signed [9:0] m200_97;
   assign m200_97 =10'b0;

   // m200_98 = W*in
   wire signed [9:0] m200_98;
   assign m200_98 =10'b0;

   // m200_99 = W*in
   wire signed [9:0] m200_99;
   assign m200_99 =10'b0;

   // m200_100 = W*in
   wire signed [9:0] m200_100;
   assign m200_100 =10'b0;

   // m200_101 = W*in
   wire signed [9:0] m200_101;
   assign m200_101 =10'b0;

   // m200_102 = W*in
   wire signed [9:0] m200_102;
   assign m200_102 =10'b0;

   // m200_103 = W*in
   wire signed [9:0] m200_103;
   assign m200_103 =10'b0;

   // m200_104 = W*in
   wire signed [9:0] m200_104;
   assign m200_104 =10'b0;

   // m200_105 = W*in
   wire signed [9:0] m200_105;
   assign m200_105 =10'b0;

   // m200_106 = W*in
   wire signed [9:0] m200_106;
   assign m200_106 =10'b0;

   // m200_107 = W*in
   wire signed [9:0] m200_107;
   assign m200_107 =10'b0;

   // m200_108 = W*in
   wire signed [9:0] m200_108;
   assign m200_108 =10'b0;

   // m200_109 = W*in
   wire signed [9:0] m200_109;
   assign m200_109 =10'b0;

   // m200_110 = W*in
   wire signed [9:0] m200_110;
   assign m200_110 =10'b0;

   // m200_111 = W*in
   wire signed [9:0] m200_111;
   assign m200_111 =10'b0;

   // m200_112 = W*in
   wire signed [9:0] m200_112;
   assign m200_112 =10'b0;

   // m200_113 = W*in
   wire signed [9:0] m200_113;
   assign m200_113 =10'b0;

   // m200_114 = W*in
   wire signed [9:0] m200_114;
   assign m200_114 =10'b0;

   // m200_115 = W*in
   wire signed [9:0] m200_115;
   assign m200_115 =10'b0;

   // m200_116 = W*in
   wire signed [9:0] m200_116;
   assign m200_116 =10'b0;

   // m200_117 = W*in
   wire signed [9:0] m200_117;
   assign m200_117 =10'b0;

   // m201_1 = W*in
   wire signed [9:0] m201_1;
   assign m201_1 =10'b0;

   // m201_2 = W*in
   wire signed [9:0] m201_2;
   assign m201_2 =10'b0;

   // m201_3 = W*in
   wire signed [9:0] m201_3;
   assign m201_3 =10'b0;

   // m201_4 = W*in
   wire signed [9:0] m201_4;
   assign m201_4 =10'b0;

   // m201_5 = W*in
   wire signed [9:0] m201_5;
   assign m201_5 =10'b0;

   // m201_6 = W*in
   wire signed [9:0] m201_6;
   assign m201_6 =10'b0;

   // m201_7 = W*in
   wire signed [9:0] m201_7;
   assign m201_7 =10'b0;

   // m201_8 = W*in
   wire signed [9:0] m201_8;
   assign m201_8 =10'b0;

   // m201_9 = W*in
   wire signed [9:0] m201_9;
   assign m201_9 =10'b0;

   // m201_10 = W*in
   wire signed [9:0] m201_10;
   assign m201_10 =10'b0;

   // m201_11 = W*in
   wire signed [9:0] m201_11;
   assign m201_11 =10'b0;

   // m201_12 = W*in
   wire signed [9:0] m201_12;
   assign m201_12 =10'b0;

   // m201_13 = W*in
   wire signed [9:0] m201_13;
   assign m201_13 =10'b0;

   // m201_14 = W*in
   wire signed [9:0] m201_14;
   assign m201_14 =10'b0;

   // m201_15 = W*in
   wire signed [9:0] m201_15;
   assign m201_15 =10'b0;

   // m201_16 = W*in
   wire signed [9:0] m201_16;
   assign m201_16 =10'b0;

   // m201_17 = W*in
   wire signed [9:0] m201_17;
   assign m201_17 =10'b0;

   // m201_18 = W*in
   wire signed [9:0] m201_18;
   assign m201_18 =10'b0;

   // m201_19 = W*in
   wire signed [9:0] m201_19;
   assign m201_19 =10'b0;

   // m201_20 = W*in
   wire signed [9:0] m201_20;
   assign m201_20 =10'b0;

   // m201_21 = W*in
   wire signed [9:0] m201_21;
   assign m201_21 =10'b0;

   // m201_22 = W*in
   wire signed [9:0] m201_22;
   assign m201_22 =10'b0;

   // m201_23 = W*in
   wire signed [9:0] m201_23;
   assign m201_23 =10'b0;

   // m201_24 = W*in
   wire signed [9:0] m201_24;
   assign m201_24 =10'b0;

   // m201_25 = W*in
   wire signed [9:0] m201_25;
   assign m201_25 =10'b0;

   // m201_26 = W*in
   wire signed [9:0] m201_26;
   assign m201_26 =10'b0;

   // m201_27 = W*in
   wire signed [9:0] m201_27;
   assign m201_27 =10'b0;

   // m201_28 = W*in
   wire signed [9:0] m201_28;
   assign m201_28 =10'b0;

   // m201_29 = W*in
   wire signed [9:0] m201_29;
   assign m201_29 =10'b0;

   // m201_30 = W*in
   wire signed [9:0] m201_30;
   assign m201_30 =10'b0;

   // m201_31 = W*in
   wire signed [9:0] m201_31;
   assign m201_31 =10'b0;

   // m201_32 = W*in
   wire signed [9:0] m201_32;
   assign m201_32 =10'b0;

   // m201_33 = W*in
   wire signed [9:0] m201_33;
   assign m201_33 =10'b0;

   // m201_34 = W*in
   wire signed [9:0] m201_34;
   assign m201_34 =10'b0;

   // m201_35 = W*in
   wire signed [9:0] m201_35;
   assign m201_35 =10'b0;

   // m201_36 = W*in
   wire signed [9:0] m201_36;
   assign m201_36 ={ {5{in201[5]}} , in201[5:1] };

   // m201_37 = W*in
   wire signed [9:0] m201_37;
   assign m201_37 =10'b0;

   // m201_38 = W*in
   wire signed [9:0] m201_38;
   assign m201_38 =10'b0;

   // m201_39 = W*in
   wire signed [9:0] m201_39;
   assign m201_39 =10'b0;

   // m201_40 = W*in
   wire signed [9:0] m201_40;
   assign m201_40 =10'b0;

   // m201_41 = W*in
   wire signed [9:0] m201_41;
   assign m201_41 =10'b0;

   // m201_42 = W*in
   wire signed [9:0] m201_42;
   assign m201_42 =10'b0;

   // m201_43 = W*in
   wire signed [9:0] m201_43;
   assign m201_43 =10'b0;

   // m201_44 = W*in
   wire signed [9:0] m201_44;
   assign m201_44 =10'b0;

   // m201_45 = W*in
   wire signed [9:0] m201_45;
   assign m201_45 =10'b0;

   // m201_46 = W*in
   wire signed [9:0] m201_46;
   assign m201_46 =10'b0;

   // m201_47 = W*in
   wire signed [9:0] m201_47;
   assign m201_47 =10'b0;

   // m201_48 = W*in
   wire signed [9:0] m201_48;
   assign m201_48 =10'b0;

   // m201_49 = W*in
   wire signed [9:0] m201_49;
   assign m201_49 =10'b0;

   // m201_50 = W*in
   wire signed [9:0] m201_50;
   assign m201_50 =10'b0;

   // m201_51 = W*in
   wire signed [9:0] m201_51;
   assign m201_51 =10'b0;

   // m201_52 = W*in
   wire signed [9:0] m201_52;
   assign m201_52 =10'b0;

   // m201_53 = W*in
   wire signed [9:0] m201_53;
   assign m201_53 =10'b0;

   // m201_54 = W*in
   wire signed [9:0] m201_54;
   assign m201_54 =10'b0;

   // m201_55 = W*in
   wire signed [9:0] m201_55;
   assign m201_55 =10'b0;

   // m201_56 = W*in
   wire signed [9:0] m201_56;
   assign m201_56 =10'b0;

   // m201_57 = W*in
   wire signed [9:0] m201_57;
   assign m201_57 =10'b0;

   // m201_58 = W*in
   wire signed [9:0] m201_58;
   assign m201_58 =10'b0;

   // m201_59 = W*in
   wire signed [9:0] m201_59;
   assign m201_59 =10'b0;

   // m201_60 = W*in
   wire signed [9:0] m201_60;
   assign m201_60 =10'b0;

   // m201_61 = W*in
   wire signed [9:0] m201_61;
   assign m201_61 =10'b0;

   // m201_62 = W*in
   wire signed [9:0] m201_62;
   assign m201_62 =10'b0;

   // m201_63 = W*in
   wire signed [9:0] m201_63;
   assign m201_63 =10'b0;

   // m201_64 = W*in
   wire signed [9:0] m201_64;
   assign m201_64 ={ {5{neg201[5]}} , neg201[5:1] };

   // m201_65 = W*in
   wire signed [9:0] m201_65;
   assign m201_65 =10'b0;

   // m201_66 = W*in
   wire signed [9:0] m201_66;
   assign m201_66 =10'b0;

   // m201_67 = W*in
   wire signed [9:0] m201_67;
   assign m201_67 =10'b0;

   // m201_68 = W*in
   wire signed [9:0] m201_68;
   assign m201_68 =10'b0;

   // m201_69 = W*in
   wire signed [9:0] m201_69;
   assign m201_69 =10'b0;

   // m201_70 = W*in
   wire signed [9:0] m201_70;
   assign m201_70 =10'b0;

   // m201_71 = W*in
   wire signed [9:0] m201_71;
   assign m201_71 =10'b0;

   // m201_72 = W*in
   wire signed [9:0] m201_72;
   assign m201_72 =10'b0;

   // m201_73 = W*in
   wire signed [9:0] m201_73;
   assign m201_73 =10'b0;

   // m201_74 = W*in
   wire signed [9:0] m201_74;
   assign m201_74 =10'b0;

   // m201_75 = W*in
   wire signed [9:0] m201_75;
   assign m201_75 =10'b0;

   // m201_76 = W*in
   wire signed [9:0] m201_76;
   assign m201_76 =10'b0;

   // m201_77 = W*in
   wire signed [9:0] m201_77;
   assign m201_77 =10'b0;

   // m201_78 = W*in
   wire signed [9:0] m201_78;
   assign m201_78 =10'b0;

   // m201_79 = W*in
   wire signed [9:0] m201_79;
   assign m201_79 =10'b0;

   // m201_80 = W*in
   wire signed [9:0] m201_80;
   assign m201_80 =10'b0;

   // m201_81 = W*in
   wire signed [9:0] m201_81;
   assign m201_81 =10'b0;

   // m201_82 = W*in
   wire signed [9:0] m201_82;
   assign m201_82 =10'b0;

   // m201_83 = W*in
   wire signed [9:0] m201_83;
   assign m201_83 =10'b0;

   // m201_84 = W*in
   wire signed [9:0] m201_84;
   assign m201_84 =10'b0;

   // m201_85 = W*in
   wire signed [9:0] m201_85;
   assign m201_85 =10'b0;

   // m201_86 = W*in
   wire signed [9:0] m201_86;
   assign m201_86 =10'b0;

   // m201_87 = W*in
   wire signed [9:0] m201_87;
   assign m201_87 =10'b0;

   // m201_88 = W*in
   wire signed [9:0] m201_88;
   assign m201_88 =10'b0;

   // m201_89 = W*in
   wire signed [9:0] m201_89;
   assign m201_89 =10'b0;

   // m201_90 = W*in
   wire signed [9:0] m201_90;
   assign m201_90 =10'b0;

   // m201_91 = W*in
   wire signed [9:0] m201_91;
   assign m201_91 =10'b0;

   // m201_92 = W*in
   wire signed [9:0] m201_92;
   assign m201_92 =10'b0;

   // m201_93 = W*in
   wire signed [9:0] m201_93;
   assign m201_93 =10'b0;

   // m201_94 = W*in
   wire signed [9:0] m201_94;
   assign m201_94 =10'b0;

   // m201_95 = W*in
   wire signed [9:0] m201_95;
   assign m201_95 =10'b0;

   // m201_96 = W*in
   wire signed [9:0] m201_96;
   assign m201_96 =10'b0;

   // m201_97 = W*in
   wire signed [9:0] m201_97;
   assign m201_97 =10'b0;

   // m201_98 = W*in
   wire signed [9:0] m201_98;
   assign m201_98 =10'b0;

   // m201_99 = W*in
   wire signed [9:0] m201_99;
   assign m201_99 =10'b0;

   // m201_100 = W*in
   wire signed [9:0] m201_100;
   assign m201_100 =10'b0;

   // m201_101 = W*in
   wire signed [9:0] m201_101;
   assign m201_101 =10'b0;

   // m201_102 = W*in
   wire signed [9:0] m201_102;
   assign m201_102 =10'b0;

   // m201_103 = W*in
   wire signed [9:0] m201_103;
   assign m201_103 =10'b0;

   // m201_104 = W*in
   wire signed [9:0] m201_104;
   assign m201_104 =10'b0;

   // m201_105 = W*in
   wire signed [9:0] m201_105;
   assign m201_105 =10'b0;

   // m201_106 = W*in
   wire signed [9:0] m201_106;
   assign m201_106 =10'b0;

   // m201_107 = W*in
   wire signed [9:0] m201_107;
   assign m201_107 =10'b0;

   // m201_108 = W*in
   wire signed [9:0] m201_108;
   assign m201_108 =10'b0;

   // m201_109 = W*in
   wire signed [9:0] m201_109;
   assign m201_109 =10'b0;

   // m201_110 = W*in
   wire signed [9:0] m201_110;
   assign m201_110 =10'b0;

   // m201_111 = W*in
   wire signed [9:0] m201_111;
   assign m201_111 =10'b0;

   // m201_112 = W*in
   wire signed [9:0] m201_112;
   assign m201_112 =10'b0;

   // m201_113 = W*in
   wire signed [9:0] m201_113;
   assign m201_113 =10'b0;

   // m201_114 = W*in
   wire signed [9:0] m201_114;
   assign m201_114 =10'b0;

   // m201_115 = W*in
   wire signed [9:0] m201_115;
   assign m201_115 =10'b0;

   // m201_116 = W*in
   wire signed [9:0] m201_116;
   assign m201_116 =10'b0;

   // m201_117 = W*in
   wire signed [9:0] m201_117;
   assign m201_117 =10'b0;

   // m202_1 = W*in
   wire signed [9:0] m202_1;
   assign m202_1 =10'b0;

   // m202_2 = W*in
   wire signed [9:0] m202_2;
   assign m202_2 =10'b0;

   // m202_3 = W*in
   wire signed [9:0] m202_3;
   assign m202_3 =10'b0;

   // m202_4 = W*in
   wire signed [9:0] m202_4;
   assign m202_4 =10'b0;

   // m202_5 = W*in
   wire signed [9:0] m202_5;
   assign m202_5 =10'b0;

   // m202_6 = W*in
   wire signed [9:0] m202_6;
   assign m202_6 =10'b0;

   // m202_7 = W*in
   wire signed [9:0] m202_7;
   assign m202_7 =10'b0;

   // m202_8 = W*in
   wire signed [9:0] m202_8;
   assign m202_8 =10'b0;

   // m202_9 = W*in
   wire signed [9:0] m202_9;
   assign m202_9 =10'b0;

   // m202_10 = W*in
   wire signed [9:0] m202_10;
   assign m202_10 =10'b0;

   // m202_11 = W*in
   wire signed [9:0] m202_11;
   assign m202_11 =10'b0;

   // m202_12 = W*in
   wire signed [9:0] m202_12;
   assign m202_12 =10'b0;

   // m202_13 = W*in
   wire signed [9:0] m202_13;
   assign m202_13 =10'b0;

   // m202_14 = W*in
   wire signed [9:0] m202_14;
   assign m202_14 =10'b0;

   // m202_15 = W*in
   wire signed [9:0] m202_15;
   assign m202_15 =10'b0;

   // m202_16 = W*in
   wire signed [9:0] m202_16;
   assign m202_16 =10'b0;

   // m202_17 = W*in
   wire signed [9:0] m202_17;
   assign m202_17 =10'b0;

   // m202_18 = W*in
   wire signed [9:0] m202_18;
   assign m202_18 =10'b0;

   // m202_19 = W*in
   wire signed [9:0] m202_19;
   assign m202_19 =10'b0;

   // m202_20 = W*in
   wire signed [9:0] m202_20;
   assign m202_20 ={ {5{in202[5]}} , in202[5:1] };

   // m202_21 = W*in
   wire signed [9:0] m202_21;
   assign m202_21 =10'b0;

   // m202_22 = W*in
   wire signed [9:0] m202_22;
   assign m202_22 ={ {5{in202[5]}} , in202[5:1] };

   // m202_23 = W*in
   wire signed [9:0] m202_23;
   assign m202_23 =10'b0;

   // m202_24 = W*in
   wire signed [9:0] m202_24;
   assign m202_24 =10'b0;

   // m202_25 = W*in
   wire signed [9:0] m202_25;
   assign m202_25 =10'b0;

   // m202_26 = W*in
   wire signed [9:0] m202_26;
   assign m202_26 =10'b0;

   // m202_27 = W*in
   wire signed [9:0] m202_27;
   assign m202_27 ={ {5{in202[5]}} , in202[5:1] };

   // m202_28 = W*in
   wire signed [9:0] m202_28;
   assign m202_28 =10'b0;

   // m202_29 = W*in
   wire signed [9:0] m202_29;
   assign m202_29 =10'b0;

   // m202_30 = W*in
   wire signed [9:0] m202_30;
   assign m202_30 =10'b0;

   // m202_31 = W*in
   wire signed [9:0] m202_31;
   assign m202_31 =10'b0;

   // m202_32 = W*in
   wire signed [9:0] m202_32;
   assign m202_32 =10'b0;

   // m202_33 = W*in
   wire signed [9:0] m202_33;
   assign m202_33 =10'b0;

   // m202_34 = W*in
   wire signed [9:0] m202_34;
   assign m202_34 =10'b0;

   // m202_35 = W*in
   wire signed [9:0] m202_35;
   assign m202_35 =10'b0;

   // m202_36 = W*in
   wire signed [9:0] m202_36;
   assign m202_36 =10'b0;

   // m202_37 = W*in
   wire signed [9:0] m202_37;
   assign m202_37 =10'b0;

   // m202_38 = W*in
   wire signed [9:0] m202_38;
   assign m202_38 =10'b0;

   // m202_39 = W*in
   wire signed [9:0] m202_39;
   assign m202_39 =10'b0;

   // m202_40 = W*in
   wire signed [9:0] m202_40;
   assign m202_40 =10'b0;

   // m202_41 = W*in
   wire signed [9:0] m202_41;
   assign m202_41 =10'b0;

   // m202_42 = W*in
   wire signed [9:0] m202_42;
   assign m202_42 =10'b0;

   // m202_43 = W*in
   wire signed [9:0] m202_43;
   assign m202_43 =10'b0;

   // m202_44 = W*in
   wire signed [9:0] m202_44;
   assign m202_44 =10'b0;

   // m202_45 = W*in
   wire signed [9:0] m202_45;
   assign m202_45 =10'b0;

   // m202_46 = W*in
   wire signed [9:0] m202_46;
   assign m202_46 =10'b0;

   // m202_47 = W*in
   wire signed [9:0] m202_47;
   assign m202_47 =10'b0;

   // m202_48 = W*in
   wire signed [9:0] m202_48;
   assign m202_48 =10'b0;

   // m202_49 = W*in
   wire signed [9:0] m202_49;
   assign m202_49 =10'b0;

   // m202_50 = W*in
   wire signed [9:0] m202_50;
   assign m202_50 =10'b0;

   // m202_51 = W*in
   wire signed [9:0] m202_51;
   assign m202_51 =10'b0;

   // m202_52 = W*in
   wire signed [9:0] m202_52;
   assign m202_52 =10'b0;

   // m202_53 = W*in
   wire signed [9:0] m202_53;
   assign m202_53 =10'b0;

   // m202_54 = W*in
   wire signed [9:0] m202_54;
   assign m202_54 =10'b0;

   // m202_55 = W*in
   wire signed [9:0] m202_55;
   assign m202_55 =10'b0;

   // m202_56 = W*in
   wire signed [9:0] m202_56;
   assign m202_56 =10'b0;

   // m202_57 = W*in
   wire signed [9:0] m202_57;
   assign m202_57 =10'b0;

   // m202_58 = W*in
   wire signed [9:0] m202_58;
   assign m202_58 =10'b0;

   // m202_59 = W*in
   wire signed [9:0] m202_59;
   assign m202_59 =10'b0;

   // m202_60 = W*in
   wire signed [9:0] m202_60;
   assign m202_60 =10'b0;

   // m202_61 = W*in
   wire signed [9:0] m202_61;
   assign m202_61 =10'b0;

   // m202_62 = W*in
   wire signed [9:0] m202_62;
   assign m202_62 =10'b0;

   // m202_63 = W*in
   wire signed [9:0] m202_63;
   assign m202_63 =10'b0;

   // m202_64 = W*in
   wire signed [9:0] m202_64;
   assign m202_64 ={ {4{in202[5]}} , in202[5:0] };

   // m202_65 = W*in
   wire signed [9:0] m202_65;
   assign m202_65 =10'b0;

   // m202_66 = W*in
   wire signed [9:0] m202_66;
   assign m202_66 =10'b0;

   // m202_67 = W*in
   wire signed [9:0] m202_67;
   assign m202_67 ={ {5{neg202[5]}} , neg202[5:1] };

   // m202_68 = W*in
   wire signed [9:0] m202_68;
   assign m202_68 =10'b0;

   // m202_69 = W*in
   wire signed [9:0] m202_69;
   assign m202_69 ={ {5{neg202[5]}} , neg202[5:1] };

   // m202_70 = W*in
   wire signed [9:0] m202_70;
   assign m202_70 =10'b0;

   // m202_71 = W*in
   wire signed [9:0] m202_71;
   assign m202_71 =10'b0;

   // m202_72 = W*in
   wire signed [9:0] m202_72;
   assign m202_72 =10'b0;

   // m202_73 = W*in
   wire signed [9:0] m202_73;
   assign m202_73 =10'b0;

   // m202_74 = W*in
   wire signed [9:0] m202_74;
   assign m202_74 =10'b0;

   // m202_75 = W*in
   wire signed [9:0] m202_75;
   assign m202_75 =10'b0;

   // m202_76 = W*in
   wire signed [9:0] m202_76;
   assign m202_76 =10'b0;

   // m202_77 = W*in
   wire signed [9:0] m202_77;
   assign m202_77 =10'b0;

   // m202_78 = W*in
   wire signed [9:0] m202_78;
   assign m202_78 =10'b0;

   // m202_79 = W*in
   wire signed [9:0] m202_79;
   assign m202_79 =10'b0;

   // m202_80 = W*in
   wire signed [9:0] m202_80;
   assign m202_80 =10'b0;

   // m202_81 = W*in
   wire signed [9:0] m202_81;
   assign m202_81 =10'b0;

   // m202_82 = W*in
   wire signed [9:0] m202_82;
   assign m202_82 =10'b0;

   // m202_83 = W*in
   wire signed [9:0] m202_83;
   assign m202_83 =10'b0;

   // m202_84 = W*in
   wire signed [9:0] m202_84;
   assign m202_84 =10'b0;

   // m202_85 = W*in
   wire signed [9:0] m202_85;
   assign m202_85 ={ {5{neg202[5]}} , neg202[5:1] };

   // m202_86 = W*in
   wire signed [9:0] m202_86;
   assign m202_86 =10'b0;

   // m202_87 = W*in
   wire signed [9:0] m202_87;
   assign m202_87 =10'b0;

   // m202_88 = W*in
   wire signed [9:0] m202_88;
   assign m202_88 =10'b0;

   // m202_89 = W*in
   wire signed [9:0] m202_89;
   assign m202_89 =10'b0;

   // m202_90 = W*in
   wire signed [9:0] m202_90;
   assign m202_90 =10'b0;

   // m202_91 = W*in
   wire signed [9:0] m202_91;
   assign m202_91 =10'b0;

   // m202_92 = W*in
   wire signed [9:0] m202_92;
   assign m202_92 =10'b0;

   // m202_93 = W*in
   wire signed [9:0] m202_93;
   assign m202_93 =10'b0;

   // m202_94 = W*in
   wire signed [9:0] m202_94;
   assign m202_94 =10'b0;

   // m202_95 = W*in
   wire signed [9:0] m202_95;
   assign m202_95 =10'b0;

   // m202_96 = W*in
   wire signed [9:0] m202_96;
   assign m202_96 =10'b0;

   // m202_97 = W*in
   wire signed [9:0] m202_97;
   assign m202_97 =10'b0;

   // m202_98 = W*in
   wire signed [9:0] m202_98;
   assign m202_98 =10'b0;

   // m202_99 = W*in
   wire signed [9:0] m202_99;
   assign m202_99 =10'b0;

   // m202_100 = W*in
   wire signed [9:0] m202_100;
   assign m202_100 =10'b0;

   // m202_101 = W*in
   wire signed [9:0] m202_101;
   assign m202_101 =10'b0;

   // m202_102 = W*in
   wire signed [9:0] m202_102;
   assign m202_102 =10'b0;

   // m202_103 = W*in
   wire signed [9:0] m202_103;
   assign m202_103 =10'b0;

   // m202_104 = W*in
   wire signed [9:0] m202_104;
   assign m202_104 =10'b0;

   // m202_105 = W*in
   wire signed [9:0] m202_105;
   assign m202_105 =10'b0;

   // m202_106 = W*in
   wire signed [9:0] m202_106;
   assign m202_106 =10'b0;

   // m202_107 = W*in
   wire signed [9:0] m202_107;
   assign m202_107 =10'b0;

   // m202_108 = W*in
   wire signed [9:0] m202_108;
   assign m202_108 =10'b0;

   // m202_109 = W*in
   wire signed [9:0] m202_109;
   assign m202_109 =10'b0;

   // m202_110 = W*in
   wire signed [9:0] m202_110;
   assign m202_110 =10'b0;

   // m202_111 = W*in
   wire signed [9:0] m202_111;
   assign m202_111 =10'b0;

   // m202_112 = W*in
   wire signed [9:0] m202_112;
   assign m202_112 =10'b0;

   // m202_113 = W*in
   wire signed [9:0] m202_113;
   assign m202_113 =10'b0;

   // m202_114 = W*in
   wire signed [9:0] m202_114;
   assign m202_114 ={ {5{in202[5]}} , in202[5:1] };

   // m202_115 = W*in
   wire signed [9:0] m202_115;
   assign m202_115 =10'b0;

   // m202_116 = W*in
   wire signed [9:0] m202_116;
   assign m202_116 =10'b0;

   // m202_117 = W*in
   wire signed [9:0] m202_117;
   assign m202_117 =10'b0;

   // m203_1 = W*in
   wire signed [9:0] m203_1;
   assign m203_1 =10'b0;

   // m203_2 = W*in
   wire signed [9:0] m203_2;
   assign m203_2 =10'b0;

   // m203_3 = W*in
   wire signed [9:0] m203_3;
   assign m203_3 =10'b0;

   // m203_4 = W*in
   wire signed [9:0] m203_4;
   assign m203_4 =10'b0;

   // m203_5 = W*in
   wire signed [9:0] m203_5;
   assign m203_5 =10'b0;

   // m203_6 = W*in
   wire signed [9:0] m203_6;
   assign m203_6 =10'b0;

   // m203_7 = W*in
   wire signed [9:0] m203_7;
   assign m203_7 =10'b0;

   // m203_8 = W*in
   wire signed [9:0] m203_8;
   assign m203_8 =10'b0;

   // m203_9 = W*in
   wire signed [9:0] m203_9;
   assign m203_9 =10'b0;

   // m203_10 = W*in
   wire signed [9:0] m203_10;
   assign m203_10 =10'b0;

   // m203_11 = W*in
   wire signed [9:0] m203_11;
   assign m203_11 =10'b0;

   // m203_12 = W*in
   wire signed [9:0] m203_12;
   assign m203_12 ={ {4{in203[5]}} , in203[5:0] };

   // m203_13 = W*in
   wire signed [9:0] m203_13;
   assign m203_13 =10'b0;

   // m203_14 = W*in
   wire signed [9:0] m203_14;
   assign m203_14 =10'b0;

   // m203_15 = W*in
   wire signed [9:0] m203_15;
   assign m203_15 =10'b0;

   // m203_16 = W*in
   wire signed [9:0] m203_16;
   assign m203_16 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_17 = W*in
   wire signed [9:0] m203_17;
   assign m203_17 ={ {5{in203[5]}} , in203[5:1] };

   // m203_18 = W*in
   wire signed [9:0] m203_18;
   assign m203_18 ={ {4{in203[5]}} , in203[5:0] };

   // m203_19 = W*in
   wire signed [9:0] m203_19;
   assign m203_19 =10'b0;

   // m203_20 = W*in
   wire signed [9:0] m203_20;
   assign m203_20 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_21 = W*in
   wire signed [9:0] m203_21;
   assign m203_21 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_22 = W*in
   wire signed [9:0] m203_22;
   assign m203_22 =10'b0;

   // m203_23 = W*in
   wire signed [9:0] m203_23;
   assign m203_23 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_24 = W*in
   wire signed [9:0] m203_24;
   assign m203_24 =10'b0;

   // m203_25 = W*in
   wire signed [9:0] m203_25;
   assign m203_25 ={ {5{in203[5]}} , in203[5:1] };

   // m203_26 = W*in
   wire signed [9:0] m203_26;
   assign m203_26 ={ {5{in203[5]}} , in203[5:1] };

   // m203_27 = W*in
   wire signed [9:0] m203_27;
   assign m203_27 ={ {4{in203[5]}} , in203[5:0] };

   // m203_28 = W*in
   wire signed [9:0] m203_28;
   assign m203_28 ={ {5{in203[5]}} , in203[5:1] };

   // m203_29 = W*in
   wire signed [9:0] m203_29;
   assign m203_29 =10'b0;

   // m203_30 = W*in
   wire signed [9:0] m203_30;
   assign m203_30 =10'b0;

   // m203_31 = W*in
   wire signed [9:0] m203_31;
   assign m203_31 =10'b0;

   // m203_32 = W*in
   wire signed [9:0] m203_32;
   assign m203_32 =10'b0;

   // m203_33 = W*in
   wire signed [9:0] m203_33;
   assign m203_33 =10'b0;

   // m203_34 = W*in
   wire signed [9:0] m203_34;
   assign m203_34 =10'b0;

   // m203_35 = W*in
   wire signed [9:0] m203_35;
   assign m203_35 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_36 = W*in
   wire signed [9:0] m203_36;
   assign m203_36 =10'b0;

   // m203_37 = W*in
   wire signed [9:0] m203_37;
   assign m203_37 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_38 = W*in
   wire signed [9:0] m203_38;
   assign m203_38 =10'b0;

   // m203_39 = W*in
   wire signed [9:0] m203_39;
   assign m203_39 =10'b0;

   // m203_40 = W*in
   wire signed [9:0] m203_40;
   assign m203_40 =10'b0;

   // m203_41 = W*in
   wire signed [9:0] m203_41;
   assign m203_41 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_42 = W*in
   wire signed [9:0] m203_42;
   assign m203_42 ={ {4{in203[5]}} , in203[5:0] };

   // m203_43 = W*in
   wire signed [9:0] m203_43;
   assign m203_43 ={ {4{in203[5]}} , in203[5:0] };

   // m203_44 = W*in
   wire signed [9:0] m203_44;
   assign m203_44 =10'b0;

   // m203_45 = W*in
   wire signed [9:0] m203_45;
   assign m203_45 =10'b0;

   // m203_46 = W*in
   wire signed [9:0] m203_46;
   assign m203_46 =10'b0;

   // m203_47 = W*in
   wire signed [9:0] m203_47;
   assign m203_47 =10'b0;

   // m203_48 = W*in
   wire signed [9:0] m203_48;
   assign m203_48 =10'b0;

   // m203_49 = W*in
   wire signed [9:0] m203_49;
   assign m203_49 =10'b0;

   // m203_50 = W*in
   wire signed [9:0] m203_50;
   assign m203_50 =10'b0;

   // m203_51 = W*in
   wire signed [9:0] m203_51;
   assign m203_51 =10'b0;

   // m203_52 = W*in
   wire signed [9:0] m203_52;
   assign m203_52 =10'b0;

   // m203_53 = W*in
   wire signed [9:0] m203_53;
   assign m203_53 =10'b0;

   // m203_54 = W*in
   wire signed [9:0] m203_54;
   assign m203_54 =10'b0;

   // m203_55 = W*in
   wire signed [9:0] m203_55;
   assign m203_55 =10'b0;

   // m203_56 = W*in
   wire signed [9:0] m203_56;
   assign m203_56 =10'b0;

   // m203_57 = W*in
   wire signed [9:0] m203_57;
   assign m203_57 =10'b0;

   // m203_58 = W*in
   wire signed [9:0] m203_58;
   assign m203_58 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_59 = W*in
   wire signed [9:0] m203_59;
   assign m203_59 =10'b0;

   // m203_60 = W*in
   wire signed [9:0] m203_60;
   assign m203_60 =10'b0;

   // m203_61 = W*in
   wire signed [9:0] m203_61;
   assign m203_61 =10'b0;

   // m203_62 = W*in
   wire signed [9:0] m203_62;
   assign m203_62 =10'b0;

   // m203_63 = W*in
   wire signed [9:0] m203_63;
   assign m203_63 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_64 = W*in
   wire signed [9:0] m203_64;
   assign m203_64 ={ {5{in203[5]}} , in203[5:1] };

   // m203_65 = W*in
   wire signed [9:0] m203_65;
   assign m203_65 =10'b0;

   // m203_66 = W*in
   wire signed [9:0] m203_66;
   assign m203_66 ={ {4{in203[5]}} , in203[5:0] };

   // m203_67 = W*in
   wire signed [9:0] m203_67;
   assign m203_67 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_68 = W*in
   wire signed [9:0] m203_68;
   assign m203_68 =10'b0;

   // m203_69 = W*in
   wire signed [9:0] m203_69;
   assign m203_69 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_70 = W*in
   wire signed [9:0] m203_70;
   assign m203_70 =10'b0;

   // m203_71 = W*in
   wire signed [9:0] m203_71;
   assign m203_71 ={ {5{in203[5]}} , in203[5:1] };

   // m203_72 = W*in
   wire signed [9:0] m203_72;
   assign m203_72 =10'b0;

   // m203_73 = W*in
   wire signed [9:0] m203_73;
   assign m203_73 =10'b0;

   // m203_74 = W*in
   wire signed [9:0] m203_74;
   assign m203_74 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_75 = W*in
   wire signed [9:0] m203_75;
   assign m203_75 =10'b0;

   // m203_76 = W*in
   wire signed [9:0] m203_76;
   assign m203_76 =10'b0;

   // m203_77 = W*in
   wire signed [9:0] m203_77;
   assign m203_77 ={ {4{in203[5]}} , in203[5:0] };

   // m203_78 = W*in
   wire signed [9:0] m203_78;
   assign m203_78 =10'b0;

   // m203_79 = W*in
   wire signed [9:0] m203_79;
   assign m203_79 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_80 = W*in
   wire signed [9:0] m203_80;
   assign m203_80 =10'b0;

   // m203_81 = W*in
   wire signed [9:0] m203_81;
   assign m203_81 =10'b0;

   // m203_82 = W*in
   wire signed [9:0] m203_82;
   assign m203_82 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_83 = W*in
   wire signed [9:0] m203_83;
   assign m203_83 =10'b0;

   // m203_84 = W*in
   wire signed [9:0] m203_84;
   assign m203_84 =10'b0;

   // m203_85 = W*in
   wire signed [9:0] m203_85;
   assign m203_85 ={ {3{neg203[5]}} , neg203 , {1{1'b0}} };

   // m203_86 = W*in
   wire signed [9:0] m203_86;
   assign m203_86 =10'b0;

   // m203_87 = W*in
   wire signed [9:0] m203_87;
   assign m203_87 =10'b0;

   // m203_88 = W*in
   wire signed [9:0] m203_88;
   assign m203_88 =10'b0;

   // m203_89 = W*in
   wire signed [9:0] m203_89;
   assign m203_89 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_90 = W*in
   wire signed [9:0] m203_90;
   assign m203_90 =10'b0;

   // m203_91 = W*in
   wire signed [9:0] m203_91;
   assign m203_91 ={ {4{in203[5]}} , in203[5:0] };

   // m203_92 = W*in
   wire signed [9:0] m203_92;
   assign m203_92 =10'b0;

   // m203_93 = W*in
   wire signed [9:0] m203_93;
   assign m203_93 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_94 = W*in
   wire signed [9:0] m203_94;
   assign m203_94 =10'b0;

   // m203_95 = W*in
   wire signed [9:0] m203_95;
   assign m203_95 =10'b0;

   // m203_96 = W*in
   wire signed [9:0] m203_96;
   assign m203_96 =10'b0;

   // m203_97 = W*in
   wire signed [9:0] m203_97;
   assign m203_97 ={ {4{in203[5]}} , in203[5:0] };

   // m203_98 = W*in
   wire signed [9:0] m203_98;
   assign m203_98 =10'b0;

   // m203_99 = W*in
   wire signed [9:0] m203_99;
   assign m203_99 =10'b0;

   // m203_100 = W*in
   wire signed [9:0] m203_100;
   assign m203_100 ={ {4{in203[5]}} , in203[5:0] };

   // m203_101 = W*in
   wire signed [9:0] m203_101;
   assign m203_101 =10'b0;

   // m203_102 = W*in
   wire signed [9:0] m203_102;
   assign m203_102 =10'b0;

   // m203_103 = W*in
   wire signed [9:0] m203_103;
   assign m203_103 =10'b0;

   // m203_104 = W*in
   wire signed [9:0] m203_104;
   assign m203_104 ={ {4{in203[5]}} , in203[5:0] };

   // m203_105 = W*in
   wire signed [9:0] m203_105;
   assign m203_105 =10'b0;

   // m203_106 = W*in
   wire signed [9:0] m203_106;
   assign m203_106 =10'b0;

   // m203_107 = W*in
   wire signed [9:0] m203_107;
   assign m203_107 =10'b0;

   // m203_108 = W*in
   wire signed [9:0] m203_108;
   assign m203_108 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_109 = W*in
   wire signed [9:0] m203_109;
   assign m203_109 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_110 = W*in
   wire signed [9:0] m203_110;
   assign m203_110 =10'b0;

   // m203_111 = W*in
   wire signed [9:0] m203_111;
   assign m203_111 =10'b0;

   // m203_112 = W*in
   wire signed [9:0] m203_112;
   assign m203_112 ={ {4{in203[5]}} , in203[5:0] };

   // m203_113 = W*in
   wire signed [9:0] m203_113;
   assign m203_113 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_114 = W*in
   wire signed [9:0] m203_114;
   assign m203_114 =10'b0;

   // m203_115 = W*in
   wire signed [9:0] m203_115;
   assign m203_115 ={ {5{neg203[5]}} , neg203[5:1] };

   // m203_116 = W*in
   wire signed [9:0] m203_116;
   assign m203_116 ={ {4{neg203[5]}} , neg203[5:0] };

   // m203_117 = W*in
   wire signed [9:0] m203_117;
   assign m203_117 =10'b0;

   // m204_1 = W*in
   wire signed [9:0] m204_1;
   assign m204_1 =10'b0;

   // m204_2 = W*in
   wire signed [9:0] m204_2;
   assign m204_2 =10'b0;

   // m204_3 = W*in
   wire signed [9:0] m204_3;
   assign m204_3 ={ {4{in204[5]}} , in204[5:0] };

   // m204_4 = W*in
   wire signed [9:0] m204_4;
   assign m204_4 =10'b0;

   // m204_5 = W*in
   wire signed [9:0] m204_5;
   assign m204_5 =10'b0;

   // m204_6 = W*in
   wire signed [9:0] m204_6;
   assign m204_6 =10'b0;

   // m204_7 = W*in
   wire signed [9:0] m204_7;
   assign m204_7 =10'b0;

   // m204_8 = W*in
   wire signed [9:0] m204_8;
   assign m204_8 =10'b0;

   // m204_9 = W*in
   wire signed [9:0] m204_9;
   assign m204_9 =10'b0;

   // m204_10 = W*in
   wire signed [9:0] m204_10;
   assign m204_10 ={ {4{neg204[5]}} , neg204[5:0] };

   // m204_11 = W*in
   wire signed [9:0] m204_11;
   assign m204_11 =10'b0;

   // m204_12 = W*in
   wire signed [9:0] m204_12;
   assign m204_12 ={ {4{in204[5]}} , in204[5:0] };

   // m204_13 = W*in
   wire signed [9:0] m204_13;
   assign m204_13 =10'b0;

   // m204_14 = W*in
   wire signed [9:0] m204_14;
   assign m204_14 =10'b0;

   // m204_15 = W*in
   wire signed [9:0] m204_15;
   assign m204_15 =10'b0;

   // m204_16 = W*in
   wire signed [9:0] m204_16;
   assign m204_16 =10'b0;

   // m204_17 = W*in
   wire signed [9:0] m204_17;
   assign m204_17 ={ {5{in204[5]}} , in204[5:1] };

   // m204_18 = W*in
   wire signed [9:0] m204_18;
   assign m204_18 ={ {5{in204[5]}} , in204[5:1] };

   // m204_19 = W*in
   wire signed [9:0] m204_19;
   assign m204_19 =10'b0;

   // m204_20 = W*in
   wire signed [9:0] m204_20;
   assign m204_20 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_21 = W*in
   wire signed [9:0] m204_21;
   assign m204_21 =10'b0;

   // m204_22 = W*in
   wire signed [9:0] m204_22;
   assign m204_22 =10'b0;

   // m204_23 = W*in
   wire signed [9:0] m204_23;
   assign m204_23 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_24 = W*in
   wire signed [9:0] m204_24;
   assign m204_24 =10'b0;

   // m204_25 = W*in
   wire signed [9:0] m204_25;
   assign m204_25 =10'b0;

   // m204_26 = W*in
   wire signed [9:0] m204_26;
   assign m204_26 =10'b0;

   // m204_27 = W*in
   wire signed [9:0] m204_27;
   assign m204_27 ={ {4{in204[5]}} , in204[5:0] };

   // m204_28 = W*in
   wire signed [9:0] m204_28;
   assign m204_28 ={ {4{in204[5]}} , in204[5:0] };

   // m204_29 = W*in
   wire signed [9:0] m204_29;
   assign m204_29 =10'b0;

   // m204_30 = W*in
   wire signed [9:0] m204_30;
   assign m204_30 =10'b0;

   // m204_31 = W*in
   wire signed [9:0] m204_31;
   assign m204_31 =10'b0;

   // m204_32 = W*in
   wire signed [9:0] m204_32;
   assign m204_32 ={ {4{neg204[5]}} , neg204[5:0] };

   // m204_33 = W*in
   wire signed [9:0] m204_33;
   assign m204_33 =10'b0;

   // m204_34 = W*in
   wire signed [9:0] m204_34;
   assign m204_34 =10'b0;

   // m204_35 = W*in
   wire signed [9:0] m204_35;
   assign m204_35 ={ {5{in204[5]}} , in204[5:1] };

   // m204_36 = W*in
   wire signed [9:0] m204_36;
   assign m204_36 =10'b0;

   // m204_37 = W*in
   wire signed [9:0] m204_37;
   assign m204_37 ={ {4{neg204[5]}} , neg204[5:0] };

   // m204_38 = W*in
   wire signed [9:0] m204_38;
   assign m204_38 =10'b0;

   // m204_39 = W*in
   wire signed [9:0] m204_39;
   assign m204_39 =10'b0;

   // m204_40 = W*in
   wire signed [9:0] m204_40;
   assign m204_40 =10'b0;

   // m204_41 = W*in
   wire signed [9:0] m204_41;
   assign m204_41 =10'b0;

   // m204_42 = W*in
   wire signed [9:0] m204_42;
   assign m204_42 =10'b0;

   // m204_43 = W*in
   wire signed [9:0] m204_43;
   assign m204_43 =10'b0;

   // m204_44 = W*in
   wire signed [9:0] m204_44;
   assign m204_44 =10'b0;

   // m204_45 = W*in
   wire signed [9:0] m204_45;
   assign m204_45 ={ {4{neg204[5]}} , neg204[5:0] };

   // m204_46 = W*in
   wire signed [9:0] m204_46;
   assign m204_46 =10'b0;

   // m204_47 = W*in
   wire signed [9:0] m204_47;
   assign m204_47 =10'b0;

   // m204_48 = W*in
   wire signed [9:0] m204_48;
   assign m204_48 =10'b0;

   // m204_49 = W*in
   wire signed [9:0] m204_49;
   assign m204_49 =10'b0;

   // m204_50 = W*in
   wire signed [9:0] m204_50;
   assign m204_50 =10'b0;

   // m204_51 = W*in
   wire signed [9:0] m204_51;
   assign m204_51 ={ {4{neg204[5]}} , neg204[5:0] };

   // m204_52 = W*in
   wire signed [9:0] m204_52;
   assign m204_52 =10'b0;

   // m204_53 = W*in
   wire signed [9:0] m204_53;
   assign m204_53 =10'b0;

   // m204_54 = W*in
   wire signed [9:0] m204_54;
   assign m204_54 =10'b0;

   // m204_55 = W*in
   wire signed [9:0] m204_55;
   assign m204_55 =10'b0;

   // m204_56 = W*in
   wire signed [9:0] m204_56;
   assign m204_56 =10'b0;

   // m204_57 = W*in
   wire signed [9:0] m204_57;
   assign m204_57 =10'b0;

   // m204_58 = W*in
   wire signed [9:0] m204_58;
   assign m204_58 =10'b0;

   // m204_59 = W*in
   wire signed [9:0] m204_59;
   assign m204_59 =10'b0;

   // m204_60 = W*in
   wire signed [9:0] m204_60;
   assign m204_60 =10'b0;

   // m204_61 = W*in
   wire signed [9:0] m204_61;
   assign m204_61 ={ {4{in204[5]}} , in204[5:0] };

   // m204_62 = W*in
   wire signed [9:0] m204_62;
   assign m204_62 =10'b0;

   // m204_63 = W*in
   wire signed [9:0] m204_63;
   assign m204_63 =10'b0;

   // m204_64 = W*in
   wire signed [9:0] m204_64;
   assign m204_64 =10'b0;

   // m204_65 = W*in
   wire signed [9:0] m204_65;
   assign m204_65 =10'b0;

   // m204_66 = W*in
   wire signed [9:0] m204_66;
   assign m204_66 ={ {4{in204[5]}} , in204[5:0] };

   // m204_67 = W*in
   wire signed [9:0] m204_67;
   assign m204_67 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_68 = W*in
   wire signed [9:0] m204_68;
   assign m204_68 =10'b0;

   // m204_69 = W*in
   wire signed [9:0] m204_69;
   assign m204_69 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_70 = W*in
   wire signed [9:0] m204_70;
   assign m204_70 =10'b0;

   // m204_71 = W*in
   wire signed [9:0] m204_71;
   assign m204_71 ={ {5{in204[5]}} , in204[5:1] };

   // m204_72 = W*in
   wire signed [9:0] m204_72;
   assign m204_72 =10'b0;

   // m204_73 = W*in
   wire signed [9:0] m204_73;
   assign m204_73 =10'b0;

   // m204_74 = W*in
   wire signed [9:0] m204_74;
   assign m204_74 =10'b0;

   // m204_75 = W*in
   wire signed [9:0] m204_75;
   assign m204_75 =10'b0;

   // m204_76 = W*in
   wire signed [9:0] m204_76;
   assign m204_76 =10'b0;

   // m204_77 = W*in
   wire signed [9:0] m204_77;
   assign m204_77 =10'b0;

   // m204_78 = W*in
   wire signed [9:0] m204_78;
   assign m204_78 =10'b0;

   // m204_79 = W*in
   wire signed [9:0] m204_79;
   assign m204_79 =10'b0;

   // m204_80 = W*in
   wire signed [9:0] m204_80;
   assign m204_80 =10'b0;

   // m204_81 = W*in
   wire signed [9:0] m204_81;
   assign m204_81 =10'b0;

   // m204_82 = W*in
   wire signed [9:0] m204_82;
   assign m204_82 =10'b0;

   // m204_83 = W*in
   wire signed [9:0] m204_83;
   assign m204_83 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_84 = W*in
   wire signed [9:0] m204_84;
   assign m204_84 =10'b0;

   // m204_85 = W*in
   wire signed [9:0] m204_85;
   assign m204_85 ={ {4{neg204[5]}} , neg204[5:0] };

   // m204_86 = W*in
   wire signed [9:0] m204_86;
   assign m204_86 =10'b0;

   // m204_87 = W*in
   wire signed [9:0] m204_87;
   assign m204_87 =10'b0;

   // m204_88 = W*in
   wire signed [9:0] m204_88;
   assign m204_88 =10'b0;

   // m204_89 = W*in
   wire signed [9:0] m204_89;
   assign m204_89 =10'b0;

   // m204_90 = W*in
   wire signed [9:0] m204_90;
   assign m204_90 =10'b0;

   // m204_91 = W*in
   wire signed [9:0] m204_91;
   assign m204_91 ={ {4{in204[5]}} , in204[5:0] };

   // m204_92 = W*in
   wire signed [9:0] m204_92;
   assign m204_92 =10'b0;

   // m204_93 = W*in
   wire signed [9:0] m204_93;
   assign m204_93 =10'b0;

   // m204_94 = W*in
   wire signed [9:0] m204_94;
   assign m204_94 =10'b0;

   // m204_95 = W*in
   wire signed [9:0] m204_95;
   assign m204_95 =10'b0;

   // m204_96 = W*in
   wire signed [9:0] m204_96;
   assign m204_96 =10'b0;

   // m204_97 = W*in
   wire signed [9:0] m204_97;
   assign m204_97 ={ {4{in204[5]}} , in204[5:0] };

   // m204_98 = W*in
   wire signed [9:0] m204_98;
   assign m204_98 =10'b0;

   // m204_99 = W*in
   wire signed [9:0] m204_99;
   assign m204_99 =10'b0;

   // m204_100 = W*in
   wire signed [9:0] m204_100;
   assign m204_100 ={ {4{in204[5]}} , in204[5:0] };

   // m204_101 = W*in
   wire signed [9:0] m204_101;
   assign m204_101 =10'b0;

   // m204_102 = W*in
   wire signed [9:0] m204_102;
   assign m204_102 =10'b0;

   // m204_103 = W*in
   wire signed [9:0] m204_103;
   assign m204_103 =10'b0;

   // m204_104 = W*in
   wire signed [9:0] m204_104;
   assign m204_104 ={ {4{in204[5]}} , in204[5:0] };

   // m204_105 = W*in
   wire signed [9:0] m204_105;
   assign m204_105 =10'b0;

   // m204_106 = W*in
   wire signed [9:0] m204_106;
   assign m204_106 =10'b0;

   // m204_107 = W*in
   wire signed [9:0] m204_107;
   assign m204_107 =10'b0;

   // m204_108 = W*in
   wire signed [9:0] m204_108;
   assign m204_108 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_109 = W*in
   wire signed [9:0] m204_109;
   assign m204_109 =10'b0;

   // m204_110 = W*in
   wire signed [9:0] m204_110;
   assign m204_110 =10'b0;

   // m204_111 = W*in
   wire signed [9:0] m204_111;
   assign m204_111 =10'b0;

   // m204_112 = W*in
   wire signed [9:0] m204_112;
   assign m204_112 ={ {4{in204[5]}} , in204[5:0] };

   // m204_113 = W*in
   wire signed [9:0] m204_113;
   assign m204_113 =10'b0;

   // m204_114 = W*in
   wire signed [9:0] m204_114;
   assign m204_114 ={ {5{neg204[5]}} , neg204[5:1] };

   // m204_115 = W*in
   wire signed [9:0] m204_115;
   assign m204_115 =10'b0;

   // m204_116 = W*in
   wire signed [9:0] m204_116;
   assign m204_116 =10'b0;

   // m204_117 = W*in
   wire signed [9:0] m204_117;
   assign m204_117 =10'b0;

   // m205_1 = W*in
   wire signed [9:0] m205_1;
   assign m205_1 =10'b0;

   // m205_2 = W*in
   wire signed [9:0] m205_2;
   assign m205_2 =10'b0;

   // m205_3 = W*in
   wire signed [9:0] m205_3;
   assign m205_3 =10'b0;

   // m205_4 = W*in
   wire signed [9:0] m205_4;
   assign m205_4 =10'b0;

   // m205_5 = W*in
   wire signed [9:0] m205_5;
   assign m205_5 =10'b0;

   // m205_6 = W*in
   wire signed [9:0] m205_6;
   assign m205_6 =10'b0;

   // m205_7 = W*in
   wire signed [9:0] m205_7;
   assign m205_7 =10'b0;

   // m205_8 = W*in
   wire signed [9:0] m205_8;
   assign m205_8 =10'b0;

   // m205_9 = W*in
   wire signed [9:0] m205_9;
   assign m205_9 =10'b0;

   // m205_10 = W*in
   wire signed [9:0] m205_10;
   assign m205_10 =10'b0;

   // m205_11 = W*in
   wire signed [9:0] m205_11;
   assign m205_11 =10'b0;

   // m205_12 = W*in
   wire signed [9:0] m205_12;
   assign m205_12 =10'b0;

   // m205_13 = W*in
   wire signed [9:0] m205_13;
   assign m205_13 =10'b0;

   // m205_14 = W*in
   wire signed [9:0] m205_14;
   assign m205_14 =10'b0;

   // m205_15 = W*in
   wire signed [9:0] m205_15;
   assign m205_15 =10'b0;

   // m205_16 = W*in
   wire signed [9:0] m205_16;
   assign m205_16 =10'b0;

   // m205_17 = W*in
   wire signed [9:0] m205_17;
   assign m205_17 =10'b0;

   // m205_18 = W*in
   wire signed [9:0] m205_18;
   assign m205_18 =10'b0;

   // m205_19 = W*in
   wire signed [9:0] m205_19;
   assign m205_19 =10'b0;

   // m205_20 = W*in
   wire signed [9:0] m205_20;
   assign m205_20 =10'b0;

   // m205_21 = W*in
   wire signed [9:0] m205_21;
   assign m205_21 =10'b0;

   // m205_22 = W*in
   wire signed [9:0] m205_22;
   assign m205_22 =10'b0;

   // m205_23 = W*in
   wire signed [9:0] m205_23;
   assign m205_23 ={ {5{neg205[5]}} , neg205[5:1] };

   // m205_24 = W*in
   wire signed [9:0] m205_24;
   assign m205_24 =10'b0;

   // m205_25 = W*in
   wire signed [9:0] m205_25;
   assign m205_25 =10'b0;

   // m205_26 = W*in
   wire signed [9:0] m205_26;
   assign m205_26 =10'b0;

   // m205_27 = W*in
   wire signed [9:0] m205_27;
   assign m205_27 =10'b0;

   // m205_28 = W*in
   wire signed [9:0] m205_28;
   assign m205_28 =10'b0;

   // m205_29 = W*in
   wire signed [9:0] m205_29;
   assign m205_29 =10'b0;

   // m205_30 = W*in
   wire signed [9:0] m205_30;
   assign m205_30 =10'b0;

   // m205_31 = W*in
   wire signed [9:0] m205_31;
   assign m205_31 =10'b0;

   // m205_32 = W*in
   wire signed [9:0] m205_32;
   assign m205_32 =10'b0;

   // m205_33 = W*in
   wire signed [9:0] m205_33;
   assign m205_33 =10'b0;

   // m205_34 = W*in
   wire signed [9:0] m205_34;
   assign m205_34 ={ {5{neg205[5]}} , neg205[5:1] };

   // m205_35 = W*in
   wire signed [9:0] m205_35;
   assign m205_35 =10'b0;

   // m205_36 = W*in
   wire signed [9:0] m205_36;
   assign m205_36 =10'b0;

   // m205_37 = W*in
   wire signed [9:0] m205_37;
   assign m205_37 =10'b0;

   // m205_38 = W*in
   wire signed [9:0] m205_38;
   assign m205_38 =10'b0;

   // m205_39 = W*in
   wire signed [9:0] m205_39;
   assign m205_39 =10'b0;

   // m205_40 = W*in
   wire signed [9:0] m205_40;
   assign m205_40 =10'b0;

   // m205_41 = W*in
   wire signed [9:0] m205_41;
   assign m205_41 =10'b0;

   // m205_42 = W*in
   wire signed [9:0] m205_42;
   assign m205_42 =10'b0;

   // m205_43 = W*in
   wire signed [9:0] m205_43;
   assign m205_43 =10'b0;

   // m205_44 = W*in
   wire signed [9:0] m205_44;
   assign m205_44 =10'b0;

   // m205_45 = W*in
   wire signed [9:0] m205_45;
   assign m205_45 =10'b0;

   // m205_46 = W*in
   wire signed [9:0] m205_46;
   assign m205_46 =10'b0;

   // m205_47 = W*in
   wire signed [9:0] m205_47;
   assign m205_47 =10'b0;

   // m205_48 = W*in
   wire signed [9:0] m205_48;
   assign m205_48 =10'b0;

   // m205_49 = W*in
   wire signed [9:0] m205_49;
   assign m205_49 =10'b0;

   // m205_50 = W*in
   wire signed [9:0] m205_50;
   assign m205_50 =10'b0;

   // m205_51 = W*in
   wire signed [9:0] m205_51;
   assign m205_51 =10'b0;

   // m205_52 = W*in
   wire signed [9:0] m205_52;
   assign m205_52 =10'b0;

   // m205_53 = W*in
   wire signed [9:0] m205_53;
   assign m205_53 =10'b0;

   // m205_54 = W*in
   wire signed [9:0] m205_54;
   assign m205_54 =10'b0;

   // m205_55 = W*in
   wire signed [9:0] m205_55;
   assign m205_55 =10'b0;

   // m205_56 = W*in
   wire signed [9:0] m205_56;
   assign m205_56 =10'b0;

   // m205_57 = W*in
   wire signed [9:0] m205_57;
   assign m205_57 =10'b0;

   // m205_58 = W*in
   wire signed [9:0] m205_58;
   assign m205_58 =10'b0;

   // m205_59 = W*in
   wire signed [9:0] m205_59;
   assign m205_59 =10'b0;

   // m205_60 = W*in
   wire signed [9:0] m205_60;
   assign m205_60 =10'b0;

   // m205_61 = W*in
   wire signed [9:0] m205_61;
   assign m205_61 =10'b0;

   // m205_62 = W*in
   wire signed [9:0] m205_62;
   assign m205_62 =10'b0;

   // m205_63 = W*in
   wire signed [9:0] m205_63;
   assign m205_63 =10'b0;

   // m205_64 = W*in
   wire signed [9:0] m205_64;
   assign m205_64 =10'b0;

   // m205_65 = W*in
   wire signed [9:0] m205_65;
   assign m205_65 =10'b0;

   // m205_66 = W*in
   wire signed [9:0] m205_66;
   assign m205_66 ={ {5{in205[5]}} , in205[5:1] };

   // m205_67 = W*in
   wire signed [9:0] m205_67;
   assign m205_67 =10'b0;

   // m205_68 = W*in
   wire signed [9:0] m205_68;
   assign m205_68 =10'b0;

   // m205_69 = W*in
   wire signed [9:0] m205_69;
   assign m205_69 ={ {5{neg205[5]}} , neg205[5:1] };

   // m205_70 = W*in
   wire signed [9:0] m205_70;
   assign m205_70 ={ {5{neg205[5]}} , neg205[5:1] };

   // m205_71 = W*in
   wire signed [9:0] m205_71;
   assign m205_71 =10'b0;

   // m205_72 = W*in
   wire signed [9:0] m205_72;
   assign m205_72 ={ {4{neg205[5]}} , neg205[5:0] };

   // m205_73 = W*in
   wire signed [9:0] m205_73;
   assign m205_73 =10'b0;

   // m205_74 = W*in
   wire signed [9:0] m205_74;
   assign m205_74 =10'b0;

   // m205_75 = W*in
   wire signed [9:0] m205_75;
   assign m205_75 =10'b0;

   // m205_76 = W*in
   wire signed [9:0] m205_76;
   assign m205_76 =10'b0;

   // m205_77 = W*in
   wire signed [9:0] m205_77;
   assign m205_77 =10'b0;

   // m205_78 = W*in
   wire signed [9:0] m205_78;
   assign m205_78 =10'b0;

   // m205_79 = W*in
   wire signed [9:0] m205_79;
   assign m205_79 =10'b0;

   // m205_80 = W*in
   wire signed [9:0] m205_80;
   assign m205_80 =10'b0;

   // m205_81 = W*in
   wire signed [9:0] m205_81;
   assign m205_81 =10'b0;

   // m205_82 = W*in
   wire signed [9:0] m205_82;
   assign m205_82 ={ {5{neg205[5]}} , neg205[5:1] };

   // m205_83 = W*in
   wire signed [9:0] m205_83;
   assign m205_83 =10'b0;

   // m205_84 = W*in
   wire signed [9:0] m205_84;
   assign m205_84 =10'b0;

   // m205_85 = W*in
   wire signed [9:0] m205_85;
   assign m205_85 ={ {5{neg205[5]}} , neg205[5:1] };

   // m205_86 = W*in
   wire signed [9:0] m205_86;
   assign m205_86 =10'b0;

   // m205_87 = W*in
   wire signed [9:0] m205_87;
   assign m205_87 ={ {4{neg205[5]}} , neg205[5:0] };

   // m205_88 = W*in
   wire signed [9:0] m205_88;
   assign m205_88 =10'b0;

   // m205_89 = W*in
   wire signed [9:0] m205_89;
   assign m205_89 ={ {4{neg205[5]}} , neg205[5:0] };

   // m205_90 = W*in
   wire signed [9:0] m205_90;
   assign m205_90 =10'b0;

   // m205_91 = W*in
   wire signed [9:0] m205_91;
   assign m205_91 =10'b0;

   // m205_92 = W*in
   wire signed [9:0] m205_92;
   assign m205_92 =10'b0;

   // m205_93 = W*in
   wire signed [9:0] m205_93;
   assign m205_93 =10'b0;

   // m205_94 = W*in
   wire signed [9:0] m205_94;
   assign m205_94 =10'b0;

   // m205_95 = W*in
   wire signed [9:0] m205_95;
   assign m205_95 =10'b0;

   // m205_96 = W*in
   wire signed [9:0] m205_96;
   assign m205_96 =10'b0;

   // m205_97 = W*in
   wire signed [9:0] m205_97;
   assign m205_97 =10'b0;

   // m205_98 = W*in
   wire signed [9:0] m205_98;
   assign m205_98 =10'b0;

   // m205_99 = W*in
   wire signed [9:0] m205_99;
   assign m205_99 =10'b0;

   // m205_100 = W*in
   wire signed [9:0] m205_100;
   assign m205_100 =10'b0;

   // m205_101 = W*in
   wire signed [9:0] m205_101;
   assign m205_101 =10'b0;

   // m205_102 = W*in
   wire signed [9:0] m205_102;
   assign m205_102 =10'b0;

   // m205_103 = W*in
   wire signed [9:0] m205_103;
   assign m205_103 =10'b0;

   // m205_104 = W*in
   wire signed [9:0] m205_104;
   assign m205_104 =10'b0;

   // m205_105 = W*in
   wire signed [9:0] m205_105;
   assign m205_105 =10'b0;

   // m205_106 = W*in
   wire signed [9:0] m205_106;
   assign m205_106 =10'b0;

   // m205_107 = W*in
   wire signed [9:0] m205_107;
   assign m205_107 =10'b0;

   // m205_108 = W*in
   wire signed [9:0] m205_108;
   assign m205_108 =10'b0;

   // m205_109 = W*in
   wire signed [9:0] m205_109;
   assign m205_109 =10'b0;

   // m205_110 = W*in
   wire signed [9:0] m205_110;
   assign m205_110 =10'b0;

   // m205_111 = W*in
   wire signed [9:0] m205_111;
   assign m205_111 =10'b0;

   // m205_112 = W*in
   wire signed [9:0] m205_112;
   assign m205_112 =10'b0;

   // m205_113 = W*in
   wire signed [9:0] m205_113;
   assign m205_113 =10'b0;

   // m205_114 = W*in
   wire signed [9:0] m205_114;
   assign m205_114 =10'b0;

   // m205_115 = W*in
   wire signed [9:0] m205_115;
   assign m205_115 =10'b0;

   // m205_116 = W*in
   wire signed [9:0] m205_116;
   assign m205_116 =10'b0;

   // m205_117 = W*in
   wire signed [9:0] m205_117;
   assign m205_117 =10'b0;

   // m206_1 = W*in
   wire signed [9:0] m206_1;
   assign m206_1 =10'b0;

   // m206_2 = W*in
   wire signed [9:0] m206_2;
   assign m206_2 =10'b0;

   // m206_3 = W*in
   wire signed [9:0] m206_3;
   assign m206_3 =10'b0;

   // m206_4 = W*in
   wire signed [9:0] m206_4;
   assign m206_4 =10'b0;

   // m206_5 = W*in
   wire signed [9:0] m206_5;
   assign m206_5 =10'b0;

   // m206_6 = W*in
   wire signed [9:0] m206_6;
   assign m206_6 =10'b0;

   // m206_7 = W*in
   wire signed [9:0] m206_7;
   assign m206_7 =10'b0;

   // m206_8 = W*in
   wire signed [9:0] m206_8;
   assign m206_8 =10'b0;

   // m206_9 = W*in
   wire signed [9:0] m206_9;
   assign m206_9 =10'b0;

   // m206_10 = W*in
   wire signed [9:0] m206_10;
   assign m206_10 =10'b0;

   // m206_11 = W*in
   wire signed [9:0] m206_11;
   assign m206_11 =10'b0;

   // m206_12 = W*in
   wire signed [9:0] m206_12;
   assign m206_12 =10'b0;

   // m206_13 = W*in
   wire signed [9:0] m206_13;
   assign m206_13 =10'b0;

   // m206_14 = W*in
   wire signed [9:0] m206_14;
   assign m206_14 =10'b0;

   // m206_15 = W*in
   wire signed [9:0] m206_15;
   assign m206_15 =10'b0;

   // m206_16 = W*in
   wire signed [9:0] m206_16;
   assign m206_16 =10'b0;

   // m206_17 = W*in
   wire signed [9:0] m206_17;
   assign m206_17 =10'b0;

   // m206_18 = W*in
   wire signed [9:0] m206_18;
   assign m206_18 =10'b0;

   // m206_19 = W*in
   wire signed [9:0] m206_19;
   assign m206_19 =10'b0;

   // m206_20 = W*in
   wire signed [9:0] m206_20;
   assign m206_20 =10'b0;

   // m206_21 = W*in
   wire signed [9:0] m206_21;
   assign m206_21 ={ {5{neg206[5]}} , neg206[5:1] };

   // m206_22 = W*in
   wire signed [9:0] m206_22;
   assign m206_22 =10'b0;

   // m206_23 = W*in
   wire signed [9:0] m206_23;
   assign m206_23 =10'b0;

   // m206_24 = W*in
   wire signed [9:0] m206_24;
   assign m206_24 =10'b0;

   // m206_25 = W*in
   wire signed [9:0] m206_25;
   assign m206_25 =10'b0;

   // m206_26 = W*in
   wire signed [9:0] m206_26;
   assign m206_26 =10'b0;

   // m206_27 = W*in
   wire signed [9:0] m206_27;
   assign m206_27 =10'b0;

   // m206_28 = W*in
   wire signed [9:0] m206_28;
   assign m206_28 =10'b0;

   // m206_29 = W*in
   wire signed [9:0] m206_29;
   assign m206_29 =10'b0;

   // m206_30 = W*in
   wire signed [9:0] m206_30;
   assign m206_30 =10'b0;

   // m206_31 = W*in
   wire signed [9:0] m206_31;
   assign m206_31 ={ {5{in206[5]}} , in206[5:1] };

   // m206_32 = W*in
   wire signed [9:0] m206_32;
   assign m206_32 =10'b0;

   // m206_33 = W*in
   wire signed [9:0] m206_33;
   assign m206_33 =10'b0;

   // m206_34 = W*in
   wire signed [9:0] m206_34;
   assign m206_34 =10'b0;

   // m206_35 = W*in
   wire signed [9:0] m206_35;
   assign m206_35 =10'b0;

   // m206_36 = W*in
   wire signed [9:0] m206_36;
   assign m206_36 =10'b0;

   // m206_37 = W*in
   wire signed [9:0] m206_37;
   assign m206_37 =10'b0;

   // m206_38 = W*in
   wire signed [9:0] m206_38;
   assign m206_38 =10'b0;

   // m206_39 = W*in
   wire signed [9:0] m206_39;
   assign m206_39 =10'b0;

   // m206_40 = W*in
   wire signed [9:0] m206_40;
   assign m206_40 =10'b0;

   // m206_41 = W*in
   wire signed [9:0] m206_41;
   assign m206_41 =10'b0;

   // m206_42 = W*in
   wire signed [9:0] m206_42;
   assign m206_42 =10'b0;

   // m206_43 = W*in
   wire signed [9:0] m206_43;
   assign m206_43 =10'b0;

   // m206_44 = W*in
   wire signed [9:0] m206_44;
   assign m206_44 =10'b0;

   // m206_45 = W*in
   wire signed [9:0] m206_45;
   assign m206_45 =10'b0;

   // m206_46 = W*in
   wire signed [9:0] m206_46;
   assign m206_46 =10'b0;

   // m206_47 = W*in
   wire signed [9:0] m206_47;
   assign m206_47 =10'b0;

   // m206_48 = W*in
   wire signed [9:0] m206_48;
   assign m206_48 =10'b0;

   // m206_49 = W*in
   wire signed [9:0] m206_49;
   assign m206_49 =10'b0;

   // m206_50 = W*in
   wire signed [9:0] m206_50;
   assign m206_50 =10'b0;

   // m206_51 = W*in
   wire signed [9:0] m206_51;
   assign m206_51 =10'b0;

   // m206_52 = W*in
   wire signed [9:0] m206_52;
   assign m206_52 =10'b0;

   // m206_53 = W*in
   wire signed [9:0] m206_53;
   assign m206_53 =10'b0;

   // m206_54 = W*in
   wire signed [9:0] m206_54;
   assign m206_54 =10'b0;

   // m206_55 = W*in
   wire signed [9:0] m206_55;
   assign m206_55 =10'b0;

   // m206_56 = W*in
   wire signed [9:0] m206_56;
   assign m206_56 =10'b0;

   // m206_57 = W*in
   wire signed [9:0] m206_57;
   assign m206_57 =10'b0;

   // m206_58 = W*in
   wire signed [9:0] m206_58;
   assign m206_58 =10'b0;

   // m206_59 = W*in
   wire signed [9:0] m206_59;
   assign m206_59 =10'b0;

   // m206_60 = W*in
   wire signed [9:0] m206_60;
   assign m206_60 =10'b0;

   // m206_61 = W*in
   wire signed [9:0] m206_61;
   assign m206_61 =10'b0;

   // m206_62 = W*in
   wire signed [9:0] m206_62;
   assign m206_62 =10'b0;

   // m206_63 = W*in
   wire signed [9:0] m206_63;
   assign m206_63 =10'b0;

   // m206_64 = W*in
   wire signed [9:0] m206_64;
   assign m206_64 =10'b0;

   // m206_65 = W*in
   wire signed [9:0] m206_65;
   assign m206_65 =10'b0;

   // m206_66 = W*in
   wire signed [9:0] m206_66;
   assign m206_66 =10'b0;

   // m206_67 = W*in
   wire signed [9:0] m206_67;
   assign m206_67 =10'b0;

   // m206_68 = W*in
   wire signed [9:0] m206_68;
   assign m206_68 =10'b0;

   // m206_69 = W*in
   wire signed [9:0] m206_69;
   assign m206_69 ={ {5{neg206[5]}} , neg206[5:1] };

   // m206_70 = W*in
   wire signed [9:0] m206_70;
   assign m206_70 =10'b0;

   // m206_71 = W*in
   wire signed [9:0] m206_71;
   assign m206_71 =10'b0;

   // m206_72 = W*in
   wire signed [9:0] m206_72;
   assign m206_72 =10'b0;

   // m206_73 = W*in
   wire signed [9:0] m206_73;
   assign m206_73 =10'b0;

   // m206_74 = W*in
   wire signed [9:0] m206_74;
   assign m206_74 =10'b0;

   // m206_75 = W*in
   wire signed [9:0] m206_75;
   assign m206_75 =10'b0;

   // m206_76 = W*in
   wire signed [9:0] m206_76;
   assign m206_76 =10'b0;

   // m206_77 = W*in
   wire signed [9:0] m206_77;
   assign m206_77 =10'b0;

   // m206_78 = W*in
   wire signed [9:0] m206_78;
   assign m206_78 =10'b0;

   // m206_79 = W*in
   wire signed [9:0] m206_79;
   assign m206_79 =10'b0;

   // m206_80 = W*in
   wire signed [9:0] m206_80;
   assign m206_80 =10'b0;

   // m206_81 = W*in
   wire signed [9:0] m206_81;
   assign m206_81 =10'b0;

   // m206_82 = W*in
   wire signed [9:0] m206_82;
   assign m206_82 =10'b0;

   // m206_83 = W*in
   wire signed [9:0] m206_83;
   assign m206_83 =10'b0;

   // m206_84 = W*in
   wire signed [9:0] m206_84;
   assign m206_84 =10'b0;

   // m206_85 = W*in
   wire signed [9:0] m206_85;
   assign m206_85 =10'b0;

   // m206_86 = W*in
   wire signed [9:0] m206_86;
   assign m206_86 =10'b0;

   // m206_87 = W*in
   wire signed [9:0] m206_87;
   assign m206_87 =10'b0;

   // m206_88 = W*in
   wire signed [9:0] m206_88;
   assign m206_88 =10'b0;

   // m206_89 = W*in
   wire signed [9:0] m206_89;
   assign m206_89 =10'b0;

   // m206_90 = W*in
   wire signed [9:0] m206_90;
   assign m206_90 =10'b0;

   // m206_91 = W*in
   wire signed [9:0] m206_91;
   assign m206_91 =10'b0;

   // m206_92 = W*in
   wire signed [9:0] m206_92;
   assign m206_92 =10'b0;

   // m206_93 = W*in
   wire signed [9:0] m206_93;
   assign m206_93 =10'b0;

   // m206_94 = W*in
   wire signed [9:0] m206_94;
   assign m206_94 =10'b0;

   // m206_95 = W*in
   wire signed [9:0] m206_95;
   assign m206_95 =10'b0;

   // m206_96 = W*in
   wire signed [9:0] m206_96;
   assign m206_96 =10'b0;

   // m206_97 = W*in
   wire signed [9:0] m206_97;
   assign m206_97 =10'b0;

   // m206_98 = W*in
   wire signed [9:0] m206_98;
   assign m206_98 =10'b0;

   // m206_99 = W*in
   wire signed [9:0] m206_99;
   assign m206_99 =10'b0;

   // m206_100 = W*in
   wire signed [9:0] m206_100;
   assign m206_100 =10'b0;

   // m206_101 = W*in
   wire signed [9:0] m206_101;
   assign m206_101 =10'b0;

   // m206_102 = W*in
   wire signed [9:0] m206_102;
   assign m206_102 =10'b0;

   // m206_103 = W*in
   wire signed [9:0] m206_103;
   assign m206_103 =10'b0;

   // m206_104 = W*in
   wire signed [9:0] m206_104;
   assign m206_104 =10'b0;

   // m206_105 = W*in
   wire signed [9:0] m206_105;
   assign m206_105 =10'b0;

   // m206_106 = W*in
   wire signed [9:0] m206_106;
   assign m206_106 =10'b0;

   // m206_107 = W*in
   wire signed [9:0] m206_107;
   assign m206_107 =10'b0;

   // m206_108 = W*in
   wire signed [9:0] m206_108;
   assign m206_108 ={ {5{neg206[5]}} , neg206[5:1] };

   // m206_109 = W*in
   wire signed [9:0] m206_109;
   assign m206_109 =10'b0;

   // m206_110 = W*in
   wire signed [9:0] m206_110;
   assign m206_110 =10'b0;

   // m206_111 = W*in
   wire signed [9:0] m206_111;
   assign m206_111 =10'b0;

   // m206_112 = W*in
   wire signed [9:0] m206_112;
   assign m206_112 =10'b0;

   // m206_113 = W*in
   wire signed [9:0] m206_113;
   assign m206_113 =10'b0;

   // m206_114 = W*in
   wire signed [9:0] m206_114;
   assign m206_114 =10'b0;

   // m206_115 = W*in
   wire signed [9:0] m206_115;
   assign m206_115 =10'b0;

   // m206_116 = W*in
   wire signed [9:0] m206_116;
   assign m206_116 =10'b0;

   // m206_117 = W*in
   wire signed [9:0] m206_117;
   assign m206_117 =10'b0;

   // m207_1 = W*in
   wire signed [9:0] m207_1;
   assign m207_1 =10'b0;

   // m207_2 = W*in
   wire signed [9:0] m207_2;
   assign m207_2 =10'b0;

   // m207_3 = W*in
   wire signed [9:0] m207_3;
   assign m207_3 =10'b0;

   // m207_4 = W*in
   wire signed [9:0] m207_4;
   assign m207_4 =10'b0;

   // m207_5 = W*in
   wire signed [9:0] m207_5;
   assign m207_5 =10'b0;

   // m207_6 = W*in
   wire signed [9:0] m207_6;
   assign m207_6 =10'b0;

   // m207_7 = W*in
   wire signed [9:0] m207_7;
   assign m207_7 =10'b0;

   // m207_8 = W*in
   wire signed [9:0] m207_8;
   assign m207_8 =10'b0;

   // m207_9 = W*in
   wire signed [9:0] m207_9;
   assign m207_9 =10'b0;

   // m207_10 = W*in
   wire signed [9:0] m207_10;
   assign m207_10 =10'b0;

   // m207_11 = W*in
   wire signed [9:0] m207_11;
   assign m207_11 =10'b0;

   // m207_12 = W*in
   wire signed [9:0] m207_12;
   assign m207_12 =10'b0;

   // m207_13 = W*in
   wire signed [9:0] m207_13;
   assign m207_13 =10'b0;

   // m207_14 = W*in
   wire signed [9:0] m207_14;
   assign m207_14 =10'b0;

   // m207_15 = W*in
   wire signed [9:0] m207_15;
   assign m207_15 =10'b0;

   // m207_16 = W*in
   wire signed [9:0] m207_16;
   assign m207_16 =10'b0;

   // m207_17 = W*in
   wire signed [9:0] m207_17;
   assign m207_17 =10'b0;

   // m207_18 = W*in
   wire signed [9:0] m207_18;
   assign m207_18 =10'b0;

   // m207_19 = W*in
   wire signed [9:0] m207_19;
   assign m207_19 =10'b0;

   // m207_20 = W*in
   wire signed [9:0] m207_20;
   assign m207_20 =10'b0;

   // m207_21 = W*in
   wire signed [9:0] m207_21;
   assign m207_21 =10'b0;

   // m207_22 = W*in
   wire signed [9:0] m207_22;
   assign m207_22 =10'b0;

   // m207_23 = W*in
   wire signed [9:0] m207_23;
   assign m207_23 =10'b0;

   // m207_24 = W*in
   wire signed [9:0] m207_24;
   assign m207_24 =10'b0;

   // m207_25 = W*in
   wire signed [9:0] m207_25;
   assign m207_25 =10'b0;

   // m207_26 = W*in
   wire signed [9:0] m207_26;
   assign m207_26 =10'b0;

   // m207_27 = W*in
   wire signed [9:0] m207_27;
   assign m207_27 =10'b0;

   // m207_28 = W*in
   wire signed [9:0] m207_28;
   assign m207_28 =10'b0;

   // m207_29 = W*in
   wire signed [9:0] m207_29;
   assign m207_29 =10'b0;

   // m207_30 = W*in
   wire signed [9:0] m207_30;
   assign m207_30 =10'b0;

   // m207_31 = W*in
   wire signed [9:0] m207_31;
   assign m207_31 =10'b0;

   // m207_32 = W*in
   wire signed [9:0] m207_32;
   assign m207_32 =10'b0;

   // m207_33 = W*in
   wire signed [9:0] m207_33;
   assign m207_33 =10'b0;

   // m207_34 = W*in
   wire signed [9:0] m207_34;
   assign m207_34 =10'b0;

   // m207_35 = W*in
   wire signed [9:0] m207_35;
   assign m207_35 =10'b0;

   // m207_36 = W*in
   wire signed [9:0] m207_36;
   assign m207_36 =10'b0;

   // m207_37 = W*in
   wire signed [9:0] m207_37;
   assign m207_37 =10'b0;

   // m207_38 = W*in
   wire signed [9:0] m207_38;
   assign m207_38 =10'b0;

   // m207_39 = W*in
   wire signed [9:0] m207_39;
   assign m207_39 =10'b0;

   // m207_40 = W*in
   wire signed [9:0] m207_40;
   assign m207_40 =10'b0;

   // m207_41 = W*in
   wire signed [9:0] m207_41;
   assign m207_41 =10'b0;

   // m207_42 = W*in
   wire signed [9:0] m207_42;
   assign m207_42 =10'b0;

   // m207_43 = W*in
   wire signed [9:0] m207_43;
   assign m207_43 =10'b0;

   // m207_44 = W*in
   wire signed [9:0] m207_44;
   assign m207_44 =10'b0;

   // m207_45 = W*in
   wire signed [9:0] m207_45;
   assign m207_45 =10'b0;

   // m207_46 = W*in
   wire signed [9:0] m207_46;
   assign m207_46 =10'b0;

   // m207_47 = W*in
   wire signed [9:0] m207_47;
   assign m207_47 =10'b0;

   // m207_48 = W*in
   wire signed [9:0] m207_48;
   assign m207_48 =10'b0;

   // m207_49 = W*in
   wire signed [9:0] m207_49;
   assign m207_49 =10'b0;

   // m207_50 = W*in
   wire signed [9:0] m207_50;
   assign m207_50 =10'b0;

   // m207_51 = W*in
   wire signed [9:0] m207_51;
   assign m207_51 =10'b0;

   // m207_52 = W*in
   wire signed [9:0] m207_52;
   assign m207_52 =10'b0;

   // m207_53 = W*in
   wire signed [9:0] m207_53;
   assign m207_53 =10'b0;

   // m207_54 = W*in
   wire signed [9:0] m207_54;
   assign m207_54 =10'b0;

   // m207_55 = W*in
   wire signed [9:0] m207_55;
   assign m207_55 =10'b0;

   // m207_56 = W*in
   wire signed [9:0] m207_56;
   assign m207_56 =10'b0;

   // m207_57 = W*in
   wire signed [9:0] m207_57;
   assign m207_57 =10'b0;

   // m207_58 = W*in
   wire signed [9:0] m207_58;
   assign m207_58 =10'b0;

   // m207_59 = W*in
   wire signed [9:0] m207_59;
   assign m207_59 =10'b0;

   // m207_60 = W*in
   wire signed [9:0] m207_60;
   assign m207_60 =10'b0;

   // m207_61 = W*in
   wire signed [9:0] m207_61;
   assign m207_61 =10'b0;

   // m207_62 = W*in
   wire signed [9:0] m207_62;
   assign m207_62 =10'b0;

   // m207_63 = W*in
   wire signed [9:0] m207_63;
   assign m207_63 =10'b0;

   // m207_64 = W*in
   wire signed [9:0] m207_64;
   assign m207_64 =10'b0;

   // m207_65 = W*in
   wire signed [9:0] m207_65;
   assign m207_65 =10'b0;

   // m207_66 = W*in
   wire signed [9:0] m207_66;
   assign m207_66 =10'b0;

   // m207_67 = W*in
   wire signed [9:0] m207_67;
   assign m207_67 =10'b0;

   // m207_68 = W*in
   wire signed [9:0] m207_68;
   assign m207_68 =10'b0;

   // m207_69 = W*in
   wire signed [9:0] m207_69;
   assign m207_69 =10'b0;

   // m207_70 = W*in
   wire signed [9:0] m207_70;
   assign m207_70 =10'b0;

   // m207_71 = W*in
   wire signed [9:0] m207_71;
   assign m207_71 =10'b0;

   // m207_72 = W*in
   wire signed [9:0] m207_72;
   assign m207_72 ={ {5{neg207[5]}} , neg207[5:1] };

   // m207_73 = W*in
   wire signed [9:0] m207_73;
   assign m207_73 =10'b0;

   // m207_74 = W*in
   wire signed [9:0] m207_74;
   assign m207_74 =10'b0;

   // m207_75 = W*in
   wire signed [9:0] m207_75;
   assign m207_75 =10'b0;

   // m207_76 = W*in
   wire signed [9:0] m207_76;
   assign m207_76 =10'b0;

   // m207_77 = W*in
   wire signed [9:0] m207_77;
   assign m207_77 =10'b0;

   // m207_78 = W*in
   wire signed [9:0] m207_78;
   assign m207_78 =10'b0;

   // m207_79 = W*in
   wire signed [9:0] m207_79;
   assign m207_79 =10'b0;

   // m207_80 = W*in
   wire signed [9:0] m207_80;
   assign m207_80 =10'b0;

   // m207_81 = W*in
   wire signed [9:0] m207_81;
   assign m207_81 =10'b0;

   // m207_82 = W*in
   wire signed [9:0] m207_82;
   assign m207_82 =10'b0;

   // m207_83 = W*in
   wire signed [9:0] m207_83;
   assign m207_83 =10'b0;

   // m207_84 = W*in
   wire signed [9:0] m207_84;
   assign m207_84 =10'b0;

   // m207_85 = W*in
   wire signed [9:0] m207_85;
   assign m207_85 =10'b0;

   // m207_86 = W*in
   wire signed [9:0] m207_86;
   assign m207_86 =10'b0;

   // m207_87 = W*in
   wire signed [9:0] m207_87;
   assign m207_87 =10'b0;

   // m207_88 = W*in
   wire signed [9:0] m207_88;
   assign m207_88 =10'b0;

   // m207_89 = W*in
   wire signed [9:0] m207_89;
   assign m207_89 =10'b0;

   // m207_90 = W*in
   wire signed [9:0] m207_90;
   assign m207_90 =10'b0;

   // m207_91 = W*in
   wire signed [9:0] m207_91;
   assign m207_91 =10'b0;

   // m207_92 = W*in
   wire signed [9:0] m207_92;
   assign m207_92 =10'b0;

   // m207_93 = W*in
   wire signed [9:0] m207_93;
   assign m207_93 =10'b0;

   // m207_94 = W*in
   wire signed [9:0] m207_94;
   assign m207_94 =10'b0;

   // m207_95 = W*in
   wire signed [9:0] m207_95;
   assign m207_95 =10'b0;

   // m207_96 = W*in
   wire signed [9:0] m207_96;
   assign m207_96 =10'b0;

   // m207_97 = W*in
   wire signed [9:0] m207_97;
   assign m207_97 =10'b0;

   // m207_98 = W*in
   wire signed [9:0] m207_98;
   assign m207_98 =10'b0;

   // m207_99 = W*in
   wire signed [9:0] m207_99;
   assign m207_99 =10'b0;

   // m207_100 = W*in
   wire signed [9:0] m207_100;
   assign m207_100 =10'b0;

   // m207_101 = W*in
   wire signed [9:0] m207_101;
   assign m207_101 =10'b0;

   // m207_102 = W*in
   wire signed [9:0] m207_102;
   assign m207_102 =10'b0;

   // m207_103 = W*in
   wire signed [9:0] m207_103;
   assign m207_103 =10'b0;

   // m207_104 = W*in
   wire signed [9:0] m207_104;
   assign m207_104 =10'b0;

   // m207_105 = W*in
   wire signed [9:0] m207_105;
   assign m207_105 =10'b0;

   // m207_106 = W*in
   wire signed [9:0] m207_106;
   assign m207_106 =10'b0;

   // m207_107 = W*in
   wire signed [9:0] m207_107;
   assign m207_107 =10'b0;

   // m207_108 = W*in
   wire signed [9:0] m207_108;
   assign m207_108 =10'b0;

   // m207_109 = W*in
   wire signed [9:0] m207_109;
   assign m207_109 =10'b0;

   // m207_110 = W*in
   wire signed [9:0] m207_110;
   assign m207_110 =10'b0;

   // m207_111 = W*in
   wire signed [9:0] m207_111;
   assign m207_111 =10'b0;

   // m207_112 = W*in
   wire signed [9:0] m207_112;
   assign m207_112 =10'b0;

   // m207_113 = W*in
   wire signed [9:0] m207_113;
   assign m207_113 =10'b0;

   // m207_114 = W*in
   wire signed [9:0] m207_114;
   assign m207_114 =10'b0;

   // m207_115 = W*in
   wire signed [9:0] m207_115;
   assign m207_115 =10'b0;

   // m207_116 = W*in
   wire signed [9:0] m207_116;
   assign m207_116 =10'b0;

   // m207_117 = W*in
   wire signed [9:0] m207_117;
   assign m207_117 =10'b0;

   // m208_1 = W*in
   wire signed [9:0] m208_1;
   assign m208_1 =10'b0;

   // m208_2 = W*in
   wire signed [9:0] m208_2;
   assign m208_2 =10'b0;

   // m208_3 = W*in
   wire signed [9:0] m208_3;
   assign m208_3 =10'b0;

   // m208_4 = W*in
   wire signed [9:0] m208_4;
   assign m208_4 =10'b0;

   // m208_5 = W*in
   wire signed [9:0] m208_5;
   assign m208_5 =10'b0;

   // m208_6 = W*in
   wire signed [9:0] m208_6;
   assign m208_6 =10'b0;

   // m208_7 = W*in
   wire signed [9:0] m208_7;
   assign m208_7 =10'b0;

   // m208_8 = W*in
   wire signed [9:0] m208_8;
   assign m208_8 =10'b0;

   // m208_9 = W*in
   wire signed [9:0] m208_9;
   assign m208_9 =10'b0;

   // m208_10 = W*in
   wire signed [9:0] m208_10;
   assign m208_10 =10'b0;

   // m208_11 = W*in
   wire signed [9:0] m208_11;
   assign m208_11 =10'b0;

   // m208_12 = W*in
   wire signed [9:0] m208_12;
   assign m208_12 =10'b0;

   // m208_13 = W*in
   wire signed [9:0] m208_13;
   assign m208_13 =10'b0;

   // m208_14 = W*in
   wire signed [9:0] m208_14;
   assign m208_14 =10'b0;

   // m208_15 = W*in
   wire signed [9:0] m208_15;
   assign m208_15 =10'b0;

   // m208_16 = W*in
   wire signed [9:0] m208_16;
   assign m208_16 =10'b0;

   // m208_17 = W*in
   wire signed [9:0] m208_17;
   assign m208_17 =10'b0;

   // m208_18 = W*in
   wire signed [9:0] m208_18;
   assign m208_18 =10'b0;

   // m208_19 = W*in
   wire signed [9:0] m208_19;
   assign m208_19 =10'b0;

   // m208_20 = W*in
   wire signed [9:0] m208_20;
   assign m208_20 =10'b0;

   // m208_21 = W*in
   wire signed [9:0] m208_21;
   assign m208_21 =10'b0;

   // m208_22 = W*in
   wire signed [9:0] m208_22;
   assign m208_22 =10'b0;

   // m208_23 = W*in
   wire signed [9:0] m208_23;
   assign m208_23 =10'b0;

   // m208_24 = W*in
   wire signed [9:0] m208_24;
   assign m208_24 =10'b0;

   // m208_25 = W*in
   wire signed [9:0] m208_25;
   assign m208_25 =10'b0;

   // m208_26 = W*in
   wire signed [9:0] m208_26;
   assign m208_26 =10'b0;

   // m208_27 = W*in
   wire signed [9:0] m208_27;
   assign m208_27 =10'b0;

   // m208_28 = W*in
   wire signed [9:0] m208_28;
   assign m208_28 =10'b0;

   // m208_29 = W*in
   wire signed [9:0] m208_29;
   assign m208_29 =10'b0;

   // m208_30 = W*in
   wire signed [9:0] m208_30;
   assign m208_30 =10'b0;

   // m208_31 = W*in
   wire signed [9:0] m208_31;
   assign m208_31 =10'b0;

   // m208_32 = W*in
   wire signed [9:0] m208_32;
   assign m208_32 =10'b0;

   // m208_33 = W*in
   wire signed [9:0] m208_33;
   assign m208_33 =10'b0;

   // m208_34 = W*in
   wire signed [9:0] m208_34;
   assign m208_34 =10'b0;

   // m208_35 = W*in
   wire signed [9:0] m208_35;
   assign m208_35 =10'b0;

   // m208_36 = W*in
   wire signed [9:0] m208_36;
   assign m208_36 =10'b0;

   // m208_37 = W*in
   wire signed [9:0] m208_37;
   assign m208_37 =10'b0;

   // m208_38 = W*in
   wire signed [9:0] m208_38;
   assign m208_38 =10'b0;

   // m208_39 = W*in
   wire signed [9:0] m208_39;
   assign m208_39 =10'b0;

   // m208_40 = W*in
   wire signed [9:0] m208_40;
   assign m208_40 =10'b0;

   // m208_41 = W*in
   wire signed [9:0] m208_41;
   assign m208_41 =10'b0;

   // m208_42 = W*in
   wire signed [9:0] m208_42;
   assign m208_42 =10'b0;

   // m208_43 = W*in
   wire signed [9:0] m208_43;
   assign m208_43 =10'b0;

   // m208_44 = W*in
   wire signed [9:0] m208_44;
   assign m208_44 =10'b0;

   // m208_45 = W*in
   wire signed [9:0] m208_45;
   assign m208_45 =10'b0;

   // m208_46 = W*in
   wire signed [9:0] m208_46;
   assign m208_46 =10'b0;

   // m208_47 = W*in
   wire signed [9:0] m208_47;
   assign m208_47 =10'b0;

   // m208_48 = W*in
   wire signed [9:0] m208_48;
   assign m208_48 =10'b0;

   // m208_49 = W*in
   wire signed [9:0] m208_49;
   assign m208_49 =10'b0;

   // m208_50 = W*in
   wire signed [9:0] m208_50;
   assign m208_50 =10'b0;

   // m208_51 = W*in
   wire signed [9:0] m208_51;
   assign m208_51 =10'b0;

   // m208_52 = W*in
   wire signed [9:0] m208_52;
   assign m208_52 =10'b0;

   // m208_53 = W*in
   wire signed [9:0] m208_53;
   assign m208_53 =10'b0;

   // m208_54 = W*in
   wire signed [9:0] m208_54;
   assign m208_54 =10'b0;

   // m208_55 = W*in
   wire signed [9:0] m208_55;
   assign m208_55 =10'b0;

   // m208_56 = W*in
   wire signed [9:0] m208_56;
   assign m208_56 =10'b0;

   // m208_57 = W*in
   wire signed [9:0] m208_57;
   assign m208_57 =10'b0;

   // m208_58 = W*in
   wire signed [9:0] m208_58;
   assign m208_58 =10'b0;

   // m208_59 = W*in
   wire signed [9:0] m208_59;
   assign m208_59 =10'b0;

   // m208_60 = W*in
   wire signed [9:0] m208_60;
   assign m208_60 =10'b0;

   // m208_61 = W*in
   wire signed [9:0] m208_61;
   assign m208_61 =10'b0;

   // m208_62 = W*in
   wire signed [9:0] m208_62;
   assign m208_62 =10'b0;

   // m208_63 = W*in
   wire signed [9:0] m208_63;
   assign m208_63 =10'b0;

   // m208_64 = W*in
   wire signed [9:0] m208_64;
   assign m208_64 =10'b0;

   // m208_65 = W*in
   wire signed [9:0] m208_65;
   assign m208_65 =10'b0;

   // m208_66 = W*in
   wire signed [9:0] m208_66;
   assign m208_66 =10'b0;

   // m208_67 = W*in
   wire signed [9:0] m208_67;
   assign m208_67 =10'b0;

   // m208_68 = W*in
   wire signed [9:0] m208_68;
   assign m208_68 =10'b0;

   // m208_69 = W*in
   wire signed [9:0] m208_69;
   assign m208_69 =10'b0;

   // m208_70 = W*in
   wire signed [9:0] m208_70;
   assign m208_70 =10'b0;

   // m208_71 = W*in
   wire signed [9:0] m208_71;
   assign m208_71 =10'b0;

   // m208_72 = W*in
   wire signed [9:0] m208_72;
   assign m208_72 =10'b0;

   // m208_73 = W*in
   wire signed [9:0] m208_73;
   assign m208_73 =10'b0;

   // m208_74 = W*in
   wire signed [9:0] m208_74;
   assign m208_74 =10'b0;

   // m208_75 = W*in
   wire signed [9:0] m208_75;
   assign m208_75 =10'b0;

   // m208_76 = W*in
   wire signed [9:0] m208_76;
   assign m208_76 =10'b0;

   // m208_77 = W*in
   wire signed [9:0] m208_77;
   assign m208_77 =10'b0;

   // m208_78 = W*in
   wire signed [9:0] m208_78;
   assign m208_78 ={ {5{neg208[5]}} , neg208[5:1] };

   // m208_79 = W*in
   wire signed [9:0] m208_79;
   assign m208_79 =10'b0;

   // m208_80 = W*in
   wire signed [9:0] m208_80;
   assign m208_80 =10'b0;

   // m208_81 = W*in
   wire signed [9:0] m208_81;
   assign m208_81 =10'b0;

   // m208_82 = W*in
   wire signed [9:0] m208_82;
   assign m208_82 =10'b0;

   // m208_83 = W*in
   wire signed [9:0] m208_83;
   assign m208_83 =10'b0;

   // m208_84 = W*in
   wire signed [9:0] m208_84;
   assign m208_84 =10'b0;

   // m208_85 = W*in
   wire signed [9:0] m208_85;
   assign m208_85 =10'b0;

   // m208_86 = W*in
   wire signed [9:0] m208_86;
   assign m208_86 =10'b0;

   // m208_87 = W*in
   wire signed [9:0] m208_87;
   assign m208_87 =10'b0;

   // m208_88 = W*in
   wire signed [9:0] m208_88;
   assign m208_88 =10'b0;

   // m208_89 = W*in
   wire signed [9:0] m208_89;
   assign m208_89 =10'b0;

   // m208_90 = W*in
   wire signed [9:0] m208_90;
   assign m208_90 =10'b0;

   // m208_91 = W*in
   wire signed [9:0] m208_91;
   assign m208_91 =10'b0;

   // m208_92 = W*in
   wire signed [9:0] m208_92;
   assign m208_92 =10'b0;

   // m208_93 = W*in
   wire signed [9:0] m208_93;
   assign m208_93 =10'b0;

   // m208_94 = W*in
   wire signed [9:0] m208_94;
   assign m208_94 =10'b0;

   // m208_95 = W*in
   wire signed [9:0] m208_95;
   assign m208_95 =10'b0;

   // m208_96 = W*in
   wire signed [9:0] m208_96;
   assign m208_96 =10'b0;

   // m208_97 = W*in
   wire signed [9:0] m208_97;
   assign m208_97 =10'b0;

   // m208_98 = W*in
   wire signed [9:0] m208_98;
   assign m208_98 =10'b0;

   // m208_99 = W*in
   wire signed [9:0] m208_99;
   assign m208_99 =10'b0;

   // m208_100 = W*in
   wire signed [9:0] m208_100;
   assign m208_100 =10'b0;

   // m208_101 = W*in
   wire signed [9:0] m208_101;
   assign m208_101 =10'b0;

   // m208_102 = W*in
   wire signed [9:0] m208_102;
   assign m208_102 =10'b0;

   // m208_103 = W*in
   wire signed [9:0] m208_103;
   assign m208_103 =10'b0;

   // m208_104 = W*in
   wire signed [9:0] m208_104;
   assign m208_104 =10'b0;

   // m208_105 = W*in
   wire signed [9:0] m208_105;
   assign m208_105 =10'b0;

   // m208_106 = W*in
   wire signed [9:0] m208_106;
   assign m208_106 =10'b0;

   // m208_107 = W*in
   wire signed [9:0] m208_107;
   assign m208_107 =10'b0;

   // m208_108 = W*in
   wire signed [9:0] m208_108;
   assign m208_108 =10'b0;

   // m208_109 = W*in
   wire signed [9:0] m208_109;
   assign m208_109 =10'b0;

   // m208_110 = W*in
   wire signed [9:0] m208_110;
   assign m208_110 =10'b0;

   // m208_111 = W*in
   wire signed [9:0] m208_111;
   assign m208_111 =10'b0;

   // m208_112 = W*in
   wire signed [9:0] m208_112;
   assign m208_112 =10'b0;

   // m208_113 = W*in
   wire signed [9:0] m208_113;
   assign m208_113 =10'b0;

   // m208_114 = W*in
   wire signed [9:0] m208_114;
   assign m208_114 =10'b0;

   // m208_115 = W*in
   wire signed [9:0] m208_115;
   assign m208_115 =10'b0;

   // m208_116 = W*in
   wire signed [9:0] m208_116;
   assign m208_116 =10'b0;

   // m208_117 = W*in
   wire signed [9:0] m208_117;
   assign m208_117 =10'b0;

   // m209_1 = W*in
   wire signed [9:0] m209_1;
   assign m209_1 =10'b0;

   // m209_2 = W*in
   wire signed [9:0] m209_2;
   assign m209_2 =10'b0;

   // m209_3 = W*in
   wire signed [9:0] m209_3;
   assign m209_3 =10'b0;

   // m209_4 = W*in
   wire signed [9:0] m209_4;
   assign m209_4 =10'b0;

   // m209_5 = W*in
   wire signed [9:0] m209_5;
   assign m209_5 =10'b0;

   // m209_6 = W*in
   wire signed [9:0] m209_6;
   assign m209_6 =10'b0;

   // m209_7 = W*in
   wire signed [9:0] m209_7;
   assign m209_7 =10'b0;

   // m209_8 = W*in
   wire signed [9:0] m209_8;
   assign m209_8 ={ {4{in209[5]}} , in209[5:0] };

   // m209_9 = W*in
   wire signed [9:0] m209_9;
   assign m209_9 =10'b0;

   // m209_10 = W*in
   wire signed [9:0] m209_10;
   assign m209_10 =10'b0;

   // m209_11 = W*in
   wire signed [9:0] m209_11;
   assign m209_11 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_12 = W*in
   wire signed [9:0] m209_12;
   assign m209_12 =10'b0;

   // m209_13 = W*in
   wire signed [9:0] m209_13;
   assign m209_13 =10'b0;

   // m209_14 = W*in
   wire signed [9:0] m209_14;
   assign m209_14 =10'b0;

   // m209_15 = W*in
   wire signed [9:0] m209_15;
   assign m209_15 =10'b0;

   // m209_16 = W*in
   wire signed [9:0] m209_16;
   assign m209_16 =10'b0;

   // m209_17 = W*in
   wire signed [9:0] m209_17;
   assign m209_17 =10'b0;

   // m209_18 = W*in
   wire signed [9:0] m209_18;
   assign m209_18 =10'b0;

   // m209_19 = W*in
   wire signed [9:0] m209_19;
   assign m209_19 =10'b0;

   // m209_20 = W*in
   wire signed [9:0] m209_20;
   assign m209_20 =10'b0;

   // m209_21 = W*in
   wire signed [9:0] m209_21;
   assign m209_21 =10'b0;

   // m209_22 = W*in
   wire signed [9:0] m209_22;
   assign m209_22 =10'b0;

   // m209_23 = W*in
   wire signed [9:0] m209_23;
   assign m209_23 =10'b0;

   // m209_24 = W*in
   wire signed [9:0] m209_24;
   assign m209_24 =10'b0;

   // m209_25 = W*in
   wire signed [9:0] m209_25;
   assign m209_25 =10'b0;

   // m209_26 = W*in
   wire signed [9:0] m209_26;
   assign m209_26 ={ {5{neg209[5]}} , neg209[5:1] };

   // m209_27 = W*in
   wire signed [9:0] m209_27;
   assign m209_27 =10'b0;

   // m209_28 = W*in
   wire signed [9:0] m209_28;
   assign m209_28 =10'b0;

   // m209_29 = W*in
   wire signed [9:0] m209_29;
   assign m209_29 =10'b0;

   // m209_30 = W*in
   wire signed [9:0] m209_30;
   assign m209_30 =10'b0;

   // m209_31 = W*in
   wire signed [9:0] m209_31;
   assign m209_31 ={ {5{in209[5]}} , in209[5:1] };

   // m209_32 = W*in
   wire signed [9:0] m209_32;
   assign m209_32 =10'b0;

   // m209_33 = W*in
   wire signed [9:0] m209_33;
   assign m209_33 =10'b0;

   // m209_34 = W*in
   wire signed [9:0] m209_34;
   assign m209_34 =10'b0;

   // m209_35 = W*in
   wire signed [9:0] m209_35;
   assign m209_35 =10'b0;

   // m209_36 = W*in
   wire signed [9:0] m209_36;
   assign m209_36 =10'b0;

   // m209_37 = W*in
   wire signed [9:0] m209_37;
   assign m209_37 =10'b0;

   // m209_38 = W*in
   wire signed [9:0] m209_38;
   assign m209_38 =10'b0;

   // m209_39 = W*in
   wire signed [9:0] m209_39;
   assign m209_39 =10'b0;

   // m209_40 = W*in
   wire signed [9:0] m209_40;
   assign m209_40 =10'b0;

   // m209_41 = W*in
   wire signed [9:0] m209_41;
   assign m209_41 =10'b0;

   // m209_42 = W*in
   wire signed [9:0] m209_42;
   assign m209_42 =10'b0;

   // m209_43 = W*in
   wire signed [9:0] m209_43;
   assign m209_43 =10'b0;

   // m209_44 = W*in
   wire signed [9:0] m209_44;
   assign m209_44 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_45 = W*in
   wire signed [9:0] m209_45;
   assign m209_45 ={ {4{in209[5]}} , in209[5:0] };

   // m209_46 = W*in
   wire signed [9:0] m209_46;
   assign m209_46 =10'b0;

   // m209_47 = W*in
   wire signed [9:0] m209_47;
   assign m209_47 =10'b0;

   // m209_48 = W*in
   wire signed [9:0] m209_48;
   assign m209_48 =10'b0;

   // m209_49 = W*in
   wire signed [9:0] m209_49;
   assign m209_49 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_50 = W*in
   wire signed [9:0] m209_50;
   assign m209_50 =10'b0;

   // m209_51 = W*in
   wire signed [9:0] m209_51;
   assign m209_51 ={ {4{in209[5]}} , in209[5:0] };

   // m209_52 = W*in
   wire signed [9:0] m209_52;
   assign m209_52 =10'b0;

   // m209_53 = W*in
   wire signed [9:0] m209_53;
   assign m209_53 =10'b0;

   // m209_54 = W*in
   wire signed [9:0] m209_54;
   assign m209_54 =10'b0;

   // m209_55 = W*in
   wire signed [9:0] m209_55;
   assign m209_55 =10'b0;

   // m209_56 = W*in
   wire signed [9:0] m209_56;
   assign m209_56 =10'b0;

   // m209_57 = W*in
   wire signed [9:0] m209_57;
   assign m209_57 =10'b0;

   // m209_58 = W*in
   wire signed [9:0] m209_58;
   assign m209_58 =10'b0;

   // m209_59 = W*in
   wire signed [9:0] m209_59;
   assign m209_59 =10'b0;

   // m209_60 = W*in
   wire signed [9:0] m209_60;
   assign m209_60 =10'b0;

   // m209_61 = W*in
   wire signed [9:0] m209_61;
   assign m209_61 =10'b0;

   // m209_62 = W*in
   wire signed [9:0] m209_62;
   assign m209_62 =10'b0;

   // m209_63 = W*in
   wire signed [9:0] m209_63;
   assign m209_63 =10'b0;

   // m209_64 = W*in
   wire signed [9:0] m209_64;
   assign m209_64 =10'b0;

   // m209_65 = W*in
   wire signed [9:0] m209_65;
   assign m209_65 =10'b0;

   // m209_66 = W*in
   wire signed [9:0] m209_66;
   assign m209_66 ={ {5{neg209[5]}} , neg209[5:1] };

   // m209_67 = W*in
   wire signed [9:0] m209_67;
   assign m209_67 =10'b0;

   // m209_68 = W*in
   wire signed [9:0] m209_68;
   assign m209_68 =10'b0;

   // m209_69 = W*in
   wire signed [9:0] m209_69;
   assign m209_69 ={ {5{neg209[5]}} , neg209[5:1] };

   // m209_70 = W*in
   wire signed [9:0] m209_70;
   assign m209_70 ={ {5{neg209[5]}} , neg209[5:1] };

   // m209_71 = W*in
   wire signed [9:0] m209_71;
   assign m209_71 ={ {5{neg209[5]}} , neg209[5:1] };

   // m209_72 = W*in
   wire signed [9:0] m209_72;
   assign m209_72 =10'b0;

   // m209_73 = W*in
   wire signed [9:0] m209_73;
   assign m209_73 ={ {4{in209[5]}} , in209[5:0] };

   // m209_74 = W*in
   wire signed [9:0] m209_74;
   assign m209_74 =10'b0;

   // m209_75 = W*in
   wire signed [9:0] m209_75;
   assign m209_75 =10'b0;

   // m209_76 = W*in
   wire signed [9:0] m209_76;
   assign m209_76 =10'b0;

   // m209_77 = W*in
   wire signed [9:0] m209_77;
   assign m209_77 =10'b0;

   // m209_78 = W*in
   wire signed [9:0] m209_78;
   assign m209_78 =10'b0;

   // m209_79 = W*in
   wire signed [9:0] m209_79;
   assign m209_79 =10'b0;

   // m209_80 = W*in
   wire signed [9:0] m209_80;
   assign m209_80 =10'b0;

   // m209_81 = W*in
   wire signed [9:0] m209_81;
   assign m209_81 =10'b0;

   // m209_82 = W*in
   wire signed [9:0] m209_82;
   assign m209_82 =10'b0;

   // m209_83 = W*in
   wire signed [9:0] m209_83;
   assign m209_83 =10'b0;

   // m209_84 = W*in
   wire signed [9:0] m209_84;
   assign m209_84 =10'b0;

   // m209_85 = W*in
   wire signed [9:0] m209_85;
   assign m209_85 =10'b0;

   // m209_86 = W*in
   wire signed [9:0] m209_86;
   assign m209_86 =10'b0;

   // m209_87 = W*in
   wire signed [9:0] m209_87;
   assign m209_87 =10'b0;

   // m209_88 = W*in
   wire signed [9:0] m209_88;
   assign m209_88 =10'b0;

   // m209_89 = W*in
   wire signed [9:0] m209_89;
   assign m209_89 =10'b0;

   // m209_90 = W*in
   wire signed [9:0] m209_90;
   assign m209_90 =10'b0;

   // m209_91 = W*in
   wire signed [9:0] m209_91;
   assign m209_91 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_92 = W*in
   wire signed [9:0] m209_92;
   assign m209_92 =10'b0;

   // m209_93 = W*in
   wire signed [9:0] m209_93;
   assign m209_93 =10'b0;

   // m209_94 = W*in
   wire signed [9:0] m209_94;
   assign m209_94 =10'b0;

   // m209_95 = W*in
   wire signed [9:0] m209_95;
   assign m209_95 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_96 = W*in
   wire signed [9:0] m209_96;
   assign m209_96 =10'b0;

   // m209_97 = W*in
   wire signed [9:0] m209_97;
   assign m209_97 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_98 = W*in
   wire signed [9:0] m209_98;
   assign m209_98 =10'b0;

   // m209_99 = W*in
   wire signed [9:0] m209_99;
   assign m209_99 =10'b0;

   // m209_100 = W*in
   wire signed [9:0] m209_100;
   assign m209_100 =10'b0;

   // m209_101 = W*in
   wire signed [9:0] m209_101;
   assign m209_101 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_102 = W*in
   wire signed [9:0] m209_102;
   assign m209_102 =10'b0;

   // m209_103 = W*in
   wire signed [9:0] m209_103;
   assign m209_103 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_104 = W*in
   wire signed [9:0] m209_104;
   assign m209_104 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_105 = W*in
   wire signed [9:0] m209_105;
   assign m209_105 =10'b0;

   // m209_106 = W*in
   wire signed [9:0] m209_106;
   assign m209_106 =10'b0;

   // m209_107 = W*in
   wire signed [9:0] m209_107;
   assign m209_107 =10'b0;

   // m209_108 = W*in
   wire signed [9:0] m209_108;
   assign m209_108 =10'b0;

   // m209_109 = W*in
   wire signed [9:0] m209_109;
   assign m209_109 =10'b0;

   // m209_110 = W*in
   wire signed [9:0] m209_110;
   assign m209_110 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_111 = W*in
   wire signed [9:0] m209_111;
   assign m209_111 =10'b0;

   // m209_112 = W*in
   wire signed [9:0] m209_112;
   assign m209_112 ={ {4{neg209[5]}} , neg209[5:0] };

   // m209_113 = W*in
   wire signed [9:0] m209_113;
   assign m209_113 =10'b0;

   // m209_114 = W*in
   wire signed [9:0] m209_114;
   assign m209_114 =10'b0;

   // m209_115 = W*in
   wire signed [9:0] m209_115;
   assign m209_115 ={ {5{in209[5]}} , in209[5:1] };

   // m209_116 = W*in
   wire signed [9:0] m209_116;
   assign m209_116 =10'b0;

   // m209_117 = W*in
   wire signed [9:0] m209_117;
   assign m209_117 =10'b0;

   // m210_1 = W*in
   wire signed [9:0] m210_1;
   assign m210_1 =10'b0;

   // m210_2 = W*in
   wire signed [9:0] m210_2;
   assign m210_2 ={ {4{in210[5]}} , in210[5:0] };

   // m210_3 = W*in
   wire signed [9:0] m210_3;
   assign m210_3 =10'b0;

   // m210_4 = W*in
   wire signed [9:0] m210_4;
   assign m210_4 =10'b0;

   // m210_5 = W*in
   wire signed [9:0] m210_5;
   assign m210_5 =10'b0;

   // m210_6 = W*in
   wire signed [9:0] m210_6;
   assign m210_6 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_7 = W*in
   wire signed [9:0] m210_7;
   assign m210_7 =10'b0;

   // m210_8 = W*in
   wire signed [9:0] m210_8;
   assign m210_8 ={ {4{in210[5]}} , in210[5:0] };

   // m210_9 = W*in
   wire signed [9:0] m210_9;
   assign m210_9 =10'b0;

   // m210_10 = W*in
   wire signed [9:0] m210_10;
   assign m210_10 =10'b0;

   // m210_11 = W*in
   wire signed [9:0] m210_11;
   assign m210_11 =10'b0;

   // m210_12 = W*in
   wire signed [9:0] m210_12;
   assign m210_12 ={ {5{in210[5]}} , in210[5:1] };

   // m210_13 = W*in
   wire signed [9:0] m210_13;
   assign m210_13 ={ {4{in210[5]}} , in210[5:0] };

   // m210_14 = W*in
   wire signed [9:0] m210_14;
   assign m210_14 =10'b0;

   // m210_15 = W*in
   wire signed [9:0] m210_15;
   assign m210_15 =10'b0;

   // m210_16 = W*in
   wire signed [9:0] m210_16;
   assign m210_16 =10'b0;

   // m210_17 = W*in
   wire signed [9:0] m210_17;
   assign m210_17 ={ {5{in210[5]}} , in210[5:1] };

   // m210_18 = W*in
   wire signed [9:0] m210_18;
   assign m210_18 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_19 = W*in
   wire signed [9:0] m210_19;
   assign m210_19 =10'b0;

   // m210_20 = W*in
   wire signed [9:0] m210_20;
   assign m210_20 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_21 = W*in
   wire signed [9:0] m210_21;
   assign m210_21 =10'b0;

   // m210_22 = W*in
   wire signed [9:0] m210_22;
   assign m210_22 =10'b0;

   // m210_23 = W*in
   wire signed [9:0] m210_23;
   assign m210_23 ={ {5{in210[5]}} , in210[5:1] };

   // m210_24 = W*in
   wire signed [9:0] m210_24;
   assign m210_24 =10'b0;

   // m210_25 = W*in
   wire signed [9:0] m210_25;
   assign m210_25 ={ {5{in210[5]}} , in210[5:1] };

   // m210_26 = W*in
   wire signed [9:0] m210_26;
   assign m210_26 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_27 = W*in
   wire signed [9:0] m210_27;
   assign m210_27 ={ {5{in210[5]}} , in210[5:1] };

   // m210_28 = W*in
   wire signed [9:0] m210_28;
   assign m210_28 ={ {5{in210[5]}} , in210[5:1] };

   // m210_29 = W*in
   wire signed [9:0] m210_29;
   assign m210_29 =10'b0;

   // m210_30 = W*in
   wire signed [9:0] m210_30;
   assign m210_30 =10'b0;

   // m210_31 = W*in
   wire signed [9:0] m210_31;
   assign m210_31 ={ {4{in210[5]}} , in210[5:0] };

   // m210_32 = W*in
   wire signed [9:0] m210_32;
   assign m210_32 =10'b0;

   // m210_33 = W*in
   wire signed [9:0] m210_33;
   assign m210_33 =10'b0;

   // m210_34 = W*in
   wire signed [9:0] m210_34;
   assign m210_34 ={ {5{in210[5]}} , in210[5:1] };

   // m210_35 = W*in
   wire signed [9:0] m210_35;
   assign m210_35 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_36 = W*in
   wire signed [9:0] m210_36;
   assign m210_36 ={ {5{in210[5]}} , in210[5:1] };

   // m210_37 = W*in
   wire signed [9:0] m210_37;
   assign m210_37 ={ {4{in210[5]}} , in210[5:0] };

   // m210_38 = W*in
   wire signed [9:0] m210_38;
   assign m210_38 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_39 = W*in
   wire signed [9:0] m210_39;
   assign m210_39 =10'b0;

   // m210_40 = W*in
   wire signed [9:0] m210_40;
   assign m210_40 =10'b0;

   // m210_41 = W*in
   wire signed [9:0] m210_41;
   assign m210_41 =10'b0;

   // m210_42 = W*in
   wire signed [9:0] m210_42;
   assign m210_42 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_43 = W*in
   wire signed [9:0] m210_43;
   assign m210_43 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_44 = W*in
   wire signed [9:0] m210_44;
   assign m210_44 =10'b0;

   // m210_45 = W*in
   wire signed [9:0] m210_45;
   assign m210_45 =10'b0;

   // m210_46 = W*in
   wire signed [9:0] m210_46;
   assign m210_46 =10'b0;

   // m210_47 = W*in
   wire signed [9:0] m210_47;
   assign m210_47 =10'b0;

   // m210_48 = W*in
   wire signed [9:0] m210_48;
   assign m210_48 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_49 = W*in
   wire signed [9:0] m210_49;
   assign m210_49 =10'b0;

   // m210_50 = W*in
   wire signed [9:0] m210_50;
   assign m210_50 =10'b0;

   // m210_51 = W*in
   wire signed [9:0] m210_51;
   assign m210_51 =10'b0;

   // m210_52 = W*in
   wire signed [9:0] m210_52;
   assign m210_52 ={ {4{in210[5]}} , in210[5:0] };

   // m210_53 = W*in
   wire signed [9:0] m210_53;
   assign m210_53 =10'b0;

   // m210_54 = W*in
   wire signed [9:0] m210_54;
   assign m210_54 =10'b0;

   // m210_55 = W*in
   wire signed [9:0] m210_55;
   assign m210_55 =10'b0;

   // m210_56 = W*in
   wire signed [9:0] m210_56;
   assign m210_56 =10'b0;

   // m210_57 = W*in
   wire signed [9:0] m210_57;
   assign m210_57 =10'b0;

   // m210_58 = W*in
   wire signed [9:0] m210_58;
   assign m210_58 =10'b0;

   // m210_59 = W*in
   wire signed [9:0] m210_59;
   assign m210_59 ={ {4{in210[5]}} , in210[5:0] };

   // m210_60 = W*in
   wire signed [9:0] m210_60;
   assign m210_60 =10'b0;

   // m210_61 = W*in
   wire signed [9:0] m210_61;
   assign m210_61 =10'b0;

   // m210_62 = W*in
   wire signed [9:0] m210_62;
   assign m210_62 =10'b0;

   // m210_63 = W*in
   wire signed [9:0] m210_63;
   assign m210_63 =10'b0;

   // m210_64 = W*in
   wire signed [9:0] m210_64;
   assign m210_64 =10'b0;

   // m210_65 = W*in
   wire signed [9:0] m210_65;
   assign m210_65 =10'b0;

   // m210_66 = W*in
   wire signed [9:0] m210_66;
   assign m210_66 ={ {5{in210[5]}} , in210[5:1] };

   // m210_67 = W*in
   wire signed [9:0] m210_67;
   assign m210_67 ={ {5{in210[5]}} , in210[5:1] };

   // m210_68 = W*in
   wire signed [9:0] m210_68;
   assign m210_68 =10'b0;

   // m210_69 = W*in
   wire signed [9:0] m210_69;
   assign m210_69 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_70 = W*in
   wire signed [9:0] m210_70;
   assign m210_70 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_71 = W*in
   wire signed [9:0] m210_71;
   assign m210_71 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_72 = W*in
   wire signed [9:0] m210_72;
   assign m210_72 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_73 = W*in
   wire signed [9:0] m210_73;
   assign m210_73 ={ {4{in210[5]}} , in210[5:0] };

   // m210_74 = W*in
   wire signed [9:0] m210_74;
   assign m210_74 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_75 = W*in
   wire signed [9:0] m210_75;
   assign m210_75 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_76 = W*in
   wire signed [9:0] m210_76;
   assign m210_76 =10'b0;

   // m210_77 = W*in
   wire signed [9:0] m210_77;
   assign m210_77 =10'b0;

   // m210_78 = W*in
   wire signed [9:0] m210_78;
   assign m210_78 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_79 = W*in
   wire signed [9:0] m210_79;
   assign m210_79 =10'b0;

   // m210_80 = W*in
   wire signed [9:0] m210_80;
   assign m210_80 ={ {4{in210[5]}} , in210[5:0] };

   // m210_81 = W*in
   wire signed [9:0] m210_81;
   assign m210_81 =10'b0;

   // m210_82 = W*in
   wire signed [9:0] m210_82;
   assign m210_82 ={ {4{in210[5]}} , in210[5:0] };

   // m210_83 = W*in
   wire signed [9:0] m210_83;
   assign m210_83 =10'b0;

   // m210_84 = W*in
   wire signed [9:0] m210_84;
   assign m210_84 =10'b0;

   // m210_85 = W*in
   wire signed [9:0] m210_85;
   assign m210_85 ={ {4{in210[5]}} , in210[5:0] };

   // m210_86 = W*in
   wire signed [9:0] m210_86;
   assign m210_86 =10'b0;

   // m210_87 = W*in
   wire signed [9:0] m210_87;
   assign m210_87 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_88 = W*in
   wire signed [9:0] m210_88;
   assign m210_88 =10'b0;

   // m210_89 = W*in
   wire signed [9:0] m210_89;
   assign m210_89 =10'b0;

   // m210_90 = W*in
   wire signed [9:0] m210_90;
   assign m210_90 =10'b0;

   // m210_91 = W*in
   wire signed [9:0] m210_91;
   assign m210_91 =10'b0;

   // m210_92 = W*in
   wire signed [9:0] m210_92;
   assign m210_92 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_93 = W*in
   wire signed [9:0] m210_93;
   assign m210_93 =10'b0;

   // m210_94 = W*in
   wire signed [9:0] m210_94;
   assign m210_94 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_95 = W*in
   wire signed [9:0] m210_95;
   assign m210_95 =10'b0;

   // m210_96 = W*in
   wire signed [9:0] m210_96;
   assign m210_96 =10'b0;

   // m210_97 = W*in
   wire signed [9:0] m210_97;
   assign m210_97 =10'b0;

   // m210_98 = W*in
   wire signed [9:0] m210_98;
   assign m210_98 ={ {4{in210[5]}} , in210[5:0] };

   // m210_99 = W*in
   wire signed [9:0] m210_99;
   assign m210_99 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_100 = W*in
   wire signed [9:0] m210_100;
   assign m210_100 =10'b0;

   // m210_101 = W*in
   wire signed [9:0] m210_101;
   assign m210_101 =10'b0;

   // m210_102 = W*in
   wire signed [9:0] m210_102;
   assign m210_102 =10'b0;

   // m210_103 = W*in
   wire signed [9:0] m210_103;
   assign m210_103 =10'b0;

   // m210_104 = W*in
   wire signed [9:0] m210_104;
   assign m210_104 =10'b0;

   // m210_105 = W*in
   wire signed [9:0] m210_105;
   assign m210_105 =10'b0;

   // m210_106 = W*in
   wire signed [9:0] m210_106;
   assign m210_106 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_107 = W*in
   wire signed [9:0] m210_107;
   assign m210_107 =10'b0;

   // m210_108 = W*in
   wire signed [9:0] m210_108;
   assign m210_108 ={ {5{in210[5]}} , in210[5:1] };

   // m210_109 = W*in
   wire signed [9:0] m210_109;
   assign m210_109 =10'b0;

   // m210_110 = W*in
   wire signed [9:0] m210_110;
   assign m210_110 =10'b0;

   // m210_111 = W*in
   wire signed [9:0] m210_111;
   assign m210_111 ={ {4{neg210[5]}} , neg210[5:0] };

   // m210_112 = W*in
   wire signed [9:0] m210_112;
   assign m210_112 =10'b0;

   // m210_113 = W*in
   wire signed [9:0] m210_113;
   assign m210_113 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_114 = W*in
   wire signed [9:0] m210_114;
   assign m210_114 =10'b0;

   // m210_115 = W*in
   wire signed [9:0] m210_115;
   assign m210_115 ={ {5{neg210[5]}} , neg210[5:1] };

   // m210_116 = W*in
   wire signed [9:0] m210_116;
   assign m210_116 =10'b0;

   // m210_117 = W*in
   wire signed [9:0] m210_117;
   assign m210_117 =10'b0;

   // m211_1 = W*in
   wire signed [9:0] m211_1;
   assign m211_1 ={ {4{in211[5]}} , in211[5:0] };

   // m211_2 = W*in
   wire signed [9:0] m211_2;
   assign m211_2 =10'b0;

   // m211_3 = W*in
   wire signed [9:0] m211_3;
   assign m211_3 =10'b0;

   // m211_4 = W*in
   wire signed [9:0] m211_4;
   assign m211_4 =10'b0;

   // m211_5 = W*in
   wire signed [9:0] m211_5;
   assign m211_5 =10'b0;

   // m211_6 = W*in
   wire signed [9:0] m211_6;
   assign m211_6 =10'b0;

   // m211_7 = W*in
   wire signed [9:0] m211_7;
   assign m211_7 =10'b0;

   // m211_8 = W*in
   wire signed [9:0] m211_8;
   assign m211_8 =10'b0;

   // m211_9 = W*in
   wire signed [9:0] m211_9;
   assign m211_9 =10'b0;

   // m211_10 = W*in
   wire signed [9:0] m211_10;
   assign m211_10 =10'b0;

   // m211_11 = W*in
   wire signed [9:0] m211_11;
   assign m211_11 =10'b0;

   // m211_12 = W*in
   wire signed [9:0] m211_12;
   assign m211_12 =10'b0;

   // m211_13 = W*in
   wire signed [9:0] m211_13;
   assign m211_13 =10'b0;

   // m211_14 = W*in
   wire signed [9:0] m211_14;
   assign m211_14 =10'b0;

   // m211_15 = W*in
   wire signed [9:0] m211_15;
   assign m211_15 =10'b0;

   // m211_16 = W*in
   wire signed [9:0] m211_16;
   assign m211_16 ={ {5{in211[5]}} , in211[5:1] };

   // m211_17 = W*in
   wire signed [9:0] m211_17;
   assign m211_17 =10'b0;

   // m211_18 = W*in
   wire signed [9:0] m211_18;
   assign m211_18 =10'b0;

   // m211_19 = W*in
   wire signed [9:0] m211_19;
   assign m211_19 ={ {5{in211[5]}} , in211[5:1] };

   // m211_20 = W*in
   wire signed [9:0] m211_20;
   assign m211_20 ={ {4{neg211[5]}} , neg211[5:0] };

   // m211_21 = W*in
   wire signed [9:0] m211_21;
   assign m211_21 ={ {5{neg211[5]}} , neg211[5:1] };

   // m211_22 = W*in
   wire signed [9:0] m211_22;
   assign m211_22 =10'b0;

   // m211_23 = W*in
   wire signed [9:0] m211_23;
   assign m211_23 =10'b0;

   // m211_24 = W*in
   wire signed [9:0] m211_24;
   assign m211_24 ={ {4{in211[5]}} , in211[5:0] };

   // m211_25 = W*in
   wire signed [9:0] m211_25;
   assign m211_25 =10'b0;

   // m211_26 = W*in
   wire signed [9:0] m211_26;
   assign m211_26 ={ {4{neg211[5]}} , neg211[5:0] };

   // m211_27 = W*in
   wire signed [9:0] m211_27;
   assign m211_27 ={ {4{in211[5]}} , in211[5:0] };

   // m211_28 = W*in
   wire signed [9:0] m211_28;
   assign m211_28 =10'b0;

   // m211_29 = W*in
   wire signed [9:0] m211_29;
   assign m211_29 =10'b0;

   // m211_30 = W*in
   wire signed [9:0] m211_30;
   assign m211_30 =10'b0;

   // m211_31 = W*in
   wire signed [9:0] m211_31;
   assign m211_31 =10'b0;

   // m211_32 = W*in
   wire signed [9:0] m211_32;
   assign m211_32 =10'b0;

   // m211_33 = W*in
   wire signed [9:0] m211_33;
   assign m211_33 =10'b0;

   // m211_34 = W*in
   wire signed [9:0] m211_34;
   assign m211_34 =10'b0;

   // m211_35 = W*in
   wire signed [9:0] m211_35;
   assign m211_35 =10'b0;

   // m211_36 = W*in
   wire signed [9:0] m211_36;
   assign m211_36 =10'b0;

   // m211_37 = W*in
   wire signed [9:0] m211_37;
   assign m211_37 =10'b0;

   // m211_38 = W*in
   wire signed [9:0] m211_38;
   assign m211_38 =10'b0;

   // m211_39 = W*in
   wire signed [9:0] m211_39;
   assign m211_39 =10'b0;

   // m211_40 = W*in
   wire signed [9:0] m211_40;
   assign m211_40 =10'b0;

   // m211_41 = W*in
   wire signed [9:0] m211_41;
   assign m211_41 =10'b0;

   // m211_42 = W*in
   wire signed [9:0] m211_42;
   assign m211_42 =10'b0;

   // m211_43 = W*in
   wire signed [9:0] m211_43;
   assign m211_43 =10'b0;

   // m211_44 = W*in
   wire signed [9:0] m211_44;
   assign m211_44 =10'b0;

   // m211_45 = W*in
   wire signed [9:0] m211_45;
   assign m211_45 =10'b0;

   // m211_46 = W*in
   wire signed [9:0] m211_46;
   assign m211_46 ={ {4{in211[5]}} , in211[5:0] };

   // m211_47 = W*in
   wire signed [9:0] m211_47;
   assign m211_47 =10'b0;

   // m211_48 = W*in
   wire signed [9:0] m211_48;
   assign m211_48 =10'b0;

   // m211_49 = W*in
   wire signed [9:0] m211_49;
   assign m211_49 =10'b0;

   // m211_50 = W*in
   wire signed [9:0] m211_50;
   assign m211_50 =10'b0;

   // m211_51 = W*in
   wire signed [9:0] m211_51;
   assign m211_51 =10'b0;

   // m211_52 = W*in
   wire signed [9:0] m211_52;
   assign m211_52 =10'b0;

   // m211_53 = W*in
   wire signed [9:0] m211_53;
   assign m211_53 =10'b0;

   // m211_54 = W*in
   wire signed [9:0] m211_54;
   assign m211_54 =10'b0;

   // m211_55 = W*in
   wire signed [9:0] m211_55;
   assign m211_55 =10'b0;

   // m211_56 = W*in
   wire signed [9:0] m211_56;
   assign m211_56 =10'b0;

   // m211_57 = W*in
   wire signed [9:0] m211_57;
   assign m211_57 =10'b0;

   // m211_58 = W*in
   wire signed [9:0] m211_58;
   assign m211_58 =10'b0;

   // m211_59 = W*in
   wire signed [9:0] m211_59;
   assign m211_59 =10'b0;

   // m211_60 = W*in
   wire signed [9:0] m211_60;
   assign m211_60 =10'b0;

   // m211_61 = W*in
   wire signed [9:0] m211_61;
   assign m211_61 ={ {4{in211[5]}} , in211[5:0] };

   // m211_62 = W*in
   wire signed [9:0] m211_62;
   assign m211_62 =10'b0;

   // m211_63 = W*in
   wire signed [9:0] m211_63;
   assign m211_63 =10'b0;

   // m211_64 = W*in
   wire signed [9:0] m211_64;
   assign m211_64 =10'b0;

   // m211_65 = W*in
   wire signed [9:0] m211_65;
   assign m211_65 =10'b0;

   // m211_66 = W*in
   wire signed [9:0] m211_66;
   assign m211_66 =10'b0;

   // m211_67 = W*in
   wire signed [9:0] m211_67;
   assign m211_67 =10'b0;

   // m211_68 = W*in
   wire signed [9:0] m211_68;
   assign m211_68 =10'b0;

   // m211_69 = W*in
   wire signed [9:0] m211_69;
   assign m211_69 ={ {4{in211[5]}} , in211[5:0] };

   // m211_70 = W*in
   wire signed [9:0] m211_70;
   assign m211_70 =10'b0;

   // m211_71 = W*in
   wire signed [9:0] m211_71;
   assign m211_71 =10'b0;

   // m211_72 = W*in
   wire signed [9:0] m211_72;
   assign m211_72 =10'b0;

   // m211_73 = W*in
   wire signed [9:0] m211_73;
   assign m211_73 ={ {4{in211[5]}} , in211[5:0] };

   // m211_74 = W*in
   wire signed [9:0] m211_74;
   assign m211_74 ={ {5{neg211[5]}} , neg211[5:1] };

   // m211_75 = W*in
   wire signed [9:0] m211_75;
   assign m211_75 =10'b0;

   // m211_76 = W*in
   wire signed [9:0] m211_76;
   assign m211_76 =10'b0;

   // m211_77 = W*in
   wire signed [9:0] m211_77;
   assign m211_77 =10'b0;

   // m211_78 = W*in
   wire signed [9:0] m211_78;
   assign m211_78 =10'b0;

   // m211_79 = W*in
   wire signed [9:0] m211_79;
   assign m211_79 =10'b0;

   // m211_80 = W*in
   wire signed [9:0] m211_80;
   assign m211_80 ={ {5{in211[5]}} , in211[5:1] };

   // m211_81 = W*in
   wire signed [9:0] m211_81;
   assign m211_81 =10'b0;

   // m211_82 = W*in
   wire signed [9:0] m211_82;
   assign m211_82 =10'b0;

   // m211_83 = W*in
   wire signed [9:0] m211_83;
   assign m211_83 =10'b0;

   // m211_84 = W*in
   wire signed [9:0] m211_84;
   assign m211_84 =10'b0;

   // m211_85 = W*in
   wire signed [9:0] m211_85;
   assign m211_85 =10'b0;

   // m211_86 = W*in
   wire signed [9:0] m211_86;
   assign m211_86 =10'b0;

   // m211_87 = W*in
   wire signed [9:0] m211_87;
   assign m211_87 =10'b0;

   // m211_88 = W*in
   wire signed [9:0] m211_88;
   assign m211_88 =10'b0;

   // m211_89 = W*in
   wire signed [9:0] m211_89;
   assign m211_89 =10'b0;

   // m211_90 = W*in
   wire signed [9:0] m211_90;
   assign m211_90 =10'b0;

   // m211_91 = W*in
   wire signed [9:0] m211_91;
   assign m211_91 =10'b0;

   // m211_92 = W*in
   wire signed [9:0] m211_92;
   assign m211_92 =10'b0;

   // m211_93 = W*in
   wire signed [9:0] m211_93;
   assign m211_93 =10'b0;

   // m211_94 = W*in
   wire signed [9:0] m211_94;
   assign m211_94 =10'b0;

   // m211_95 = W*in
   wire signed [9:0] m211_95;
   assign m211_95 =10'b0;

   // m211_96 = W*in
   wire signed [9:0] m211_96;
   assign m211_96 =10'b0;

   // m211_97 = W*in
   wire signed [9:0] m211_97;
   assign m211_97 ={ {5{in211[5]}} , in211[5:1] };

   // m211_98 = W*in
   wire signed [9:0] m211_98;
   assign m211_98 =10'b0;

   // m211_99 = W*in
   wire signed [9:0] m211_99;
   assign m211_99 ={ {4{neg211[5]}} , neg211[5:0] };

   // m211_100 = W*in
   wire signed [9:0] m211_100;
   assign m211_100 =10'b0;

   // m211_101 = W*in
   wire signed [9:0] m211_101;
   assign m211_101 =10'b0;

   // m211_102 = W*in
   wire signed [9:0] m211_102;
   assign m211_102 =10'b0;

   // m211_103 = W*in
   wire signed [9:0] m211_103;
   assign m211_103 =10'b0;

   // m211_104 = W*in
   wire signed [9:0] m211_104;
   assign m211_104 =10'b0;

   // m211_105 = W*in
   wire signed [9:0] m211_105;
   assign m211_105 =10'b0;

   // m211_106 = W*in
   wire signed [9:0] m211_106;
   assign m211_106 ={ {5{neg211[5]}} , neg211[5:1] };

   // m211_107 = W*in
   wire signed [9:0] m211_107;
   assign m211_107 ={ {4{in211[5]}} , in211[5:0] };

   // m211_108 = W*in
   wire signed [9:0] m211_108;
   assign m211_108 =10'b0;

   // m211_109 = W*in
   wire signed [9:0] m211_109;
   assign m211_109 =10'b0;

   // m211_110 = W*in
   wire signed [9:0] m211_110;
   assign m211_110 =10'b0;

   // m211_111 = W*in
   wire signed [9:0] m211_111;
   assign m211_111 =10'b0;

   // m211_112 = W*in
   wire signed [9:0] m211_112;
   assign m211_112 =10'b0;

   // m211_113 = W*in
   wire signed [9:0] m211_113;
   assign m211_113 =10'b0;

   // m211_114 = W*in
   wire signed [9:0] m211_114;
   assign m211_114 =10'b0;

   // m211_115 = W*in
   wire signed [9:0] m211_115;
   assign m211_115 =10'b0;

   // m211_116 = W*in
   wire signed [9:0] m211_116;
   assign m211_116 =10'b0;

   // m211_117 = W*in
   wire signed [9:0] m211_117;
   assign m211_117 =10'b0;

   // m212_1 = W*in
   wire signed [9:0] m212_1;
   assign m212_1 =10'b0;

   // m212_2 = W*in
   wire signed [9:0] m212_2;
   assign m212_2 =10'b0;

   // m212_3 = W*in
   wire signed [9:0] m212_3;
   assign m212_3 =10'b0;

   // m212_4 = W*in
   wire signed [9:0] m212_4;
   assign m212_4 =10'b0;

   // m212_5 = W*in
   wire signed [9:0] m212_5;
   assign m212_5 =10'b0;

   // m212_6 = W*in
   wire signed [9:0] m212_6;
   assign m212_6 =10'b0;

   // m212_7 = W*in
   wire signed [9:0] m212_7;
   assign m212_7 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_8 = W*in
   wire signed [9:0] m212_8;
   assign m212_8 =10'b0;

   // m212_9 = W*in
   wire signed [9:0] m212_9;
   assign m212_9 =10'b0;

   // m212_10 = W*in
   wire signed [9:0] m212_10;
   assign m212_10 =10'b0;

   // m212_11 = W*in
   wire signed [9:0] m212_11;
   assign m212_11 ={ {4{in212[5]}} , in212[5:0] };

   // m212_12 = W*in
   wire signed [9:0] m212_12;
   assign m212_12 =10'b0;

   // m212_13 = W*in
   wire signed [9:0] m212_13;
   assign m212_13 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_14 = W*in
   wire signed [9:0] m212_14;
   assign m212_14 =10'b0;

   // m212_15 = W*in
   wire signed [9:0] m212_15;
   assign m212_15 =10'b0;

   // m212_16 = W*in
   wire signed [9:0] m212_16;
   assign m212_16 ={ {5{neg212[5]}} , neg212[5:1] };

   // m212_17 = W*in
   wire signed [9:0] m212_17;
   assign m212_17 =10'b0;

   // m212_18 = W*in
   wire signed [9:0] m212_18;
   assign m212_18 =10'b0;

   // m212_19 = W*in
   wire signed [9:0] m212_19;
   assign m212_19 =10'b0;

   // m212_20 = W*in
   wire signed [9:0] m212_20;
   assign m212_20 =10'b0;

   // m212_21 = W*in
   wire signed [9:0] m212_21;
   assign m212_21 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_22 = W*in
   wire signed [9:0] m212_22;
   assign m212_22 =10'b0;

   // m212_23 = W*in
   wire signed [9:0] m212_23;
   assign m212_23 ={ {5{neg212[5]}} , neg212[5:1] };

   // m212_24 = W*in
   wire signed [9:0] m212_24;
   assign m212_24 =10'b0;

   // m212_25 = W*in
   wire signed [9:0] m212_25;
   assign m212_25 =10'b0;

   // m212_26 = W*in
   wire signed [9:0] m212_26;
   assign m212_26 =10'b0;

   // m212_27 = W*in
   wire signed [9:0] m212_27;
   assign m212_27 ={ {5{in212[5]}} , in212[5:1] };

   // m212_28 = W*in
   wire signed [9:0] m212_28;
   assign m212_28 =10'b0;

   // m212_29 = W*in
   wire signed [9:0] m212_29;
   assign m212_29 =10'b0;

   // m212_30 = W*in
   wire signed [9:0] m212_30;
   assign m212_30 =10'b0;

   // m212_31 = W*in
   wire signed [9:0] m212_31;
   assign m212_31 =10'b0;

   // m212_32 = W*in
   wire signed [9:0] m212_32;
   assign m212_32 =10'b0;

   // m212_33 = W*in
   wire signed [9:0] m212_33;
   assign m212_33 =10'b0;

   // m212_34 = W*in
   wire signed [9:0] m212_34;
   assign m212_34 =10'b0;

   // m212_35 = W*in
   wire signed [9:0] m212_35;
   assign m212_35 =10'b0;

   // m212_36 = W*in
   wire signed [9:0] m212_36;
   assign m212_36 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_37 = W*in
   wire signed [9:0] m212_37;
   assign m212_37 =10'b0;

   // m212_38 = W*in
   wire signed [9:0] m212_38;
   assign m212_38 =10'b0;

   // m212_39 = W*in
   wire signed [9:0] m212_39;
   assign m212_39 =10'b0;

   // m212_40 = W*in
   wire signed [9:0] m212_40;
   assign m212_40 =10'b0;

   // m212_41 = W*in
   wire signed [9:0] m212_41;
   assign m212_41 =10'b0;

   // m212_42 = W*in
   wire signed [9:0] m212_42;
   assign m212_42 =10'b0;

   // m212_43 = W*in
   wire signed [9:0] m212_43;
   assign m212_43 =10'b0;

   // m212_44 = W*in
   wire signed [9:0] m212_44;
   assign m212_44 =10'b0;

   // m212_45 = W*in
   wire signed [9:0] m212_45;
   assign m212_45 =10'b0;

   // m212_46 = W*in
   wire signed [9:0] m212_46;
   assign m212_46 =10'b0;

   // m212_47 = W*in
   wire signed [9:0] m212_47;
   assign m212_47 =10'b0;

   // m212_48 = W*in
   wire signed [9:0] m212_48;
   assign m212_48 =10'b0;

   // m212_49 = W*in
   wire signed [9:0] m212_49;
   assign m212_49 =10'b0;

   // m212_50 = W*in
   wire signed [9:0] m212_50;
   assign m212_50 =10'b0;

   // m212_51 = W*in
   wire signed [9:0] m212_51;
   assign m212_51 =10'b0;

   // m212_52 = W*in
   wire signed [9:0] m212_52;
   assign m212_52 =10'b0;

   // m212_53 = W*in
   wire signed [9:0] m212_53;
   assign m212_53 =10'b0;

   // m212_54 = W*in
   wire signed [9:0] m212_54;
   assign m212_54 =10'b0;

   // m212_55 = W*in
   wire signed [9:0] m212_55;
   assign m212_55 =10'b0;

   // m212_56 = W*in
   wire signed [9:0] m212_56;
   assign m212_56 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_57 = W*in
   wire signed [9:0] m212_57;
   assign m212_57 =10'b0;

   // m212_58 = W*in
   wire signed [9:0] m212_58;
   assign m212_58 =10'b0;

   // m212_59 = W*in
   wire signed [9:0] m212_59;
   assign m212_59 =10'b0;

   // m212_60 = W*in
   wire signed [9:0] m212_60;
   assign m212_60 =10'b0;

   // m212_61 = W*in
   wire signed [9:0] m212_61;
   assign m212_61 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_62 = W*in
   wire signed [9:0] m212_62;
   assign m212_62 =10'b0;

   // m212_63 = W*in
   wire signed [9:0] m212_63;
   assign m212_63 =10'b0;

   // m212_64 = W*in
   wire signed [9:0] m212_64;
   assign m212_64 =10'b0;

   // m212_65 = W*in
   wire signed [9:0] m212_65;
   assign m212_65 =10'b0;

   // m212_66 = W*in
   wire signed [9:0] m212_66;
   assign m212_66 =10'b0;

   // m212_67 = W*in
   wire signed [9:0] m212_67;
   assign m212_67 =10'b0;

   // m212_68 = W*in
   wire signed [9:0] m212_68;
   assign m212_68 =10'b0;

   // m212_69 = W*in
   wire signed [9:0] m212_69;
   assign m212_69 =10'b0;

   // m212_70 = W*in
   wire signed [9:0] m212_70;
   assign m212_70 ={ {5{neg212[5]}} , neg212[5:1] };

   // m212_71 = W*in
   wire signed [9:0] m212_71;
   assign m212_71 =10'b0;

   // m212_72 = W*in
   wire signed [9:0] m212_72;
   assign m212_72 =10'b0;

   // m212_73 = W*in
   wire signed [9:0] m212_73;
   assign m212_73 ={ {5{neg212[5]}} , neg212[5:1] };

   // m212_74 = W*in
   wire signed [9:0] m212_74;
   assign m212_74 =10'b0;

   // m212_75 = W*in
   wire signed [9:0] m212_75;
   assign m212_75 ={ {5{in212[5]}} , in212[5:1] };

   // m212_76 = W*in
   wire signed [9:0] m212_76;
   assign m212_76 =10'b0;

   // m212_77 = W*in
   wire signed [9:0] m212_77;
   assign m212_77 =10'b0;

   // m212_78 = W*in
   wire signed [9:0] m212_78;
   assign m212_78 =10'b0;

   // m212_79 = W*in
   wire signed [9:0] m212_79;
   assign m212_79 =10'b0;

   // m212_80 = W*in
   wire signed [9:0] m212_80;
   assign m212_80 =10'b0;

   // m212_81 = W*in
   wire signed [9:0] m212_81;
   assign m212_81 =10'b0;

   // m212_82 = W*in
   wire signed [9:0] m212_82;
   assign m212_82 =10'b0;

   // m212_83 = W*in
   wire signed [9:0] m212_83;
   assign m212_83 =10'b0;

   // m212_84 = W*in
   wire signed [9:0] m212_84;
   assign m212_84 =10'b0;

   // m212_85 = W*in
   wire signed [9:0] m212_85;
   assign m212_85 ={ {5{neg212[5]}} , neg212[5:1] };

   // m212_86 = W*in
   wire signed [9:0] m212_86;
   assign m212_86 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_87 = W*in
   wire signed [9:0] m212_87;
   assign m212_87 =10'b0;

   // m212_88 = W*in
   wire signed [9:0] m212_88;
   assign m212_88 =10'b0;

   // m212_89 = W*in
   wire signed [9:0] m212_89;
   assign m212_89 =10'b0;

   // m212_90 = W*in
   wire signed [9:0] m212_90;
   assign m212_90 =10'b0;

   // m212_91 = W*in
   wire signed [9:0] m212_91;
   assign m212_91 =10'b0;

   // m212_92 = W*in
   wire signed [9:0] m212_92;
   assign m212_92 =10'b0;

   // m212_93 = W*in
   wire signed [9:0] m212_93;
   assign m212_93 =10'b0;

   // m212_94 = W*in
   wire signed [9:0] m212_94;
   assign m212_94 =10'b0;

   // m212_95 = W*in
   wire signed [9:0] m212_95;
   assign m212_95 =10'b0;

   // m212_96 = W*in
   wire signed [9:0] m212_96;
   assign m212_96 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_97 = W*in
   wire signed [9:0] m212_97;
   assign m212_97 ={ {4{in212[5]}} , in212[5:0] };

   // m212_98 = W*in
   wire signed [9:0] m212_98;
   assign m212_98 =10'b0;

   // m212_99 = W*in
   wire signed [9:0] m212_99;
   assign m212_99 =10'b0;

   // m212_100 = W*in
   wire signed [9:0] m212_100;
   assign m212_100 =10'b0;

   // m212_101 = W*in
   wire signed [9:0] m212_101;
   assign m212_101 =10'b0;

   // m212_102 = W*in
   wire signed [9:0] m212_102;
   assign m212_102 =10'b0;

   // m212_103 = W*in
   wire signed [9:0] m212_103;
   assign m212_103 =10'b0;

   // m212_104 = W*in
   wire signed [9:0] m212_104;
   assign m212_104 =10'b0;

   // m212_105 = W*in
   wire signed [9:0] m212_105;
   assign m212_105 =10'b0;

   // m212_106 = W*in
   wire signed [9:0] m212_106;
   assign m212_106 =10'b0;

   // m212_107 = W*in
   wire signed [9:0] m212_107;
   assign m212_107 =10'b0;

   // m212_108 = W*in
   wire signed [9:0] m212_108;
   assign m212_108 =10'b0;

   // m212_109 = W*in
   wire signed [9:0] m212_109;
   assign m212_109 =10'b0;

   // m212_110 = W*in
   wire signed [9:0] m212_110;
   assign m212_110 =10'b0;

   // m212_111 = W*in
   wire signed [9:0] m212_111;
   assign m212_111 =10'b0;

   // m212_112 = W*in
   wire signed [9:0] m212_112;
   assign m212_112 =10'b0;

   // m212_113 = W*in
   wire signed [9:0] m212_113;
   assign m212_113 =10'b0;

   // m212_114 = W*in
   wire signed [9:0] m212_114;
   assign m212_114 =10'b0;

   // m212_115 = W*in
   wire signed [9:0] m212_115;
   assign m212_115 =10'b0;

   // m212_116 = W*in
   wire signed [9:0] m212_116;
   assign m212_116 ={ {4{neg212[5]}} , neg212[5:0] };

   // m212_117 = W*in
   wire signed [9:0] m212_117;
   assign m212_117 =10'b0;

   // m213_1 = W*in
   wire signed [9:0] m213_1;
   assign m213_1 =10'b0;

   // m213_2 = W*in
   wire signed [9:0] m213_2;
   assign m213_2 =10'b0;

   // m213_3 = W*in
   wire signed [9:0] m213_3;
   assign m213_3 =10'b0;

   // m213_4 = W*in
   wire signed [9:0] m213_4;
   assign m213_4 =10'b0;

   // m213_5 = W*in
   wire signed [9:0] m213_5;
   assign m213_5 =10'b0;

   // m213_6 = W*in
   wire signed [9:0] m213_6;
   assign m213_6 =10'b0;

   // m213_7 = W*in
   wire signed [9:0] m213_7;
   assign m213_7 =10'b0;

   // m213_8 = W*in
   wire signed [9:0] m213_8;
   assign m213_8 =10'b0;

   // m213_9 = W*in
   wire signed [9:0] m213_9;
   assign m213_9 =10'b0;

   // m213_10 = W*in
   wire signed [9:0] m213_10;
   assign m213_10 =10'b0;

   // m213_11 = W*in
   wire signed [9:0] m213_11;
   assign m213_11 =10'b0;

   // m213_12 = W*in
   wire signed [9:0] m213_12;
   assign m213_12 =10'b0;

   // m213_13 = W*in
   wire signed [9:0] m213_13;
   assign m213_13 =10'b0;

   // m213_14 = W*in
   wire signed [9:0] m213_14;
   assign m213_14 =10'b0;

   // m213_15 = W*in
   wire signed [9:0] m213_15;
   assign m213_15 =10'b0;

   // m213_16 = W*in
   wire signed [9:0] m213_16;
   assign m213_16 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_17 = W*in
   wire signed [9:0] m213_17;
   assign m213_17 =10'b0;

   // m213_18 = W*in
   wire signed [9:0] m213_18;
   assign m213_18 ={ {5{in213[5]}} , in213[5:1] };

   // m213_19 = W*in
   wire signed [9:0] m213_19;
   assign m213_19 =10'b0;

   // m213_20 = W*in
   wire signed [9:0] m213_20;
   assign m213_20 =10'b0;

   // m213_21 = W*in
   wire signed [9:0] m213_21;
   assign m213_21 =10'b0;

   // m213_22 = W*in
   wire signed [9:0] m213_22;
   assign m213_22 =10'b0;

   // m213_23 = W*in
   wire signed [9:0] m213_23;
   assign m213_23 ={ {5{in213[5]}} , in213[5:1] };

   // m213_24 = W*in
   wire signed [9:0] m213_24;
   assign m213_24 =10'b0;

   // m213_25 = W*in
   wire signed [9:0] m213_25;
   assign m213_25 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_26 = W*in
   wire signed [9:0] m213_26;
   assign m213_26 ={ {5{in213[5]}} , in213[5:1] };

   // m213_27 = W*in
   wire signed [9:0] m213_27;
   assign m213_27 =10'b0;

   // m213_28 = W*in
   wire signed [9:0] m213_28;
   assign m213_28 ={ {4{neg213[5]}} , neg213[5:0] };

   // m213_29 = W*in
   wire signed [9:0] m213_29;
   assign m213_29 =10'b0;

   // m213_30 = W*in
   wire signed [9:0] m213_30;
   assign m213_30 =10'b0;

   // m213_31 = W*in
   wire signed [9:0] m213_31;
   assign m213_31 =10'b0;

   // m213_32 = W*in
   wire signed [9:0] m213_32;
   assign m213_32 =10'b0;

   // m213_33 = W*in
   wire signed [9:0] m213_33;
   assign m213_33 =10'b0;

   // m213_34 = W*in
   wire signed [9:0] m213_34;
   assign m213_34 ={ {5{in213[5]}} , in213[5:1] };

   // m213_35 = W*in
   wire signed [9:0] m213_35;
   assign m213_35 =10'b0;

   // m213_36 = W*in
   wire signed [9:0] m213_36;
   assign m213_36 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_37 = W*in
   wire signed [9:0] m213_37;
   assign m213_37 =10'b0;

   // m213_38 = W*in
   wire signed [9:0] m213_38;
   assign m213_38 ={ {4{in213[5]}} , in213[5:0] };

   // m213_39 = W*in
   wire signed [9:0] m213_39;
   assign m213_39 =10'b0;

   // m213_40 = W*in
   wire signed [9:0] m213_40;
   assign m213_40 =10'b0;

   // m213_41 = W*in
   wire signed [9:0] m213_41;
   assign m213_41 ={ {4{neg213[5]}} , neg213[5:0] };

   // m213_42 = W*in
   wire signed [9:0] m213_42;
   assign m213_42 =10'b0;

   // m213_43 = W*in
   wire signed [9:0] m213_43;
   assign m213_43 =10'b0;

   // m213_44 = W*in
   wire signed [9:0] m213_44;
   assign m213_44 =10'b0;

   // m213_45 = W*in
   wire signed [9:0] m213_45;
   assign m213_45 =10'b0;

   // m213_46 = W*in
   wire signed [9:0] m213_46;
   assign m213_46 =10'b0;

   // m213_47 = W*in
   wire signed [9:0] m213_47;
   assign m213_47 =10'b0;

   // m213_48 = W*in
   wire signed [9:0] m213_48;
   assign m213_48 =10'b0;

   // m213_49 = W*in
   wire signed [9:0] m213_49;
   assign m213_49 =10'b0;

   // m213_50 = W*in
   wire signed [9:0] m213_50;
   assign m213_50 =10'b0;

   // m213_51 = W*in
   wire signed [9:0] m213_51;
   assign m213_51 =10'b0;

   // m213_52 = W*in
   wire signed [9:0] m213_52;
   assign m213_52 =10'b0;

   // m213_53 = W*in
   wire signed [9:0] m213_53;
   assign m213_53 =10'b0;

   // m213_54 = W*in
   wire signed [9:0] m213_54;
   assign m213_54 =10'b0;

   // m213_55 = W*in
   wire signed [9:0] m213_55;
   assign m213_55 =10'b0;

   // m213_56 = W*in
   wire signed [9:0] m213_56;
   assign m213_56 =10'b0;

   // m213_57 = W*in
   wire signed [9:0] m213_57;
   assign m213_57 =10'b0;

   // m213_58 = W*in
   wire signed [9:0] m213_58;
   assign m213_58 =10'b0;

   // m213_59 = W*in
   wire signed [9:0] m213_59;
   assign m213_59 =10'b0;

   // m213_60 = W*in
   wire signed [9:0] m213_60;
   assign m213_60 =10'b0;

   // m213_61 = W*in
   wire signed [9:0] m213_61;
   assign m213_61 =10'b0;

   // m213_62 = W*in
   wire signed [9:0] m213_62;
   assign m213_62 =10'b0;

   // m213_63 = W*in
   wire signed [9:0] m213_63;
   assign m213_63 =10'b0;

   // m213_64 = W*in
   wire signed [9:0] m213_64;
   assign m213_64 ={ {4{in213[5]}} , in213[5:0] };

   // m213_65 = W*in
   wire signed [9:0] m213_65;
   assign m213_65 =10'b0;

   // m213_66 = W*in
   wire signed [9:0] m213_66;
   assign m213_66 =10'b0;

   // m213_67 = W*in
   wire signed [9:0] m213_67;
   assign m213_67 =10'b0;

   // m213_68 = W*in
   wire signed [9:0] m213_68;
   assign m213_68 =10'b0;

   // m213_69 = W*in
   wire signed [9:0] m213_69;
   assign m213_69 =10'b0;

   // m213_70 = W*in
   wire signed [9:0] m213_70;
   assign m213_70 =10'b0;

   // m213_71 = W*in
   wire signed [9:0] m213_71;
   assign m213_71 =10'b0;

   // m213_72 = W*in
   wire signed [9:0] m213_72;
   assign m213_72 =10'b0;

   // m213_73 = W*in
   wire signed [9:0] m213_73;
   assign m213_73 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_74 = W*in
   wire signed [9:0] m213_74;
   assign m213_74 =10'b0;

   // m213_75 = W*in
   wire signed [9:0] m213_75;
   assign m213_75 =10'b0;

   // m213_76 = W*in
   wire signed [9:0] m213_76;
   assign m213_76 =10'b0;

   // m213_77 = W*in
   wire signed [9:0] m213_77;
   assign m213_77 =10'b0;

   // m213_78 = W*in
   wire signed [9:0] m213_78;
   assign m213_78 =10'b0;

   // m213_79 = W*in
   wire signed [9:0] m213_79;
   assign m213_79 ={ {4{neg213[5]}} , neg213[5:0] };

   // m213_80 = W*in
   wire signed [9:0] m213_80;
   assign m213_80 =10'b0;

   // m213_81 = W*in
   wire signed [9:0] m213_81;
   assign m213_81 =10'b0;

   // m213_82 = W*in
   wire signed [9:0] m213_82;
   assign m213_82 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_83 = W*in
   wire signed [9:0] m213_83;
   assign m213_83 =10'b0;

   // m213_84 = W*in
   wire signed [9:0] m213_84;
   assign m213_84 =10'b0;

   // m213_85 = W*in
   wire signed [9:0] m213_85;
   assign m213_85 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_86 = W*in
   wire signed [9:0] m213_86;
   assign m213_86 =10'b0;

   // m213_87 = W*in
   wire signed [9:0] m213_87;
   assign m213_87 =10'b0;

   // m213_88 = W*in
   wire signed [9:0] m213_88;
   assign m213_88 =10'b0;

   // m213_89 = W*in
   wire signed [9:0] m213_89;
   assign m213_89 =10'b0;

   // m213_90 = W*in
   wire signed [9:0] m213_90;
   assign m213_90 =10'b0;

   // m213_91 = W*in
   wire signed [9:0] m213_91;
   assign m213_91 ={ {4{in213[5]}} , in213[5:0] };

   // m213_92 = W*in
   wire signed [9:0] m213_92;
   assign m213_92 =10'b0;

   // m213_93 = W*in
   wire signed [9:0] m213_93;
   assign m213_93 =10'b0;

   // m213_94 = W*in
   wire signed [9:0] m213_94;
   assign m213_94 =10'b0;

   // m213_95 = W*in
   wire signed [9:0] m213_95;
   assign m213_95 =10'b0;

   // m213_96 = W*in
   wire signed [9:0] m213_96;
   assign m213_96 =10'b0;

   // m213_97 = W*in
   wire signed [9:0] m213_97;
   assign m213_97 ={ {4{in213[5]}} , in213[5:0] };

   // m213_98 = W*in
   wire signed [9:0] m213_98;
   assign m213_98 =10'b0;

   // m213_99 = W*in
   wire signed [9:0] m213_99;
   assign m213_99 =10'b0;

   // m213_100 = W*in
   wire signed [9:0] m213_100;
   assign m213_100 =10'b0;

   // m213_101 = W*in
   wire signed [9:0] m213_101;
   assign m213_101 =10'b0;

   // m213_102 = W*in
   wire signed [9:0] m213_102;
   assign m213_102 =10'b0;

   // m213_103 = W*in
   wire signed [9:0] m213_103;
   assign m213_103 =10'b0;

   // m213_104 = W*in
   wire signed [9:0] m213_104;
   assign m213_104 =10'b0;

   // m213_105 = W*in
   wire signed [9:0] m213_105;
   assign m213_105 =10'b0;

   // m213_106 = W*in
   wire signed [9:0] m213_106;
   assign m213_106 =10'b0;

   // m213_107 = W*in
   wire signed [9:0] m213_107;
   assign m213_107 =10'b0;

   // m213_108 = W*in
   wire signed [9:0] m213_108;
   assign m213_108 ={ {4{neg213[5]}} , neg213[5:0] };

   // m213_109 = W*in
   wire signed [9:0] m213_109;
   assign m213_109 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_110 = W*in
   wire signed [9:0] m213_110;
   assign m213_110 ={ {4{in213[5]}} , in213[5:0] };

   // m213_111 = W*in
   wire signed [9:0] m213_111;
   assign m213_111 =10'b0;

   // m213_112 = W*in
   wire signed [9:0] m213_112;
   assign m213_112 =10'b0;

   // m213_113 = W*in
   wire signed [9:0] m213_113;
   assign m213_113 ={ {5{neg213[5]}} , neg213[5:1] };

   // m213_114 = W*in
   wire signed [9:0] m213_114;
   assign m213_114 ={ {5{in213[5]}} , in213[5:1] };

   // m213_115 = W*in
   wire signed [9:0] m213_115;
   assign m213_115 =10'b0;

   // m213_116 = W*in
   wire signed [9:0] m213_116;
   assign m213_116 ={ {4{neg213[5]}} , neg213[5:0] };

   // m213_117 = W*in
   wire signed [9:0] m213_117;
   assign m213_117 =10'b0;

   // m214_1 = W*in
   wire signed [9:0] m214_1;
   assign m214_1 =10'b0;

   // m214_2 = W*in
   wire signed [9:0] m214_2;
   assign m214_2 =10'b0;

   // m214_3 = W*in
   wire signed [9:0] m214_3;
   assign m214_3 =10'b0;

   // m214_4 = W*in
   wire signed [9:0] m214_4;
   assign m214_4 =10'b0;

   // m214_5 = W*in
   wire signed [9:0] m214_5;
   assign m214_5 =10'b0;

   // m214_6 = W*in
   wire signed [9:0] m214_6;
   assign m214_6 =10'b0;

   // m214_7 = W*in
   wire signed [9:0] m214_7;
   assign m214_7 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_8 = W*in
   wire signed [9:0] m214_8;
   assign m214_8 =10'b0;

   // m214_9 = W*in
   wire signed [9:0] m214_9;
   assign m214_9 =10'b0;

   // m214_10 = W*in
   wire signed [9:0] m214_10;
   assign m214_10 =10'b0;

   // m214_11 = W*in
   wire signed [9:0] m214_11;
   assign m214_11 =10'b0;

   // m214_12 = W*in
   wire signed [9:0] m214_12;
   assign m214_12 =10'b0;

   // m214_13 = W*in
   wire signed [9:0] m214_13;
   assign m214_13 =10'b0;

   // m214_14 = W*in
   wire signed [9:0] m214_14;
   assign m214_14 ={ {4{in214[5]}} , in214[5:0] };

   // m214_15 = W*in
   wire signed [9:0] m214_15;
   assign m214_15 =10'b0;

   // m214_16 = W*in
   wire signed [9:0] m214_16;
   assign m214_16 =10'b0;

   // m214_17 = W*in
   wire signed [9:0] m214_17;
   assign m214_17 =10'b0;

   // m214_18 = W*in
   wire signed [9:0] m214_18;
   assign m214_18 ={ {4{in214[5]}} , in214[5:0] };

   // m214_19 = W*in
   wire signed [9:0] m214_19;
   assign m214_19 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_20 = W*in
   wire signed [9:0] m214_20;
   assign m214_20 ={ {5{neg214[5]}} , neg214[5:1] };

   // m214_21 = W*in
   wire signed [9:0] m214_21;
   assign m214_21 =10'b0;

   // m214_22 = W*in
   wire signed [9:0] m214_22;
   assign m214_22 =10'b0;

   // m214_23 = W*in
   wire signed [9:0] m214_23;
   assign m214_23 =10'b0;

   // m214_24 = W*in
   wire signed [9:0] m214_24;
   assign m214_24 =10'b0;

   // m214_25 = W*in
   wire signed [9:0] m214_25;
   assign m214_25 =10'b0;

   // m214_26 = W*in
   wire signed [9:0] m214_26;
   assign m214_26 ={ {4{in214[5]}} , in214[5:0] };

   // m214_27 = W*in
   wire signed [9:0] m214_27;
   assign m214_27 ={ {5{neg214[5]}} , neg214[5:1] };

   // m214_28 = W*in
   wire signed [9:0] m214_28;
   assign m214_28 =10'b0;

   // m214_29 = W*in
   wire signed [9:0] m214_29;
   assign m214_29 =10'b0;

   // m214_30 = W*in
   wire signed [9:0] m214_30;
   assign m214_30 =10'b0;

   // m214_31 = W*in
   wire signed [9:0] m214_31;
   assign m214_31 =10'b0;

   // m214_32 = W*in
   wire signed [9:0] m214_32;
   assign m214_32 =10'b0;

   // m214_33 = W*in
   wire signed [9:0] m214_33;
   assign m214_33 =10'b0;

   // m214_34 = W*in
   wire signed [9:0] m214_34;
   assign m214_34 =10'b0;

   // m214_35 = W*in
   wire signed [9:0] m214_35;
   assign m214_35 ={ {5{neg214[5]}} , neg214[5:1] };

   // m214_36 = W*in
   wire signed [9:0] m214_36;
   assign m214_36 =10'b0;

   // m214_37 = W*in
   wire signed [9:0] m214_37;
   assign m214_37 =10'b0;

   // m214_38 = W*in
   wire signed [9:0] m214_38;
   assign m214_38 =10'b0;

   // m214_39 = W*in
   wire signed [9:0] m214_39;
   assign m214_39 =10'b0;

   // m214_40 = W*in
   wire signed [9:0] m214_40;
   assign m214_40 =10'b0;

   // m214_41 = W*in
   wire signed [9:0] m214_41;
   assign m214_41 =10'b0;

   // m214_42 = W*in
   wire signed [9:0] m214_42;
   assign m214_42 ={ {4{in214[5]}} , in214[5:0] };

   // m214_43 = W*in
   wire signed [9:0] m214_43;
   assign m214_43 =10'b0;

   // m214_44 = W*in
   wire signed [9:0] m214_44;
   assign m214_44 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_45 = W*in
   wire signed [9:0] m214_45;
   assign m214_45 =10'b0;

   // m214_46 = W*in
   wire signed [9:0] m214_46;
   assign m214_46 =10'b0;

   // m214_47 = W*in
   wire signed [9:0] m214_47;
   assign m214_47 =10'b0;

   // m214_48 = W*in
   wire signed [9:0] m214_48;
   assign m214_48 =10'b0;

   // m214_49 = W*in
   wire signed [9:0] m214_49;
   assign m214_49 ={ {5{neg214[5]}} , neg214[5:1] };

   // m214_50 = W*in
   wire signed [9:0] m214_50;
   assign m214_50 =10'b0;

   // m214_51 = W*in
   wire signed [9:0] m214_51;
   assign m214_51 =10'b0;

   // m214_52 = W*in
   wire signed [9:0] m214_52;
   assign m214_52 =10'b0;

   // m214_53 = W*in
   wire signed [9:0] m214_53;
   assign m214_53 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_54 = W*in
   wire signed [9:0] m214_54;
   assign m214_54 =10'b0;

   // m214_55 = W*in
   wire signed [9:0] m214_55;
   assign m214_55 =10'b0;

   // m214_56 = W*in
   wire signed [9:0] m214_56;
   assign m214_56 =10'b0;

   // m214_57 = W*in
   wire signed [9:0] m214_57;
   assign m214_57 =10'b0;

   // m214_58 = W*in
   wire signed [9:0] m214_58;
   assign m214_58 =10'b0;

   // m214_59 = W*in
   wire signed [9:0] m214_59;
   assign m214_59 =10'b0;

   // m214_60 = W*in
   wire signed [9:0] m214_60;
   assign m214_60 =10'b0;

   // m214_61 = W*in
   wire signed [9:0] m214_61;
   assign m214_61 =10'b0;

   // m214_62 = W*in
   wire signed [9:0] m214_62;
   assign m214_62 =10'b0;

   // m214_63 = W*in
   wire signed [9:0] m214_63;
   assign m214_63 =10'b0;

   // m214_64 = W*in
   wire signed [9:0] m214_64;
   assign m214_64 ={ {4{in214[5]}} , in214[5:0] };

   // m214_65 = W*in
   wire signed [9:0] m214_65;
   assign m214_65 =10'b0;

   // m214_66 = W*in
   wire signed [9:0] m214_66;
   assign m214_66 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_67 = W*in
   wire signed [9:0] m214_67;
   assign m214_67 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_68 = W*in
   wire signed [9:0] m214_68;
   assign m214_68 =10'b0;

   // m214_69 = W*in
   wire signed [9:0] m214_69;
   assign m214_69 =10'b0;

   // m214_70 = W*in
   wire signed [9:0] m214_70;
   assign m214_70 =10'b0;

   // m214_71 = W*in
   wire signed [9:0] m214_71;
   assign m214_71 =10'b0;

   // m214_72 = W*in
   wire signed [9:0] m214_72;
   assign m214_72 =10'b0;

   // m214_73 = W*in
   wire signed [9:0] m214_73;
   assign m214_73 =10'b0;

   // m214_74 = W*in
   wire signed [9:0] m214_74;
   assign m214_74 =10'b0;

   // m214_75 = W*in
   wire signed [9:0] m214_75;
   assign m214_75 =10'b0;

   // m214_76 = W*in
   wire signed [9:0] m214_76;
   assign m214_76 =10'b0;

   // m214_77 = W*in
   wire signed [9:0] m214_77;
   assign m214_77 =10'b0;

   // m214_78 = W*in
   wire signed [9:0] m214_78;
   assign m214_78 =10'b0;

   // m214_79 = W*in
   wire signed [9:0] m214_79;
   assign m214_79 =10'b0;

   // m214_80 = W*in
   wire signed [9:0] m214_80;
   assign m214_80 =10'b0;

   // m214_81 = W*in
   wire signed [9:0] m214_81;
   assign m214_81 =10'b0;

   // m214_82 = W*in
   wire signed [9:0] m214_82;
   assign m214_82 =10'b0;

   // m214_83 = W*in
   wire signed [9:0] m214_83;
   assign m214_83 =10'b0;

   // m214_84 = W*in
   wire signed [9:0] m214_84;
   assign m214_84 =10'b0;

   // m214_85 = W*in
   wire signed [9:0] m214_85;
   assign m214_85 =10'b0;

   // m214_86 = W*in
   wire signed [9:0] m214_86;
   assign m214_86 =10'b0;

   // m214_87 = W*in
   wire signed [9:0] m214_87;
   assign m214_87 =10'b0;

   // m214_88 = W*in
   wire signed [9:0] m214_88;
   assign m214_88 =10'b0;

   // m214_89 = W*in
   wire signed [9:0] m214_89;
   assign m214_89 ={ {4{in214[5]}} , in214[5:0] };

   // m214_90 = W*in
   wire signed [9:0] m214_90;
   assign m214_90 =10'b0;

   // m214_91 = W*in
   wire signed [9:0] m214_91;
   assign m214_91 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_92 = W*in
   wire signed [9:0] m214_92;
   assign m214_92 =10'b0;

   // m214_93 = W*in
   wire signed [9:0] m214_93;
   assign m214_93 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_94 = W*in
   wire signed [9:0] m214_94;
   assign m214_94 ={ {4{in214[5]}} , in214[5:0] };

   // m214_95 = W*in
   wire signed [9:0] m214_95;
   assign m214_95 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_96 = W*in
   wire signed [9:0] m214_96;
   assign m214_96 =10'b0;

   // m214_97 = W*in
   wire signed [9:0] m214_97;
   assign m214_97 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_98 = W*in
   wire signed [9:0] m214_98;
   assign m214_98 ={ {4{neg214[5]}} , neg214[5:0] };

   // m214_99 = W*in
   wire signed [9:0] m214_99;
   assign m214_99 =10'b0;

   // m214_100 = W*in
   wire signed [9:0] m214_100;
   assign m214_100 =10'b0;

   // m214_101 = W*in
   wire signed [9:0] m214_101;
   assign m214_101 =10'b0;

   // m214_102 = W*in
   wire signed [9:0] m214_102;
   assign m214_102 ={ {4{in214[5]}} , in214[5:0] };

   // m214_103 = W*in
   wire signed [9:0] m214_103;
   assign m214_103 =10'b0;

   // m214_104 = W*in
   wire signed [9:0] m214_104;
   assign m214_104 =10'b0;

   // m214_105 = W*in
   wire signed [9:0] m214_105;
   assign m214_105 =10'b0;

   // m214_106 = W*in
   wire signed [9:0] m214_106;
   assign m214_106 =10'b0;

   // m214_107 = W*in
   wire signed [9:0] m214_107;
   assign m214_107 =10'b0;

   // m214_108 = W*in
   wire signed [9:0] m214_108;
   assign m214_108 =10'b0;

   // m214_109 = W*in
   wire signed [9:0] m214_109;
   assign m214_109 =10'b0;

   // m214_110 = W*in
   wire signed [9:0] m214_110;
   assign m214_110 =10'b0;

   // m214_111 = W*in
   wire signed [9:0] m214_111;
   assign m214_111 =10'b0;

   // m214_112 = W*in
   wire signed [9:0] m214_112;
   assign m214_112 =10'b0;

   // m214_113 = W*in
   wire signed [9:0] m214_113;
   assign m214_113 =10'b0;

   // m214_114 = W*in
   wire signed [9:0] m214_114;
   assign m214_114 =10'b0;

   // m214_115 = W*in
   wire signed [9:0] m214_115;
   assign m214_115 ={ {5{neg214[5]}} , neg214[5:1] };

   // m214_116 = W*in
   wire signed [9:0] m214_116;
   assign m214_116 =10'b0;

   // m214_117 = W*in
   wire signed [9:0] m214_117;
   assign m214_117 =10'b0;

   // m215_1 = W*in
   wire signed [9:0] m215_1;
   assign m215_1 =10'b0;

   // m215_2 = W*in
   wire signed [9:0] m215_2;
   assign m215_2 =10'b0;

   // m215_3 = W*in
   wire signed [9:0] m215_3;
   assign m215_3 =10'b0;

   // m215_4 = W*in
   wire signed [9:0] m215_4;
   assign m215_4 =10'b0;

   // m215_5 = W*in
   wire signed [9:0] m215_5;
   assign m215_5 =10'b0;

   // m215_6 = W*in
   wire signed [9:0] m215_6;
   assign m215_6 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_7 = W*in
   wire signed [9:0] m215_7;
   assign m215_7 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_8 = W*in
   wire signed [9:0] m215_8;
   assign m215_8 =10'b0;

   // m215_9 = W*in
   wire signed [9:0] m215_9;
   assign m215_9 =10'b0;

   // m215_10 = W*in
   wire signed [9:0] m215_10;
   assign m215_10 ={ {4{in215[5]}} , in215[5:0] };

   // m215_11 = W*in
   wire signed [9:0] m215_11;
   assign m215_11 =10'b0;

   // m215_12 = W*in
   wire signed [9:0] m215_12;
   assign m215_12 =10'b0;

   // m215_13 = W*in
   wire signed [9:0] m215_13;
   assign m215_13 =10'b0;

   // m215_14 = W*in
   wire signed [9:0] m215_14;
   assign m215_14 ={ {4{in215[5]}} , in215[5:0] };

   // m215_15 = W*in
   wire signed [9:0] m215_15;
   assign m215_15 =10'b0;

   // m215_16 = W*in
   wire signed [9:0] m215_16;
   assign m215_16 =10'b0;

   // m215_17 = W*in
   wire signed [9:0] m215_17;
   assign m215_17 =10'b0;

   // m215_18 = W*in
   wire signed [9:0] m215_18;
   assign m215_18 ={ {3{in215[5]}} , in215 , {1{1'b0}} };

   // m215_19 = W*in
   wire signed [9:0] m215_19;
   assign m215_19 ={ {3{neg215[5]}} , neg215 , {1{1'b0}} };

   // m215_20 = W*in
   wire signed [9:0] m215_20;
   assign m215_20 ={ {3{neg215[5]}} , neg215 , {1{1'b0}} };

   // m215_21 = W*in
   wire signed [9:0] m215_21;
   assign m215_21 =10'b0;

   // m215_22 = W*in
   wire signed [9:0] m215_22;
   assign m215_22 =10'b0;

   // m215_23 = W*in
   wire signed [9:0] m215_23;
   assign m215_23 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_24 = W*in
   wire signed [9:0] m215_24;
   assign m215_24 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_25 = W*in
   wire signed [9:0] m215_25;
   assign m215_25 ={ {5{in215[5]}} , in215[5:1] };

   // m215_26 = W*in
   wire signed [9:0] m215_26;
   assign m215_26 ={ {3{in215[5]}} , in215 , {1{1'b0}} };

   // m215_27 = W*in
   wire signed [9:0] m215_27;
   assign m215_27 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_28 = W*in
   wire signed [9:0] m215_28;
   assign m215_28 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_29 = W*in
   wire signed [9:0] m215_29;
   assign m215_29 =10'b0;

   // m215_30 = W*in
   wire signed [9:0] m215_30;
   assign m215_30 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_31 = W*in
   wire signed [9:0] m215_31;
   assign m215_31 =10'b0;

   // m215_32 = W*in
   wire signed [9:0] m215_32;
   assign m215_32 =10'b0;

   // m215_33 = W*in
   wire signed [9:0] m215_33;
   assign m215_33 ={ {5{in215[5]}} , in215[5:1] };

   // m215_34 = W*in
   wire signed [9:0] m215_34;
   assign m215_34 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_35 = W*in
   wire signed [9:0] m215_35;
   assign m215_35 ={ {3{neg215[5]}} , neg215 , {1{1'b0}} };

   // m215_36 = W*in
   wire signed [9:0] m215_36;
   assign m215_36 =10'b0;

   // m215_37 = W*in
   wire signed [9:0] m215_37;
   assign m215_37 =10'b0;

   // m215_38 = W*in
   wire signed [9:0] m215_38;
   assign m215_38 ={ {4{in215[5]}} , in215[5:0] };

   // m215_39 = W*in
   wire signed [9:0] m215_39;
   assign m215_39 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_40 = W*in
   wire signed [9:0] m215_40;
   assign m215_40 =10'b0;

   // m215_41 = W*in
   wire signed [9:0] m215_41;
   assign m215_41 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_42 = W*in
   wire signed [9:0] m215_42;
   assign m215_42 ={ {4{in215[5]}} , in215[5:0] };

   // m215_43 = W*in
   wire signed [9:0] m215_43;
   assign m215_43 ={ {4{in215[5]}} , in215[5:0] };

   // m215_44 = W*in
   wire signed [9:0] m215_44;
   assign m215_44 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_45 = W*in
   wire signed [9:0] m215_45;
   assign m215_45 =10'b0;

   // m215_46 = W*in
   wire signed [9:0] m215_46;
   assign m215_46 =10'b0;

   // m215_47 = W*in
   wire signed [9:0] m215_47;
   assign m215_47 =10'b0;

   // m215_48 = W*in
   wire signed [9:0] m215_48;
   assign m215_48 =10'b0;

   // m215_49 = W*in
   wire signed [9:0] m215_49;
   assign m215_49 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_50 = W*in
   wire signed [9:0] m215_50;
   assign m215_50 =10'b0;

   // m215_51 = W*in
   wire signed [9:0] m215_51;
   assign m215_51 =10'b0;

   // m215_52 = W*in
   wire signed [9:0] m215_52;
   assign m215_52 =10'b0;

   // m215_53 = W*in
   wire signed [9:0] m215_53;
   assign m215_53 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_54 = W*in
   wire signed [9:0] m215_54;
   assign m215_54 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_55 = W*in
   wire signed [9:0] m215_55;
   assign m215_55 =10'b0;

   // m215_56 = W*in
   wire signed [9:0] m215_56;
   assign m215_56 =10'b0;

   // m215_57 = W*in
   wire signed [9:0] m215_57;
   assign m215_57 =10'b0;

   // m215_58 = W*in
   wire signed [9:0] m215_58;
   assign m215_58 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_59 = W*in
   wire signed [9:0] m215_59;
   assign m215_59 =10'b0;

   // m215_60 = W*in
   wire signed [9:0] m215_60;
   assign m215_60 ={ {3{neg215[5]}} , neg215 , {1{1'b0}} };

   // m215_61 = W*in
   wire signed [9:0] m215_61;
   assign m215_61 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_62 = W*in
   wire signed [9:0] m215_62;
   assign m215_62 =10'b0;

   // m215_63 = W*in
   wire signed [9:0] m215_63;
   assign m215_63 =10'b0;

   // m215_64 = W*in
   wire signed [9:0] m215_64;
   assign m215_64 ={ {4{in215[5]}} , in215[5:0] };

   // m215_65 = W*in
   wire signed [9:0] m215_65;
   assign m215_65 =10'b0;

   // m215_66 = W*in
   wire signed [9:0] m215_66;
   assign m215_66 =10'b0;

   // m215_67 = W*in
   wire signed [9:0] m215_67;
   assign m215_67 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_68 = W*in
   wire signed [9:0] m215_68;
   assign m215_68 =10'b0;

   // m215_69 = W*in
   wire signed [9:0] m215_69;
   assign m215_69 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_70 = W*in
   wire signed [9:0] m215_70;
   assign m215_70 ={ {3{in215[5]}} , in215 , {1{1'b0}} };

   // m215_71 = W*in
   wire signed [9:0] m215_71;
   assign m215_71 ={ {4{in215[5]}} , in215[5:0] };

   // m215_72 = W*in
   wire signed [9:0] m215_72;
   assign m215_72 ={ {3{in215[5]}} , in215 , {1{1'b0}} };

   // m215_73 = W*in
   wire signed [9:0] m215_73;
   assign m215_73 =10'b0;

   // m215_74 = W*in
   wire signed [9:0] m215_74;
   assign m215_74 =10'b0;

   // m215_75 = W*in
   wire signed [9:0] m215_75;
   assign m215_75 =10'b0;

   // m215_76 = W*in
   wire signed [9:0] m215_76;
   assign m215_76 =10'b0;

   // m215_77 = W*in
   wire signed [9:0] m215_77;
   assign m215_77 ={ {4{in215[5]}} , in215[5:0] };

   // m215_78 = W*in
   wire signed [9:0] m215_78;
   assign m215_78 =10'b0;

   // m215_79 = W*in
   wire signed [9:0] m215_79;
   assign m215_79 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_80 = W*in
   wire signed [9:0] m215_80;
   assign m215_80 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_81 = W*in
   wire signed [9:0] m215_81;
   assign m215_81 ={ {4{in215[5]}} , in215[5:0] };

   // m215_82 = W*in
   wire signed [9:0] m215_82;
   assign m215_82 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_83 = W*in
   wire signed [9:0] m215_83;
   assign m215_83 =10'b0;

   // m215_84 = W*in
   wire signed [9:0] m215_84;
   assign m215_84 ={ {3{in215[5]}} , in215 , {1{1'b0}} };

   // m215_85 = W*in
   wire signed [9:0] m215_85;
   assign m215_85 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_86 = W*in
   wire signed [9:0] m215_86;
   assign m215_86 ={ {4{in215[5]}} , in215[5:0] };

   // m215_87 = W*in
   wire signed [9:0] m215_87;
   assign m215_87 ={ {4{in215[5]}} , in215[5:0] };

   // m215_88 = W*in
   wire signed [9:0] m215_88;
   assign m215_88 =10'b0;

   // m215_89 = W*in
   wire signed [9:0] m215_89;
   assign m215_89 =10'b0;

   // m215_90 = W*in
   wire signed [9:0] m215_90;
   assign m215_90 =10'b0;

   // m215_91 = W*in
   wire signed [9:0] m215_91;
   assign m215_91 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_92 = W*in
   wire signed [9:0] m215_92;
   assign m215_92 =10'b0;

   // m215_93 = W*in
   wire signed [9:0] m215_93;
   assign m215_93 ={ {3{neg215[5]}} , neg215 , {1{1'b0}} };

   // m215_94 = W*in
   wire signed [9:0] m215_94;
   assign m215_94 ={ {4{in215[5]}} , in215[5:0] };

   // m215_95 = W*in
   wire signed [9:0] m215_95;
   assign m215_95 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_96 = W*in
   wire signed [9:0] m215_96;
   assign m215_96 ={ {4{in215[5]}} , in215[5:0] };

   // m215_97 = W*in
   wire signed [9:0] m215_97;
   assign m215_97 =10'b0;

   // m215_98 = W*in
   wire signed [9:0] m215_98;
   assign m215_98 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_99 = W*in
   wire signed [9:0] m215_99;
   assign m215_99 ={ {3{in215[5]}} , in215 , {1{1'b0}} };

   // m215_100 = W*in
   wire signed [9:0] m215_100;
   assign m215_100 ={ {4{in215[5]}} , in215[5:0] };

   // m215_101 = W*in
   wire signed [9:0] m215_101;
   assign m215_101 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_102 = W*in
   wire signed [9:0] m215_102;
   assign m215_102 =10'b0;

   // m215_103 = W*in
   wire signed [9:0] m215_103;
   assign m215_103 =10'b0;

   // m215_104 = W*in
   wire signed [9:0] m215_104;
   assign m215_104 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_105 = W*in
   wire signed [9:0] m215_105;
   assign m215_105 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_106 = W*in
   wire signed [9:0] m215_106;
   assign m215_106 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_107 = W*in
   wire signed [9:0] m215_107;
   assign m215_107 =10'b0;

   // m215_108 = W*in
   wire signed [9:0] m215_108;
   assign m215_108 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_109 = W*in
   wire signed [9:0] m215_109;
   assign m215_109 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_110 = W*in
   wire signed [9:0] m215_110;
   assign m215_110 =10'b0;

   // m215_111 = W*in
   wire signed [9:0] m215_111;
   assign m215_111 =10'b0;

   // m215_112 = W*in
   wire signed [9:0] m215_112;
   assign m215_112 ={ {4{in215[5]}} , in215[5:0] };

   // m215_113 = W*in
   wire signed [9:0] m215_113;
   assign m215_113 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_114 = W*in
   wire signed [9:0] m215_114;
   assign m215_114 ={ {5{neg215[5]}} , neg215[5:1] };

   // m215_115 = W*in
   wire signed [9:0] m215_115;
   assign m215_115 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_116 = W*in
   wire signed [9:0] m215_116;
   assign m215_116 ={ {4{neg215[5]}} , neg215[5:0] };

   // m215_117 = W*in
   wire signed [9:0] m215_117;
   assign m215_117 ={ {3{neg215[5]}} , neg215 , {1{1'b0}} };

   // m216_1 = W*in
   wire signed [9:0] m216_1;
   assign m216_1 =10'b0;

   // m216_2 = W*in
   wire signed [9:0] m216_2;
   assign m216_2 =10'b0;

   // m216_3 = W*in
   wire signed [9:0] m216_3;
   assign m216_3 ={ {4{in216[5]}} , in216[5:0] };

   // m216_4 = W*in
   wire signed [9:0] m216_4;
   assign m216_4 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_5 = W*in
   wire signed [9:0] m216_5;
   assign m216_5 =10'b0;

   // m216_6 = W*in
   wire signed [9:0] m216_6;
   assign m216_6 =10'b0;

   // m216_7 = W*in
   wire signed [9:0] m216_7;
   assign m216_7 =10'b0;

   // m216_8 = W*in
   wire signed [9:0] m216_8;
   assign m216_8 =10'b0;

   // m216_9 = W*in
   wire signed [9:0] m216_9;
   assign m216_9 =10'b0;

   // m216_10 = W*in
   wire signed [9:0] m216_10;
   assign m216_10 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_11 = W*in
   wire signed [9:0] m216_11;
   assign m216_11 =10'b0;

   // m216_12 = W*in
   wire signed [9:0] m216_12;
   assign m216_12 ={ {4{in216[5]}} , in216[5:0] };

   // m216_13 = W*in
   wire signed [9:0] m216_13;
   assign m216_13 =10'b0;

   // m216_14 = W*in
   wire signed [9:0] m216_14;
   assign m216_14 ={ {4{in216[5]}} , in216[5:0] };

   // m216_15 = W*in
   wire signed [9:0] m216_15;
   assign m216_15 =10'b0;

   // m216_16 = W*in
   wire signed [9:0] m216_16;
   assign m216_16 =10'b0;

   // m216_17 = W*in
   wire signed [9:0] m216_17;
   assign m216_17 ={ {3{neg216[5]}} , neg216 , {1{1'b0}} };

   // m216_18 = W*in
   wire signed [9:0] m216_18;
   assign m216_18 ={ {3{in216[5]}} , in216 , {1{1'b0}} };

   // m216_19 = W*in
   wire signed [9:0] m216_19;
   assign m216_19 ={ {5{neg216[5]}} , neg216[5:1] };

   // m216_20 = W*in
   wire signed [9:0] m216_20;
   assign m216_20 =10'b0;

   // m216_21 = W*in
   wire signed [9:0] m216_21;
   assign m216_21 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_22 = W*in
   wire signed [9:0] m216_22;
   assign m216_22 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_23 = W*in
   wire signed [9:0] m216_23;
   assign m216_23 =10'b0;

   // m216_24 = W*in
   wire signed [9:0] m216_24;
   assign m216_24 ={ {4{in216[5]}} , in216[5:0] };

   // m216_25 = W*in
   wire signed [9:0] m216_25;
   assign m216_25 ={ {5{neg216[5]}} , neg216[5:1] };

   // m216_26 = W*in
   wire signed [9:0] m216_26;
   assign m216_26 ={ {4{in216[5]}} , in216[5:0] };

   // m216_27 = W*in
   wire signed [9:0] m216_27;
   assign m216_27 ={ {4{in216[5]}} , in216[5:0] };

   // m216_28 = W*in
   wire signed [9:0] m216_28;
   assign m216_28 =10'b0;

   // m216_29 = W*in
   wire signed [9:0] m216_29;
   assign m216_29 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_30 = W*in
   wire signed [9:0] m216_30;
   assign m216_30 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_31 = W*in
   wire signed [9:0] m216_31;
   assign m216_31 =10'b0;

   // m216_32 = W*in
   wire signed [9:0] m216_32;
   assign m216_32 =10'b0;

   // m216_33 = W*in
   wire signed [9:0] m216_33;
   assign m216_33 =10'b0;

   // m216_34 = W*in
   wire signed [9:0] m216_34;
   assign m216_34 ={ {5{in216[5]}} , in216[5:1] };

   // m216_35 = W*in
   wire signed [9:0] m216_35;
   assign m216_35 =10'b0;

   // m216_36 = W*in
   wire signed [9:0] m216_36;
   assign m216_36 =10'b0;

   // m216_37 = W*in
   wire signed [9:0] m216_37;
   assign m216_37 =10'b0;

   // m216_38 = W*in
   wire signed [9:0] m216_38;
   assign m216_38 ={ {4{in216[5]}} , in216[5:0] };

   // m216_39 = W*in
   wire signed [9:0] m216_39;
   assign m216_39 =10'b0;

   // m216_40 = W*in
   wire signed [9:0] m216_40;
   assign m216_40 =10'b0;

   // m216_41 = W*in
   wire signed [9:0] m216_41;
   assign m216_41 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_42 = W*in
   wire signed [9:0] m216_42;
   assign m216_42 ={ {4{in216[5]}} , in216[5:0] };

   // m216_43 = W*in
   wire signed [9:0] m216_43;
   assign m216_43 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_44 = W*in
   wire signed [9:0] m216_44;
   assign m216_44 =10'b0;

   // m216_45 = W*in
   wire signed [9:0] m216_45;
   assign m216_45 =10'b0;

   // m216_46 = W*in
   wire signed [9:0] m216_46;
   assign m216_46 =10'b0;

   // m216_47 = W*in
   wire signed [9:0] m216_47;
   assign m216_47 =10'b0;

   // m216_48 = W*in
   wire signed [9:0] m216_48;
   assign m216_48 =10'b0;

   // m216_49 = W*in
   wire signed [9:0] m216_49;
   assign m216_49 =10'b0;

   // m216_50 = W*in
   wire signed [9:0] m216_50;
   assign m216_50 =10'b0;

   // m216_51 = W*in
   wire signed [9:0] m216_51;
   assign m216_51 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_52 = W*in
   wire signed [9:0] m216_52;
   assign m216_52 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_53 = W*in
   wire signed [9:0] m216_53;
   assign m216_53 =10'b0;

   // m216_54 = W*in
   wire signed [9:0] m216_54;
   assign m216_54 =10'b0;

   // m216_55 = W*in
   wire signed [9:0] m216_55;
   assign m216_55 =10'b0;

   // m216_56 = W*in
   wire signed [9:0] m216_56;
   assign m216_56 =10'b0;

   // m216_57 = W*in
   wire signed [9:0] m216_57;
   assign m216_57 =10'b0;

   // m216_58 = W*in
   wire signed [9:0] m216_58;
   assign m216_58 ={ {5{in216[5]}} , in216[5:1] };

   // m216_59 = W*in
   wire signed [9:0] m216_59;
   assign m216_59 =10'b0;

   // m216_60 = W*in
   wire signed [9:0] m216_60;
   assign m216_60 =10'b0;

   // m216_61 = W*in
   wire signed [9:0] m216_61;
   assign m216_61 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_62 = W*in
   wire signed [9:0] m216_62;
   assign m216_62 =10'b0;

   // m216_63 = W*in
   wire signed [9:0] m216_63;
   assign m216_63 =10'b0;

   // m216_64 = W*in
   wire signed [9:0] m216_64;
   assign m216_64 ={ {4{in216[5]}} , in216[5:0] };

   // m216_65 = W*in
   wire signed [9:0] m216_65;
   assign m216_65 =10'b0;

   // m216_66 = W*in
   wire signed [9:0] m216_66;
   assign m216_66 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_67 = W*in
   wire signed [9:0] m216_67;
   assign m216_67 =10'b0;

   // m216_68 = W*in
   wire signed [9:0] m216_68;
   assign m216_68 =10'b0;

   // m216_69 = W*in
   wire signed [9:0] m216_69;
   assign m216_69 =10'b0;

   // m216_70 = W*in
   wire signed [9:0] m216_70;
   assign m216_70 ={ {4{in216[5]}} , in216[5:0] };

   // m216_71 = W*in
   wire signed [9:0] m216_71;
   assign m216_71 ={ {5{in216[5]}} , in216[5:1] };

   // m216_72 = W*in
   wire signed [9:0] m216_72;
   assign m216_72 =10'b0;

   // m216_73 = W*in
   wire signed [9:0] m216_73;
   assign m216_73 ={ {4{in216[5]}} , in216[5:0] };

   // m216_74 = W*in
   wire signed [9:0] m216_74;
   assign m216_74 =10'b0;

   // m216_75 = W*in
   wire signed [9:0] m216_75;
   assign m216_75 =10'b0;

   // m216_76 = W*in
   wire signed [9:0] m216_76;
   assign m216_76 =10'b0;

   // m216_77 = W*in
   wire signed [9:0] m216_77;
   assign m216_77 ={ {4{in216[5]}} , in216[5:0] };

   // m216_78 = W*in
   wire signed [9:0] m216_78;
   assign m216_78 ={ {5{neg216[5]}} , neg216[5:1] };

   // m216_79 = W*in
   wire signed [9:0] m216_79;
   assign m216_79 ={ {3{neg216[5]}} , neg216 , {1{1'b0}} };

   // m216_80 = W*in
   wire signed [9:0] m216_80;
   assign m216_80 ={ {4{in216[5]}} , in216[5:0] };

   // m216_81 = W*in
   wire signed [9:0] m216_81;
   assign m216_81 ={ {4{in216[5]}} , in216[5:0] };

   // m216_82 = W*in
   wire signed [9:0] m216_82;
   assign m216_82 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_83 = W*in
   wire signed [9:0] m216_83;
   assign m216_83 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_84 = W*in
   wire signed [9:0] m216_84;
   assign m216_84 ={ {4{in216[5]}} , in216[5:0] };

   // m216_85 = W*in
   wire signed [9:0] m216_85;
   assign m216_85 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_86 = W*in
   wire signed [9:0] m216_86;
   assign m216_86 ={ {4{in216[5]}} , in216[5:0] };

   // m216_87 = W*in
   wire signed [9:0] m216_87;
   assign m216_87 =10'b0;

   // m216_88 = W*in
   wire signed [9:0] m216_88;
   assign m216_88 ={ {4{in216[5]}} , in216[5:0] };

   // m216_89 = W*in
   wire signed [9:0] m216_89;
   assign m216_89 =10'b0;

   // m216_90 = W*in
   wire signed [9:0] m216_90;
   assign m216_90 =10'b0;

   // m216_91 = W*in
   wire signed [9:0] m216_91;
   assign m216_91 =10'b0;

   // m216_92 = W*in
   wire signed [9:0] m216_92;
   assign m216_92 =10'b0;

   // m216_93 = W*in
   wire signed [9:0] m216_93;
   assign m216_93 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_94 = W*in
   wire signed [9:0] m216_94;
   assign m216_94 =10'b0;

   // m216_95 = W*in
   wire signed [9:0] m216_95;
   assign m216_95 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_96 = W*in
   wire signed [9:0] m216_96;
   assign m216_96 =10'b0;

   // m216_97 = W*in
   wire signed [9:0] m216_97;
   assign m216_97 =10'b0;

   // m216_98 = W*in
   wire signed [9:0] m216_98;
   assign m216_98 =10'b0;

   // m216_99 = W*in
   wire signed [9:0] m216_99;
   assign m216_99 =10'b0;

   // m216_100 = W*in
   wire signed [9:0] m216_100;
   assign m216_100 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_101 = W*in
   wire signed [9:0] m216_101;
   assign m216_101 =10'b0;

   // m216_102 = W*in
   wire signed [9:0] m216_102;
   assign m216_102 =10'b0;

   // m216_103 = W*in
   wire signed [9:0] m216_103;
   assign m216_103 =10'b0;

   // m216_104 = W*in
   wire signed [9:0] m216_104;
   assign m216_104 =10'b0;

   // m216_105 = W*in
   wire signed [9:0] m216_105;
   assign m216_105 ={ {4{in216[5]}} , in216[5:0] };

   // m216_106 = W*in
   wire signed [9:0] m216_106;
   assign m216_106 ={ {5{neg216[5]}} , neg216[5:1] };

   // m216_107 = W*in
   wire signed [9:0] m216_107;
   assign m216_107 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_108 = W*in
   wire signed [9:0] m216_108;
   assign m216_108 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_109 = W*in
   wire signed [9:0] m216_109;
   assign m216_109 =10'b0;

   // m216_110 = W*in
   wire signed [9:0] m216_110;
   assign m216_110 ={ {4{in216[5]}} , in216[5:0] };

   // m216_111 = W*in
   wire signed [9:0] m216_111;
   assign m216_111 =10'b0;

   // m216_112 = W*in
   wire signed [9:0] m216_112;
   assign m216_112 =10'b0;

   // m216_113 = W*in
   wire signed [9:0] m216_113;
   assign m216_113 =10'b0;

   // m216_114 = W*in
   wire signed [9:0] m216_114;
   assign m216_114 =10'b0;

   // m216_115 = W*in
   wire signed [9:0] m216_115;
   assign m216_115 ={ {5{neg216[5]}} , neg216[5:1] };

   // m216_116 = W*in
   wire signed [9:0] m216_116;
   assign m216_116 ={ {4{neg216[5]}} , neg216[5:0] };

   // m216_117 = W*in
   wire signed [9:0] m216_117;
   assign m216_117 =10'b0;

   // m217_1 = W*in
   wire signed [9:0] m217_1;
   assign m217_1 =10'b0;

   // m217_2 = W*in
   wire signed [9:0] m217_2;
   assign m217_2 =10'b0;

   // m217_3 = W*in
   wire signed [9:0] m217_3;
   assign m217_3 =10'b0;

   // m217_4 = W*in
   wire signed [9:0] m217_4;
   assign m217_4 =10'b0;

   // m217_5 = W*in
   wire signed [9:0] m217_5;
   assign m217_5 =10'b0;

   // m217_6 = W*in
   wire signed [9:0] m217_6;
   assign m217_6 =10'b0;

   // m217_7 = W*in
   wire signed [9:0] m217_7;
   assign m217_7 =10'b0;

   // m217_8 = W*in
   wire signed [9:0] m217_8;
   assign m217_8 =10'b0;

   // m217_9 = W*in
   wire signed [9:0] m217_9;
   assign m217_9 =10'b0;

   // m217_10 = W*in
   wire signed [9:0] m217_10;
   assign m217_10 =10'b0;

   // m217_11 = W*in
   wire signed [9:0] m217_11;
   assign m217_11 =10'b0;

   // m217_12 = W*in
   wire signed [9:0] m217_12;
   assign m217_12 =10'b0;

   // m217_13 = W*in
   wire signed [9:0] m217_13;
   assign m217_13 =10'b0;

   // m217_14 = W*in
   wire signed [9:0] m217_14;
   assign m217_14 =10'b0;

   // m217_15 = W*in
   wire signed [9:0] m217_15;
   assign m217_15 =10'b0;

   // m217_16 = W*in
   wire signed [9:0] m217_16;
   assign m217_16 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_17 = W*in
   wire signed [9:0] m217_17;
   assign m217_17 =10'b0;

   // m217_18 = W*in
   wire signed [9:0] m217_18;
   assign m217_18 =10'b0;

   // m217_19 = W*in
   wire signed [9:0] m217_19;
   assign m217_19 =10'b0;

   // m217_20 = W*in
   wire signed [9:0] m217_20;
   assign m217_20 =10'b0;

   // m217_21 = W*in
   wire signed [9:0] m217_21;
   assign m217_21 =10'b0;

   // m217_22 = W*in
   wire signed [9:0] m217_22;
   assign m217_22 ={ {4{in217[5]}} , in217[5:0] };

   // m217_23 = W*in
   wire signed [9:0] m217_23;
   assign m217_23 ={ {4{in217[5]}} , in217[5:0] };

   // m217_24 = W*in
   wire signed [9:0] m217_24;
   assign m217_24 =10'b0;

   // m217_25 = W*in
   wire signed [9:0] m217_25;
   assign m217_25 =10'b0;

   // m217_26 = W*in
   wire signed [9:0] m217_26;
   assign m217_26 =10'b0;

   // m217_27 = W*in
   wire signed [9:0] m217_27;
   assign m217_27 =10'b0;

   // m217_28 = W*in
   wire signed [9:0] m217_28;
   assign m217_28 =10'b0;

   // m217_29 = W*in
   wire signed [9:0] m217_29;
   assign m217_29 =10'b0;

   // m217_30 = W*in
   wire signed [9:0] m217_30;
   assign m217_30 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_31 = W*in
   wire signed [9:0] m217_31;
   assign m217_31 =10'b0;

   // m217_32 = W*in
   wire signed [9:0] m217_32;
   assign m217_32 =10'b0;

   // m217_33 = W*in
   wire signed [9:0] m217_33;
   assign m217_33 =10'b0;

   // m217_34 = W*in
   wire signed [9:0] m217_34;
   assign m217_34 ={ {5{in217[5]}} , in217[5:1] };

   // m217_35 = W*in
   wire signed [9:0] m217_35;
   assign m217_35 =10'b0;

   // m217_36 = W*in
   wire signed [9:0] m217_36;
   assign m217_36 ={ {5{neg217[5]}} , neg217[5:1] };

   // m217_37 = W*in
   wire signed [9:0] m217_37;
   assign m217_37 =10'b0;

   // m217_38 = W*in
   wire signed [9:0] m217_38;
   assign m217_38 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_39 = W*in
   wire signed [9:0] m217_39;
   assign m217_39 =10'b0;

   // m217_40 = W*in
   wire signed [9:0] m217_40;
   assign m217_40 =10'b0;

   // m217_41 = W*in
   wire signed [9:0] m217_41;
   assign m217_41 =10'b0;

   // m217_42 = W*in
   wire signed [9:0] m217_42;
   assign m217_42 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_43 = W*in
   wire signed [9:0] m217_43;
   assign m217_43 =10'b0;

   // m217_44 = W*in
   wire signed [9:0] m217_44;
   assign m217_44 =10'b0;

   // m217_45 = W*in
   wire signed [9:0] m217_45;
   assign m217_45 =10'b0;

   // m217_46 = W*in
   wire signed [9:0] m217_46;
   assign m217_46 =10'b0;

   // m217_47 = W*in
   wire signed [9:0] m217_47;
   assign m217_47 =10'b0;

   // m217_48 = W*in
   wire signed [9:0] m217_48;
   assign m217_48 =10'b0;

   // m217_49 = W*in
   wire signed [9:0] m217_49;
   assign m217_49 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_50 = W*in
   wire signed [9:0] m217_50;
   assign m217_50 =10'b0;

   // m217_51 = W*in
   wire signed [9:0] m217_51;
   assign m217_51 =10'b0;

   // m217_52 = W*in
   wire signed [9:0] m217_52;
   assign m217_52 =10'b0;

   // m217_53 = W*in
   wire signed [9:0] m217_53;
   assign m217_53 =10'b0;

   // m217_54 = W*in
   wire signed [9:0] m217_54;
   assign m217_54 =10'b0;

   // m217_55 = W*in
   wire signed [9:0] m217_55;
   assign m217_55 =10'b0;

   // m217_56 = W*in
   wire signed [9:0] m217_56;
   assign m217_56 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_57 = W*in
   wire signed [9:0] m217_57;
   assign m217_57 =10'b0;

   // m217_58 = W*in
   wire signed [9:0] m217_58;
   assign m217_58 ={ {5{in217[5]}} , in217[5:1] };

   // m217_59 = W*in
   wire signed [9:0] m217_59;
   assign m217_59 =10'b0;

   // m217_60 = W*in
   wire signed [9:0] m217_60;
   assign m217_60 =10'b0;

   // m217_61 = W*in
   wire signed [9:0] m217_61;
   assign m217_61 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_62 = W*in
   wire signed [9:0] m217_62;
   assign m217_62 =10'b0;

   // m217_63 = W*in
   wire signed [9:0] m217_63;
   assign m217_63 =10'b0;

   // m217_64 = W*in
   wire signed [9:0] m217_64;
   assign m217_64 =10'b0;

   // m217_65 = W*in
   wire signed [9:0] m217_65;
   assign m217_65 =10'b0;

   // m217_66 = W*in
   wire signed [9:0] m217_66;
   assign m217_66 =10'b0;

   // m217_67 = W*in
   wire signed [9:0] m217_67;
   assign m217_67 =10'b0;

   // m217_68 = W*in
   wire signed [9:0] m217_68;
   assign m217_68 =10'b0;

   // m217_69 = W*in
   wire signed [9:0] m217_69;
   assign m217_69 =10'b0;

   // m217_70 = W*in
   wire signed [9:0] m217_70;
   assign m217_70 =10'b0;

   // m217_71 = W*in
   wire signed [9:0] m217_71;
   assign m217_71 ={ {5{neg217[5]}} , neg217[5:1] };

   // m217_72 = W*in
   wire signed [9:0] m217_72;
   assign m217_72 =10'b0;

   // m217_73 = W*in
   wire signed [9:0] m217_73;
   assign m217_73 =10'b0;

   // m217_74 = W*in
   wire signed [9:0] m217_74;
   assign m217_74 =10'b0;

   // m217_75 = W*in
   wire signed [9:0] m217_75;
   assign m217_75 =10'b0;

   // m217_76 = W*in
   wire signed [9:0] m217_76;
   assign m217_76 ={ {4{in217[5]}} , in217[5:0] };

   // m217_77 = W*in
   wire signed [9:0] m217_77;
   assign m217_77 =10'b0;

   // m217_78 = W*in
   wire signed [9:0] m217_78;
   assign m217_78 =10'b0;

   // m217_79 = W*in
   wire signed [9:0] m217_79;
   assign m217_79 =10'b0;

   // m217_80 = W*in
   wire signed [9:0] m217_80;
   assign m217_80 =10'b0;

   // m217_81 = W*in
   wire signed [9:0] m217_81;
   assign m217_81 =10'b0;

   // m217_82 = W*in
   wire signed [9:0] m217_82;
   assign m217_82 =10'b0;

   // m217_83 = W*in
   wire signed [9:0] m217_83;
   assign m217_83 =10'b0;

   // m217_84 = W*in
   wire signed [9:0] m217_84;
   assign m217_84 =10'b0;

   // m217_85 = W*in
   wire signed [9:0] m217_85;
   assign m217_85 =10'b0;

   // m217_86 = W*in
   wire signed [9:0] m217_86;
   assign m217_86 =10'b0;

   // m217_87 = W*in
   wire signed [9:0] m217_87;
   assign m217_87 =10'b0;

   // m217_88 = W*in
   wire signed [9:0] m217_88;
   assign m217_88 =10'b0;

   // m217_89 = W*in
   wire signed [9:0] m217_89;
   assign m217_89 ={ {4{in217[5]}} , in217[5:0] };

   // m217_90 = W*in
   wire signed [9:0] m217_90;
   assign m217_90 =10'b0;

   // m217_91 = W*in
   wire signed [9:0] m217_91;
   assign m217_91 =10'b0;

   // m217_92 = W*in
   wire signed [9:0] m217_92;
   assign m217_92 =10'b0;

   // m217_93 = W*in
   wire signed [9:0] m217_93;
   assign m217_93 ={ {4{in217[5]}} , in217[5:0] };

   // m217_94 = W*in
   wire signed [9:0] m217_94;
   assign m217_94 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_95 = W*in
   wire signed [9:0] m217_95;
   assign m217_95 ={ {4{in217[5]}} , in217[5:0] };

   // m217_96 = W*in
   wire signed [9:0] m217_96;
   assign m217_96 ={ {4{in217[5]}} , in217[5:0] };

   // m217_97 = W*in
   wire signed [9:0] m217_97;
   assign m217_97 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_98 = W*in
   wire signed [9:0] m217_98;
   assign m217_98 ={ {4{in217[5]}} , in217[5:0] };

   // m217_99 = W*in
   wire signed [9:0] m217_99;
   assign m217_99 ={ {4{in217[5]}} , in217[5:0] };

   // m217_100 = W*in
   wire signed [9:0] m217_100;
   assign m217_100 =10'b0;

   // m217_101 = W*in
   wire signed [9:0] m217_101;
   assign m217_101 =10'b0;

   // m217_102 = W*in
   wire signed [9:0] m217_102;
   assign m217_102 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_103 = W*in
   wire signed [9:0] m217_103;
   assign m217_103 =10'b0;

   // m217_104 = W*in
   wire signed [9:0] m217_104;
   assign m217_104 =10'b0;

   // m217_105 = W*in
   wire signed [9:0] m217_105;
   assign m217_105 =10'b0;

   // m217_106 = W*in
   wire signed [9:0] m217_106;
   assign m217_106 ={ {4{neg217[5]}} , neg217[5:0] };

   // m217_107 = W*in
   wire signed [9:0] m217_107;
   assign m217_107 =10'b0;

   // m217_108 = W*in
   wire signed [9:0] m217_108;
   assign m217_108 ={ {4{in217[5]}} , in217[5:0] };

   // m217_109 = W*in
   wire signed [9:0] m217_109;
   assign m217_109 ={ {4{in217[5]}} , in217[5:0] };

   // m217_110 = W*in
   wire signed [9:0] m217_110;
   assign m217_110 =10'b0;

   // m217_111 = W*in
   wire signed [9:0] m217_111;
   assign m217_111 =10'b0;

   // m217_112 = W*in
   wire signed [9:0] m217_112;
   assign m217_112 =10'b0;

   // m217_113 = W*in
   wire signed [9:0] m217_113;
   assign m217_113 =10'b0;

   // m217_114 = W*in
   wire signed [9:0] m217_114;
   assign m217_114 ={ {5{in217[5]}} , in217[5:1] };

   // m217_115 = W*in
   wire signed [9:0] m217_115;
   assign m217_115 ={ {5{in217[5]}} , in217[5:1] };

   // m217_116 = W*in
   wire signed [9:0] m217_116;
   assign m217_116 =10'b0;

   // m217_117 = W*in
   wire signed [9:0] m217_117;
   assign m217_117 =10'b0;

   // m218_1 = W*in
   wire signed [9:0] m218_1;
   assign m218_1 =10'b0;

   // m218_2 = W*in
   wire signed [9:0] m218_2;
   assign m218_2 =10'b0;

   // m218_3 = W*in
   wire signed [9:0] m218_3;
   assign m218_3 =10'b0;

   // m218_4 = W*in
   wire signed [9:0] m218_4;
   assign m218_4 =10'b0;

   // m218_5 = W*in
   wire signed [9:0] m218_5;
   assign m218_5 =10'b0;

   // m218_6 = W*in
   wire signed [9:0] m218_6;
   assign m218_6 =10'b0;

   // m218_7 = W*in
   wire signed [9:0] m218_7;
   assign m218_7 =10'b0;

   // m218_8 = W*in
   wire signed [9:0] m218_8;
   assign m218_8 =10'b0;

   // m218_9 = W*in
   wire signed [9:0] m218_9;
   assign m218_9 =10'b0;

   // m218_10 = W*in
   wire signed [9:0] m218_10;
   assign m218_10 =10'b0;

   // m218_11 = W*in
   wire signed [9:0] m218_11;
   assign m218_11 =10'b0;

   // m218_12 = W*in
   wire signed [9:0] m218_12;
   assign m218_12 =10'b0;

   // m218_13 = W*in
   wire signed [9:0] m218_13;
   assign m218_13 =10'b0;

   // m218_14 = W*in
   wire signed [9:0] m218_14;
   assign m218_14 =10'b0;

   // m218_15 = W*in
   wire signed [9:0] m218_15;
   assign m218_15 =10'b0;

   // m218_16 = W*in
   wire signed [9:0] m218_16;
   assign m218_16 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_17 = W*in
   wire signed [9:0] m218_17;
   assign m218_17 =10'b0;

   // m218_18 = W*in
   wire signed [9:0] m218_18;
   assign m218_18 =10'b0;

   // m218_19 = W*in
   wire signed [9:0] m218_19;
   assign m218_19 =10'b0;

   // m218_20 = W*in
   wire signed [9:0] m218_20;
   assign m218_20 =10'b0;

   // m218_21 = W*in
   wire signed [9:0] m218_21;
   assign m218_21 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_22 = W*in
   wire signed [9:0] m218_22;
   assign m218_22 =10'b0;

   // m218_23 = W*in
   wire signed [9:0] m218_23;
   assign m218_23 ={ {4{in218[5]}} , in218[5:0] };

   // m218_24 = W*in
   wire signed [9:0] m218_24;
   assign m218_24 =10'b0;

   // m218_25 = W*in
   wire signed [9:0] m218_25;
   assign m218_25 =10'b0;

   // m218_26 = W*in
   wire signed [9:0] m218_26;
   assign m218_26 =10'b0;

   // m218_27 = W*in
   wire signed [9:0] m218_27;
   assign m218_27 ={ {4{in218[5]}} , in218[5:0] };

   // m218_28 = W*in
   wire signed [9:0] m218_28;
   assign m218_28 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_29 = W*in
   wire signed [9:0] m218_29;
   assign m218_29 =10'b0;

   // m218_30 = W*in
   wire signed [9:0] m218_30;
   assign m218_30 =10'b0;

   // m218_31 = W*in
   wire signed [9:0] m218_31;
   assign m218_31 =10'b0;

   // m218_32 = W*in
   wire signed [9:0] m218_32;
   assign m218_32 =10'b0;

   // m218_33 = W*in
   wire signed [9:0] m218_33;
   assign m218_33 =10'b0;

   // m218_34 = W*in
   wire signed [9:0] m218_34;
   assign m218_34 ={ {4{in218[5]}} , in218[5:0] };

   // m218_35 = W*in
   wire signed [9:0] m218_35;
   assign m218_35 =10'b0;

   // m218_36 = W*in
   wire signed [9:0] m218_36;
   assign m218_36 =10'b0;

   // m218_37 = W*in
   wire signed [9:0] m218_37;
   assign m218_37 =10'b0;

   // m218_38 = W*in
   wire signed [9:0] m218_38;
   assign m218_38 =10'b0;

   // m218_39 = W*in
   wire signed [9:0] m218_39;
   assign m218_39 ={ {4{in218[5]}} , in218[5:0] };

   // m218_40 = W*in
   wire signed [9:0] m218_40;
   assign m218_40 =10'b0;

   // m218_41 = W*in
   wire signed [9:0] m218_41;
   assign m218_41 =10'b0;

   // m218_42 = W*in
   wire signed [9:0] m218_42;
   assign m218_42 =10'b0;

   // m218_43 = W*in
   wire signed [9:0] m218_43;
   assign m218_43 =10'b0;

   // m218_44 = W*in
   wire signed [9:0] m218_44;
   assign m218_44 =10'b0;

   // m218_45 = W*in
   wire signed [9:0] m218_45;
   assign m218_45 =10'b0;

   // m218_46 = W*in
   wire signed [9:0] m218_46;
   assign m218_46 =10'b0;

   // m218_47 = W*in
   wire signed [9:0] m218_47;
   assign m218_47 ={ {4{in218[5]}} , in218[5:0] };

   // m218_48 = W*in
   wire signed [9:0] m218_48;
   assign m218_48 =10'b0;

   // m218_49 = W*in
   wire signed [9:0] m218_49;
   assign m218_49 =10'b0;

   // m218_50 = W*in
   wire signed [9:0] m218_50;
   assign m218_50 =10'b0;

   // m218_51 = W*in
   wire signed [9:0] m218_51;
   assign m218_51 =10'b0;

   // m218_52 = W*in
   wire signed [9:0] m218_52;
   assign m218_52 =10'b0;

   // m218_53 = W*in
   wire signed [9:0] m218_53;
   assign m218_53 =10'b0;

   // m218_54 = W*in
   wire signed [9:0] m218_54;
   assign m218_54 =10'b0;

   // m218_55 = W*in
   wire signed [9:0] m218_55;
   assign m218_55 =10'b0;

   // m218_56 = W*in
   wire signed [9:0] m218_56;
   assign m218_56 =10'b0;

   // m218_57 = W*in
   wire signed [9:0] m218_57;
   assign m218_57 =10'b0;

   // m218_58 = W*in
   wire signed [9:0] m218_58;
   assign m218_58 =10'b0;

   // m218_59 = W*in
   wire signed [9:0] m218_59;
   assign m218_59 =10'b0;

   // m218_60 = W*in
   wire signed [9:0] m218_60;
   assign m218_60 ={ {4{in218[5]}} , in218[5:0] };

   // m218_61 = W*in
   wire signed [9:0] m218_61;
   assign m218_61 =10'b0;

   // m218_62 = W*in
   wire signed [9:0] m218_62;
   assign m218_62 =10'b0;

   // m218_63 = W*in
   wire signed [9:0] m218_63;
   assign m218_63 =10'b0;

   // m218_64 = W*in
   wire signed [9:0] m218_64;
   assign m218_64 ={ {4{in218[5]}} , in218[5:0] };

   // m218_65 = W*in
   wire signed [9:0] m218_65;
   assign m218_65 =10'b0;

   // m218_66 = W*in
   wire signed [9:0] m218_66;
   assign m218_66 =10'b0;

   // m218_67 = W*in
   wire signed [9:0] m218_67;
   assign m218_67 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_68 = W*in
   wire signed [9:0] m218_68;
   assign m218_68 =10'b0;

   // m218_69 = W*in
   wire signed [9:0] m218_69;
   assign m218_69 ={ {4{neg218[5]}} , neg218[5:0] };

   // m218_70 = W*in
   wire signed [9:0] m218_70;
   assign m218_70 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_71 = W*in
   wire signed [9:0] m218_71;
   assign m218_71 ={ {5{in218[5]}} , in218[5:1] };

   // m218_72 = W*in
   wire signed [9:0] m218_72;
   assign m218_72 =10'b0;

   // m218_73 = W*in
   wire signed [9:0] m218_73;
   assign m218_73 =10'b0;

   // m218_74 = W*in
   wire signed [9:0] m218_74;
   assign m218_74 =10'b0;

   // m218_75 = W*in
   wire signed [9:0] m218_75;
   assign m218_75 =10'b0;

   // m218_76 = W*in
   wire signed [9:0] m218_76;
   assign m218_76 =10'b0;

   // m218_77 = W*in
   wire signed [9:0] m218_77;
   assign m218_77 =10'b0;

   // m218_78 = W*in
   wire signed [9:0] m218_78;
   assign m218_78 =10'b0;

   // m218_79 = W*in
   wire signed [9:0] m218_79;
   assign m218_79 =10'b0;

   // m218_80 = W*in
   wire signed [9:0] m218_80;
   assign m218_80 =10'b0;

   // m218_81 = W*in
   wire signed [9:0] m218_81;
   assign m218_81 =10'b0;

   // m218_82 = W*in
   wire signed [9:0] m218_82;
   assign m218_82 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_83 = W*in
   wire signed [9:0] m218_83;
   assign m218_83 =10'b0;

   // m218_84 = W*in
   wire signed [9:0] m218_84;
   assign m218_84 =10'b0;

   // m218_85 = W*in
   wire signed [9:0] m218_85;
   assign m218_85 ={ {5{neg218[5]}} , neg218[5:1] };

   // m218_86 = W*in
   wire signed [9:0] m218_86;
   assign m218_86 =10'b0;

   // m218_87 = W*in
   wire signed [9:0] m218_87;
   assign m218_87 =10'b0;

   // m218_88 = W*in
   wire signed [9:0] m218_88;
   assign m218_88 ={ {4{neg218[5]}} , neg218[5:0] };

   // m218_89 = W*in
   wire signed [9:0] m218_89;
   assign m218_89 ={ {4{in218[5]}} , in218[5:0] };

   // m218_90 = W*in
   wire signed [9:0] m218_90;
   assign m218_90 =10'b0;

   // m218_91 = W*in
   wire signed [9:0] m218_91;
   assign m218_91 =10'b0;

   // m218_92 = W*in
   wire signed [9:0] m218_92;
   assign m218_92 =10'b0;

   // m218_93 = W*in
   wire signed [9:0] m218_93;
   assign m218_93 =10'b0;

   // m218_94 = W*in
   wire signed [9:0] m218_94;
   assign m218_94 =10'b0;

   // m218_95 = W*in
   wire signed [9:0] m218_95;
   assign m218_95 =10'b0;

   // m218_96 = W*in
   wire signed [9:0] m218_96;
   assign m218_96 =10'b0;

   // m218_97 = W*in
   wire signed [9:0] m218_97;
   assign m218_97 =10'b0;

   // m218_98 = W*in
   wire signed [9:0] m218_98;
   assign m218_98 =10'b0;

   // m218_99 = W*in
   wire signed [9:0] m218_99;
   assign m218_99 =10'b0;

   // m218_100 = W*in
   wire signed [9:0] m218_100;
   assign m218_100 =10'b0;

   // m218_101 = W*in
   wire signed [9:0] m218_101;
   assign m218_101 =10'b0;

   // m218_102 = W*in
   wire signed [9:0] m218_102;
   assign m218_102 =10'b0;

   // m218_103 = W*in
   wire signed [9:0] m218_103;
   assign m218_103 =10'b0;

   // m218_104 = W*in
   wire signed [9:0] m218_104;
   assign m218_104 =10'b0;

   // m218_105 = W*in
   wire signed [9:0] m218_105;
   assign m218_105 =10'b0;

   // m218_106 = W*in
   wire signed [9:0] m218_106;
   assign m218_106 =10'b0;

   // m218_107 = W*in
   wire signed [9:0] m218_107;
   assign m218_107 =10'b0;

   // m218_108 = W*in
   wire signed [9:0] m218_108;
   assign m218_108 ={ {5{in218[5]}} , in218[5:1] };

   // m218_109 = W*in
   wire signed [9:0] m218_109;
   assign m218_109 ={ {4{in218[5]}} , in218[5:0] };

   // m218_110 = W*in
   wire signed [9:0] m218_110;
   assign m218_110 =10'b0;

   // m218_111 = W*in
   wire signed [9:0] m218_111;
   assign m218_111 =10'b0;

   // m218_112 = W*in
   wire signed [9:0] m218_112;
   assign m218_112 =10'b0;

   // m218_113 = W*in
   wire signed [9:0] m218_113;
   assign m218_113 =10'b0;

   // m218_114 = W*in
   wire signed [9:0] m218_114;
   assign m218_114 ={ {4{in218[5]}} , in218[5:0] };

   // m218_115 = W*in
   wire signed [9:0] m218_115;
   assign m218_115 =10'b0;

   // m218_116 = W*in
   wire signed [9:0] m218_116;
   assign m218_116 =10'b0;

   // m218_117 = W*in
   wire signed [9:0] m218_117;
   assign m218_117 =10'b0;

   // m219_1 = W*in
   wire signed [9:0] m219_1;
   assign m219_1 =10'b0;

   // m219_2 = W*in
   wire signed [9:0] m219_2;
   assign m219_2 =10'b0;

   // m219_3 = W*in
   wire signed [9:0] m219_3;
   assign m219_3 =10'b0;

   // m219_4 = W*in
   wire signed [9:0] m219_4;
   assign m219_4 =10'b0;

   // m219_5 = W*in
   wire signed [9:0] m219_5;
   assign m219_5 =10'b0;

   // m219_6 = W*in
   wire signed [9:0] m219_6;
   assign m219_6 =10'b0;

   // m219_7 = W*in
   wire signed [9:0] m219_7;
   assign m219_7 ={ {4{in219[5]}} , in219[5:0] };

   // m219_8 = W*in
   wire signed [9:0] m219_8;
   assign m219_8 =10'b0;

   // m219_9 = W*in
   wire signed [9:0] m219_9;
   assign m219_9 =10'b0;

   // m219_10 = W*in
   wire signed [9:0] m219_10;
   assign m219_10 ={ {4{in219[5]}} , in219[5:0] };

   // m219_11 = W*in
   wire signed [9:0] m219_11;
   assign m219_11 =10'b0;

   // m219_12 = W*in
   wire signed [9:0] m219_12;
   assign m219_12 =10'b0;

   // m219_13 = W*in
   wire signed [9:0] m219_13;
   assign m219_13 =10'b0;

   // m219_14 = W*in
   wire signed [9:0] m219_14;
   assign m219_14 =10'b0;

   // m219_15 = W*in
   wire signed [9:0] m219_15;
   assign m219_15 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_16 = W*in
   wire signed [9:0] m219_16;
   assign m219_16 ={ {4{in219[5]}} , in219[5:0] };

   // m219_17 = W*in
   wire signed [9:0] m219_17;
   assign m219_17 ={ {5{neg219[5]}} , neg219[5:1] };

   // m219_18 = W*in
   wire signed [9:0] m219_18;
   assign m219_18 ={ {4{in219[5]}} , in219[5:0] };

   // m219_19 = W*in
   wire signed [9:0] m219_19;
   assign m219_19 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_20 = W*in
   wire signed [9:0] m219_20;
   assign m219_20 =10'b0;

   // m219_21 = W*in
   wire signed [9:0] m219_21;
   assign m219_21 =10'b0;

   // m219_22 = W*in
   wire signed [9:0] m219_22;
   assign m219_22 =10'b0;

   // m219_23 = W*in
   wire signed [9:0] m219_23;
   assign m219_23 =10'b0;

   // m219_24 = W*in
   wire signed [9:0] m219_24;
   assign m219_24 =10'b0;

   // m219_25 = W*in
   wire signed [9:0] m219_25;
   assign m219_25 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_26 = W*in
   wire signed [9:0] m219_26;
   assign m219_26 ={ {3{in219[5]}} , in219 , {1{1'b0}} };

   // m219_27 = W*in
   wire signed [9:0] m219_27;
   assign m219_27 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_28 = W*in
   wire signed [9:0] m219_28;
   assign m219_28 ={ {5{neg219[5]}} , neg219[5:1] };

   // m219_29 = W*in
   wire signed [9:0] m219_29;
   assign m219_29 =10'b0;

   // m219_30 = W*in
   wire signed [9:0] m219_30;
   assign m219_30 =10'b0;

   // m219_31 = W*in
   wire signed [9:0] m219_31;
   assign m219_31 ={ {5{neg219[5]}} , neg219[5:1] };

   // m219_32 = W*in
   wire signed [9:0] m219_32;
   assign m219_32 =10'b0;

   // m219_33 = W*in
   wire signed [9:0] m219_33;
   assign m219_33 =10'b0;

   // m219_34 = W*in
   wire signed [9:0] m219_34;
   assign m219_34 =10'b0;

   // m219_35 = W*in
   wire signed [9:0] m219_35;
   assign m219_35 =10'b0;

   // m219_36 = W*in
   wire signed [9:0] m219_36;
   assign m219_36 =10'b0;

   // m219_37 = W*in
   wire signed [9:0] m219_37;
   assign m219_37 =10'b0;

   // m219_38 = W*in
   wire signed [9:0] m219_38;
   assign m219_38 =10'b0;

   // m219_39 = W*in
   wire signed [9:0] m219_39;
   assign m219_39 =10'b0;

   // m219_40 = W*in
   wire signed [9:0] m219_40;
   assign m219_40 =10'b0;

   // m219_41 = W*in
   wire signed [9:0] m219_41;
   assign m219_41 =10'b0;

   // m219_42 = W*in
   wire signed [9:0] m219_42;
   assign m219_42 =10'b0;

   // m219_43 = W*in
   wire signed [9:0] m219_43;
   assign m219_43 =10'b0;

   // m219_44 = W*in
   wire signed [9:0] m219_44;
   assign m219_44 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_45 = W*in
   wire signed [9:0] m219_45;
   assign m219_45 =10'b0;

   // m219_46 = W*in
   wire signed [9:0] m219_46;
   assign m219_46 =10'b0;

   // m219_47 = W*in
   wire signed [9:0] m219_47;
   assign m219_47 =10'b0;

   // m219_48 = W*in
   wire signed [9:0] m219_48;
   assign m219_48 =10'b0;

   // m219_49 = W*in
   wire signed [9:0] m219_49;
   assign m219_49 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_50 = W*in
   wire signed [9:0] m219_50;
   assign m219_50 =10'b0;

   // m219_51 = W*in
   wire signed [9:0] m219_51;
   assign m219_51 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_52 = W*in
   wire signed [9:0] m219_52;
   assign m219_52 =10'b0;

   // m219_53 = W*in
   wire signed [9:0] m219_53;
   assign m219_53 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_54 = W*in
   wire signed [9:0] m219_54;
   assign m219_54 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_55 = W*in
   wire signed [9:0] m219_55;
   assign m219_55 ={ {4{in219[5]}} , in219[5:0] };

   // m219_56 = W*in
   wire signed [9:0] m219_56;
   assign m219_56 =10'b0;

   // m219_57 = W*in
   wire signed [9:0] m219_57;
   assign m219_57 =10'b0;

   // m219_58 = W*in
   wire signed [9:0] m219_58;
   assign m219_58 =10'b0;

   // m219_59 = W*in
   wire signed [9:0] m219_59;
   assign m219_59 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_60 = W*in
   wire signed [9:0] m219_60;
   assign m219_60 =10'b0;

   // m219_61 = W*in
   wire signed [9:0] m219_61;
   assign m219_61 =10'b0;

   // m219_62 = W*in
   wire signed [9:0] m219_62;
   assign m219_62 =10'b0;

   // m219_63 = W*in
   wire signed [9:0] m219_63;
   assign m219_63 =10'b0;

   // m219_64 = W*in
   wire signed [9:0] m219_64;
   assign m219_64 ={ {5{in219[5]}} , in219[5:1] };

   // m219_65 = W*in
   wire signed [9:0] m219_65;
   assign m219_65 =10'b0;

   // m219_66 = W*in
   wire signed [9:0] m219_66;
   assign m219_66 =10'b0;

   // m219_67 = W*in
   wire signed [9:0] m219_67;
   assign m219_67 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_68 = W*in
   wire signed [9:0] m219_68;
   assign m219_68 =10'b0;

   // m219_69 = W*in
   wire signed [9:0] m219_69;
   assign m219_69 ={ {4{in219[5]}} , in219[5:0] };

   // m219_70 = W*in
   wire signed [9:0] m219_70;
   assign m219_70 ={ {4{in219[5]}} , in219[5:0] };

   // m219_71 = W*in
   wire signed [9:0] m219_71;
   assign m219_71 ={ {5{in219[5]}} , in219[5:1] };

   // m219_72 = W*in
   wire signed [9:0] m219_72;
   assign m219_72 ={ {4{in219[5]}} , in219[5:0] };

   // m219_73 = W*in
   wire signed [9:0] m219_73;
   assign m219_73 ={ {5{neg219[5]}} , neg219[5:1] };

   // m219_74 = W*in
   wire signed [9:0] m219_74;
   assign m219_74 ={ {4{in219[5]}} , in219[5:0] };

   // m219_75 = W*in
   wire signed [9:0] m219_75;
   assign m219_75 =10'b0;

   // m219_76 = W*in
   wire signed [9:0] m219_76;
   assign m219_76 =10'b0;

   // m219_77 = W*in
   wire signed [9:0] m219_77;
   assign m219_77 =10'b0;

   // m219_78 = W*in
   wire signed [9:0] m219_78;
   assign m219_78 ={ {4{in219[5]}} , in219[5:0] };

   // m219_79 = W*in
   wire signed [9:0] m219_79;
   assign m219_79 =10'b0;

   // m219_80 = W*in
   wire signed [9:0] m219_80;
   assign m219_80 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_81 = W*in
   wire signed [9:0] m219_81;
   assign m219_81 =10'b0;

   // m219_82 = W*in
   wire signed [9:0] m219_82;
   assign m219_82 =10'b0;

   // m219_83 = W*in
   wire signed [9:0] m219_83;
   assign m219_83 =10'b0;

   // m219_84 = W*in
   wire signed [9:0] m219_84;
   assign m219_84 ={ {4{in219[5]}} , in219[5:0] };

   // m219_85 = W*in
   wire signed [9:0] m219_85;
   assign m219_85 =10'b0;

   // m219_86 = W*in
   wire signed [9:0] m219_86;
   assign m219_86 ={ {4{in219[5]}} , in219[5:0] };

   // m219_87 = W*in
   wire signed [9:0] m219_87;
   assign m219_87 =10'b0;

   // m219_88 = W*in
   wire signed [9:0] m219_88;
   assign m219_88 =10'b0;

   // m219_89 = W*in
   wire signed [9:0] m219_89;
   assign m219_89 =10'b0;

   // m219_90 = W*in
   wire signed [9:0] m219_90;
   assign m219_90 =10'b0;

   // m219_91 = W*in
   wire signed [9:0] m219_91;
   assign m219_91 =10'b0;

   // m219_92 = W*in
   wire signed [9:0] m219_92;
   assign m219_92 =10'b0;

   // m219_93 = W*in
   wire signed [9:0] m219_93;
   assign m219_93 =10'b0;

   // m219_94 = W*in
   wire signed [9:0] m219_94;
   assign m219_94 ={ {4{in219[5]}} , in219[5:0] };

   // m219_95 = W*in
   wire signed [9:0] m219_95;
   assign m219_95 =10'b0;

   // m219_96 = W*in
   wire signed [9:0] m219_96;
   assign m219_96 =10'b0;

   // m219_97 = W*in
   wire signed [9:0] m219_97;
   assign m219_97 ={ {4{neg219[5]}} , neg219[5:0] };

   // m219_98 = W*in
   wire signed [9:0] m219_98;
   assign m219_98 =10'b0;

   // m219_99 = W*in
   wire signed [9:0] m219_99;
   assign m219_99 ={ {4{in219[5]}} , in219[5:0] };

   // m219_100 = W*in
   wire signed [9:0] m219_100;
   assign m219_100 =10'b0;

   // m219_101 = W*in
   wire signed [9:0] m219_101;
   assign m219_101 =10'b0;

   // m219_102 = W*in
   wire signed [9:0] m219_102;
   assign m219_102 ={ {4{in219[5]}} , in219[5:0] };

   // m219_103 = W*in
   wire signed [9:0] m219_103;
   assign m219_103 =10'b0;

   // m219_104 = W*in
   wire signed [9:0] m219_104;
   assign m219_104 =10'b0;

   // m219_105 = W*in
   wire signed [9:0] m219_105;
   assign m219_105 =10'b0;

   // m219_106 = W*in
   wire signed [9:0] m219_106;
   assign m219_106 =10'b0;

   // m219_107 = W*in
   wire signed [9:0] m219_107;
   assign m219_107 =10'b0;

   // m219_108 = W*in
   wire signed [9:0] m219_108;
   assign m219_108 =10'b0;

   // m219_109 = W*in
   wire signed [9:0] m219_109;
   assign m219_109 =10'b0;

   // m219_110 = W*in
   wire signed [9:0] m219_110;
   assign m219_110 =10'b0;

   // m219_111 = W*in
   wire signed [9:0] m219_111;
   assign m219_111 =10'b0;

   // m219_112 = W*in
   wire signed [9:0] m219_112;
   assign m219_112 =10'b0;

   // m219_113 = W*in
   wire signed [9:0] m219_113;
   assign m219_113 =10'b0;

   // m219_114 = W*in
   wire signed [9:0] m219_114;
   assign m219_114 =10'b0;

   // m219_115 = W*in
   wire signed [9:0] m219_115;
   assign m219_115 ={ {5{neg219[5]}} , neg219[5:1] };

   // m219_116 = W*in
   wire signed [9:0] m219_116;
   assign m219_116 =10'b0;

   // m219_117 = W*in
   wire signed [9:0] m219_117;
   assign m219_117 =10'b0;

   // m220_1 = W*in
   wire signed [9:0] m220_1;
   assign m220_1 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_2 = W*in
   wire signed [9:0] m220_2;
   assign m220_2 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_3 = W*in
   wire signed [9:0] m220_3;
   assign m220_3 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_4 = W*in
   wire signed [9:0] m220_4;
   assign m220_4 =10'b0;

   // m220_5 = W*in
   wire signed [9:0] m220_5;
   assign m220_5 =10'b0;

   // m220_6 = W*in
   wire signed [9:0] m220_6;
   assign m220_6 ={ {4{in220[5]}} , in220[5:0] };

   // m220_7 = W*in
   wire signed [9:0] m220_7;
   assign m220_7 =10'b0;

   // m220_8 = W*in
   wire signed [9:0] m220_8;
   assign m220_8 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_9 = W*in
   wire signed [9:0] m220_9;
   assign m220_9 =10'b0;

   // m220_10 = W*in
   wire signed [9:0] m220_10;
   assign m220_10 =10'b0;

   // m220_11 = W*in
   wire signed [9:0] m220_11;
   assign m220_11 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_12 = W*in
   wire signed [9:0] m220_12;
   assign m220_12 =10'b0;

   // m220_13 = W*in
   wire signed [9:0] m220_13;
   assign m220_13 =10'b0;

   // m220_14 = W*in
   wire signed [9:0] m220_14;
   assign m220_14 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_15 = W*in
   wire signed [9:0] m220_15;
   assign m220_15 =10'b0;

   // m220_16 = W*in
   wire signed [9:0] m220_16;
   assign m220_16 =10'b0;

   // m220_17 = W*in
   wire signed [9:0] m220_17;
   assign m220_17 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_18 = W*in
   wire signed [9:0] m220_18;
   assign m220_18 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_19 = W*in
   wire signed [9:0] m220_19;
   assign m220_19 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_20 = W*in
   wire signed [9:0] m220_20;
   assign m220_20 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_21 = W*in
   wire signed [9:0] m220_21;
   assign m220_21 ={ {4{in220[5]}} , in220[5:0] };

   // m220_22 = W*in
   wire signed [9:0] m220_22;
   assign m220_22 =10'b0;

   // m220_23 = W*in
   wire signed [9:0] m220_23;
   assign m220_23 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_24 = W*in
   wire signed [9:0] m220_24;
   assign m220_24 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_25 = W*in
   wire signed [9:0] m220_25;
   assign m220_25 =10'b0;

   // m220_26 = W*in
   wire signed [9:0] m220_26;
   assign m220_26 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_27 = W*in
   wire signed [9:0] m220_27;
   assign m220_27 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_28 = W*in
   wire signed [9:0] m220_28;
   assign m220_28 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_29 = W*in
   wire signed [9:0] m220_29;
   assign m220_29 ={ {4{in220[5]}} , in220[5:0] };

   // m220_30 = W*in
   wire signed [9:0] m220_30;
   assign m220_30 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_31 = W*in
   wire signed [9:0] m220_31;
   assign m220_31 ={ {5{neg220[5]}} , neg220[5:1] };

   // m220_32 = W*in
   wire signed [9:0] m220_32;
   assign m220_32 ={ {5{in220[5]}} , in220[5:1] };

   // m220_33 = W*in
   wire signed [9:0] m220_33;
   assign m220_33 ={ {4{in220[5]}} , in220[5:0] };

   // m220_34 = W*in
   wire signed [9:0] m220_34;
   assign m220_34 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_35 = W*in
   wire signed [9:0] m220_35;
   assign m220_35 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_36 = W*in
   wire signed [9:0] m220_36;
   assign m220_36 =10'b0;

   // m220_37 = W*in
   wire signed [9:0] m220_37;
   assign m220_37 =10'b0;

   // m220_38 = W*in
   wire signed [9:0] m220_38;
   assign m220_38 ={ {4{in220[5]}} , in220[5:0] };

   // m220_39 = W*in
   wire signed [9:0] m220_39;
   assign m220_39 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_40 = W*in
   wire signed [9:0] m220_40;
   assign m220_40 =10'b0;

   // m220_41 = W*in
   wire signed [9:0] m220_41;
   assign m220_41 =10'b0;

   // m220_42 = W*in
   wire signed [9:0] m220_42;
   assign m220_42 =10'b0;

   // m220_43 = W*in
   wire signed [9:0] m220_43;
   assign m220_43 ={ {4{in220[5]}} , in220[5:0] };

   // m220_44 = W*in
   wire signed [9:0] m220_44;
   assign m220_44 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_45 = W*in
   wire signed [9:0] m220_45;
   assign m220_45 =10'b0;

   // m220_46 = W*in
   wire signed [9:0] m220_46;
   assign m220_46 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_47 = W*in
   wire signed [9:0] m220_47;
   assign m220_47 =10'b0;

   // m220_48 = W*in
   wire signed [9:0] m220_48;
   assign m220_48 ={ {4{in220[5]}} , in220[5:0] };

   // m220_49 = W*in
   wire signed [9:0] m220_49;
   assign m220_49 =10'b0;

   // m220_50 = W*in
   wire signed [9:0] m220_50;
   assign m220_50 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_51 = W*in
   wire signed [9:0] m220_51;
   assign m220_51 =10'b0;

   // m220_52 = W*in
   wire signed [9:0] m220_52;
   assign m220_52 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_53 = W*in
   wire signed [9:0] m220_53;
   assign m220_53 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_54 = W*in
   wire signed [9:0] m220_54;
   assign m220_54 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_55 = W*in
   wire signed [9:0] m220_55;
   assign m220_55 ={ {4{in220[5]}} , in220[5:0] };

   // m220_56 = W*in
   wire signed [9:0] m220_56;
   assign m220_56 =10'b0;

   // m220_57 = W*in
   wire signed [9:0] m220_57;
   assign m220_57 =10'b0;

   // m220_58 = W*in
   wire signed [9:0] m220_58;
   assign m220_58 =10'b0;

   // m220_59 = W*in
   wire signed [9:0] m220_59;
   assign m220_59 =10'b0;

   // m220_60 = W*in
   wire signed [9:0] m220_60;
   assign m220_60 ={ {3{neg220[5]}} , neg220 , {1{1'b0}} };

   // m220_61 = W*in
   wire signed [9:0] m220_61;
   assign m220_61 ={ {3{neg220[5]}} , neg220 , {1{1'b0}} };

   // m220_62 = W*in
   wire signed [9:0] m220_62;
   assign m220_62 =10'b0;

   // m220_63 = W*in
   wire signed [9:0] m220_63;
   assign m220_63 ={ {4{in220[5]}} , in220[5:0] };

   // m220_64 = W*in
   wire signed [9:0] m220_64;
   assign m220_64 ={ {4{in220[5]}} , in220[5:0] };

   // m220_65 = W*in
   wire signed [9:0] m220_65;
   assign m220_65 ={ {4{in220[5]}} , in220[5:0] };

   // m220_66 = W*in
   wire signed [9:0] m220_66;
   assign m220_66 =10'b0;

   // m220_67 = W*in
   wire signed [9:0] m220_67;
   assign m220_67 =10'b0;

   // m220_68 = W*in
   wire signed [9:0] m220_68;
   assign m220_68 =10'b0;

   // m220_69 = W*in
   wire signed [9:0] m220_69;
   assign m220_69 =10'b0;

   // m220_70 = W*in
   wire signed [9:0] m220_70;
   assign m220_70 ={ {4{in220[5]}} , in220[5:0] };

   // m220_71 = W*in
   wire signed [9:0] m220_71;
   assign m220_71 =10'b0;

   // m220_72 = W*in
   wire signed [9:0] m220_72;
   assign m220_72 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_73 = W*in
   wire signed [9:0] m220_73;
   assign m220_73 =10'b0;

   // m220_74 = W*in
   wire signed [9:0] m220_74;
   assign m220_74 ={ {4{in220[5]}} , in220[5:0] };

   // m220_75 = W*in
   wire signed [9:0] m220_75;
   assign m220_75 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_76 = W*in
   wire signed [9:0] m220_76;
   assign m220_76 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_77 = W*in
   wire signed [9:0] m220_77;
   assign m220_77 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_78 = W*in
   wire signed [9:0] m220_78;
   assign m220_78 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_79 = W*in
   wire signed [9:0] m220_79;
   assign m220_79 =10'b0;

   // m220_80 = W*in
   wire signed [9:0] m220_80;
   assign m220_80 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_81 = W*in
   wire signed [9:0] m220_81;
   assign m220_81 =10'b0;

   // m220_82 = W*in
   wire signed [9:0] m220_82;
   assign m220_82 ={ {5{neg220[5]}} , neg220[5:1] };

   // m220_83 = W*in
   wire signed [9:0] m220_83;
   assign m220_83 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_84 = W*in
   wire signed [9:0] m220_84;
   assign m220_84 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_85 = W*in
   wire signed [9:0] m220_85;
   assign m220_85 ={ {5{neg220[5]}} , neg220[5:1] };

   // m220_86 = W*in
   wire signed [9:0] m220_86;
   assign m220_86 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_87 = W*in
   wire signed [9:0] m220_87;
   assign m220_87 ={ {4{in220[5]}} , in220[5:0] };

   // m220_88 = W*in
   wire signed [9:0] m220_88;
   assign m220_88 =10'b0;

   // m220_89 = W*in
   wire signed [9:0] m220_89;
   assign m220_89 ={ {4{in220[5]}} , in220[5:0] };

   // m220_90 = W*in
   wire signed [9:0] m220_90;
   assign m220_90 =10'b0;

   // m220_91 = W*in
   wire signed [9:0] m220_91;
   assign m220_91 =10'b0;

   // m220_92 = W*in
   wire signed [9:0] m220_92;
   assign m220_92 =10'b0;

   // m220_93 = W*in
   wire signed [9:0] m220_93;
   assign m220_93 =10'b0;

   // m220_94 = W*in
   wire signed [9:0] m220_94;
   assign m220_94 ={ {3{in220[5]}} , in220 , {1{1'b0}} };

   // m220_95 = W*in
   wire signed [9:0] m220_95;
   assign m220_95 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_96 = W*in
   wire signed [9:0] m220_96;
   assign m220_96 =10'b0;

   // m220_97 = W*in
   wire signed [9:0] m220_97;
   assign m220_97 =10'b0;

   // m220_98 = W*in
   wire signed [9:0] m220_98;
   assign m220_98 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_99 = W*in
   wire signed [9:0] m220_99;
   assign m220_99 ={ {4{in220[5]}} , in220[5:0] };

   // m220_100 = W*in
   wire signed [9:0] m220_100;
   assign m220_100 =10'b0;

   // m220_101 = W*in
   wire signed [9:0] m220_101;
   assign m220_101 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_102 = W*in
   wire signed [9:0] m220_102;
   assign m220_102 =10'b0;

   // m220_103 = W*in
   wire signed [9:0] m220_103;
   assign m220_103 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_104 = W*in
   wire signed [9:0] m220_104;
   assign m220_104 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_105 = W*in
   wire signed [9:0] m220_105;
   assign m220_105 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_106 = W*in
   wire signed [9:0] m220_106;
   assign m220_106 =10'b0;

   // m220_107 = W*in
   wire signed [9:0] m220_107;
   assign m220_107 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_108 = W*in
   wire signed [9:0] m220_108;
   assign m220_108 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_109 = W*in
   wire signed [9:0] m220_109;
   assign m220_109 =10'b0;

   // m220_110 = W*in
   wire signed [9:0] m220_110;
   assign m220_110 =10'b0;

   // m220_111 = W*in
   wire signed [9:0] m220_111;
   assign m220_111 ={ {4{in220[5]}} , in220[5:0] };

   // m220_112 = W*in
   wire signed [9:0] m220_112;
   assign m220_112 ={ {4{in220[5]}} , in220[5:0] };

   // m220_113 = W*in
   wire signed [9:0] m220_113;
   assign m220_113 =10'b0;

   // m220_114 = W*in
   wire signed [9:0] m220_114;
   assign m220_114 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_115 = W*in
   wire signed [9:0] m220_115;
   assign m220_115 ={ {4{neg220[5]}} , neg220[5:0] };

   // m220_116 = W*in
   wire signed [9:0] m220_116;
   assign m220_116 =10'b0;

   // m220_117 = W*in
   wire signed [9:0] m220_117;
   assign m220_117 ={ {3{neg220[5]}} , neg220 , {1{1'b0}} };

   // m221_1 = W*in
   wire signed [9:0] m221_1;
   assign m221_1 =10'b0;

   // m221_2 = W*in
   wire signed [9:0] m221_2;
   assign m221_2 =10'b0;

   // m221_3 = W*in
   wire signed [9:0] m221_3;
   assign m221_3 =10'b0;

   // m221_4 = W*in
   wire signed [9:0] m221_4;
   assign m221_4 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_5 = W*in
   wire signed [9:0] m221_5;
   assign m221_5 ={ {4{in221[5]}} , in221[5:0] };

   // m221_6 = W*in
   wire signed [9:0] m221_6;
   assign m221_6 =10'b0;

   // m221_7 = W*in
   wire signed [9:0] m221_7;
   assign m221_7 =10'b0;

   // m221_8 = W*in
   wire signed [9:0] m221_8;
   assign m221_8 =10'b0;

   // m221_9 = W*in
   wire signed [9:0] m221_9;
   assign m221_9 =10'b0;

   // m221_10 = W*in
   wire signed [9:0] m221_10;
   assign m221_10 =10'b0;

   // m221_11 = W*in
   wire signed [9:0] m221_11;
   assign m221_11 =10'b0;

   // m221_12 = W*in
   wire signed [9:0] m221_12;
   assign m221_12 ={ {4{in221[5]}} , in221[5:0] };

   // m221_13 = W*in
   wire signed [9:0] m221_13;
   assign m221_13 =10'b0;

   // m221_14 = W*in
   wire signed [9:0] m221_14;
   assign m221_14 =10'b0;

   // m221_15 = W*in
   wire signed [9:0] m221_15;
   assign m221_15 =10'b0;

   // m221_16 = W*in
   wire signed [9:0] m221_16;
   assign m221_16 =10'b0;

   // m221_17 = W*in
   wire signed [9:0] m221_17;
   assign m221_17 ={ {5{neg221[5]}} , neg221[5:1] };

   // m221_18 = W*in
   wire signed [9:0] m221_18;
   assign m221_18 ={ {5{in221[5]}} , in221[5:1] };

   // m221_19 = W*in
   wire signed [9:0] m221_19;
   assign m221_19 =10'b0;

   // m221_20 = W*in
   wire signed [9:0] m221_20;
   assign m221_20 =10'b0;

   // m221_21 = W*in
   wire signed [9:0] m221_21;
   assign m221_21 =10'b0;

   // m221_22 = W*in
   wire signed [9:0] m221_22;
   assign m221_22 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_23 = W*in
   wire signed [9:0] m221_23;
   assign m221_23 =10'b0;

   // m221_24 = W*in
   wire signed [9:0] m221_24;
   assign m221_24 =10'b0;

   // m221_25 = W*in
   wire signed [9:0] m221_25;
   assign m221_25 ={ {4{in221[5]}} , in221[5:0] };

   // m221_26 = W*in
   wire signed [9:0] m221_26;
   assign m221_26 ={ {4{in221[5]}} , in221[5:0] };

   // m221_27 = W*in
   wire signed [9:0] m221_27;
   assign m221_27 =10'b0;

   // m221_28 = W*in
   wire signed [9:0] m221_28;
   assign m221_28 ={ {4{in221[5]}} , in221[5:0] };

   // m221_29 = W*in
   wire signed [9:0] m221_29;
   assign m221_29 =10'b0;

   // m221_30 = W*in
   wire signed [9:0] m221_30;
   assign m221_30 =10'b0;

   // m221_31 = W*in
   wire signed [9:0] m221_31;
   assign m221_31 =10'b0;

   // m221_32 = W*in
   wire signed [9:0] m221_32;
   assign m221_32 ={ {4{in221[5]}} , in221[5:0] };

   // m221_33 = W*in
   wire signed [9:0] m221_33;
   assign m221_33 ={ {4{in221[5]}} , in221[5:0] };

   // m221_34 = W*in
   wire signed [9:0] m221_34;
   assign m221_34 =10'b0;

   // m221_35 = W*in
   wire signed [9:0] m221_35;
   assign m221_35 =10'b0;

   // m221_36 = W*in
   wire signed [9:0] m221_36;
   assign m221_36 =10'b0;

   // m221_37 = W*in
   wire signed [9:0] m221_37;
   assign m221_37 =10'b0;

   // m221_38 = W*in
   wire signed [9:0] m221_38;
   assign m221_38 =10'b0;

   // m221_39 = W*in
   wire signed [9:0] m221_39;
   assign m221_39 =10'b0;

   // m221_40 = W*in
   wire signed [9:0] m221_40;
   assign m221_40 =10'b0;

   // m221_41 = W*in
   wire signed [9:0] m221_41;
   assign m221_41 =10'b0;

   // m221_42 = W*in
   wire signed [9:0] m221_42;
   assign m221_42 =10'b0;

   // m221_43 = W*in
   wire signed [9:0] m221_43;
   assign m221_43 =10'b0;

   // m221_44 = W*in
   wire signed [9:0] m221_44;
   assign m221_44 =10'b0;

   // m221_45 = W*in
   wire signed [9:0] m221_45;
   assign m221_45 =10'b0;

   // m221_46 = W*in
   wire signed [9:0] m221_46;
   assign m221_46 =10'b0;

   // m221_47 = W*in
   wire signed [9:0] m221_47;
   assign m221_47 =10'b0;

   // m221_48 = W*in
   wire signed [9:0] m221_48;
   assign m221_48 =10'b0;

   // m221_49 = W*in
   wire signed [9:0] m221_49;
   assign m221_49 ={ {4{in221[5]}} , in221[5:0] };

   // m221_50 = W*in
   wire signed [9:0] m221_50;
   assign m221_50 =10'b0;

   // m221_51 = W*in
   wire signed [9:0] m221_51;
   assign m221_51 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_52 = W*in
   wire signed [9:0] m221_52;
   assign m221_52 =10'b0;

   // m221_53 = W*in
   wire signed [9:0] m221_53;
   assign m221_53 ={ {4{in221[5]}} , in221[5:0] };

   // m221_54 = W*in
   wire signed [9:0] m221_54;
   assign m221_54 =10'b0;

   // m221_55 = W*in
   wire signed [9:0] m221_55;
   assign m221_55 =10'b0;

   // m221_56 = W*in
   wire signed [9:0] m221_56;
   assign m221_56 =10'b0;

   // m221_57 = W*in
   wire signed [9:0] m221_57;
   assign m221_57 =10'b0;

   // m221_58 = W*in
   wire signed [9:0] m221_58;
   assign m221_58 =10'b0;

   // m221_59 = W*in
   wire signed [9:0] m221_59;
   assign m221_59 ={ {4{in221[5]}} , in221[5:0] };

   // m221_60 = W*in
   wire signed [9:0] m221_60;
   assign m221_60 =10'b0;

   // m221_61 = W*in
   wire signed [9:0] m221_61;
   assign m221_61 =10'b0;

   // m221_62 = W*in
   wire signed [9:0] m221_62;
   assign m221_62 =10'b0;

   // m221_63 = W*in
   wire signed [9:0] m221_63;
   assign m221_63 =10'b0;

   // m221_64 = W*in
   wire signed [9:0] m221_64;
   assign m221_64 ={ {5{in221[5]}} , in221[5:1] };

   // m221_65 = W*in
   wire signed [9:0] m221_65;
   assign m221_65 ={ {4{in221[5]}} , in221[5:0] };

   // m221_66 = W*in
   wire signed [9:0] m221_66;
   assign m221_66 =10'b0;

   // m221_67 = W*in
   wire signed [9:0] m221_67;
   assign m221_67 =10'b0;

   // m221_68 = W*in
   wire signed [9:0] m221_68;
   assign m221_68 =10'b0;

   // m221_69 = W*in
   wire signed [9:0] m221_69;
   assign m221_69 =10'b0;

   // m221_70 = W*in
   wire signed [9:0] m221_70;
   assign m221_70 =10'b0;

   // m221_71 = W*in
   wire signed [9:0] m221_71;
   assign m221_71 =10'b0;

   // m221_72 = W*in
   wire signed [9:0] m221_72;
   assign m221_72 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_73 = W*in
   wire signed [9:0] m221_73;
   assign m221_73 =10'b0;

   // m221_74 = W*in
   wire signed [9:0] m221_74;
   assign m221_74 =10'b0;

   // m221_75 = W*in
   wire signed [9:0] m221_75;
   assign m221_75 =10'b0;

   // m221_76 = W*in
   wire signed [9:0] m221_76;
   assign m221_76 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_77 = W*in
   wire signed [9:0] m221_77;
   assign m221_77 =10'b0;

   // m221_78 = W*in
   wire signed [9:0] m221_78;
   assign m221_78 ={ {5{in221[5]}} , in221[5:1] };

   // m221_79 = W*in
   wire signed [9:0] m221_79;
   assign m221_79 =10'b0;

   // m221_80 = W*in
   wire signed [9:0] m221_80;
   assign m221_80 =10'b0;

   // m221_81 = W*in
   wire signed [9:0] m221_81;
   assign m221_81 =10'b0;

   // m221_82 = W*in
   wire signed [9:0] m221_82;
   assign m221_82 ={ {5{neg221[5]}} , neg221[5:1] };

   // m221_83 = W*in
   wire signed [9:0] m221_83;
   assign m221_83 =10'b0;

   // m221_84 = W*in
   wire signed [9:0] m221_84;
   assign m221_84 =10'b0;

   // m221_85 = W*in
   wire signed [9:0] m221_85;
   assign m221_85 =10'b0;

   // m221_86 = W*in
   wire signed [9:0] m221_86;
   assign m221_86 =10'b0;

   // m221_87 = W*in
   wire signed [9:0] m221_87;
   assign m221_87 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_88 = W*in
   wire signed [9:0] m221_88;
   assign m221_88 =10'b0;

   // m221_89 = W*in
   wire signed [9:0] m221_89;
   assign m221_89 =10'b0;

   // m221_90 = W*in
   wire signed [9:0] m221_90;
   assign m221_90 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_91 = W*in
   wire signed [9:0] m221_91;
   assign m221_91 ={ {4{in221[5]}} , in221[5:0] };

   // m221_92 = W*in
   wire signed [9:0] m221_92;
   assign m221_92 =10'b0;

   // m221_93 = W*in
   wire signed [9:0] m221_93;
   assign m221_93 =10'b0;

   // m221_94 = W*in
   wire signed [9:0] m221_94;
   assign m221_94 ={ {4{in221[5]}} , in221[5:0] };

   // m221_95 = W*in
   wire signed [9:0] m221_95;
   assign m221_95 =10'b0;

   // m221_96 = W*in
   wire signed [9:0] m221_96;
   assign m221_96 =10'b0;

   // m221_97 = W*in
   wire signed [9:0] m221_97;
   assign m221_97 =10'b0;

   // m221_98 = W*in
   wire signed [9:0] m221_98;
   assign m221_98 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_99 = W*in
   wire signed [9:0] m221_99;
   assign m221_99 =10'b0;

   // m221_100 = W*in
   wire signed [9:0] m221_100;
   assign m221_100 =10'b0;

   // m221_101 = W*in
   wire signed [9:0] m221_101;
   assign m221_101 =10'b0;

   // m221_102 = W*in
   wire signed [9:0] m221_102;
   assign m221_102 ={ {4{in221[5]}} , in221[5:0] };

   // m221_103 = W*in
   wire signed [9:0] m221_103;
   assign m221_103 =10'b0;

   // m221_104 = W*in
   wire signed [9:0] m221_104;
   assign m221_104 =10'b0;

   // m221_105 = W*in
   wire signed [9:0] m221_105;
   assign m221_105 =10'b0;

   // m221_106 = W*in
   wire signed [9:0] m221_106;
   assign m221_106 =10'b0;

   // m221_107 = W*in
   wire signed [9:0] m221_107;
   assign m221_107 ={ {4{neg221[5]}} , neg221[5:0] };

   // m221_108 = W*in
   wire signed [9:0] m221_108;
   assign m221_108 =10'b0;

   // m221_109 = W*in
   wire signed [9:0] m221_109;
   assign m221_109 =10'b0;

   // m221_110 = W*in
   wire signed [9:0] m221_110;
   assign m221_110 =10'b0;

   // m221_111 = W*in
   wire signed [9:0] m221_111;
   assign m221_111 ={ {4{in221[5]}} , in221[5:0] };

   // m221_112 = W*in
   wire signed [9:0] m221_112;
   assign m221_112 =10'b0;

   // m221_113 = W*in
   wire signed [9:0] m221_113;
   assign m221_113 =10'b0;

   // m221_114 = W*in
   wire signed [9:0] m221_114;
   assign m221_114 =10'b0;

   // m221_115 = W*in
   wire signed [9:0] m221_115;
   assign m221_115 =10'b0;

   // m221_116 = W*in
   wire signed [9:0] m221_116;
   assign m221_116 ={ {5{neg221[5]}} , neg221[5:1] };

   // m221_117 = W*in
   wire signed [9:0] m221_117;
   assign m221_117 =10'b0;

   // m222_1 = W*in
   wire signed [9:0] m222_1;
   assign m222_1 =10'b0;

   // m222_2 = W*in
   wire signed [9:0] m222_2;
   assign m222_2 =10'b0;

   // m222_3 = W*in
   wire signed [9:0] m222_3;
   assign m222_3 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_4 = W*in
   wire signed [9:0] m222_4;
   assign m222_4 =10'b0;

   // m222_5 = W*in
   wire signed [9:0] m222_5;
   assign m222_5 =10'b0;

   // m222_6 = W*in
   wire signed [9:0] m222_6;
   assign m222_6 ={ {5{in222[5]}} , in222[5:1] };

   // m222_7 = W*in
   wire signed [9:0] m222_7;
   assign m222_7 =10'b0;

   // m222_8 = W*in
   wire signed [9:0] m222_8;
   assign m222_8 =10'b0;

   // m222_9 = W*in
   wire signed [9:0] m222_9;
   assign m222_9 =10'b0;

   // m222_10 = W*in
   wire signed [9:0] m222_10;
   assign m222_10 ={ {4{in222[5]}} , in222[5:0] };

   // m222_11 = W*in
   wire signed [9:0] m222_11;
   assign m222_11 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_12 = W*in
   wire signed [9:0] m222_12;
   assign m222_12 =10'b0;

   // m222_13 = W*in
   wire signed [9:0] m222_13;
   assign m222_13 =10'b0;

   // m222_14 = W*in
   wire signed [9:0] m222_14;
   assign m222_14 =10'b0;

   // m222_15 = W*in
   wire signed [9:0] m222_15;
   assign m222_15 =10'b0;

   // m222_16 = W*in
   wire signed [9:0] m222_16;
   assign m222_16 =10'b0;

   // m222_17 = W*in
   wire signed [9:0] m222_17;
   assign m222_17 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_18 = W*in
   wire signed [9:0] m222_18;
   assign m222_18 =10'b0;

   // m222_19 = W*in
   wire signed [9:0] m222_19;
   assign m222_19 =10'b0;

   // m222_20 = W*in
   wire signed [9:0] m222_20;
   assign m222_20 =10'b0;

   // m222_21 = W*in
   wire signed [9:0] m222_21;
   assign m222_21 =10'b0;

   // m222_22 = W*in
   wire signed [9:0] m222_22;
   assign m222_22 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_23 = W*in
   wire signed [9:0] m222_23;
   assign m222_23 ={ {5{neg222[5]}} , neg222[5:1] };

   // m222_24 = W*in
   wire signed [9:0] m222_24;
   assign m222_24 =10'b0;

   // m222_25 = W*in
   wire signed [9:0] m222_25;
   assign m222_25 ={ {5{neg222[5]}} , neg222[5:1] };

   // m222_26 = W*in
   wire signed [9:0] m222_26;
   assign m222_26 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_27 = W*in
   wire signed [9:0] m222_27;
   assign m222_27 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_28 = W*in
   wire signed [9:0] m222_28;
   assign m222_28 =10'b0;

   // m222_29 = W*in
   wire signed [9:0] m222_29;
   assign m222_29 ={ {4{in222[5]}} , in222[5:0] };

   // m222_30 = W*in
   wire signed [9:0] m222_30;
   assign m222_30 =10'b0;

   // m222_31 = W*in
   wire signed [9:0] m222_31;
   assign m222_31 =10'b0;

   // m222_32 = W*in
   wire signed [9:0] m222_32;
   assign m222_32 ={ {4{in222[5]}} , in222[5:0] };

   // m222_33 = W*in
   wire signed [9:0] m222_33;
   assign m222_33 =10'b0;

   // m222_34 = W*in
   wire signed [9:0] m222_34;
   assign m222_34 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_35 = W*in
   wire signed [9:0] m222_35;
   assign m222_35 =10'b0;

   // m222_36 = W*in
   wire signed [9:0] m222_36;
   assign m222_36 ={ {5{neg222[5]}} , neg222[5:1] };

   // m222_37 = W*in
   wire signed [9:0] m222_37;
   assign m222_37 =10'b0;

   // m222_38 = W*in
   wire signed [9:0] m222_38;
   assign m222_38 =10'b0;

   // m222_39 = W*in
   wire signed [9:0] m222_39;
   assign m222_39 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_40 = W*in
   wire signed [9:0] m222_40;
   assign m222_40 =10'b0;

   // m222_41 = W*in
   wire signed [9:0] m222_41;
   assign m222_41 =10'b0;

   // m222_42 = W*in
   wire signed [9:0] m222_42;
   assign m222_42 =10'b0;

   // m222_43 = W*in
   wire signed [9:0] m222_43;
   assign m222_43 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_44 = W*in
   wire signed [9:0] m222_44;
   assign m222_44 =10'b0;

   // m222_45 = W*in
   wire signed [9:0] m222_45;
   assign m222_45 =10'b0;

   // m222_46 = W*in
   wire signed [9:0] m222_46;
   assign m222_46 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_47 = W*in
   wire signed [9:0] m222_47;
   assign m222_47 =10'b0;

   // m222_48 = W*in
   wire signed [9:0] m222_48;
   assign m222_48 =10'b0;

   // m222_49 = W*in
   wire signed [9:0] m222_49;
   assign m222_49 =10'b0;

   // m222_50 = W*in
   wire signed [9:0] m222_50;
   assign m222_50 =10'b0;

   // m222_51 = W*in
   wire signed [9:0] m222_51;
   assign m222_51 =10'b0;

   // m222_52 = W*in
   wire signed [9:0] m222_52;
   assign m222_52 =10'b0;

   // m222_53 = W*in
   wire signed [9:0] m222_53;
   assign m222_53 =10'b0;

   // m222_54 = W*in
   wire signed [9:0] m222_54;
   assign m222_54 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_55 = W*in
   wire signed [9:0] m222_55;
   assign m222_55 =10'b0;

   // m222_56 = W*in
   wire signed [9:0] m222_56;
   assign m222_56 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_57 = W*in
   wire signed [9:0] m222_57;
   assign m222_57 =10'b0;

   // m222_58 = W*in
   wire signed [9:0] m222_58;
   assign m222_58 =10'b0;

   // m222_59 = W*in
   wire signed [9:0] m222_59;
   assign m222_59 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_60 = W*in
   wire signed [9:0] m222_60;
   assign m222_60 =10'b0;

   // m222_61 = W*in
   wire signed [9:0] m222_61;
   assign m222_61 =10'b0;

   // m222_62 = W*in
   wire signed [9:0] m222_62;
   assign m222_62 =10'b0;

   // m222_63 = W*in
   wire signed [9:0] m222_63;
   assign m222_63 ={ {4{in222[5]}} , in222[5:0] };

   // m222_64 = W*in
   wire signed [9:0] m222_64;
   assign m222_64 =10'b0;

   // m222_65 = W*in
   wire signed [9:0] m222_65;
   assign m222_65 =10'b0;

   // m222_66 = W*in
   wire signed [9:0] m222_66;
   assign m222_66 =10'b0;

   // m222_67 = W*in
   wire signed [9:0] m222_67;
   assign m222_67 ={ {4{in222[5]}} , in222[5:0] };

   // m222_68 = W*in
   wire signed [9:0] m222_68;
   assign m222_68 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_69 = W*in
   wire signed [9:0] m222_69;
   assign m222_69 =10'b0;

   // m222_70 = W*in
   wire signed [9:0] m222_70;
   assign m222_70 =10'b0;

   // m222_71 = W*in
   wire signed [9:0] m222_71;
   assign m222_71 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_72 = W*in
   wire signed [9:0] m222_72;
   assign m222_72 =10'b0;

   // m222_73 = W*in
   wire signed [9:0] m222_73;
   assign m222_73 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_74 = W*in
   wire signed [9:0] m222_74;
   assign m222_74 =10'b0;

   // m222_75 = W*in
   wire signed [9:0] m222_75;
   assign m222_75 =10'b0;

   // m222_76 = W*in
   wire signed [9:0] m222_76;
   assign m222_76 =10'b0;

   // m222_77 = W*in
   wire signed [9:0] m222_77;
   assign m222_77 =10'b0;

   // m222_78 = W*in
   wire signed [9:0] m222_78;
   assign m222_78 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_79 = W*in
   wire signed [9:0] m222_79;
   assign m222_79 =10'b0;

   // m222_80 = W*in
   wire signed [9:0] m222_80;
   assign m222_80 =10'b0;

   // m222_81 = W*in
   wire signed [9:0] m222_81;
   assign m222_81 =10'b0;

   // m222_82 = W*in
   wire signed [9:0] m222_82;
   assign m222_82 =10'b0;

   // m222_83 = W*in
   wire signed [9:0] m222_83;
   assign m222_83 =10'b0;

   // m222_84 = W*in
   wire signed [9:0] m222_84;
   assign m222_84 =10'b0;

   // m222_85 = W*in
   wire signed [9:0] m222_85;
   assign m222_85 ={ {5{in222[5]}} , in222[5:1] };

   // m222_86 = W*in
   wire signed [9:0] m222_86;
   assign m222_86 =10'b0;

   // m222_87 = W*in
   wire signed [9:0] m222_87;
   assign m222_87 =10'b0;

   // m222_88 = W*in
   wire signed [9:0] m222_88;
   assign m222_88 ={ {5{neg222[5]}} , neg222[5:1] };

   // m222_89 = W*in
   wire signed [9:0] m222_89;
   assign m222_89 =10'b0;

   // m222_90 = W*in
   wire signed [9:0] m222_90;
   assign m222_90 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_91 = W*in
   wire signed [9:0] m222_91;
   assign m222_91 =10'b0;

   // m222_92 = W*in
   wire signed [9:0] m222_92;
   assign m222_92 =10'b0;

   // m222_93 = W*in
   wire signed [9:0] m222_93;
   assign m222_93 ={ {4{in222[5]}} , in222[5:0] };

   // m222_94 = W*in
   wire signed [9:0] m222_94;
   assign m222_94 =10'b0;

   // m222_95 = W*in
   wire signed [9:0] m222_95;
   assign m222_95 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_96 = W*in
   wire signed [9:0] m222_96;
   assign m222_96 =10'b0;

   // m222_97 = W*in
   wire signed [9:0] m222_97;
   assign m222_97 =10'b0;

   // m222_98 = W*in
   wire signed [9:0] m222_98;
   assign m222_98 =10'b0;

   // m222_99 = W*in
   wire signed [9:0] m222_99;
   assign m222_99 =10'b0;

   // m222_100 = W*in
   wire signed [9:0] m222_100;
   assign m222_100 =10'b0;

   // m222_101 = W*in
   wire signed [9:0] m222_101;
   assign m222_101 =10'b0;

   // m222_102 = W*in
   wire signed [9:0] m222_102;
   assign m222_102 =10'b0;

   // m222_103 = W*in
   wire signed [9:0] m222_103;
   assign m222_103 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_104 = W*in
   wire signed [9:0] m222_104;
   assign m222_104 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_105 = W*in
   wire signed [9:0] m222_105;
   assign m222_105 =10'b0;

   // m222_106 = W*in
   wire signed [9:0] m222_106;
   assign m222_106 =10'b0;

   // m222_107 = W*in
   wire signed [9:0] m222_107;
   assign m222_107 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_108 = W*in
   wire signed [9:0] m222_108;
   assign m222_108 =10'b0;

   // m222_109 = W*in
   wire signed [9:0] m222_109;
   assign m222_109 =10'b0;

   // m222_110 = W*in
   wire signed [9:0] m222_110;
   assign m222_110 =10'b0;

   // m222_111 = W*in
   wire signed [9:0] m222_111;
   assign m222_111 ={ {4{neg222[5]}} , neg222[5:0] };

   // m222_112 = W*in
   wire signed [9:0] m222_112;
   assign m222_112 =10'b0;

   // m222_113 = W*in
   wire signed [9:0] m222_113;
   assign m222_113 =10'b0;

   // m222_114 = W*in
   wire signed [9:0] m222_114;
   assign m222_114 ={ {5{neg222[5]}} , neg222[5:1] };

   // m222_115 = W*in
   wire signed [9:0] m222_115;
   assign m222_115 =10'b0;

   // m222_116 = W*in
   wire signed [9:0] m222_116;
   assign m222_116 =10'b0;

   // m222_117 = W*in
   wire signed [9:0] m222_117;
   assign m222_117 =10'b0;

   // m223_1 = W*in
   wire signed [9:0] m223_1;
   assign m223_1 =10'b0;

   // m223_2 = W*in
   wire signed [9:0] m223_2;
   assign m223_2 =10'b0;

   // m223_3 = W*in
   wire signed [9:0] m223_3;
   assign m223_3 =10'b0;

   // m223_4 = W*in
   wire signed [9:0] m223_4;
   assign m223_4 =10'b0;

   // m223_5 = W*in
   wire signed [9:0] m223_5;
   assign m223_5 =10'b0;

   // m223_6 = W*in
   wire signed [9:0] m223_6;
   assign m223_6 =10'b0;

   // m223_7 = W*in
   wire signed [9:0] m223_7;
   assign m223_7 =10'b0;

   // m223_8 = W*in
   wire signed [9:0] m223_8;
   assign m223_8 =10'b0;

   // m223_9 = W*in
   wire signed [9:0] m223_9;
   assign m223_9 =10'b0;

   // m223_10 = W*in
   wire signed [9:0] m223_10;
   assign m223_10 =10'b0;

   // m223_11 = W*in
   wire signed [9:0] m223_11;
   assign m223_11 =10'b0;

   // m223_12 = W*in
   wire signed [9:0] m223_12;
   assign m223_12 =10'b0;

   // m223_13 = W*in
   wire signed [9:0] m223_13;
   assign m223_13 =10'b0;

   // m223_14 = W*in
   wire signed [9:0] m223_14;
   assign m223_14 =10'b0;

   // m223_15 = W*in
   wire signed [9:0] m223_15;
   assign m223_15 =10'b0;

   // m223_16 = W*in
   wire signed [9:0] m223_16;
   assign m223_16 =10'b0;

   // m223_17 = W*in
   wire signed [9:0] m223_17;
   assign m223_17 =10'b0;

   // m223_18 = W*in
   wire signed [9:0] m223_18;
   assign m223_18 =10'b0;

   // m223_19 = W*in
   wire signed [9:0] m223_19;
   assign m223_19 =10'b0;

   // m223_20 = W*in
   wire signed [9:0] m223_20;
   assign m223_20 ={ {5{in223[5]}} , in223[5:1] };

   // m223_21 = W*in
   wire signed [9:0] m223_21;
   assign m223_21 =10'b0;

   // m223_22 = W*in
   wire signed [9:0] m223_22;
   assign m223_22 =10'b0;

   // m223_23 = W*in
   wire signed [9:0] m223_23;
   assign m223_23 ={ {4{in223[5]}} , in223[5:0] };

   // m223_24 = W*in
   wire signed [9:0] m223_24;
   assign m223_24 =10'b0;

   // m223_25 = W*in
   wire signed [9:0] m223_25;
   assign m223_25 =10'b0;

   // m223_26 = W*in
   wire signed [9:0] m223_26;
   assign m223_26 =10'b0;

   // m223_27 = W*in
   wire signed [9:0] m223_27;
   assign m223_27 ={ {5{in223[5]}} , in223[5:1] };

   // m223_28 = W*in
   wire signed [9:0] m223_28;
   assign m223_28 ={ {5{in223[5]}} , in223[5:1] };

   // m223_29 = W*in
   wire signed [9:0] m223_29;
   assign m223_29 =10'b0;

   // m223_30 = W*in
   wire signed [9:0] m223_30;
   assign m223_30 =10'b0;

   // m223_31 = W*in
   wire signed [9:0] m223_31;
   assign m223_31 =10'b0;

   // m223_32 = W*in
   wire signed [9:0] m223_32;
   assign m223_32 =10'b0;

   // m223_33 = W*in
   wire signed [9:0] m223_33;
   assign m223_33 =10'b0;

   // m223_34 = W*in
   wire signed [9:0] m223_34;
   assign m223_34 ={ {4{in223[5]}} , in223[5:0] };

   // m223_35 = W*in
   wire signed [9:0] m223_35;
   assign m223_35 ={ {5{in223[5]}} , in223[5:1] };

   // m223_36 = W*in
   wire signed [9:0] m223_36;
   assign m223_36 =10'b0;

   // m223_37 = W*in
   wire signed [9:0] m223_37;
   assign m223_37 =10'b0;

   // m223_38 = W*in
   wire signed [9:0] m223_38;
   assign m223_38 =10'b0;

   // m223_39 = W*in
   wire signed [9:0] m223_39;
   assign m223_39 =10'b0;

   // m223_40 = W*in
   wire signed [9:0] m223_40;
   assign m223_40 =10'b0;

   // m223_41 = W*in
   wire signed [9:0] m223_41;
   assign m223_41 =10'b0;

   // m223_42 = W*in
   wire signed [9:0] m223_42;
   assign m223_42 =10'b0;

   // m223_43 = W*in
   wire signed [9:0] m223_43;
   assign m223_43 =10'b0;

   // m223_44 = W*in
   wire signed [9:0] m223_44;
   assign m223_44 =10'b0;

   // m223_45 = W*in
   wire signed [9:0] m223_45;
   assign m223_45 =10'b0;

   // m223_46 = W*in
   wire signed [9:0] m223_46;
   assign m223_46 =10'b0;

   // m223_47 = W*in
   wire signed [9:0] m223_47;
   assign m223_47 =10'b0;

   // m223_48 = W*in
   wire signed [9:0] m223_48;
   assign m223_48 =10'b0;

   // m223_49 = W*in
   wire signed [9:0] m223_49;
   assign m223_49 =10'b0;

   // m223_50 = W*in
   wire signed [9:0] m223_50;
   assign m223_50 =10'b0;

   // m223_51 = W*in
   wire signed [9:0] m223_51;
   assign m223_51 =10'b0;

   // m223_52 = W*in
   wire signed [9:0] m223_52;
   assign m223_52 =10'b0;

   // m223_53 = W*in
   wire signed [9:0] m223_53;
   assign m223_53 =10'b0;

   // m223_54 = W*in
   wire signed [9:0] m223_54;
   assign m223_54 =10'b0;

   // m223_55 = W*in
   wire signed [9:0] m223_55;
   assign m223_55 =10'b0;

   // m223_56 = W*in
   wire signed [9:0] m223_56;
   assign m223_56 =10'b0;

   // m223_57 = W*in
   wire signed [9:0] m223_57;
   assign m223_57 =10'b0;

   // m223_58 = W*in
   wire signed [9:0] m223_58;
   assign m223_58 =10'b0;

   // m223_59 = W*in
   wire signed [9:0] m223_59;
   assign m223_59 =10'b0;

   // m223_60 = W*in
   wire signed [9:0] m223_60;
   assign m223_60 =10'b0;

   // m223_61 = W*in
   wire signed [9:0] m223_61;
   assign m223_61 =10'b0;

   // m223_62 = W*in
   wire signed [9:0] m223_62;
   assign m223_62 =10'b0;

   // m223_63 = W*in
   wire signed [9:0] m223_63;
   assign m223_63 =10'b0;

   // m223_64 = W*in
   wire signed [9:0] m223_64;
   assign m223_64 ={ {4{in223[5]}} , in223[5:0] };

   // m223_65 = W*in
   wire signed [9:0] m223_65;
   assign m223_65 ={ {5{in223[5]}} , in223[5:1] };

   // m223_66 = W*in
   wire signed [9:0] m223_66;
   assign m223_66 =10'b0;

   // m223_67 = W*in
   wire signed [9:0] m223_67;
   assign m223_67 ={ {5{in223[5]}} , in223[5:1] };

   // m223_68 = W*in
   wire signed [9:0] m223_68;
   assign m223_68 =10'b0;

   // m223_69 = W*in
   wire signed [9:0] m223_69;
   assign m223_69 =10'b0;

   // m223_70 = W*in
   wire signed [9:0] m223_70;
   assign m223_70 ={ {5{in223[5]}} , in223[5:1] };

   // m223_71 = W*in
   wire signed [9:0] m223_71;
   assign m223_71 ={ {5{neg223[5]}} , neg223[5:1] };

   // m223_72 = W*in
   wire signed [9:0] m223_72;
   assign m223_72 ={ {5{neg223[5]}} , neg223[5:1] };

   // m223_73 = W*in
   wire signed [9:0] m223_73;
   assign m223_73 =10'b0;

   // m223_74 = W*in
   wire signed [9:0] m223_74;
   assign m223_74 =10'b0;

   // m223_75 = W*in
   wire signed [9:0] m223_75;
   assign m223_75 =10'b0;

   // m223_76 = W*in
   wire signed [9:0] m223_76;
   assign m223_76 =10'b0;

   // m223_77 = W*in
   wire signed [9:0] m223_77;
   assign m223_77 =10'b0;

   // m223_78 = W*in
   wire signed [9:0] m223_78;
   assign m223_78 =10'b0;

   // m223_79 = W*in
   wire signed [9:0] m223_79;
   assign m223_79 =10'b0;

   // m223_80 = W*in
   wire signed [9:0] m223_80;
   assign m223_80 =10'b0;

   // m223_81 = W*in
   wire signed [9:0] m223_81;
   assign m223_81 =10'b0;

   // m223_82 = W*in
   wire signed [9:0] m223_82;
   assign m223_82 =10'b0;

   // m223_83 = W*in
   wire signed [9:0] m223_83;
   assign m223_83 =10'b0;

   // m223_84 = W*in
   wire signed [9:0] m223_84;
   assign m223_84 =10'b0;

   // m223_85 = W*in
   wire signed [9:0] m223_85;
   assign m223_85 =10'b0;

   // m223_86 = W*in
   wire signed [9:0] m223_86;
   assign m223_86 =10'b0;

   // m223_87 = W*in
   wire signed [9:0] m223_87;
   assign m223_87 =10'b0;

   // m223_88 = W*in
   wire signed [9:0] m223_88;
   assign m223_88 =10'b0;

   // m223_89 = W*in
   wire signed [9:0] m223_89;
   assign m223_89 =10'b0;

   // m223_90 = W*in
   wire signed [9:0] m223_90;
   assign m223_90 =10'b0;

   // m223_91 = W*in
   wire signed [9:0] m223_91;
   assign m223_91 =10'b0;

   // m223_92 = W*in
   wire signed [9:0] m223_92;
   assign m223_92 =10'b0;

   // m223_93 = W*in
   wire signed [9:0] m223_93;
   assign m223_93 =10'b0;

   // m223_94 = W*in
   wire signed [9:0] m223_94;
   assign m223_94 =10'b0;

   // m223_95 = W*in
   wire signed [9:0] m223_95;
   assign m223_95 =10'b0;

   // m223_96 = W*in
   wire signed [9:0] m223_96;
   assign m223_96 =10'b0;

   // m223_97 = W*in
   wire signed [9:0] m223_97;
   assign m223_97 =10'b0;

   // m223_98 = W*in
   wire signed [9:0] m223_98;
   assign m223_98 =10'b0;

   // m223_99 = W*in
   wire signed [9:0] m223_99;
   assign m223_99 =10'b0;

   // m223_100 = W*in
   wire signed [9:0] m223_100;
   assign m223_100 ={ {4{in223[5]}} , in223[5:0] };

   // m223_101 = W*in
   wire signed [9:0] m223_101;
   assign m223_101 =10'b0;

   // m223_102 = W*in
   wire signed [9:0] m223_102;
   assign m223_102 =10'b0;

   // m223_103 = W*in
   wire signed [9:0] m223_103;
   assign m223_103 =10'b0;

   // m223_104 = W*in
   wire signed [9:0] m223_104;
   assign m223_104 =10'b0;

   // m223_105 = W*in
   wire signed [9:0] m223_105;
   assign m223_105 =10'b0;

   // m223_106 = W*in
   wire signed [9:0] m223_106;
   assign m223_106 =10'b0;

   // m223_107 = W*in
   wire signed [9:0] m223_107;
   assign m223_107 =10'b0;

   // m223_108 = W*in
   wire signed [9:0] m223_108;
   assign m223_108 =10'b0;

   // m223_109 = W*in
   wire signed [9:0] m223_109;
   assign m223_109 =10'b0;

   // m223_110 = W*in
   wire signed [9:0] m223_110;
   assign m223_110 =10'b0;

   // m223_111 = W*in
   wire signed [9:0] m223_111;
   assign m223_111 =10'b0;

   // m223_112 = W*in
   wire signed [9:0] m223_112;
   assign m223_112 =10'b0;

   // m223_113 = W*in
   wire signed [9:0] m223_113;
   assign m223_113 =10'b0;

   // m223_114 = W*in
   wire signed [9:0] m223_114;
   assign m223_114 ={ {5{in223[5]}} , in223[5:1] };

   // m223_115 = W*in
   wire signed [9:0] m223_115;
   assign m223_115 ={ {5{in223[5]}} , in223[5:1] };

   // m223_116 = W*in
   wire signed [9:0] m223_116;
   assign m223_116 =10'b0;

   // m223_117 = W*in
   wire signed [9:0] m223_117;
   assign m223_117 =10'b0;

   // m224_1 = W*in
   wire signed [9:0] m224_1;
   assign m224_1 =10'b0;

   // m224_2 = W*in
   wire signed [9:0] m224_2;
   assign m224_2 =10'b0;

   // m224_3 = W*in
   wire signed [9:0] m224_3;
   assign m224_3 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_4 = W*in
   wire signed [9:0] m224_4;
   assign m224_4 =10'b0;

   // m224_5 = W*in
   wire signed [9:0] m224_5;
   assign m224_5 =10'b0;

   // m224_6 = W*in
   wire signed [9:0] m224_6;
   assign m224_6 =10'b0;

   // m224_7 = W*in
   wire signed [9:0] m224_7;
   assign m224_7 =10'b0;

   // m224_8 = W*in
   wire signed [9:0] m224_8;
   assign m224_8 =10'b0;

   // m224_9 = W*in
   wire signed [9:0] m224_9;
   assign m224_9 =10'b0;

   // m224_10 = W*in
   wire signed [9:0] m224_10;
   assign m224_10 =10'b0;

   // m224_11 = W*in
   wire signed [9:0] m224_11;
   assign m224_11 =10'b0;

   // m224_12 = W*in
   wire signed [9:0] m224_12;
   assign m224_12 =10'b0;

   // m224_13 = W*in
   wire signed [9:0] m224_13;
   assign m224_13 =10'b0;

   // m224_14 = W*in
   wire signed [9:0] m224_14;
   assign m224_14 =10'b0;

   // m224_15 = W*in
   wire signed [9:0] m224_15;
   assign m224_15 =10'b0;

   // m224_16 = W*in
   wire signed [9:0] m224_16;
   assign m224_16 =10'b0;

   // m224_17 = W*in
   wire signed [9:0] m224_17;
   assign m224_17 =10'b0;

   // m224_18 = W*in
   wire signed [9:0] m224_18;
   assign m224_18 =10'b0;

   // m224_19 = W*in
   wire signed [9:0] m224_19;
   assign m224_19 =10'b0;

   // m224_20 = W*in
   wire signed [9:0] m224_20;
   assign m224_20 ={ {5{in224[5]}} , in224[5:1] };

   // m224_21 = W*in
   wire signed [9:0] m224_21;
   assign m224_21 ={ {5{neg224[5]}} , neg224[5:1] };

   // m224_22 = W*in
   wire signed [9:0] m224_22;
   assign m224_22 =10'b0;

   // m224_23 = W*in
   wire signed [9:0] m224_23;
   assign m224_23 =10'b0;

   // m224_24 = W*in
   wire signed [9:0] m224_24;
   assign m224_24 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_25 = W*in
   wire signed [9:0] m224_25;
   assign m224_25 ={ {4{in224[5]}} , in224[5:0] };

   // m224_26 = W*in
   wire signed [9:0] m224_26;
   assign m224_26 =10'b0;

   // m224_27 = W*in
   wire signed [9:0] m224_27;
   assign m224_27 =10'b0;

   // m224_28 = W*in
   wire signed [9:0] m224_28;
   assign m224_28 =10'b0;

   // m224_29 = W*in
   wire signed [9:0] m224_29;
   assign m224_29 =10'b0;

   // m224_30 = W*in
   wire signed [9:0] m224_30;
   assign m224_30 ={ {4{in224[5]}} , in224[5:0] };

   // m224_31 = W*in
   wire signed [9:0] m224_31;
   assign m224_31 ={ {5{neg224[5]}} , neg224[5:1] };

   // m224_32 = W*in
   wire signed [9:0] m224_32;
   assign m224_32 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_33 = W*in
   wire signed [9:0] m224_33;
   assign m224_33 =10'b0;

   // m224_34 = W*in
   wire signed [9:0] m224_34;
   assign m224_34 =10'b0;

   // m224_35 = W*in
   wire signed [9:0] m224_35;
   assign m224_35 =10'b0;

   // m224_36 = W*in
   wire signed [9:0] m224_36;
   assign m224_36 =10'b0;

   // m224_37 = W*in
   wire signed [9:0] m224_37;
   assign m224_37 =10'b0;

   // m224_38 = W*in
   wire signed [9:0] m224_38;
   assign m224_38 =10'b0;

   // m224_39 = W*in
   wire signed [9:0] m224_39;
   assign m224_39 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_40 = W*in
   wire signed [9:0] m224_40;
   assign m224_40 =10'b0;

   // m224_41 = W*in
   wire signed [9:0] m224_41;
   assign m224_41 =10'b0;

   // m224_42 = W*in
   wire signed [9:0] m224_42;
   assign m224_42 ={ {4{in224[5]}} , in224[5:0] };

   // m224_43 = W*in
   wire signed [9:0] m224_43;
   assign m224_43 =10'b0;

   // m224_44 = W*in
   wire signed [9:0] m224_44;
   assign m224_44 ={ {5{in224[5]}} , in224[5:1] };

   // m224_45 = W*in
   wire signed [9:0] m224_45;
   assign m224_45 =10'b0;

   // m224_46 = W*in
   wire signed [9:0] m224_46;
   assign m224_46 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_47 = W*in
   wire signed [9:0] m224_47;
   assign m224_47 =10'b0;

   // m224_48 = W*in
   wire signed [9:0] m224_48;
   assign m224_48 =10'b0;

   // m224_49 = W*in
   wire signed [9:0] m224_49;
   assign m224_49 =10'b0;

   // m224_50 = W*in
   wire signed [9:0] m224_50;
   assign m224_50 =10'b0;

   // m224_51 = W*in
   wire signed [9:0] m224_51;
   assign m224_51 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_52 = W*in
   wire signed [9:0] m224_52;
   assign m224_52 =10'b0;

   // m224_53 = W*in
   wire signed [9:0] m224_53;
   assign m224_53 ={ {4{in224[5]}} , in224[5:0] };

   // m224_54 = W*in
   wire signed [9:0] m224_54;
   assign m224_54 =10'b0;

   // m224_55 = W*in
   wire signed [9:0] m224_55;
   assign m224_55 =10'b0;

   // m224_56 = W*in
   wire signed [9:0] m224_56;
   assign m224_56 =10'b0;

   // m224_57 = W*in
   wire signed [9:0] m224_57;
   assign m224_57 =10'b0;

   // m224_58 = W*in
   wire signed [9:0] m224_58;
   assign m224_58 =10'b0;

   // m224_59 = W*in
   wire signed [9:0] m224_59;
   assign m224_59 =10'b0;

   // m224_60 = W*in
   wire signed [9:0] m224_60;
   assign m224_60 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_61 = W*in
   wire signed [9:0] m224_61;
   assign m224_61 =10'b0;

   // m224_62 = W*in
   wire signed [9:0] m224_62;
   assign m224_62 =10'b0;

   // m224_63 = W*in
   wire signed [9:0] m224_63;
   assign m224_63 =10'b0;

   // m224_64 = W*in
   wire signed [9:0] m224_64;
   assign m224_64 ={ {4{in224[5]}} , in224[5:0] };

   // m224_65 = W*in
   wire signed [9:0] m224_65;
   assign m224_65 =10'b0;

   // m224_66 = W*in
   wire signed [9:0] m224_66;
   assign m224_66 =10'b0;

   // m224_67 = W*in
   wire signed [9:0] m224_67;
   assign m224_67 =10'b0;

   // m224_68 = W*in
   wire signed [9:0] m224_68;
   assign m224_68 =10'b0;

   // m224_69 = W*in
   wire signed [9:0] m224_69;
   assign m224_69 =10'b0;

   // m224_70 = W*in
   wire signed [9:0] m224_70;
   assign m224_70 =10'b0;

   // m224_71 = W*in
   wire signed [9:0] m224_71;
   assign m224_71 =10'b0;

   // m224_72 = W*in
   wire signed [9:0] m224_72;
   assign m224_72 =10'b0;

   // m224_73 = W*in
   wire signed [9:0] m224_73;
   assign m224_73 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_74 = W*in
   wire signed [9:0] m224_74;
   assign m224_74 ={ {5{in224[5]}} , in224[5:1] };

   // m224_75 = W*in
   wire signed [9:0] m224_75;
   assign m224_75 =10'b0;

   // m224_76 = W*in
   wire signed [9:0] m224_76;
   assign m224_76 ={ {4{in224[5]}} , in224[5:0] };

   // m224_77 = W*in
   wire signed [9:0] m224_77;
   assign m224_77 ={ {4{in224[5]}} , in224[5:0] };

   // m224_78 = W*in
   wire signed [9:0] m224_78;
   assign m224_78 ={ {4{in224[5]}} , in224[5:0] };

   // m224_79 = W*in
   wire signed [9:0] m224_79;
   assign m224_79 ={ {4{in224[5]}} , in224[5:0] };

   // m224_80 = W*in
   wire signed [9:0] m224_80;
   assign m224_80 =10'b0;

   // m224_81 = W*in
   wire signed [9:0] m224_81;
   assign m224_81 =10'b0;

   // m224_82 = W*in
   wire signed [9:0] m224_82;
   assign m224_82 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_83 = W*in
   wire signed [9:0] m224_83;
   assign m224_83 =10'b0;

   // m224_84 = W*in
   wire signed [9:0] m224_84;
   assign m224_84 =10'b0;

   // m224_85 = W*in
   wire signed [9:0] m224_85;
   assign m224_85 =10'b0;

   // m224_86 = W*in
   wire signed [9:0] m224_86;
   assign m224_86 =10'b0;

   // m224_87 = W*in
   wire signed [9:0] m224_87;
   assign m224_87 =10'b0;

   // m224_88 = W*in
   wire signed [9:0] m224_88;
   assign m224_88 =10'b0;

   // m224_89 = W*in
   wire signed [9:0] m224_89;
   assign m224_89 =10'b0;

   // m224_90 = W*in
   wire signed [9:0] m224_90;
   assign m224_90 =10'b0;

   // m224_91 = W*in
   wire signed [9:0] m224_91;
   assign m224_91 =10'b0;

   // m224_92 = W*in
   wire signed [9:0] m224_92;
   assign m224_92 =10'b0;

   // m224_93 = W*in
   wire signed [9:0] m224_93;
   assign m224_93 =10'b0;

   // m224_94 = W*in
   wire signed [9:0] m224_94;
   assign m224_94 =10'b0;

   // m224_95 = W*in
   wire signed [9:0] m224_95;
   assign m224_95 =10'b0;

   // m224_96 = W*in
   wire signed [9:0] m224_96;
   assign m224_96 =10'b0;

   // m224_97 = W*in
   wire signed [9:0] m224_97;
   assign m224_97 =10'b0;

   // m224_98 = W*in
   wire signed [9:0] m224_98;
   assign m224_98 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_99 = W*in
   wire signed [9:0] m224_99;
   assign m224_99 =10'b0;

   // m224_100 = W*in
   wire signed [9:0] m224_100;
   assign m224_100 =10'b0;

   // m224_101 = W*in
   wire signed [9:0] m224_101;
   assign m224_101 =10'b0;

   // m224_102 = W*in
   wire signed [9:0] m224_102;
   assign m224_102 ={ {4{in224[5]}} , in224[5:0] };

   // m224_103 = W*in
   wire signed [9:0] m224_103;
   assign m224_103 =10'b0;

   // m224_104 = W*in
   wire signed [9:0] m224_104;
   assign m224_104 =10'b0;

   // m224_105 = W*in
   wire signed [9:0] m224_105;
   assign m224_105 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_106 = W*in
   wire signed [9:0] m224_106;
   assign m224_106 =10'b0;

   // m224_107 = W*in
   wire signed [9:0] m224_107;
   assign m224_107 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_108 = W*in
   wire signed [9:0] m224_108;
   assign m224_108 =10'b0;

   // m224_109 = W*in
   wire signed [9:0] m224_109;
   assign m224_109 =10'b0;

   // m224_110 = W*in
   wire signed [9:0] m224_110;
   assign m224_110 =10'b0;

   // m224_111 = W*in
   wire signed [9:0] m224_111;
   assign m224_111 =10'b0;

   // m224_112 = W*in
   wire signed [9:0] m224_112;
   assign m224_112 ={ {4{neg224[5]}} , neg224[5:0] };

   // m224_113 = W*in
   wire signed [9:0] m224_113;
   assign m224_113 =10'b0;

   // m224_114 = W*in
   wire signed [9:0] m224_114;
   assign m224_114 =10'b0;

   // m224_115 = W*in
   wire signed [9:0] m224_115;
   assign m224_115 =10'b0;

   // m224_116 = W*in
   wire signed [9:0] m224_116;
   assign m224_116 =10'b0;

   // m224_117 = W*in
   wire signed [9:0] m224_117;
   assign m224_117 ={ {5{in224[5]}} , in224[5:1] };

   // m225_1 = W*in
   wire signed [9:0] m225_1;
   assign m225_1 =10'b0;

   // m225_2 = W*in
   wire signed [9:0] m225_2;
   assign m225_2 =10'b0;

   // m225_3 = W*in
   wire signed [9:0] m225_3;
   assign m225_3 =10'b0;

   // m225_4 = W*in
   wire signed [9:0] m225_4;
   assign m225_4 =10'b0;

   // m225_5 = W*in
   wire signed [9:0] m225_5;
   assign m225_5 =10'b0;

   // m225_6 = W*in
   wire signed [9:0] m225_6;
   assign m225_6 =10'b0;

   // m225_7 = W*in
   wire signed [9:0] m225_7;
   assign m225_7 =10'b0;

   // m225_8 = W*in
   wire signed [9:0] m225_8;
   assign m225_8 =10'b0;

   // m225_9 = W*in
   wire signed [9:0] m225_9;
   assign m225_9 =10'b0;

   // m225_10 = W*in
   wire signed [9:0] m225_10;
   assign m225_10 ={ {5{neg225[5]}} , neg225[5:1] };

   // m225_11 = W*in
   wire signed [9:0] m225_11;
   assign m225_11 =10'b0;

   // m225_12 = W*in
   wire signed [9:0] m225_12;
   assign m225_12 =10'b0;

   // m225_13 = W*in
   wire signed [9:0] m225_13;
   assign m225_13 ={ {4{in225[5]}} , in225[5:0] };

   // m225_14 = W*in
   wire signed [9:0] m225_14;
   assign m225_14 =10'b0;

   // m225_15 = W*in
   wire signed [9:0] m225_15;
   assign m225_15 =10'b0;

   // m225_16 = W*in
   wire signed [9:0] m225_16;
   assign m225_16 =10'b0;

   // m225_17 = W*in
   wire signed [9:0] m225_17;
   assign m225_17 =10'b0;

   // m225_18 = W*in
   wire signed [9:0] m225_18;
   assign m225_18 =10'b0;

   // m225_19 = W*in
   wire signed [9:0] m225_19;
   assign m225_19 =10'b0;

   // m225_20 = W*in
   wire signed [9:0] m225_20;
   assign m225_20 ={ {4{in225[5]}} , in225[5:0] };

   // m225_21 = W*in
   wire signed [9:0] m225_21;
   assign m225_21 =10'b0;

   // m225_22 = W*in
   wire signed [9:0] m225_22;
   assign m225_22 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_23 = W*in
   wire signed [9:0] m225_23;
   assign m225_23 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_24 = W*in
   wire signed [9:0] m225_24;
   assign m225_24 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_25 = W*in
   wire signed [9:0] m225_25;
   assign m225_25 =10'b0;

   // m225_26 = W*in
   wire signed [9:0] m225_26;
   assign m225_26 =10'b0;

   // m225_27 = W*in
   wire signed [9:0] m225_27;
   assign m225_27 =10'b0;

   // m225_28 = W*in
   wire signed [9:0] m225_28;
   assign m225_28 ={ {5{in225[5]}} , in225[5:1] };

   // m225_29 = W*in
   wire signed [9:0] m225_29;
   assign m225_29 ={ {4{in225[5]}} , in225[5:0] };

   // m225_30 = W*in
   wire signed [9:0] m225_30;
   assign m225_30 ={ {4{in225[5]}} , in225[5:0] };

   // m225_31 = W*in
   wire signed [9:0] m225_31;
   assign m225_31 ={ {5{neg225[5]}} , neg225[5:1] };

   // m225_32 = W*in
   wire signed [9:0] m225_32;
   assign m225_32 =10'b0;

   // m225_33 = W*in
   wire signed [9:0] m225_33;
   assign m225_33 ={ {4{in225[5]}} , in225[5:0] };

   // m225_34 = W*in
   wire signed [9:0] m225_34;
   assign m225_34 =10'b0;

   // m225_35 = W*in
   wire signed [9:0] m225_35;
   assign m225_35 ={ {4{in225[5]}} , in225[5:0] };

   // m225_36 = W*in
   wire signed [9:0] m225_36;
   assign m225_36 ={ {4{in225[5]}} , in225[5:0] };

   // m225_37 = W*in
   wire signed [9:0] m225_37;
   assign m225_37 =10'b0;

   // m225_38 = W*in
   wire signed [9:0] m225_38;
   assign m225_38 =10'b0;

   // m225_39 = W*in
   wire signed [9:0] m225_39;
   assign m225_39 =10'b0;

   // m225_40 = W*in
   wire signed [9:0] m225_40;
   assign m225_40 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_41 = W*in
   wire signed [9:0] m225_41;
   assign m225_41 =10'b0;

   // m225_42 = W*in
   wire signed [9:0] m225_42;
   assign m225_42 =10'b0;

   // m225_43 = W*in
   wire signed [9:0] m225_43;
   assign m225_43 =10'b0;

   // m225_44 = W*in
   wire signed [9:0] m225_44;
   assign m225_44 =10'b0;

   // m225_45 = W*in
   wire signed [9:0] m225_45;
   assign m225_45 =10'b0;

   // m225_46 = W*in
   wire signed [9:0] m225_46;
   assign m225_46 =10'b0;

   // m225_47 = W*in
   wire signed [9:0] m225_47;
   assign m225_47 =10'b0;

   // m225_48 = W*in
   wire signed [9:0] m225_48;
   assign m225_48 ={ {4{in225[5]}} , in225[5:0] };

   // m225_49 = W*in
   wire signed [9:0] m225_49;
   assign m225_49 =10'b0;

   // m225_50 = W*in
   wire signed [9:0] m225_50;
   assign m225_50 =10'b0;

   // m225_51 = W*in
   wire signed [9:0] m225_51;
   assign m225_51 =10'b0;

   // m225_52 = W*in
   wire signed [9:0] m225_52;
   assign m225_52 =10'b0;

   // m225_53 = W*in
   wire signed [9:0] m225_53;
   assign m225_53 ={ {5{in225[5]}} , in225[5:1] };

   // m225_54 = W*in
   wire signed [9:0] m225_54;
   assign m225_54 =10'b0;

   // m225_55 = W*in
   wire signed [9:0] m225_55;
   assign m225_55 ={ {4{in225[5]}} , in225[5:0] };

   // m225_56 = W*in
   wire signed [9:0] m225_56;
   assign m225_56 ={ {4{in225[5]}} , in225[5:0] };

   // m225_57 = W*in
   wire signed [9:0] m225_57;
   assign m225_57 =10'b0;

   // m225_58 = W*in
   wire signed [9:0] m225_58;
   assign m225_58 =10'b0;

   // m225_59 = W*in
   wire signed [9:0] m225_59;
   assign m225_59 =10'b0;

   // m225_60 = W*in
   wire signed [9:0] m225_60;
   assign m225_60 =10'b0;

   // m225_61 = W*in
   wire signed [9:0] m225_61;
   assign m225_61 =10'b0;

   // m225_62 = W*in
   wire signed [9:0] m225_62;
   assign m225_62 =10'b0;

   // m225_63 = W*in
   wire signed [9:0] m225_63;
   assign m225_63 =10'b0;

   // m225_64 = W*in
   wire signed [9:0] m225_64;
   assign m225_64 =10'b0;

   // m225_65 = W*in
   wire signed [9:0] m225_65;
   assign m225_65 =10'b0;

   // m225_66 = W*in
   wire signed [9:0] m225_66;
   assign m225_66 ={ {5{in225[5]}} , in225[5:1] };

   // m225_67 = W*in
   wire signed [9:0] m225_67;
   assign m225_67 ={ {5{in225[5]}} , in225[5:1] };

   // m225_68 = W*in
   wire signed [9:0] m225_68;
   assign m225_68 =10'b0;

   // m225_69 = W*in
   wire signed [9:0] m225_69;
   assign m225_69 =10'b0;

   // m225_70 = W*in
   wire signed [9:0] m225_70;
   assign m225_70 ={ {4{in225[5]}} , in225[5:0] };

   // m225_71 = W*in
   wire signed [9:0] m225_71;
   assign m225_71 ={ {5{in225[5]}} , in225[5:1] };

   // m225_72 = W*in
   wire signed [9:0] m225_72;
   assign m225_72 ={ {4{in225[5]}} , in225[5:0] };

   // m225_73 = W*in
   wire signed [9:0] m225_73;
   assign m225_73 =10'b0;

   // m225_74 = W*in
   wire signed [9:0] m225_74;
   assign m225_74 ={ {4{in225[5]}} , in225[5:0] };

   // m225_75 = W*in
   wire signed [9:0] m225_75;
   assign m225_75 =10'b0;

   // m225_76 = W*in
   wire signed [9:0] m225_76;
   assign m225_76 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_77 = W*in
   wire signed [9:0] m225_77;
   assign m225_77 =10'b0;

   // m225_78 = W*in
   wire signed [9:0] m225_78;
   assign m225_78 =10'b0;

   // m225_79 = W*in
   wire signed [9:0] m225_79;
   assign m225_79 =10'b0;

   // m225_80 = W*in
   wire signed [9:0] m225_80;
   assign m225_80 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_81 = W*in
   wire signed [9:0] m225_81;
   assign m225_81 =10'b0;

   // m225_82 = W*in
   wire signed [9:0] m225_82;
   assign m225_82 =10'b0;

   // m225_83 = W*in
   wire signed [9:0] m225_83;
   assign m225_83 =10'b0;

   // m225_84 = W*in
   wire signed [9:0] m225_84;
   assign m225_84 =10'b0;

   // m225_85 = W*in
   wire signed [9:0] m225_85;
   assign m225_85 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_86 = W*in
   wire signed [9:0] m225_86;
   assign m225_86 =10'b0;

   // m225_87 = W*in
   wire signed [9:0] m225_87;
   assign m225_87 =10'b0;

   // m225_88 = W*in
   wire signed [9:0] m225_88;
   assign m225_88 =10'b0;

   // m225_89 = W*in
   wire signed [9:0] m225_89;
   assign m225_89 =10'b0;

   // m225_90 = W*in
   wire signed [9:0] m225_90;
   assign m225_90 =10'b0;

   // m225_91 = W*in
   wire signed [9:0] m225_91;
   assign m225_91 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_92 = W*in
   wire signed [9:0] m225_92;
   assign m225_92 =10'b0;

   // m225_93 = W*in
   wire signed [9:0] m225_93;
   assign m225_93 =10'b0;

   // m225_94 = W*in
   wire signed [9:0] m225_94;
   assign m225_94 ={ {4{in225[5]}} , in225[5:0] };

   // m225_95 = W*in
   wire signed [9:0] m225_95;
   assign m225_95 =10'b0;

   // m225_96 = W*in
   wire signed [9:0] m225_96;
   assign m225_96 =10'b0;

   // m225_97 = W*in
   wire signed [9:0] m225_97;
   assign m225_97 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_98 = W*in
   wire signed [9:0] m225_98;
   assign m225_98 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_99 = W*in
   wire signed [9:0] m225_99;
   assign m225_99 =10'b0;

   // m225_100 = W*in
   wire signed [9:0] m225_100;
   assign m225_100 =10'b0;

   // m225_101 = W*in
   wire signed [9:0] m225_101;
   assign m225_101 =10'b0;

   // m225_102 = W*in
   wire signed [9:0] m225_102;
   assign m225_102 ={ {4{in225[5]}} , in225[5:0] };

   // m225_103 = W*in
   wire signed [9:0] m225_103;
   assign m225_103 =10'b0;

   // m225_104 = W*in
   wire signed [9:0] m225_104;
   assign m225_104 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_105 = W*in
   wire signed [9:0] m225_105;
   assign m225_105 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_106 = W*in
   wire signed [9:0] m225_106;
   assign m225_106 ={ {4{in225[5]}} , in225[5:0] };

   // m225_107 = W*in
   wire signed [9:0] m225_107;
   assign m225_107 =10'b0;

   // m225_108 = W*in
   wire signed [9:0] m225_108;
   assign m225_108 =10'b0;

   // m225_109 = W*in
   wire signed [9:0] m225_109;
   assign m225_109 ={ {4{neg225[5]}} , neg225[5:0] };

   // m225_110 = W*in
   wire signed [9:0] m225_110;
   assign m225_110 =10'b0;

   // m225_111 = W*in
   wire signed [9:0] m225_111;
   assign m225_111 =10'b0;

   // m225_112 = W*in
   wire signed [9:0] m225_112;
   assign m225_112 =10'b0;

   // m225_113 = W*in
   wire signed [9:0] m225_113;
   assign m225_113 ={ {4{in225[5]}} , in225[5:0] };

   // m225_114 = W*in
   wire signed [9:0] m225_114;
   assign m225_114 =10'b0;

   // m225_115 = W*in
   wire signed [9:0] m225_115;
   assign m225_115 =10'b0;

   // m225_116 = W*in
   wire signed [9:0] m225_116;
   assign m225_116 =10'b0;

   // m225_117 = W*in
   wire signed [9:0] m225_117;
   assign m225_117 ={ {4{in225[5]}} , in225[5:0] };

   // m226_1 = W*in
   wire signed [9:0] m226_1;
   assign m226_1 ={ {4{in226[5]}} , in226[5:0] };

   // m226_2 = W*in
   wire signed [9:0] m226_2;
   assign m226_2 =10'b0;

   // m226_3 = W*in
   wire signed [9:0] m226_3;
   assign m226_3 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_4 = W*in
   wire signed [9:0] m226_4;
   assign m226_4 =10'b0;

   // m226_5 = W*in
   wire signed [9:0] m226_5;
   assign m226_5 ={ {4{in226[5]}} , in226[5:0] };

   // m226_6 = W*in
   wire signed [9:0] m226_6;
   assign m226_6 =10'b0;

   // m226_7 = W*in
   wire signed [9:0] m226_7;
   assign m226_7 ={ {4{in226[5]}} , in226[5:0] };

   // m226_8 = W*in
   wire signed [9:0] m226_8;
   assign m226_8 =10'b0;

   // m226_9 = W*in
   wire signed [9:0] m226_9;
   assign m226_9 =10'b0;

   // m226_10 = W*in
   wire signed [9:0] m226_10;
   assign m226_10 =10'b0;

   // m226_11 = W*in
   wire signed [9:0] m226_11;
   assign m226_11 ={ {4{in226[5]}} , in226[5:0] };

   // m226_12 = W*in
   wire signed [9:0] m226_12;
   assign m226_12 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_13 = W*in
   wire signed [9:0] m226_13;
   assign m226_13 =10'b0;

   // m226_14 = W*in
   wire signed [9:0] m226_14;
   assign m226_14 =10'b0;

   // m226_15 = W*in
   wire signed [9:0] m226_15;
   assign m226_15 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_16 = W*in
   wire signed [9:0] m226_16;
   assign m226_16 ={ {5{in226[5]}} , in226[5:1] };

   // m226_17 = W*in
   wire signed [9:0] m226_17;
   assign m226_17 =10'b0;

   // m226_18 = W*in
   wire signed [9:0] m226_18;
   assign m226_18 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_19 = W*in
   wire signed [9:0] m226_19;
   assign m226_19 ={ {4{in226[5]}} , in226[5:0] };

   // m226_20 = W*in
   wire signed [9:0] m226_20;
   assign m226_20 =10'b0;

   // m226_21 = W*in
   wire signed [9:0] m226_21;
   assign m226_21 ={ {4{in226[5]}} , in226[5:0] };

   // m226_22 = W*in
   wire signed [9:0] m226_22;
   assign m226_22 =10'b0;

   // m226_23 = W*in
   wire signed [9:0] m226_23;
   assign m226_23 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_24 = W*in
   wire signed [9:0] m226_24;
   assign m226_24 =10'b0;

   // m226_25 = W*in
   wire signed [9:0] m226_25;
   assign m226_25 =10'b0;

   // m226_26 = W*in
   wire signed [9:0] m226_26;
   assign m226_26 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_27 = W*in
   wire signed [9:0] m226_27;
   assign m226_27 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_28 = W*in
   wire signed [9:0] m226_28;
   assign m226_28 =10'b0;

   // m226_29 = W*in
   wire signed [9:0] m226_29;
   assign m226_29 =10'b0;

   // m226_30 = W*in
   wire signed [9:0] m226_30;
   assign m226_30 =10'b0;

   // m226_31 = W*in
   wire signed [9:0] m226_31;
   assign m226_31 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_32 = W*in
   wire signed [9:0] m226_32;
   assign m226_32 =10'b0;

   // m226_33 = W*in
   wire signed [9:0] m226_33;
   assign m226_33 =10'b0;

   // m226_34 = W*in
   wire signed [9:0] m226_34;
   assign m226_34 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_35 = W*in
   wire signed [9:0] m226_35;
   assign m226_35 ={ {4{in226[5]}} , in226[5:0] };

   // m226_36 = W*in
   wire signed [9:0] m226_36;
   assign m226_36 ={ {5{in226[5]}} , in226[5:1] };

   // m226_37 = W*in
   wire signed [9:0] m226_37;
   assign m226_37 =10'b0;

   // m226_38 = W*in
   wire signed [9:0] m226_38;
   assign m226_38 =10'b0;

   // m226_39 = W*in
   wire signed [9:0] m226_39;
   assign m226_39 =10'b0;

   // m226_40 = W*in
   wire signed [9:0] m226_40;
   assign m226_40 =10'b0;

   // m226_41 = W*in
   wire signed [9:0] m226_41;
   assign m226_41 =10'b0;

   // m226_42 = W*in
   wire signed [9:0] m226_42;
   assign m226_42 =10'b0;

   // m226_43 = W*in
   wire signed [9:0] m226_43;
   assign m226_43 =10'b0;

   // m226_44 = W*in
   wire signed [9:0] m226_44;
   assign m226_44 ={ {3{in226[5]}} , in226 , {1{1'b0}} };

   // m226_45 = W*in
   wire signed [9:0] m226_45;
   assign m226_45 =10'b0;

   // m226_46 = W*in
   wire signed [9:0] m226_46;
   assign m226_46 =10'b0;

   // m226_47 = W*in
   wire signed [9:0] m226_47;
   assign m226_47 =10'b0;

   // m226_48 = W*in
   wire signed [9:0] m226_48;
   assign m226_48 =10'b0;

   // m226_49 = W*in
   wire signed [9:0] m226_49;
   assign m226_49 ={ {4{in226[5]}} , in226[5:0] };

   // m226_50 = W*in
   wire signed [9:0] m226_50;
   assign m226_50 =10'b0;

   // m226_51 = W*in
   wire signed [9:0] m226_51;
   assign m226_51 =10'b0;

   // m226_52 = W*in
   wire signed [9:0] m226_52;
   assign m226_52 =10'b0;

   // m226_53 = W*in
   wire signed [9:0] m226_53;
   assign m226_53 =10'b0;

   // m226_54 = W*in
   wire signed [9:0] m226_54;
   assign m226_54 =10'b0;

   // m226_55 = W*in
   wire signed [9:0] m226_55;
   assign m226_55 =10'b0;

   // m226_56 = W*in
   wire signed [9:0] m226_56;
   assign m226_56 ={ {4{in226[5]}} , in226[5:0] };

   // m226_57 = W*in
   wire signed [9:0] m226_57;
   assign m226_57 =10'b0;

   // m226_58 = W*in
   wire signed [9:0] m226_58;
   assign m226_58 =10'b0;

   // m226_59 = W*in
   wire signed [9:0] m226_59;
   assign m226_59 =10'b0;

   // m226_60 = W*in
   wire signed [9:0] m226_60;
   assign m226_60 =10'b0;

   // m226_61 = W*in
   wire signed [9:0] m226_61;
   assign m226_61 =10'b0;

   // m226_62 = W*in
   wire signed [9:0] m226_62;
   assign m226_62 =10'b0;

   // m226_63 = W*in
   wire signed [9:0] m226_63;
   assign m226_63 ={ {4{in226[5]}} , in226[5:0] };

   // m226_64 = W*in
   wire signed [9:0] m226_64;
   assign m226_64 =10'b0;

   // m226_65 = W*in
   wire signed [9:0] m226_65;
   assign m226_65 =10'b0;

   // m226_66 = W*in
   wire signed [9:0] m226_66;
   assign m226_66 =10'b0;

   // m226_67 = W*in
   wire signed [9:0] m226_67;
   assign m226_67 ={ {4{in226[5]}} , in226[5:0] };

   // m226_68 = W*in
   wire signed [9:0] m226_68;
   assign m226_68 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_69 = W*in
   wire signed [9:0] m226_69;
   assign m226_69 =10'b0;

   // m226_70 = W*in
   wire signed [9:0] m226_70;
   assign m226_70 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_71 = W*in
   wire signed [9:0] m226_71;
   assign m226_71 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_72 = W*in
   wire signed [9:0] m226_72;
   assign m226_72 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_73 = W*in
   wire signed [9:0] m226_73;
   assign m226_73 =10'b0;

   // m226_74 = W*in
   wire signed [9:0] m226_74;
   assign m226_74 =10'b0;

   // m226_75 = W*in
   wire signed [9:0] m226_75;
   assign m226_75 =10'b0;

   // m226_76 = W*in
   wire signed [9:0] m226_76;
   assign m226_76 =10'b0;

   // m226_77 = W*in
   wire signed [9:0] m226_77;
   assign m226_77 =10'b0;

   // m226_78 = W*in
   wire signed [9:0] m226_78;
   assign m226_78 ={ {5{neg226[5]}} , neg226[5:1] };

   // m226_79 = W*in
   wire signed [9:0] m226_79;
   assign m226_79 =10'b0;

   // m226_80 = W*in
   wire signed [9:0] m226_80;
   assign m226_80 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_81 = W*in
   wire signed [9:0] m226_81;
   assign m226_81 =10'b0;

   // m226_82 = W*in
   wire signed [9:0] m226_82;
   assign m226_82 ={ {4{in226[5]}} , in226[5:0] };

   // m226_83 = W*in
   wire signed [9:0] m226_83;
   assign m226_83 =10'b0;

   // m226_84 = W*in
   wire signed [9:0] m226_84;
   assign m226_84 =10'b0;

   // m226_85 = W*in
   wire signed [9:0] m226_85;
   assign m226_85 =10'b0;

   // m226_86 = W*in
   wire signed [9:0] m226_86;
   assign m226_86 =10'b0;

   // m226_87 = W*in
   wire signed [9:0] m226_87;
   assign m226_87 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_88 = W*in
   wire signed [9:0] m226_88;
   assign m226_88 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_89 = W*in
   wire signed [9:0] m226_89;
   assign m226_89 =10'b0;

   // m226_90 = W*in
   wire signed [9:0] m226_90;
   assign m226_90 =10'b0;

   // m226_91 = W*in
   wire signed [9:0] m226_91;
   assign m226_91 ={ {4{in226[5]}} , in226[5:0] };

   // m226_92 = W*in
   wire signed [9:0] m226_92;
   assign m226_92 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_93 = W*in
   wire signed [9:0] m226_93;
   assign m226_93 ={ {3{in226[5]}} , in226 , {1{1'b0}} };

   // m226_94 = W*in
   wire signed [9:0] m226_94;
   assign m226_94 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_95 = W*in
   wire signed [9:0] m226_95;
   assign m226_95 =10'b0;

   // m226_96 = W*in
   wire signed [9:0] m226_96;
   assign m226_96 =10'b0;

   // m226_97 = W*in
   wire signed [9:0] m226_97;
   assign m226_97 ={ {4{in226[5]}} , in226[5:0] };

   // m226_98 = W*in
   wire signed [9:0] m226_98;
   assign m226_98 ={ {5{in226[5]}} , in226[5:1] };

   // m226_99 = W*in
   wire signed [9:0] m226_99;
   assign m226_99 =10'b0;

   // m226_100 = W*in
   wire signed [9:0] m226_100;
   assign m226_100 =10'b0;

   // m226_101 = W*in
   wire signed [9:0] m226_101;
   assign m226_101 =10'b0;

   // m226_102 = W*in
   wire signed [9:0] m226_102;
   assign m226_102 =10'b0;

   // m226_103 = W*in
   wire signed [9:0] m226_103;
   assign m226_103 =10'b0;

   // m226_104 = W*in
   wire signed [9:0] m226_104;
   assign m226_104 =10'b0;

   // m226_105 = W*in
   wire signed [9:0] m226_105;
   assign m226_105 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_106 = W*in
   wire signed [9:0] m226_106;
   assign m226_106 ={ {4{in226[5]}} , in226[5:0] };

   // m226_107 = W*in
   wire signed [9:0] m226_107;
   assign m226_107 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_108 = W*in
   wire signed [9:0] m226_108;
   assign m226_108 =10'b0;

   // m226_109 = W*in
   wire signed [9:0] m226_109;
   assign m226_109 =10'b0;

   // m226_110 = W*in
   wire signed [9:0] m226_110;
   assign m226_110 ={ {4{in226[5]}} , in226[5:0] };

   // m226_111 = W*in
   wire signed [9:0] m226_111;
   assign m226_111 =10'b0;

   // m226_112 = W*in
   wire signed [9:0] m226_112;
   assign m226_112 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_113 = W*in
   wire signed [9:0] m226_113;
   assign m226_113 =10'b0;

   // m226_114 = W*in
   wire signed [9:0] m226_114;
   assign m226_114 =10'b0;

   // m226_115 = W*in
   wire signed [9:0] m226_115;
   assign m226_115 =10'b0;

   // m226_116 = W*in
   wire signed [9:0] m226_116;
   assign m226_116 ={ {4{neg226[5]}} , neg226[5:0] };

   // m226_117 = W*in
   wire signed [9:0] m226_117;
   assign m226_117 =10'b0;

   // m227_1 = W*in
   wire signed [9:0] m227_1;
   assign m227_1 =10'b0;

   // m227_2 = W*in
   wire signed [9:0] m227_2;
   assign m227_2 =10'b0;

   // m227_3 = W*in
   wire signed [9:0] m227_3;
   assign m227_3 =10'b0;

   // m227_4 = W*in
   wire signed [9:0] m227_4;
   assign m227_4 =10'b0;

   // m227_5 = W*in
   wire signed [9:0] m227_5;
   assign m227_5 =10'b0;

   // m227_6 = W*in
   wire signed [9:0] m227_6;
   assign m227_6 =10'b0;

   // m227_7 = W*in
   wire signed [9:0] m227_7;
   assign m227_7 =10'b0;

   // m227_8 = W*in
   wire signed [9:0] m227_8;
   assign m227_8 =10'b0;

   // m227_9 = W*in
   wire signed [9:0] m227_9;
   assign m227_9 =10'b0;

   // m227_10 = W*in
   wire signed [9:0] m227_10;
   assign m227_10 =10'b0;

   // m227_11 = W*in
   wire signed [9:0] m227_11;
   assign m227_11 ={ {4{in227[5]}} , in227[5:0] };

   // m227_12 = W*in
   wire signed [9:0] m227_12;
   assign m227_12 =10'b0;

   // m227_13 = W*in
   wire signed [9:0] m227_13;
   assign m227_13 =10'b0;

   // m227_14 = W*in
   wire signed [9:0] m227_14;
   assign m227_14 ={ {5{neg227[5]}} , neg227[5:1] };

   // m227_15 = W*in
   wire signed [9:0] m227_15;
   assign m227_15 =10'b0;

   // m227_16 = W*in
   wire signed [9:0] m227_16;
   assign m227_16 =10'b0;

   // m227_17 = W*in
   wire signed [9:0] m227_17;
   assign m227_17 =10'b0;

   // m227_18 = W*in
   wire signed [9:0] m227_18;
   assign m227_18 =10'b0;

   // m227_19 = W*in
   wire signed [9:0] m227_19;
   assign m227_19 =10'b0;

   // m227_20 = W*in
   wire signed [9:0] m227_20;
   assign m227_20 ={ {5{in227[5]}} , in227[5:1] };

   // m227_21 = W*in
   wire signed [9:0] m227_21;
   assign m227_21 =10'b0;

   // m227_22 = W*in
   wire signed [9:0] m227_22;
   assign m227_22 =10'b0;

   // m227_23 = W*in
   wire signed [9:0] m227_23;
   assign m227_23 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_24 = W*in
   wire signed [9:0] m227_24;
   assign m227_24 =10'b0;

   // m227_25 = W*in
   wire signed [9:0] m227_25;
   assign m227_25 =10'b0;

   // m227_26 = W*in
   wire signed [9:0] m227_26;
   assign m227_26 =10'b0;

   // m227_27 = W*in
   wire signed [9:0] m227_27;
   assign m227_27 =10'b0;

   // m227_28 = W*in
   wire signed [9:0] m227_28;
   assign m227_28 ={ {4{in227[5]}} , in227[5:0] };

   // m227_29 = W*in
   wire signed [9:0] m227_29;
   assign m227_29 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_30 = W*in
   wire signed [9:0] m227_30;
   assign m227_30 =10'b0;

   // m227_31 = W*in
   wire signed [9:0] m227_31;
   assign m227_31 ={ {5{neg227[5]}} , neg227[5:1] };

   // m227_32 = W*in
   wire signed [9:0] m227_32;
   assign m227_32 =10'b0;

   // m227_33 = W*in
   wire signed [9:0] m227_33;
   assign m227_33 =10'b0;

   // m227_34 = W*in
   wire signed [9:0] m227_34;
   assign m227_34 ={ {5{neg227[5]}} , neg227[5:1] };

   // m227_35 = W*in
   wire signed [9:0] m227_35;
   assign m227_35 ={ {4{in227[5]}} , in227[5:0] };

   // m227_36 = W*in
   wire signed [9:0] m227_36;
   assign m227_36 =10'b0;

   // m227_37 = W*in
   wire signed [9:0] m227_37;
   assign m227_37 =10'b0;

   // m227_38 = W*in
   wire signed [9:0] m227_38;
   assign m227_38 ={ {4{in227[5]}} , in227[5:0] };

   // m227_39 = W*in
   wire signed [9:0] m227_39;
   assign m227_39 =10'b0;

   // m227_40 = W*in
   wire signed [9:0] m227_40;
   assign m227_40 =10'b0;

   // m227_41 = W*in
   wire signed [9:0] m227_41;
   assign m227_41 =10'b0;

   // m227_42 = W*in
   wire signed [9:0] m227_42;
   assign m227_42 =10'b0;

   // m227_43 = W*in
   wire signed [9:0] m227_43;
   assign m227_43 =10'b0;

   // m227_44 = W*in
   wire signed [9:0] m227_44;
   assign m227_44 ={ {4{in227[5]}} , in227[5:0] };

   // m227_45 = W*in
   wire signed [9:0] m227_45;
   assign m227_45 =10'b0;

   // m227_46 = W*in
   wire signed [9:0] m227_46;
   assign m227_46 =10'b0;

   // m227_47 = W*in
   wire signed [9:0] m227_47;
   assign m227_47 =10'b0;

   // m227_48 = W*in
   wire signed [9:0] m227_48;
   assign m227_48 =10'b0;

   // m227_49 = W*in
   wire signed [9:0] m227_49;
   assign m227_49 =10'b0;

   // m227_50 = W*in
   wire signed [9:0] m227_50;
   assign m227_50 =10'b0;

   // m227_51 = W*in
   wire signed [9:0] m227_51;
   assign m227_51 =10'b0;

   // m227_52 = W*in
   wire signed [9:0] m227_52;
   assign m227_52 =10'b0;

   // m227_53 = W*in
   wire signed [9:0] m227_53;
   assign m227_53 =10'b0;

   // m227_54 = W*in
   wire signed [9:0] m227_54;
   assign m227_54 ={ {4{in227[5]}} , in227[5:0] };

   // m227_55 = W*in
   wire signed [9:0] m227_55;
   assign m227_55 =10'b0;

   // m227_56 = W*in
   wire signed [9:0] m227_56;
   assign m227_56 =10'b0;

   // m227_57 = W*in
   wire signed [9:0] m227_57;
   assign m227_57 =10'b0;

   // m227_58 = W*in
   wire signed [9:0] m227_58;
   assign m227_58 =10'b0;

   // m227_59 = W*in
   wire signed [9:0] m227_59;
   assign m227_59 ={ {4{in227[5]}} , in227[5:0] };

   // m227_60 = W*in
   wire signed [9:0] m227_60;
   assign m227_60 ={ {4{in227[5]}} , in227[5:0] };

   // m227_61 = W*in
   wire signed [9:0] m227_61;
   assign m227_61 =10'b0;

   // m227_62 = W*in
   wire signed [9:0] m227_62;
   assign m227_62 =10'b0;

   // m227_63 = W*in
   wire signed [9:0] m227_63;
   assign m227_63 ={ {4{in227[5]}} , in227[5:0] };

   // m227_64 = W*in
   wire signed [9:0] m227_64;
   assign m227_64 =10'b0;

   // m227_65 = W*in
   wire signed [9:0] m227_65;
   assign m227_65 =10'b0;

   // m227_66 = W*in
   wire signed [9:0] m227_66;
   assign m227_66 =10'b0;

   // m227_67 = W*in
   wire signed [9:0] m227_67;
   assign m227_67 ={ {4{in227[5]}} , in227[5:0] };

   // m227_68 = W*in
   wire signed [9:0] m227_68;
   assign m227_68 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_69 = W*in
   wire signed [9:0] m227_69;
   assign m227_69 =10'b0;

   // m227_70 = W*in
   wire signed [9:0] m227_70;
   assign m227_70 =10'b0;

   // m227_71 = W*in
   wire signed [9:0] m227_71;
   assign m227_71 =10'b0;

   // m227_72 = W*in
   wire signed [9:0] m227_72;
   assign m227_72 =10'b0;

   // m227_73 = W*in
   wire signed [9:0] m227_73;
   assign m227_73 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_74 = W*in
   wire signed [9:0] m227_74;
   assign m227_74 =10'b0;

   // m227_75 = W*in
   wire signed [9:0] m227_75;
   assign m227_75 ={ {4{in227[5]}} , in227[5:0] };

   // m227_76 = W*in
   wire signed [9:0] m227_76;
   assign m227_76 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_77 = W*in
   wire signed [9:0] m227_77;
   assign m227_77 ={ {4{in227[5]}} , in227[5:0] };

   // m227_78 = W*in
   wire signed [9:0] m227_78;
   assign m227_78 =10'b0;

   // m227_79 = W*in
   wire signed [9:0] m227_79;
   assign m227_79 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_80 = W*in
   wire signed [9:0] m227_80;
   assign m227_80 =10'b0;

   // m227_81 = W*in
   wire signed [9:0] m227_81;
   assign m227_81 =10'b0;

   // m227_82 = W*in
   wire signed [9:0] m227_82;
   assign m227_82 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_83 = W*in
   wire signed [9:0] m227_83;
   assign m227_83 =10'b0;

   // m227_84 = W*in
   wire signed [9:0] m227_84;
   assign m227_84 =10'b0;

   // m227_85 = W*in
   wire signed [9:0] m227_85;
   assign m227_85 =10'b0;

   // m227_86 = W*in
   wire signed [9:0] m227_86;
   assign m227_86 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_87 = W*in
   wire signed [9:0] m227_87;
   assign m227_87 =10'b0;

   // m227_88 = W*in
   wire signed [9:0] m227_88;
   assign m227_88 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_89 = W*in
   wire signed [9:0] m227_89;
   assign m227_89 =10'b0;

   // m227_90 = W*in
   wire signed [9:0] m227_90;
   assign m227_90 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_91 = W*in
   wire signed [9:0] m227_91;
   assign m227_91 =10'b0;

   // m227_92 = W*in
   wire signed [9:0] m227_92;
   assign m227_92 =10'b0;

   // m227_93 = W*in
   wire signed [9:0] m227_93;
   assign m227_93 =10'b0;

   // m227_94 = W*in
   wire signed [9:0] m227_94;
   assign m227_94 =10'b0;

   // m227_95 = W*in
   wire signed [9:0] m227_95;
   assign m227_95 ={ {4{in227[5]}} , in227[5:0] };

   // m227_96 = W*in
   wire signed [9:0] m227_96;
   assign m227_96 =10'b0;

   // m227_97 = W*in
   wire signed [9:0] m227_97;
   assign m227_97 =10'b0;

   // m227_98 = W*in
   wire signed [9:0] m227_98;
   assign m227_98 =10'b0;

   // m227_99 = W*in
   wire signed [9:0] m227_99;
   assign m227_99 =10'b0;

   // m227_100 = W*in
   wire signed [9:0] m227_100;
   assign m227_100 =10'b0;

   // m227_101 = W*in
   wire signed [9:0] m227_101;
   assign m227_101 =10'b0;

   // m227_102 = W*in
   wire signed [9:0] m227_102;
   assign m227_102 =10'b0;

   // m227_103 = W*in
   wire signed [9:0] m227_103;
   assign m227_103 =10'b0;

   // m227_104 = W*in
   wire signed [9:0] m227_104;
   assign m227_104 =10'b0;

   // m227_105 = W*in
   wire signed [9:0] m227_105;
   assign m227_105 =10'b0;

   // m227_106 = W*in
   wire signed [9:0] m227_106;
   assign m227_106 =10'b0;

   // m227_107 = W*in
   wire signed [9:0] m227_107;
   assign m227_107 ={ {4{neg227[5]}} , neg227[5:0] };

   // m227_108 = W*in
   wire signed [9:0] m227_108;
   assign m227_108 =10'b0;

   // m227_109 = W*in
   wire signed [9:0] m227_109;
   assign m227_109 =10'b0;

   // m227_110 = W*in
   wire signed [9:0] m227_110;
   assign m227_110 =10'b0;

   // m227_111 = W*in
   wire signed [9:0] m227_111;
   assign m227_111 =10'b0;

   // m227_112 = W*in
   wire signed [9:0] m227_112;
   assign m227_112 =10'b0;

   // m227_113 = W*in
   wire signed [9:0] m227_113;
   assign m227_113 =10'b0;

   // m227_114 = W*in
   wire signed [9:0] m227_114;
   assign m227_114 =10'b0;

   // m227_115 = W*in
   wire signed [9:0] m227_115;
   assign m227_115 =10'b0;

   // m227_116 = W*in
   wire signed [9:0] m227_116;
   assign m227_116 =10'b0;

   // m227_117 = W*in
   wire signed [9:0] m227_117;
   assign m227_117 ={ {4{in227[5]}} , in227[5:0] };

   // m228_1 = W*in
   wire signed [9:0] m228_1;
   assign m228_1 =10'b0;

   // m228_2 = W*in
   wire signed [9:0] m228_2;
   assign m228_2 =10'b0;

   // m228_3 = W*in
   wire signed [9:0] m228_3;
   assign m228_3 =10'b0;

   // m228_4 = W*in
   wire signed [9:0] m228_4;
   assign m228_4 =10'b0;

   // m228_5 = W*in
   wire signed [9:0] m228_5;
   assign m228_5 =10'b0;

   // m228_6 = W*in
   wire signed [9:0] m228_6;
   assign m228_6 =10'b0;

   // m228_7 = W*in
   wire signed [9:0] m228_7;
   assign m228_7 =10'b0;

   // m228_8 = W*in
   wire signed [9:0] m228_8;
   assign m228_8 =10'b0;

   // m228_9 = W*in
   wire signed [9:0] m228_9;
   assign m228_9 =10'b0;

   // m228_10 = W*in
   wire signed [9:0] m228_10;
   assign m228_10 =10'b0;

   // m228_11 = W*in
   wire signed [9:0] m228_11;
   assign m228_11 =10'b0;

   // m228_12 = W*in
   wire signed [9:0] m228_12;
   assign m228_12 =10'b0;

   // m228_13 = W*in
   wire signed [9:0] m228_13;
   assign m228_13 =10'b0;

   // m228_14 = W*in
   wire signed [9:0] m228_14;
   assign m228_14 =10'b0;

   // m228_15 = W*in
   wire signed [9:0] m228_15;
   assign m228_15 =10'b0;

   // m228_16 = W*in
   wire signed [9:0] m228_16;
   assign m228_16 =10'b0;

   // m228_17 = W*in
   wire signed [9:0] m228_17;
   assign m228_17 =10'b0;

   // m228_18 = W*in
   wire signed [9:0] m228_18;
   assign m228_18 =10'b0;

   // m228_19 = W*in
   wire signed [9:0] m228_19;
   assign m228_19 =10'b0;

   // m228_20 = W*in
   wire signed [9:0] m228_20;
   assign m228_20 ={ {5{neg228[5]}} , neg228[5:1] };

   // m228_21 = W*in
   wire signed [9:0] m228_21;
   assign m228_21 =10'b0;

   // m228_22 = W*in
   wire signed [9:0] m228_22;
   assign m228_22 =10'b0;

   // m228_23 = W*in
   wire signed [9:0] m228_23;
   assign m228_23 =10'b0;

   // m228_24 = W*in
   wire signed [9:0] m228_24;
   assign m228_24 =10'b0;

   // m228_25 = W*in
   wire signed [9:0] m228_25;
   assign m228_25 ={ {5{in228[5]}} , in228[5:1] };

   // m228_26 = W*in
   wire signed [9:0] m228_26;
   assign m228_26 ={ {5{in228[5]}} , in228[5:1] };

   // m228_27 = W*in
   wire signed [9:0] m228_27;
   assign m228_27 ={ {5{in228[5]}} , in228[5:1] };

   // m228_28 = W*in
   wire signed [9:0] m228_28;
   assign m228_28 =10'b0;

   // m228_29 = W*in
   wire signed [9:0] m228_29;
   assign m228_29 =10'b0;

   // m228_30 = W*in
   wire signed [9:0] m228_30;
   assign m228_30 =10'b0;

   // m228_31 = W*in
   wire signed [9:0] m228_31;
   assign m228_31 =10'b0;

   // m228_32 = W*in
   wire signed [9:0] m228_32;
   assign m228_32 =10'b0;

   // m228_33 = W*in
   wire signed [9:0] m228_33;
   assign m228_33 =10'b0;

   // m228_34 = W*in
   wire signed [9:0] m228_34;
   assign m228_34 =10'b0;

   // m228_35 = W*in
   wire signed [9:0] m228_35;
   assign m228_35 =10'b0;

   // m228_36 = W*in
   wire signed [9:0] m228_36;
   assign m228_36 =10'b0;

   // m228_37 = W*in
   wire signed [9:0] m228_37;
   assign m228_37 =10'b0;

   // m228_38 = W*in
   wire signed [9:0] m228_38;
   assign m228_38 =10'b0;

   // m228_39 = W*in
   wire signed [9:0] m228_39;
   assign m228_39 =10'b0;

   // m228_40 = W*in
   wire signed [9:0] m228_40;
   assign m228_40 =10'b0;

   // m228_41 = W*in
   wire signed [9:0] m228_41;
   assign m228_41 =10'b0;

   // m228_42 = W*in
   wire signed [9:0] m228_42;
   assign m228_42 =10'b0;

   // m228_43 = W*in
   wire signed [9:0] m228_43;
   assign m228_43 =10'b0;

   // m228_44 = W*in
   wire signed [9:0] m228_44;
   assign m228_44 =10'b0;

   // m228_45 = W*in
   wire signed [9:0] m228_45;
   assign m228_45 =10'b0;

   // m228_46 = W*in
   wire signed [9:0] m228_46;
   assign m228_46 =10'b0;

   // m228_47 = W*in
   wire signed [9:0] m228_47;
   assign m228_47 =10'b0;

   // m228_48 = W*in
   wire signed [9:0] m228_48;
   assign m228_48 =10'b0;

   // m228_49 = W*in
   wire signed [9:0] m228_49;
   assign m228_49 =10'b0;

   // m228_50 = W*in
   wire signed [9:0] m228_50;
   assign m228_50 =10'b0;

   // m228_51 = W*in
   wire signed [9:0] m228_51;
   assign m228_51 =10'b0;

   // m228_52 = W*in
   wire signed [9:0] m228_52;
   assign m228_52 =10'b0;

   // m228_53 = W*in
   wire signed [9:0] m228_53;
   assign m228_53 =10'b0;

   // m228_54 = W*in
   wire signed [9:0] m228_54;
   assign m228_54 =10'b0;

   // m228_55 = W*in
   wire signed [9:0] m228_55;
   assign m228_55 =10'b0;

   // m228_56 = W*in
   wire signed [9:0] m228_56;
   assign m228_56 =10'b0;

   // m228_57 = W*in
   wire signed [9:0] m228_57;
   assign m228_57 =10'b0;

   // m228_58 = W*in
   wire signed [9:0] m228_58;
   assign m228_58 =10'b0;

   // m228_59 = W*in
   wire signed [9:0] m228_59;
   assign m228_59 =10'b0;

   // m228_60 = W*in
   wire signed [9:0] m228_60;
   assign m228_60 =10'b0;

   // m228_61 = W*in
   wire signed [9:0] m228_61;
   assign m228_61 =10'b0;

   // m228_62 = W*in
   wire signed [9:0] m228_62;
   assign m228_62 =10'b0;

   // m228_63 = W*in
   wire signed [9:0] m228_63;
   assign m228_63 =10'b0;

   // m228_64 = W*in
   wire signed [9:0] m228_64;
   assign m228_64 =10'b0;

   // m228_65 = W*in
   wire signed [9:0] m228_65;
   assign m228_65 =10'b0;

   // m228_66 = W*in
   wire signed [9:0] m228_66;
   assign m228_66 =10'b0;

   // m228_67 = W*in
   wire signed [9:0] m228_67;
   assign m228_67 ={ {5{neg228[5]}} , neg228[5:1] };

   // m228_68 = W*in
   wire signed [9:0] m228_68;
   assign m228_68 =10'b0;

   // m228_69 = W*in
   wire signed [9:0] m228_69;
   assign m228_69 =10'b0;

   // m228_70 = W*in
   wire signed [9:0] m228_70;
   assign m228_70 =10'b0;

   // m228_71 = W*in
   wire signed [9:0] m228_71;
   assign m228_71 ={ {5{in228[5]}} , in228[5:1] };

   // m228_72 = W*in
   wire signed [9:0] m228_72;
   assign m228_72 =10'b0;

   // m228_73 = W*in
   wire signed [9:0] m228_73;
   assign m228_73 =10'b0;

   // m228_74 = W*in
   wire signed [9:0] m228_74;
   assign m228_74 =10'b0;

   // m228_75 = W*in
   wire signed [9:0] m228_75;
   assign m228_75 =10'b0;

   // m228_76 = W*in
   wire signed [9:0] m228_76;
   assign m228_76 =10'b0;

   // m228_77 = W*in
   wire signed [9:0] m228_77;
   assign m228_77 =10'b0;

   // m228_78 = W*in
   wire signed [9:0] m228_78;
   assign m228_78 =10'b0;

   // m228_79 = W*in
   wire signed [9:0] m228_79;
   assign m228_79 =10'b0;

   // m228_80 = W*in
   wire signed [9:0] m228_80;
   assign m228_80 =10'b0;

   // m228_81 = W*in
   wire signed [9:0] m228_81;
   assign m228_81 =10'b0;

   // m228_82 = W*in
   wire signed [9:0] m228_82;
   assign m228_82 ={ {5{in228[5]}} , in228[5:1] };

   // m228_83 = W*in
   wire signed [9:0] m228_83;
   assign m228_83 =10'b0;

   // m228_84 = W*in
   wire signed [9:0] m228_84;
   assign m228_84 =10'b0;

   // m228_85 = W*in
   wire signed [9:0] m228_85;
   assign m228_85 =10'b0;

   // m228_86 = W*in
   wire signed [9:0] m228_86;
   assign m228_86 =10'b0;

   // m228_87 = W*in
   wire signed [9:0] m228_87;
   assign m228_87 =10'b0;

   // m228_88 = W*in
   wire signed [9:0] m228_88;
   assign m228_88 =10'b0;

   // m228_89 = W*in
   wire signed [9:0] m228_89;
   assign m228_89 =10'b0;

   // m228_90 = W*in
   wire signed [9:0] m228_90;
   assign m228_90 =10'b0;

   // m228_91 = W*in
   wire signed [9:0] m228_91;
   assign m228_91 =10'b0;

   // m228_92 = W*in
   wire signed [9:0] m228_92;
   assign m228_92 =10'b0;

   // m228_93 = W*in
   wire signed [9:0] m228_93;
   assign m228_93 =10'b0;

   // m228_94 = W*in
   wire signed [9:0] m228_94;
   assign m228_94 =10'b0;

   // m228_95 = W*in
   wire signed [9:0] m228_95;
   assign m228_95 =10'b0;

   // m228_96 = W*in
   wire signed [9:0] m228_96;
   assign m228_96 =10'b0;

   // m228_97 = W*in
   wire signed [9:0] m228_97;
   assign m228_97 ={ {4{in228[5]}} , in228[5:0] };

   // m228_98 = W*in
   wire signed [9:0] m228_98;
   assign m228_98 =10'b0;

   // m228_99 = W*in
   wire signed [9:0] m228_99;
   assign m228_99 =10'b0;

   // m228_100 = W*in
   wire signed [9:0] m228_100;
   assign m228_100 =10'b0;

   // m228_101 = W*in
   wire signed [9:0] m228_101;
   assign m228_101 =10'b0;

   // m228_102 = W*in
   wire signed [9:0] m228_102;
   assign m228_102 =10'b0;

   // m228_103 = W*in
   wire signed [9:0] m228_103;
   assign m228_103 =10'b0;

   // m228_104 = W*in
   wire signed [9:0] m228_104;
   assign m228_104 =10'b0;

   // m228_105 = W*in
   wire signed [9:0] m228_105;
   assign m228_105 =10'b0;

   // m228_106 = W*in
   wire signed [9:0] m228_106;
   assign m228_106 =10'b0;

   // m228_107 = W*in
   wire signed [9:0] m228_107;
   assign m228_107 =10'b0;

   // m228_108 = W*in
   wire signed [9:0] m228_108;
   assign m228_108 ={ {5{neg228[5]}} , neg228[5:1] };

   // m228_109 = W*in
   wire signed [9:0] m228_109;
   assign m228_109 =10'b0;

   // m228_110 = W*in
   wire signed [9:0] m228_110;
   assign m228_110 =10'b0;

   // m228_111 = W*in
   wire signed [9:0] m228_111;
   assign m228_111 =10'b0;

   // m228_112 = W*in
   wire signed [9:0] m228_112;
   assign m228_112 =10'b0;

   // m228_113 = W*in
   wire signed [9:0] m228_113;
   assign m228_113 =10'b0;

   // m228_114 = W*in
   wire signed [9:0] m228_114;
   assign m228_114 =10'b0;

   // m228_115 = W*in
   wire signed [9:0] m228_115;
   assign m228_115 =10'b0;

   // m228_116 = W*in
   wire signed [9:0] m228_116;
   assign m228_116 =10'b0;

   // m228_117 = W*in
   wire signed [9:0] m228_117;
   assign m228_117 =10'b0;

   // m229_1 = W*in
   wire signed [9:0] m229_1;
   assign m229_1 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_2 = W*in
   wire signed [9:0] m229_2;
   assign m229_2 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_3 = W*in
   wire signed [9:0] m229_3;
   assign m229_3 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_4 = W*in
   wire signed [9:0] m229_4;
   assign m229_4 =10'b0;

   // m229_5 = W*in
   wire signed [9:0] m229_5;
   assign m229_5 =10'b0;

   // m229_6 = W*in
   wire signed [9:0] m229_6;
   assign m229_6 ={ {5{in229[5]}} , in229[5:1] };

   // m229_7 = W*in
   wire signed [9:0] m229_7;
   assign m229_7 =10'b0;

   // m229_8 = W*in
   wire signed [9:0] m229_8;
   assign m229_8 =10'b0;

   // m229_9 = W*in
   wire signed [9:0] m229_9;
   assign m229_9 =10'b0;

   // m229_10 = W*in
   wire signed [9:0] m229_10;
   assign m229_10 =10'b0;

   // m229_11 = W*in
   wire signed [9:0] m229_11;
   assign m229_11 =10'b0;

   // m229_12 = W*in
   wire signed [9:0] m229_12;
   assign m229_12 =10'b0;

   // m229_13 = W*in
   wire signed [9:0] m229_13;
   assign m229_13 =10'b0;

   // m229_14 = W*in
   wire signed [9:0] m229_14;
   assign m229_14 =10'b0;

   // m229_15 = W*in
   wire signed [9:0] m229_15;
   assign m229_15 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_16 = W*in
   wire signed [9:0] m229_16;
   assign m229_16 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_17 = W*in
   wire signed [9:0] m229_17;
   assign m229_17 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_18 = W*in
   wire signed [9:0] m229_18;
   assign m229_18 ={ {4{in229[5]}} , in229[5:0] };

   // m229_19 = W*in
   wire signed [9:0] m229_19;
   assign m229_19 =10'b0;

   // m229_20 = W*in
   wire signed [9:0] m229_20;
   assign m229_20 =10'b0;

   // m229_21 = W*in
   wire signed [9:0] m229_21;
   assign m229_21 =10'b0;

   // m229_22 = W*in
   wire signed [9:0] m229_22;
   assign m229_22 =10'b0;

   // m229_23 = W*in
   wire signed [9:0] m229_23;
   assign m229_23 =10'b0;

   // m229_24 = W*in
   wire signed [9:0] m229_24;
   assign m229_24 =10'b0;

   // m229_25 = W*in
   wire signed [9:0] m229_25;
   assign m229_25 =10'b0;

   // m229_26 = W*in
   wire signed [9:0] m229_26;
   assign m229_26 ={ {4{in229[5]}} , in229[5:0] };

   // m229_27 = W*in
   wire signed [9:0] m229_27;
   assign m229_27 ={ {5{neg229[5]}} , neg229[5:1] };

   // m229_28 = W*in
   wire signed [9:0] m229_28;
   assign m229_28 =10'b0;

   // m229_29 = W*in
   wire signed [9:0] m229_29;
   assign m229_29 ={ {5{in229[5]}} , in229[5:1] };

   // m229_30 = W*in
   wire signed [9:0] m229_30;
   assign m229_30 =10'b0;

   // m229_31 = W*in
   wire signed [9:0] m229_31;
   assign m229_31 ={ {5{neg229[5]}} , neg229[5:1] };

   // m229_32 = W*in
   wire signed [9:0] m229_32;
   assign m229_32 =10'b0;

   // m229_33 = W*in
   wire signed [9:0] m229_33;
   assign m229_33 =10'b0;

   // m229_34 = W*in
   wire signed [9:0] m229_34;
   assign m229_34 =10'b0;

   // m229_35 = W*in
   wire signed [9:0] m229_35;
   assign m229_35 =10'b0;

   // m229_36 = W*in
   wire signed [9:0] m229_36;
   assign m229_36 =10'b0;

   // m229_37 = W*in
   wire signed [9:0] m229_37;
   assign m229_37 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_38 = W*in
   wire signed [9:0] m229_38;
   assign m229_38 ={ {3{in229[5]}} , in229 , {1{1'b0}} };

   // m229_39 = W*in
   wire signed [9:0] m229_39;
   assign m229_39 =10'b0;

   // m229_40 = W*in
   wire signed [9:0] m229_40;
   assign m229_40 =10'b0;

   // m229_41 = W*in
   wire signed [9:0] m229_41;
   assign m229_41 =10'b0;

   // m229_42 = W*in
   wire signed [9:0] m229_42;
   assign m229_42 ={ {4{in229[5]}} , in229[5:0] };

   // m229_43 = W*in
   wire signed [9:0] m229_43;
   assign m229_43 =10'b0;

   // m229_44 = W*in
   wire signed [9:0] m229_44;
   assign m229_44 ={ {4{in229[5]}} , in229[5:0] };

   // m229_45 = W*in
   wire signed [9:0] m229_45;
   assign m229_45 =10'b0;

   // m229_46 = W*in
   wire signed [9:0] m229_46;
   assign m229_46 =10'b0;

   // m229_47 = W*in
   wire signed [9:0] m229_47;
   assign m229_47 =10'b0;

   // m229_48 = W*in
   wire signed [9:0] m229_48;
   assign m229_48 =10'b0;

   // m229_49 = W*in
   wire signed [9:0] m229_49;
   assign m229_49 =10'b0;

   // m229_50 = W*in
   wire signed [9:0] m229_50;
   assign m229_50 =10'b0;

   // m229_51 = W*in
   wire signed [9:0] m229_51;
   assign m229_51 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_52 = W*in
   wire signed [9:0] m229_52;
   assign m229_52 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_53 = W*in
   wire signed [9:0] m229_53;
   assign m229_53 ={ {4{in229[5]}} , in229[5:0] };

   // m229_54 = W*in
   wire signed [9:0] m229_54;
   assign m229_54 ={ {4{in229[5]}} , in229[5:0] };

   // m229_55 = W*in
   wire signed [9:0] m229_55;
   assign m229_55 =10'b0;

   // m229_56 = W*in
   wire signed [9:0] m229_56;
   assign m229_56 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_57 = W*in
   wire signed [9:0] m229_57;
   assign m229_57 =10'b0;

   // m229_58 = W*in
   wire signed [9:0] m229_58;
   assign m229_58 =10'b0;

   // m229_59 = W*in
   wire signed [9:0] m229_59;
   assign m229_59 =10'b0;

   // m229_60 = W*in
   wire signed [9:0] m229_60;
   assign m229_60 =10'b0;

   // m229_61 = W*in
   wire signed [9:0] m229_61;
   assign m229_61 =10'b0;

   // m229_62 = W*in
   wire signed [9:0] m229_62;
   assign m229_62 =10'b0;

   // m229_63 = W*in
   wire signed [9:0] m229_63;
   assign m229_63 =10'b0;

   // m229_64 = W*in
   wire signed [9:0] m229_64;
   assign m229_64 ={ {4{in229[5]}} , in229[5:0] };

   // m229_65 = W*in
   wire signed [9:0] m229_65;
   assign m229_65 ={ {4{in229[5]}} , in229[5:0] };

   // m229_66 = W*in
   wire signed [9:0] m229_66;
   assign m229_66 ={ {4{in229[5]}} , in229[5:0] };

   // m229_67 = W*in
   wire signed [9:0] m229_67;
   assign m229_67 ={ {4{in229[5]}} , in229[5:0] };

   // m229_68 = W*in
   wire signed [9:0] m229_68;
   assign m229_68 =10'b0;

   // m229_69 = W*in
   wire signed [9:0] m229_69;
   assign m229_69 =10'b0;

   // m229_70 = W*in
   wire signed [9:0] m229_70;
   assign m229_70 ={ {5{in229[5]}} , in229[5:1] };

   // m229_71 = W*in
   wire signed [9:0] m229_71;
   assign m229_71 =10'b0;

   // m229_72 = W*in
   wire signed [9:0] m229_72;
   assign m229_72 =10'b0;

   // m229_73 = W*in
   wire signed [9:0] m229_73;
   assign m229_73 ={ {5{neg229[5]}} , neg229[5:1] };

   // m229_74 = W*in
   wire signed [9:0] m229_74;
   assign m229_74 =10'b0;

   // m229_75 = W*in
   wire signed [9:0] m229_75;
   assign m229_75 ={ {5{neg229[5]}} , neg229[5:1] };

   // m229_76 = W*in
   wire signed [9:0] m229_76;
   assign m229_76 =10'b0;

   // m229_77 = W*in
   wire signed [9:0] m229_77;
   assign m229_77 ={ {4{in229[5]}} , in229[5:0] };

   // m229_78 = W*in
   wire signed [9:0] m229_78;
   assign m229_78 =10'b0;

   // m229_79 = W*in
   wire signed [9:0] m229_79;
   assign m229_79 =10'b0;

   // m229_80 = W*in
   wire signed [9:0] m229_80;
   assign m229_80 =10'b0;

   // m229_81 = W*in
   wire signed [9:0] m229_81;
   assign m229_81 =10'b0;

   // m229_82 = W*in
   wire signed [9:0] m229_82;
   assign m229_82 =10'b0;

   // m229_83 = W*in
   wire signed [9:0] m229_83;
   assign m229_83 ={ {5{neg229[5]}} , neg229[5:1] };

   // m229_84 = W*in
   wire signed [9:0] m229_84;
   assign m229_84 =10'b0;

   // m229_85 = W*in
   wire signed [9:0] m229_85;
   assign m229_85 =10'b0;

   // m229_86 = W*in
   wire signed [9:0] m229_86;
   assign m229_86 =10'b0;

   // m229_87 = W*in
   wire signed [9:0] m229_87;
   assign m229_87 =10'b0;

   // m229_88 = W*in
   wire signed [9:0] m229_88;
   assign m229_88 =10'b0;

   // m229_89 = W*in
   wire signed [9:0] m229_89;
   assign m229_89 =10'b0;

   // m229_90 = W*in
   wire signed [9:0] m229_90;
   assign m229_90 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_91 = W*in
   wire signed [9:0] m229_91;
   assign m229_91 ={ {3{in229[5]}} , in229 , {1{1'b0}} };

   // m229_92 = W*in
   wire signed [9:0] m229_92;
   assign m229_92 =10'b0;

   // m229_93 = W*in
   wire signed [9:0] m229_93;
   assign m229_93 =10'b0;

   // m229_94 = W*in
   wire signed [9:0] m229_94;
   assign m229_94 =10'b0;

   // m229_95 = W*in
   wire signed [9:0] m229_95;
   assign m229_95 =10'b0;

   // m229_96 = W*in
   wire signed [9:0] m229_96;
   assign m229_96 =10'b0;

   // m229_97 = W*in
   wire signed [9:0] m229_97;
   assign m229_97 ={ {4{in229[5]}} , in229[5:0] };

   // m229_98 = W*in
   wire signed [9:0] m229_98;
   assign m229_98 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_99 = W*in
   wire signed [9:0] m229_99;
   assign m229_99 ={ {4{in229[5]}} , in229[5:0] };

   // m229_100 = W*in
   wire signed [9:0] m229_100;
   assign m229_100 =10'b0;

   // m229_101 = W*in
   wire signed [9:0] m229_101;
   assign m229_101 =10'b0;

   // m229_102 = W*in
   wire signed [9:0] m229_102;
   assign m229_102 =10'b0;

   // m229_103 = W*in
   wire signed [9:0] m229_103;
   assign m229_103 =10'b0;

   // m229_104 = W*in
   wire signed [9:0] m229_104;
   assign m229_104 =10'b0;

   // m229_105 = W*in
   wire signed [9:0] m229_105;
   assign m229_105 =10'b0;

   // m229_106 = W*in
   wire signed [9:0] m229_106;
   assign m229_106 =10'b0;

   // m229_107 = W*in
   wire signed [9:0] m229_107;
   assign m229_107 ={ {4{neg229[5]}} , neg229[5:0] };

   // m229_108 = W*in
   wire signed [9:0] m229_108;
   assign m229_108 =10'b0;

   // m229_109 = W*in
   wire signed [9:0] m229_109;
   assign m229_109 =10'b0;

   // m229_110 = W*in
   wire signed [9:0] m229_110;
   assign m229_110 ={ {3{in229[5]}} , in229 , {1{1'b0}} };

   // m229_111 = W*in
   wire signed [9:0] m229_111;
   assign m229_111 =10'b0;

   // m229_112 = W*in
   wire signed [9:0] m229_112;
   assign m229_112 =10'b0;

   // m229_113 = W*in
   wire signed [9:0] m229_113;
   assign m229_113 ={ {5{neg229[5]}} , neg229[5:1] };

   // m229_114 = W*in
   wire signed [9:0] m229_114;
   assign m229_114 =10'b0;

   // m229_115 = W*in
   wire signed [9:0] m229_115;
   assign m229_115 =10'b0;

   // m229_116 = W*in
   wire signed [9:0] m229_116;
   assign m229_116 =10'b0;

   // m229_117 = W*in
   wire signed [9:0] m229_117;
   assign m229_117 =10'b0;

   // m230_1 = W*in
   wire signed [9:0] m230_1;
   assign m230_1 =10'b0;

   // m230_2 = W*in
   wire signed [9:0] m230_2;
   assign m230_2 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_3 = W*in
   wire signed [9:0] m230_3;
   assign m230_3 =10'b0;

   // m230_4 = W*in
   wire signed [9:0] m230_4;
   assign m230_4 =10'b0;

   // m230_5 = W*in
   wire signed [9:0] m230_5;
   assign m230_5 =10'b0;

   // m230_6 = W*in
   wire signed [9:0] m230_6;
   assign m230_6 =10'b0;

   // m230_7 = W*in
   wire signed [9:0] m230_7;
   assign m230_7 =10'b0;

   // m230_8 = W*in
   wire signed [9:0] m230_8;
   assign m230_8 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_9 = W*in
   wire signed [9:0] m230_9;
   assign m230_9 =10'b0;

   // m230_10 = W*in
   wire signed [9:0] m230_10;
   assign m230_10 ={ {4{in230[5]}} , in230[5:0] };

   // m230_11 = W*in
   wire signed [9:0] m230_11;
   assign m230_11 =10'b0;

   // m230_12 = W*in
   wire signed [9:0] m230_12;
   assign m230_12 =10'b0;

   // m230_13 = W*in
   wire signed [9:0] m230_13;
   assign m230_13 =10'b0;

   // m230_14 = W*in
   wire signed [9:0] m230_14;
   assign m230_14 =10'b0;

   // m230_15 = W*in
   wire signed [9:0] m230_15;
   assign m230_15 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_16 = W*in
   wire signed [9:0] m230_16;
   assign m230_16 =10'b0;

   // m230_17 = W*in
   wire signed [9:0] m230_17;
   assign m230_17 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_18 = W*in
   wire signed [9:0] m230_18;
   assign m230_18 =10'b0;

   // m230_19 = W*in
   wire signed [9:0] m230_19;
   assign m230_19 =10'b0;

   // m230_20 = W*in
   wire signed [9:0] m230_20;
   assign m230_20 =10'b0;

   // m230_21 = W*in
   wire signed [9:0] m230_21;
   assign m230_21 ={ {4{in230[5]}} , in230[5:0] };

   // m230_22 = W*in
   wire signed [9:0] m230_22;
   assign m230_22 =10'b0;

   // m230_23 = W*in
   wire signed [9:0] m230_23;
   assign m230_23 ={ {5{in230[5]}} , in230[5:1] };

   // m230_24 = W*in
   wire signed [9:0] m230_24;
   assign m230_24 =10'b0;

   // m230_25 = W*in
   wire signed [9:0] m230_25;
   assign m230_25 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_26 = W*in
   wire signed [9:0] m230_26;
   assign m230_26 =10'b0;

   // m230_27 = W*in
   wire signed [9:0] m230_27;
   assign m230_27 =10'b0;

   // m230_28 = W*in
   wire signed [9:0] m230_28;
   assign m230_28 ={ {5{in230[5]}} , in230[5:1] };

   // m230_29 = W*in
   wire signed [9:0] m230_29;
   assign m230_29 =10'b0;

   // m230_30 = W*in
   wire signed [9:0] m230_30;
   assign m230_30 =10'b0;

   // m230_31 = W*in
   wire signed [9:0] m230_31;
   assign m230_31 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_32 = W*in
   wire signed [9:0] m230_32;
   assign m230_32 =10'b0;

   // m230_33 = W*in
   wire signed [9:0] m230_33;
   assign m230_33 =10'b0;

   // m230_34 = W*in
   wire signed [9:0] m230_34;
   assign m230_34 =10'b0;

   // m230_35 = W*in
   wire signed [9:0] m230_35;
   assign m230_35 =10'b0;

   // m230_36 = W*in
   wire signed [9:0] m230_36;
   assign m230_36 =10'b0;

   // m230_37 = W*in
   wire signed [9:0] m230_37;
   assign m230_37 =10'b0;

   // m230_38 = W*in
   wire signed [9:0] m230_38;
   assign m230_38 =10'b0;

   // m230_39 = W*in
   wire signed [9:0] m230_39;
   assign m230_39 =10'b0;

   // m230_40 = W*in
   wire signed [9:0] m230_40;
   assign m230_40 =10'b0;

   // m230_41 = W*in
   wire signed [9:0] m230_41;
   assign m230_41 =10'b0;

   // m230_42 = W*in
   wire signed [9:0] m230_42;
   assign m230_42 =10'b0;

   // m230_43 = W*in
   wire signed [9:0] m230_43;
   assign m230_43 =10'b0;

   // m230_44 = W*in
   wire signed [9:0] m230_44;
   assign m230_44 =10'b0;

   // m230_45 = W*in
   wire signed [9:0] m230_45;
   assign m230_45 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_46 = W*in
   wire signed [9:0] m230_46;
   assign m230_46 ={ {4{in230[5]}} , in230[5:0] };

   // m230_47 = W*in
   wire signed [9:0] m230_47;
   assign m230_47 ={ {4{in230[5]}} , in230[5:0] };

   // m230_48 = W*in
   wire signed [9:0] m230_48;
   assign m230_48 =10'b0;

   // m230_49 = W*in
   wire signed [9:0] m230_49;
   assign m230_49 =10'b0;

   // m230_50 = W*in
   wire signed [9:0] m230_50;
   assign m230_50 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_51 = W*in
   wire signed [9:0] m230_51;
   assign m230_51 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_52 = W*in
   wire signed [9:0] m230_52;
   assign m230_52 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_53 = W*in
   wire signed [9:0] m230_53;
   assign m230_53 =10'b0;

   // m230_54 = W*in
   wire signed [9:0] m230_54;
   assign m230_54 =10'b0;

   // m230_55 = W*in
   wire signed [9:0] m230_55;
   assign m230_55 =10'b0;

   // m230_56 = W*in
   wire signed [9:0] m230_56;
   assign m230_56 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_57 = W*in
   wire signed [9:0] m230_57;
   assign m230_57 =10'b0;

   // m230_58 = W*in
   wire signed [9:0] m230_58;
   assign m230_58 =10'b0;

   // m230_59 = W*in
   wire signed [9:0] m230_59;
   assign m230_59 =10'b0;

   // m230_60 = W*in
   wire signed [9:0] m230_60;
   assign m230_60 ={ {4{in230[5]}} , in230[5:0] };

   // m230_61 = W*in
   wire signed [9:0] m230_61;
   assign m230_61 =10'b0;

   // m230_62 = W*in
   wire signed [9:0] m230_62;
   assign m230_62 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_63 = W*in
   wire signed [9:0] m230_63;
   assign m230_63 ={ {3{in230[5]}} , in230 , {1{1'b0}} };

   // m230_64 = W*in
   wire signed [9:0] m230_64;
   assign m230_64 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_65 = W*in
   wire signed [9:0] m230_65;
   assign m230_65 =10'b0;

   // m230_66 = W*in
   wire signed [9:0] m230_66;
   assign m230_66 =10'b0;

   // m230_67 = W*in
   wire signed [9:0] m230_67;
   assign m230_67 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_68 = W*in
   wire signed [9:0] m230_68;
   assign m230_68 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_69 = W*in
   wire signed [9:0] m230_69;
   assign m230_69 ={ {5{in230[5]}} , in230[5:1] };

   // m230_70 = W*in
   wire signed [9:0] m230_70;
   assign m230_70 =10'b0;

   // m230_71 = W*in
   wire signed [9:0] m230_71;
   assign m230_71 ={ {5{in230[5]}} , in230[5:1] };

   // m230_72 = W*in
   wire signed [9:0] m230_72;
   assign m230_72 =10'b0;

   // m230_73 = W*in
   wire signed [9:0] m230_73;
   assign m230_73 =10'b0;

   // m230_74 = W*in
   wire signed [9:0] m230_74;
   assign m230_74 =10'b0;

   // m230_75 = W*in
   wire signed [9:0] m230_75;
   assign m230_75 =10'b0;

   // m230_76 = W*in
   wire signed [9:0] m230_76;
   assign m230_76 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_77 = W*in
   wire signed [9:0] m230_77;
   assign m230_77 =10'b0;

   // m230_78 = W*in
   wire signed [9:0] m230_78;
   assign m230_78 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_79 = W*in
   wire signed [9:0] m230_79;
   assign m230_79 =10'b0;

   // m230_80 = W*in
   wire signed [9:0] m230_80;
   assign m230_80 =10'b0;

   // m230_81 = W*in
   wire signed [9:0] m230_81;
   assign m230_81 =10'b0;

   // m230_82 = W*in
   wire signed [9:0] m230_82;
   assign m230_82 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_83 = W*in
   wire signed [9:0] m230_83;
   assign m230_83 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_84 = W*in
   wire signed [9:0] m230_84;
   assign m230_84 =10'b0;

   // m230_85 = W*in
   wire signed [9:0] m230_85;
   assign m230_85 =10'b0;

   // m230_86 = W*in
   wire signed [9:0] m230_86;
   assign m230_86 =10'b0;

   // m230_87 = W*in
   wire signed [9:0] m230_87;
   assign m230_87 =10'b0;

   // m230_88 = W*in
   wire signed [9:0] m230_88;
   assign m230_88 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_89 = W*in
   wire signed [9:0] m230_89;
   assign m230_89 ={ {4{in230[5]}} , in230[5:0] };

   // m230_90 = W*in
   wire signed [9:0] m230_90;
   assign m230_90 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_91 = W*in
   wire signed [9:0] m230_91;
   assign m230_91 =10'b0;

   // m230_92 = W*in
   wire signed [9:0] m230_92;
   assign m230_92 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_93 = W*in
   wire signed [9:0] m230_93;
   assign m230_93 =10'b0;

   // m230_94 = W*in
   wire signed [9:0] m230_94;
   assign m230_94 ={ {4{in230[5]}} , in230[5:0] };

   // m230_95 = W*in
   wire signed [9:0] m230_95;
   assign m230_95 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_96 = W*in
   wire signed [9:0] m230_96;
   assign m230_96 =10'b0;

   // m230_97 = W*in
   wire signed [9:0] m230_97;
   assign m230_97 =10'b0;

   // m230_98 = W*in
   wire signed [9:0] m230_98;
   assign m230_98 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_99 = W*in
   wire signed [9:0] m230_99;
   assign m230_99 ={ {4{in230[5]}} , in230[5:0] };

   // m230_100 = W*in
   wire signed [9:0] m230_100;
   assign m230_100 =10'b0;

   // m230_101 = W*in
   wire signed [9:0] m230_101;
   assign m230_101 =10'b0;

   // m230_102 = W*in
   wire signed [9:0] m230_102;
   assign m230_102 =10'b0;

   // m230_103 = W*in
   wire signed [9:0] m230_103;
   assign m230_103 =10'b0;

   // m230_104 = W*in
   wire signed [9:0] m230_104;
   assign m230_104 =10'b0;

   // m230_105 = W*in
   wire signed [9:0] m230_105;
   assign m230_105 =10'b0;

   // m230_106 = W*in
   wire signed [9:0] m230_106;
   assign m230_106 =10'b0;

   // m230_107 = W*in
   wire signed [9:0] m230_107;
   assign m230_107 ={ {4{neg230[5]}} , neg230[5:0] };

   // m230_108 = W*in
   wire signed [9:0] m230_108;
   assign m230_108 ={ {4{in230[5]}} , in230[5:0] };

   // m230_109 = W*in
   wire signed [9:0] m230_109;
   assign m230_109 ={ {4{in230[5]}} , in230[5:0] };

   // m230_110 = W*in
   wire signed [9:0] m230_110;
   assign m230_110 ={ {4{in230[5]}} , in230[5:0] };

   // m230_111 = W*in
   wire signed [9:0] m230_111;
   assign m230_111 =10'b0;

   // m230_112 = W*in
   wire signed [9:0] m230_112;
   assign m230_112 =10'b0;

   // m230_113 = W*in
   wire signed [9:0] m230_113;
   assign m230_113 ={ {5{neg230[5]}} , neg230[5:1] };

   // m230_114 = W*in
   wire signed [9:0] m230_114;
   assign m230_114 ={ {4{in230[5]}} , in230[5:0] };

   // m230_115 = W*in
   wire signed [9:0] m230_115;
   assign m230_115 =10'b0;

   // m230_116 = W*in
   wire signed [9:0] m230_116;
   assign m230_116 =10'b0;

   // m230_117 = W*in
   wire signed [9:0] m230_117;
   assign m230_117 ={ {4{in230[5]}} , in230[5:0] };

   // m231_1 = W*in
   wire signed [9:0] m231_1;
   assign m231_1 =10'b0;

   // m231_2 = W*in
   wire signed [9:0] m231_2;
   assign m231_2 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_3 = W*in
   wire signed [9:0] m231_3;
   assign m231_3 =10'b0;

   // m231_4 = W*in
   wire signed [9:0] m231_4;
   assign m231_4 =10'b0;

   // m231_5 = W*in
   wire signed [9:0] m231_5;
   assign m231_5 =10'b0;

   // m231_6 = W*in
   wire signed [9:0] m231_6;
   assign m231_6 =10'b0;

   // m231_7 = W*in
   wire signed [9:0] m231_7;
   assign m231_7 =10'b0;

   // m231_8 = W*in
   wire signed [9:0] m231_8;
   assign m231_8 =10'b0;

   // m231_9 = W*in
   wire signed [9:0] m231_9;
   assign m231_9 =10'b0;

   // m231_10 = W*in
   wire signed [9:0] m231_10;
   assign m231_10 =10'b0;

   // m231_11 = W*in
   wire signed [9:0] m231_11;
   assign m231_11 =10'b0;

   // m231_12 = W*in
   wire signed [9:0] m231_12;
   assign m231_12 =10'b0;

   // m231_13 = W*in
   wire signed [9:0] m231_13;
   assign m231_13 =10'b0;

   // m231_14 = W*in
   wire signed [9:0] m231_14;
   assign m231_14 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_15 = W*in
   wire signed [9:0] m231_15;
   assign m231_15 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_16 = W*in
   wire signed [9:0] m231_16;
   assign m231_16 =10'b0;

   // m231_17 = W*in
   wire signed [9:0] m231_17;
   assign m231_17 ={ {5{neg231[5]}} , neg231[5:1] };

   // m231_18 = W*in
   wire signed [9:0] m231_18;
   assign m231_18 =10'b0;

   // m231_19 = W*in
   wire signed [9:0] m231_19;
   assign m231_19 =10'b0;

   // m231_20 = W*in
   wire signed [9:0] m231_20;
   assign m231_20 ={ {4{in231[5]}} , in231[5:0] };

   // m231_21 = W*in
   wire signed [9:0] m231_21;
   assign m231_21 =10'b0;

   // m231_22 = W*in
   wire signed [9:0] m231_22;
   assign m231_22 =10'b0;

   // m231_23 = W*in
   wire signed [9:0] m231_23;
   assign m231_23 =10'b0;

   // m231_24 = W*in
   wire signed [9:0] m231_24;
   assign m231_24 =10'b0;

   // m231_25 = W*in
   wire signed [9:0] m231_25;
   assign m231_25 ={ {5{neg231[5]}} , neg231[5:1] };

   // m231_26 = W*in
   wire signed [9:0] m231_26;
   assign m231_26 =10'b0;

   // m231_27 = W*in
   wire signed [9:0] m231_27;
   assign m231_27 =10'b0;

   // m231_28 = W*in
   wire signed [9:0] m231_28;
   assign m231_28 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_29 = W*in
   wire signed [9:0] m231_29;
   assign m231_29 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_30 = W*in
   wire signed [9:0] m231_30;
   assign m231_30 ={ {4{in231[5]}} , in231[5:0] };

   // m231_31 = W*in
   wire signed [9:0] m231_31;
   assign m231_31 ={ {5{neg231[5]}} , neg231[5:1] };

   // m231_32 = W*in
   wire signed [9:0] m231_32;
   assign m231_32 =10'b0;

   // m231_33 = W*in
   wire signed [9:0] m231_33;
   assign m231_33 =10'b0;

   // m231_34 = W*in
   wire signed [9:0] m231_34;
   assign m231_34 ={ {5{neg231[5]}} , neg231[5:1] };

   // m231_35 = W*in
   wire signed [9:0] m231_35;
   assign m231_35 ={ {4{in231[5]}} , in231[5:0] };

   // m231_36 = W*in
   wire signed [9:0] m231_36;
   assign m231_36 =10'b0;

   // m231_37 = W*in
   wire signed [9:0] m231_37;
   assign m231_37 =10'b0;

   // m231_38 = W*in
   wire signed [9:0] m231_38;
   assign m231_38 ={ {4{in231[5]}} , in231[5:0] };

   // m231_39 = W*in
   wire signed [9:0] m231_39;
   assign m231_39 ={ {4{in231[5]}} , in231[5:0] };

   // m231_40 = W*in
   wire signed [9:0] m231_40;
   assign m231_40 =10'b0;

   // m231_41 = W*in
   wire signed [9:0] m231_41;
   assign m231_41 =10'b0;

   // m231_42 = W*in
   wire signed [9:0] m231_42;
   assign m231_42 =10'b0;

   // m231_43 = W*in
   wire signed [9:0] m231_43;
   assign m231_43 =10'b0;

   // m231_44 = W*in
   wire signed [9:0] m231_44;
   assign m231_44 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_45 = W*in
   wire signed [9:0] m231_45;
   assign m231_45 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_46 = W*in
   wire signed [9:0] m231_46;
   assign m231_46 ={ {3{in231[5]}} , in231 , {1{1'b0}} };

   // m231_47 = W*in
   wire signed [9:0] m231_47;
   assign m231_47 =10'b0;

   // m231_48 = W*in
   wire signed [9:0] m231_48;
   assign m231_48 =10'b0;

   // m231_49 = W*in
   wire signed [9:0] m231_49;
   assign m231_49 =10'b0;

   // m231_50 = W*in
   wire signed [9:0] m231_50;
   assign m231_50 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_51 = W*in
   wire signed [9:0] m231_51;
   assign m231_51 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_52 = W*in
   wire signed [9:0] m231_52;
   assign m231_52 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_53 = W*in
   wire signed [9:0] m231_53;
   assign m231_53 =10'b0;

   // m231_54 = W*in
   wire signed [9:0] m231_54;
   assign m231_54 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_55 = W*in
   wire signed [9:0] m231_55;
   assign m231_55 =10'b0;

   // m231_56 = W*in
   wire signed [9:0] m231_56;
   assign m231_56 =10'b0;

   // m231_57 = W*in
   wire signed [9:0] m231_57;
   assign m231_57 =10'b0;

   // m231_58 = W*in
   wire signed [9:0] m231_58;
   assign m231_58 =10'b0;

   // m231_59 = W*in
   wire signed [9:0] m231_59;
   assign m231_59 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_60 = W*in
   wire signed [9:0] m231_60;
   assign m231_60 ={ {4{in231[5]}} , in231[5:0] };

   // m231_61 = W*in
   wire signed [9:0] m231_61;
   assign m231_61 =10'b0;

   // m231_62 = W*in
   wire signed [9:0] m231_62;
   assign m231_62 =10'b0;

   // m231_63 = W*in
   wire signed [9:0] m231_63;
   assign m231_63 =10'b0;

   // m231_64 = W*in
   wire signed [9:0] m231_64;
   assign m231_64 =10'b0;

   // m231_65 = W*in
   wire signed [9:0] m231_65;
   assign m231_65 =10'b0;

   // m231_66 = W*in
   wire signed [9:0] m231_66;
   assign m231_66 ={ {4{in231[5]}} , in231[5:0] };

   // m231_67 = W*in
   wire signed [9:0] m231_67;
   assign m231_67 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_68 = W*in
   wire signed [9:0] m231_68;
   assign m231_68 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_69 = W*in
   wire signed [9:0] m231_69;
   assign m231_69 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_70 = W*in
   wire signed [9:0] m231_70;
   assign m231_70 =10'b0;

   // m231_71 = W*in
   wire signed [9:0] m231_71;
   assign m231_71 ={ {5{in231[5]}} , in231[5:1] };

   // m231_72 = W*in
   wire signed [9:0] m231_72;
   assign m231_72 =10'b0;

   // m231_73 = W*in
   wire signed [9:0] m231_73;
   assign m231_73 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_74 = W*in
   wire signed [9:0] m231_74;
   assign m231_74 ={ {4{in231[5]}} , in231[5:0] };

   // m231_75 = W*in
   wire signed [9:0] m231_75;
   assign m231_75 ={ {4{in231[5]}} , in231[5:0] };

   // m231_76 = W*in
   wire signed [9:0] m231_76;
   assign m231_76 =10'b0;

   // m231_77 = W*in
   wire signed [9:0] m231_77;
   assign m231_77 =10'b0;

   // m231_78 = W*in
   wire signed [9:0] m231_78;
   assign m231_78 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_79 = W*in
   wire signed [9:0] m231_79;
   assign m231_79 =10'b0;

   // m231_80 = W*in
   wire signed [9:0] m231_80;
   assign m231_80 =10'b0;

   // m231_81 = W*in
   wire signed [9:0] m231_81;
   assign m231_81 ={ {5{in231[5]}} , in231[5:1] };

   // m231_82 = W*in
   wire signed [9:0] m231_82;
   assign m231_82 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_83 = W*in
   wire signed [9:0] m231_83;
   assign m231_83 ={ {5{neg231[5]}} , neg231[5:1] };

   // m231_84 = W*in
   wire signed [9:0] m231_84;
   assign m231_84 =10'b0;

   // m231_85 = W*in
   wire signed [9:0] m231_85;
   assign m231_85 =10'b0;

   // m231_86 = W*in
   wire signed [9:0] m231_86;
   assign m231_86 =10'b0;

   // m231_87 = W*in
   wire signed [9:0] m231_87;
   assign m231_87 =10'b0;

   // m231_88 = W*in
   wire signed [9:0] m231_88;
   assign m231_88 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_89 = W*in
   wire signed [9:0] m231_89;
   assign m231_89 =10'b0;

   // m231_90 = W*in
   wire signed [9:0] m231_90;
   assign m231_90 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_91 = W*in
   wire signed [9:0] m231_91;
   assign m231_91 ={ {4{in231[5]}} , in231[5:0] };

   // m231_92 = W*in
   wire signed [9:0] m231_92;
   assign m231_92 =10'b0;

   // m231_93 = W*in
   wire signed [9:0] m231_93;
   assign m231_93 =10'b0;

   // m231_94 = W*in
   wire signed [9:0] m231_94;
   assign m231_94 ={ {4{in231[5]}} , in231[5:0] };

   // m231_95 = W*in
   wire signed [9:0] m231_95;
   assign m231_95 =10'b0;

   // m231_96 = W*in
   wire signed [9:0] m231_96;
   assign m231_96 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_97 = W*in
   wire signed [9:0] m231_97;
   assign m231_97 =10'b0;

   // m231_98 = W*in
   wire signed [9:0] m231_98;
   assign m231_98 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_99 = W*in
   wire signed [9:0] m231_99;
   assign m231_99 =10'b0;

   // m231_100 = W*in
   wire signed [9:0] m231_100;
   assign m231_100 =10'b0;

   // m231_101 = W*in
   wire signed [9:0] m231_101;
   assign m231_101 =10'b0;

   // m231_102 = W*in
   wire signed [9:0] m231_102;
   assign m231_102 =10'b0;

   // m231_103 = W*in
   wire signed [9:0] m231_103;
   assign m231_103 ={ {4{in231[5]}} , in231[5:0] };

   // m231_104 = W*in
   wire signed [9:0] m231_104;
   assign m231_104 =10'b0;

   // m231_105 = W*in
   wire signed [9:0] m231_105;
   assign m231_105 =10'b0;

   // m231_106 = W*in
   wire signed [9:0] m231_106;
   assign m231_106 =10'b0;

   // m231_107 = W*in
   wire signed [9:0] m231_107;
   assign m231_107 =10'b0;

   // m231_108 = W*in
   wire signed [9:0] m231_108;
   assign m231_108 =10'b0;

   // m231_109 = W*in
   wire signed [9:0] m231_109;
   assign m231_109 ={ {4{in231[5]}} , in231[5:0] };

   // m231_110 = W*in
   wire signed [9:0] m231_110;
   assign m231_110 ={ {5{in231[5]}} , in231[5:1] };

   // m231_111 = W*in
   wire signed [9:0] m231_111;
   assign m231_111 ={ {4{neg231[5]}} , neg231[5:0] };

   // m231_112 = W*in
   wire signed [9:0] m231_112;
   assign m231_112 =10'b0;

   // m231_113 = W*in
   wire signed [9:0] m231_113;
   assign m231_113 =10'b0;

   // m231_114 = W*in
   wire signed [9:0] m231_114;
   assign m231_114 =10'b0;

   // m231_115 = W*in
   wire signed [9:0] m231_115;
   assign m231_115 ={ {4{in231[5]}} , in231[5:0] };

   // m231_116 = W*in
   wire signed [9:0] m231_116;
   assign m231_116 =10'b0;

   // m231_117 = W*in
   wire signed [9:0] m231_117;
   assign m231_117 ={ {4{in231[5]}} , in231[5:0] };

   // m232_1 = W*in
   wire signed [9:0] m232_1;
   assign m232_1 =10'b0;

   // m232_2 = W*in
   wire signed [9:0] m232_2;
   assign m232_2 =10'b0;

   // m232_3 = W*in
   wire signed [9:0] m232_3;
   assign m232_3 ={ {4{in232[5]}} , in232[5:0] };

   // m232_4 = W*in
   wire signed [9:0] m232_4;
   assign m232_4 =10'b0;

   // m232_5 = W*in
   wire signed [9:0] m232_5;
   assign m232_5 =10'b0;

   // m232_6 = W*in
   wire signed [9:0] m232_6;
   assign m232_6 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_7 = W*in
   wire signed [9:0] m232_7;
   assign m232_7 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_8 = W*in
   wire signed [9:0] m232_8;
   assign m232_8 =10'b0;

   // m232_9 = W*in
   wire signed [9:0] m232_9;
   assign m232_9 =10'b0;

   // m232_10 = W*in
   wire signed [9:0] m232_10;
   assign m232_10 =10'b0;

   // m232_11 = W*in
   wire signed [9:0] m232_11;
   assign m232_11 =10'b0;

   // m232_12 = W*in
   wire signed [9:0] m232_12;
   assign m232_12 ={ {4{in232[5]}} , in232[5:0] };

   // m232_13 = W*in
   wire signed [9:0] m232_13;
   assign m232_13 =10'b0;

   // m232_14 = W*in
   wire signed [9:0] m232_14;
   assign m232_14 =10'b0;

   // m232_15 = W*in
   wire signed [9:0] m232_15;
   assign m232_15 ={ {4{in232[5]}} , in232[5:0] };

   // m232_16 = W*in
   wire signed [9:0] m232_16;
   assign m232_16 =10'b0;

   // m232_17 = W*in
   wire signed [9:0] m232_17;
   assign m232_17 ={ {5{in232[5]}} , in232[5:1] };

   // m232_18 = W*in
   wire signed [9:0] m232_18;
   assign m232_18 =10'b0;

   // m232_19 = W*in
   wire signed [9:0] m232_19;
   assign m232_19 =10'b0;

   // m232_20 = W*in
   wire signed [9:0] m232_20;
   assign m232_20 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_21 = W*in
   wire signed [9:0] m232_21;
   assign m232_21 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_22 = W*in
   wire signed [9:0] m232_22;
   assign m232_22 =10'b0;

   // m232_23 = W*in
   wire signed [9:0] m232_23;
   assign m232_23 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_24 = W*in
   wire signed [9:0] m232_24;
   assign m232_24 =10'b0;

   // m232_25 = W*in
   wire signed [9:0] m232_25;
   assign m232_25 =10'b0;

   // m232_26 = W*in
   wire signed [9:0] m232_26;
   assign m232_26 =10'b0;

   // m232_27 = W*in
   wire signed [9:0] m232_27;
   assign m232_27 ={ {5{in232[5]}} , in232[5:1] };

   // m232_28 = W*in
   wire signed [9:0] m232_28;
   assign m232_28 ={ {5{in232[5]}} , in232[5:1] };

   // m232_29 = W*in
   wire signed [9:0] m232_29;
   assign m232_29 =10'b0;

   // m232_30 = W*in
   wire signed [9:0] m232_30;
   assign m232_30 =10'b0;

   // m232_31 = W*in
   wire signed [9:0] m232_31;
   assign m232_31 ={ {5{in232[5]}} , in232[5:1] };

   // m232_32 = W*in
   wire signed [9:0] m232_32;
   assign m232_32 =10'b0;

   // m232_33 = W*in
   wire signed [9:0] m232_33;
   assign m232_33 =10'b0;

   // m232_34 = W*in
   wire signed [9:0] m232_34;
   assign m232_34 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_35 = W*in
   wire signed [9:0] m232_35;
   assign m232_35 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_36 = W*in
   wire signed [9:0] m232_36;
   assign m232_36 =10'b0;

   // m232_37 = W*in
   wire signed [9:0] m232_37;
   assign m232_37 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_38 = W*in
   wire signed [9:0] m232_38;
   assign m232_38 ={ {4{in232[5]}} , in232[5:0] };

   // m232_39 = W*in
   wire signed [9:0] m232_39;
   assign m232_39 =10'b0;

   // m232_40 = W*in
   wire signed [9:0] m232_40;
   assign m232_40 =10'b0;

   // m232_41 = W*in
   wire signed [9:0] m232_41;
   assign m232_41 =10'b0;

   // m232_42 = W*in
   wire signed [9:0] m232_42;
   assign m232_42 =10'b0;

   // m232_43 = W*in
   wire signed [9:0] m232_43;
   assign m232_43 ={ {4{in232[5]}} , in232[5:0] };

   // m232_44 = W*in
   wire signed [9:0] m232_44;
   assign m232_44 =10'b0;

   // m232_45 = W*in
   wire signed [9:0] m232_45;
   assign m232_45 =10'b0;

   // m232_46 = W*in
   wire signed [9:0] m232_46;
   assign m232_46 =10'b0;

   // m232_47 = W*in
   wire signed [9:0] m232_47;
   assign m232_47 =10'b0;

   // m232_48 = W*in
   wire signed [9:0] m232_48;
   assign m232_48 =10'b0;

   // m232_49 = W*in
   wire signed [9:0] m232_49;
   assign m232_49 =10'b0;

   // m232_50 = W*in
   wire signed [9:0] m232_50;
   assign m232_50 =10'b0;

   // m232_51 = W*in
   wire signed [9:0] m232_51;
   assign m232_51 =10'b0;

   // m232_52 = W*in
   wire signed [9:0] m232_52;
   assign m232_52 =10'b0;

   // m232_53 = W*in
   wire signed [9:0] m232_53;
   assign m232_53 =10'b0;

   // m232_54 = W*in
   wire signed [9:0] m232_54;
   assign m232_54 =10'b0;

   // m232_55 = W*in
   wire signed [9:0] m232_55;
   assign m232_55 =10'b0;

   // m232_56 = W*in
   wire signed [9:0] m232_56;
   assign m232_56 =10'b0;

   // m232_57 = W*in
   wire signed [9:0] m232_57;
   assign m232_57 =10'b0;

   // m232_58 = W*in
   wire signed [9:0] m232_58;
   assign m232_58 =10'b0;

   // m232_59 = W*in
   wire signed [9:0] m232_59;
   assign m232_59 ={ {4{in232[5]}} , in232[5:0] };

   // m232_60 = W*in
   wire signed [9:0] m232_60;
   assign m232_60 =10'b0;

   // m232_61 = W*in
   wire signed [9:0] m232_61;
   assign m232_61 =10'b0;

   // m232_62 = W*in
   wire signed [9:0] m232_62;
   assign m232_62 =10'b0;

   // m232_63 = W*in
   wire signed [9:0] m232_63;
   assign m232_63 =10'b0;

   // m232_64 = W*in
   wire signed [9:0] m232_64;
   assign m232_64 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_65 = W*in
   wire signed [9:0] m232_65;
   assign m232_65 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_66 = W*in
   wire signed [9:0] m232_66;
   assign m232_66 =10'b0;

   // m232_67 = W*in
   wire signed [9:0] m232_67;
   assign m232_67 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_68 = W*in
   wire signed [9:0] m232_68;
   assign m232_68 =10'b0;

   // m232_69 = W*in
   wire signed [9:0] m232_69;
   assign m232_69 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_70 = W*in
   wire signed [9:0] m232_70;
   assign m232_70 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_71 = W*in
   wire signed [9:0] m232_71;
   assign m232_71 ={ {4{in232[5]}} , in232[5:0] };

   // m232_72 = W*in
   wire signed [9:0] m232_72;
   assign m232_72 =10'b0;

   // m232_73 = W*in
   wire signed [9:0] m232_73;
   assign m232_73 =10'b0;

   // m232_74 = W*in
   wire signed [9:0] m232_74;
   assign m232_74 =10'b0;

   // m232_75 = W*in
   wire signed [9:0] m232_75;
   assign m232_75 ={ {5{in232[5]}} , in232[5:1] };

   // m232_76 = W*in
   wire signed [9:0] m232_76;
   assign m232_76 =10'b0;

   // m232_77 = W*in
   wire signed [9:0] m232_77;
   assign m232_77 =10'b0;

   // m232_78 = W*in
   wire signed [9:0] m232_78;
   assign m232_78 =10'b0;

   // m232_79 = W*in
   wire signed [9:0] m232_79;
   assign m232_79 =10'b0;

   // m232_80 = W*in
   wire signed [9:0] m232_80;
   assign m232_80 =10'b0;

   // m232_81 = W*in
   wire signed [9:0] m232_81;
   assign m232_81 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_82 = W*in
   wire signed [9:0] m232_82;
   assign m232_82 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_83 = W*in
   wire signed [9:0] m232_83;
   assign m232_83 ={ {5{in232[5]}} , in232[5:1] };

   // m232_84 = W*in
   wire signed [9:0] m232_84;
   assign m232_84 =10'b0;

   // m232_85 = W*in
   wire signed [9:0] m232_85;
   assign m232_85 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_86 = W*in
   wire signed [9:0] m232_86;
   assign m232_86 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_87 = W*in
   wire signed [9:0] m232_87;
   assign m232_87 =10'b0;

   // m232_88 = W*in
   wire signed [9:0] m232_88;
   assign m232_88 ={ {4{in232[5]}} , in232[5:0] };

   // m232_89 = W*in
   wire signed [9:0] m232_89;
   assign m232_89 =10'b0;

   // m232_90 = W*in
   wire signed [9:0] m232_90;
   assign m232_90 =10'b0;

   // m232_91 = W*in
   wire signed [9:0] m232_91;
   assign m232_91 =10'b0;

   // m232_92 = W*in
   wire signed [9:0] m232_92;
   assign m232_92 ={ {4{in232[5]}} , in232[5:0] };

   // m232_93 = W*in
   wire signed [9:0] m232_93;
   assign m232_93 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_94 = W*in
   wire signed [9:0] m232_94;
   assign m232_94 =10'b0;

   // m232_95 = W*in
   wire signed [9:0] m232_95;
   assign m232_95 =10'b0;

   // m232_96 = W*in
   wire signed [9:0] m232_96;
   assign m232_96 =10'b0;

   // m232_97 = W*in
   wire signed [9:0] m232_97;
   assign m232_97 =10'b0;

   // m232_98 = W*in
   wire signed [9:0] m232_98;
   assign m232_98 =10'b0;

   // m232_99 = W*in
   wire signed [9:0] m232_99;
   assign m232_99 ={ {4{neg232[5]}} , neg232[5:0] };

   // m232_100 = W*in
   wire signed [9:0] m232_100;
   assign m232_100 =10'b0;

   // m232_101 = W*in
   wire signed [9:0] m232_101;
   assign m232_101 ={ {4{in232[5]}} , in232[5:0] };

   // m232_102 = W*in
   wire signed [9:0] m232_102;
   assign m232_102 =10'b0;

   // m232_103 = W*in
   wire signed [9:0] m232_103;
   assign m232_103 ={ {4{in232[5]}} , in232[5:0] };

   // m232_104 = W*in
   wire signed [9:0] m232_104;
   assign m232_104 ={ {4{in232[5]}} , in232[5:0] };

   // m232_105 = W*in
   wire signed [9:0] m232_105;
   assign m232_105 =10'b0;

   // m232_106 = W*in
   wire signed [9:0] m232_106;
   assign m232_106 =10'b0;

   // m232_107 = W*in
   wire signed [9:0] m232_107;
   assign m232_107 =10'b0;

   // m232_108 = W*in
   wire signed [9:0] m232_108;
   assign m232_108 =10'b0;

   // m232_109 = W*in
   wire signed [9:0] m232_109;
   assign m232_109 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_110 = W*in
   wire signed [9:0] m232_110;
   assign m232_110 =10'b0;

   // m232_111 = W*in
   wire signed [9:0] m232_111;
   assign m232_111 =10'b0;

   // m232_112 = W*in
   wire signed [9:0] m232_112;
   assign m232_112 =10'b0;

   // m232_113 = W*in
   wire signed [9:0] m232_113;
   assign m232_113 =10'b0;

   // m232_114 = W*in
   wire signed [9:0] m232_114;
   assign m232_114 ={ {5{neg232[5]}} , neg232[5:1] };

   // m232_115 = W*in
   wire signed [9:0] m232_115;
   assign m232_115 =10'b0;

   // m232_116 = W*in
   wire signed [9:0] m232_116;
   assign m232_116 =10'b0;

   // m232_117 = W*in
   wire signed [9:0] m232_117;
   assign m232_117 =10'b0;

   // m233_1 = W*in
   wire signed [9:0] m233_1;
   assign m233_1 =10'b0;

   // m233_2 = W*in
   wire signed [9:0] m233_2;
   assign m233_2 =10'b0;

   // m233_3 = W*in
   wire signed [9:0] m233_3;
   assign m233_3 =10'b0;

   // m233_4 = W*in
   wire signed [9:0] m233_4;
   assign m233_4 =10'b0;

   // m233_5 = W*in
   wire signed [9:0] m233_5;
   assign m233_5 =10'b0;

   // m233_6 = W*in
   wire signed [9:0] m233_6;
   assign m233_6 =10'b0;

   // m233_7 = W*in
   wire signed [9:0] m233_7;
   assign m233_7 =10'b0;

   // m233_8 = W*in
   wire signed [9:0] m233_8;
   assign m233_8 =10'b0;

   // m233_9 = W*in
   wire signed [9:0] m233_9;
   assign m233_9 =10'b0;

   // m233_10 = W*in
   wire signed [9:0] m233_10;
   assign m233_10 =10'b0;

   // m233_11 = W*in
   wire signed [9:0] m233_11;
   assign m233_11 =10'b0;

   // m233_12 = W*in
   wire signed [9:0] m233_12;
   assign m233_12 =10'b0;

   // m233_13 = W*in
   wire signed [9:0] m233_13;
   assign m233_13 =10'b0;

   // m233_14 = W*in
   wire signed [9:0] m233_14;
   assign m233_14 =10'b0;

   // m233_15 = W*in
   wire signed [9:0] m233_15;
   assign m233_15 =10'b0;

   // m233_16 = W*in
   wire signed [9:0] m233_16;
   assign m233_16 =10'b0;

   // m233_17 = W*in
   wire signed [9:0] m233_17;
   assign m233_17 =10'b0;

   // m233_18 = W*in
   wire signed [9:0] m233_18;
   assign m233_18 =10'b0;

   // m233_19 = W*in
   wire signed [9:0] m233_19;
   assign m233_19 =10'b0;

   // m233_20 = W*in
   wire signed [9:0] m233_20;
   assign m233_20 =10'b0;

   // m233_21 = W*in
   wire signed [9:0] m233_21;
   assign m233_21 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_22 = W*in
   wire signed [9:0] m233_22;
   assign m233_22 =10'b0;

   // m233_23 = W*in
   wire signed [9:0] m233_23;
   assign m233_23 =10'b0;

   // m233_24 = W*in
   wire signed [9:0] m233_24;
   assign m233_24 =10'b0;

   // m233_25 = W*in
   wire signed [9:0] m233_25;
   assign m233_25 ={ {5{in233[5]}} , in233[5:1] };

   // m233_26 = W*in
   wire signed [9:0] m233_26;
   assign m233_26 =10'b0;

   // m233_27 = W*in
   wire signed [9:0] m233_27;
   assign m233_27 ={ {5{in233[5]}} , in233[5:1] };

   // m233_28 = W*in
   wire signed [9:0] m233_28;
   assign m233_28 ={ {4{in233[5]}} , in233[5:0] };

   // m233_29 = W*in
   wire signed [9:0] m233_29;
   assign m233_29 =10'b0;

   // m233_30 = W*in
   wire signed [9:0] m233_30;
   assign m233_30 =10'b0;

   // m233_31 = W*in
   wire signed [9:0] m233_31;
   assign m233_31 =10'b0;

   // m233_32 = W*in
   wire signed [9:0] m233_32;
   assign m233_32 =10'b0;

   // m233_33 = W*in
   wire signed [9:0] m233_33;
   assign m233_33 =10'b0;

   // m233_34 = W*in
   wire signed [9:0] m233_34;
   assign m233_34 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_35 = W*in
   wire signed [9:0] m233_35;
   assign m233_35 =10'b0;

   // m233_36 = W*in
   wire signed [9:0] m233_36;
   assign m233_36 =10'b0;

   // m233_37 = W*in
   wire signed [9:0] m233_37;
   assign m233_37 =10'b0;

   // m233_38 = W*in
   wire signed [9:0] m233_38;
   assign m233_38 =10'b0;

   // m233_39 = W*in
   wire signed [9:0] m233_39;
   assign m233_39 =10'b0;

   // m233_40 = W*in
   wire signed [9:0] m233_40;
   assign m233_40 =10'b0;

   // m233_41 = W*in
   wire signed [9:0] m233_41;
   assign m233_41 =10'b0;

   // m233_42 = W*in
   wire signed [9:0] m233_42;
   assign m233_42 =10'b0;

   // m233_43 = W*in
   wire signed [9:0] m233_43;
   assign m233_43 ={ {4{in233[5]}} , in233[5:0] };

   // m233_44 = W*in
   wire signed [9:0] m233_44;
   assign m233_44 =10'b0;

   // m233_45 = W*in
   wire signed [9:0] m233_45;
   assign m233_45 =10'b0;

   // m233_46 = W*in
   wire signed [9:0] m233_46;
   assign m233_46 =10'b0;

   // m233_47 = W*in
   wire signed [9:0] m233_47;
   assign m233_47 =10'b0;

   // m233_48 = W*in
   wire signed [9:0] m233_48;
   assign m233_48 ={ {4{in233[5]}} , in233[5:0] };

   // m233_49 = W*in
   wire signed [9:0] m233_49;
   assign m233_49 =10'b0;

   // m233_50 = W*in
   wire signed [9:0] m233_50;
   assign m233_50 =10'b0;

   // m233_51 = W*in
   wire signed [9:0] m233_51;
   assign m233_51 =10'b0;

   // m233_52 = W*in
   wire signed [9:0] m233_52;
   assign m233_52 =10'b0;

   // m233_53 = W*in
   wire signed [9:0] m233_53;
   assign m233_53 =10'b0;

   // m233_54 = W*in
   wire signed [9:0] m233_54;
   assign m233_54 =10'b0;

   // m233_55 = W*in
   wire signed [9:0] m233_55;
   assign m233_55 =10'b0;

   // m233_56 = W*in
   wire signed [9:0] m233_56;
   assign m233_56 =10'b0;

   // m233_57 = W*in
   wire signed [9:0] m233_57;
   assign m233_57 =10'b0;

   // m233_58 = W*in
   wire signed [9:0] m233_58;
   assign m233_58 =10'b0;

   // m233_59 = W*in
   wire signed [9:0] m233_59;
   assign m233_59 =10'b0;

   // m233_60 = W*in
   wire signed [9:0] m233_60;
   assign m233_60 =10'b0;

   // m233_61 = W*in
   wire signed [9:0] m233_61;
   assign m233_61 =10'b0;

   // m233_62 = W*in
   wire signed [9:0] m233_62;
   assign m233_62 =10'b0;

   // m233_63 = W*in
   wire signed [9:0] m233_63;
   assign m233_63 =10'b0;

   // m233_64 = W*in
   wire signed [9:0] m233_64;
   assign m233_64 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_65 = W*in
   wire signed [9:0] m233_65;
   assign m233_65 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_66 = W*in
   wire signed [9:0] m233_66;
   assign m233_66 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_67 = W*in
   wire signed [9:0] m233_67;
   assign m233_67 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_68 = W*in
   wire signed [9:0] m233_68;
   assign m233_68 =10'b0;

   // m233_69 = W*in
   wire signed [9:0] m233_69;
   assign m233_69 =10'b0;

   // m233_70 = W*in
   wire signed [9:0] m233_70;
   assign m233_70 =10'b0;

   // m233_71 = W*in
   wire signed [9:0] m233_71;
   assign m233_71 ={ {5{in233[5]}} , in233[5:1] };

   // m233_72 = W*in
   wire signed [9:0] m233_72;
   assign m233_72 ={ {5{in233[5]}} , in233[5:1] };

   // m233_73 = W*in
   wire signed [9:0] m233_73;
   assign m233_73 =10'b0;

   // m233_74 = W*in
   wire signed [9:0] m233_74;
   assign m233_74 =10'b0;

   // m233_75 = W*in
   wire signed [9:0] m233_75;
   assign m233_75 =10'b0;

   // m233_76 = W*in
   wire signed [9:0] m233_76;
   assign m233_76 =10'b0;

   // m233_77 = W*in
   wire signed [9:0] m233_77;
   assign m233_77 =10'b0;

   // m233_78 = W*in
   wire signed [9:0] m233_78;
   assign m233_78 ={ {5{in233[5]}} , in233[5:1] };

   // m233_79 = W*in
   wire signed [9:0] m233_79;
   assign m233_79 =10'b0;

   // m233_80 = W*in
   wire signed [9:0] m233_80;
   assign m233_80 =10'b0;

   // m233_81 = W*in
   wire signed [9:0] m233_81;
   assign m233_81 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_82 = W*in
   wire signed [9:0] m233_82;
   assign m233_82 =10'b0;

   // m233_83 = W*in
   wire signed [9:0] m233_83;
   assign m233_83 =10'b0;

   // m233_84 = W*in
   wire signed [9:0] m233_84;
   assign m233_84 =10'b0;

   // m233_85 = W*in
   wire signed [9:0] m233_85;
   assign m233_85 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_86 = W*in
   wire signed [9:0] m233_86;
   assign m233_86 =10'b0;

   // m233_87 = W*in
   wire signed [9:0] m233_87;
   assign m233_87 =10'b0;

   // m233_88 = W*in
   wire signed [9:0] m233_88;
   assign m233_88 =10'b0;

   // m233_89 = W*in
   wire signed [9:0] m233_89;
   assign m233_89 =10'b0;

   // m233_90 = W*in
   wire signed [9:0] m233_90;
   assign m233_90 =10'b0;

   // m233_91 = W*in
   wire signed [9:0] m233_91;
   assign m233_91 =10'b0;

   // m233_92 = W*in
   wire signed [9:0] m233_92;
   assign m233_92 =10'b0;

   // m233_93 = W*in
   wire signed [9:0] m233_93;
   assign m233_93 =10'b0;

   // m233_94 = W*in
   wire signed [9:0] m233_94;
   assign m233_94 =10'b0;

   // m233_95 = W*in
   wire signed [9:0] m233_95;
   assign m233_95 =10'b0;

   // m233_96 = W*in
   wire signed [9:0] m233_96;
   assign m233_96 =10'b0;

   // m233_97 = W*in
   wire signed [9:0] m233_97;
   assign m233_97 =10'b0;

   // m233_98 = W*in
   wire signed [9:0] m233_98;
   assign m233_98 =10'b0;

   // m233_99 = W*in
   wire signed [9:0] m233_99;
   assign m233_99 =10'b0;

   // m233_100 = W*in
   wire signed [9:0] m233_100;
   assign m233_100 =10'b0;

   // m233_101 = W*in
   wire signed [9:0] m233_101;
   assign m233_101 =10'b0;

   // m233_102 = W*in
   wire signed [9:0] m233_102;
   assign m233_102 =10'b0;

   // m233_103 = W*in
   wire signed [9:0] m233_103;
   assign m233_103 =10'b0;

   // m233_104 = W*in
   wire signed [9:0] m233_104;
   assign m233_104 =10'b0;

   // m233_105 = W*in
   wire signed [9:0] m233_105;
   assign m233_105 =10'b0;

   // m233_106 = W*in
   wire signed [9:0] m233_106;
   assign m233_106 =10'b0;

   // m233_107 = W*in
   wire signed [9:0] m233_107;
   assign m233_107 =10'b0;

   // m233_108 = W*in
   wire signed [9:0] m233_108;
   assign m233_108 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_109 = W*in
   wire signed [9:0] m233_109;
   assign m233_109 ={ {5{neg233[5]}} , neg233[5:1] };

   // m233_110 = W*in
   wire signed [9:0] m233_110;
   assign m233_110 =10'b0;

   // m233_111 = W*in
   wire signed [9:0] m233_111;
   assign m233_111 =10'b0;

   // m233_112 = W*in
   wire signed [9:0] m233_112;
   assign m233_112 =10'b0;

   // m233_113 = W*in
   wire signed [9:0] m233_113;
   assign m233_113 =10'b0;

   // m233_114 = W*in
   wire signed [9:0] m233_114;
   assign m233_114 =10'b0;

   // m233_115 = W*in
   wire signed [9:0] m233_115;
   assign m233_115 =10'b0;

   // m233_116 = W*in
   wire signed [9:0] m233_116;
   assign m233_116 =10'b0;

   // m233_117 = W*in
   wire signed [9:0] m233_117;
   assign m233_117 =10'b0;

   // m234_1 = W*in
   wire signed [9:0] m234_1;
   assign m234_1 =10'b0;

   // m234_2 = W*in
   wire signed [9:0] m234_2;
   assign m234_2 =10'b0;

   // m234_3 = W*in
   wire signed [9:0] m234_3;
   assign m234_3 =10'b0;

   // m234_4 = W*in
   wire signed [9:0] m234_4;
   assign m234_4 =10'b0;

   // m234_5 = W*in
   wire signed [9:0] m234_5;
   assign m234_5 ={ {4{in234[5]}} , in234[5:0] };

   // m234_6 = W*in
   wire signed [9:0] m234_6;
   assign m234_6 =10'b0;

   // m234_7 = W*in
   wire signed [9:0] m234_7;
   assign m234_7 =10'b0;

   // m234_8 = W*in
   wire signed [9:0] m234_8;
   assign m234_8 =10'b0;

   // m234_9 = W*in
   wire signed [9:0] m234_9;
   assign m234_9 =10'b0;

   // m234_10 = W*in
   wire signed [9:0] m234_10;
   assign m234_10 =10'b0;

   // m234_11 = W*in
   wire signed [9:0] m234_11;
   assign m234_11 =10'b0;

   // m234_12 = W*in
   wire signed [9:0] m234_12;
   assign m234_12 =10'b0;

   // m234_13 = W*in
   wire signed [9:0] m234_13;
   assign m234_13 =10'b0;

   // m234_14 = W*in
   wire signed [9:0] m234_14;
   assign m234_14 =10'b0;

   // m234_15 = W*in
   wire signed [9:0] m234_15;
   assign m234_15 =10'b0;

   // m234_16 = W*in
   wire signed [9:0] m234_16;
   assign m234_16 =10'b0;

   // m234_17 = W*in
   wire signed [9:0] m234_17;
   assign m234_17 =10'b0;

   // m234_18 = W*in
   wire signed [9:0] m234_18;
   assign m234_18 =10'b0;

   // m234_19 = W*in
   wire signed [9:0] m234_19;
   assign m234_19 ={ {5{in234[5]}} , in234[5:1] };

   // m234_20 = W*in
   wire signed [9:0] m234_20;
   assign m234_20 =10'b0;

   // m234_21 = W*in
   wire signed [9:0] m234_21;
   assign m234_21 =10'b0;

   // m234_22 = W*in
   wire signed [9:0] m234_22;
   assign m234_22 =10'b0;

   // m234_23 = W*in
   wire signed [9:0] m234_23;
   assign m234_23 =10'b0;

   // m234_24 = W*in
   wire signed [9:0] m234_24;
   assign m234_24 =10'b0;

   // m234_25 = W*in
   wire signed [9:0] m234_25;
   assign m234_25 =10'b0;

   // m234_26 = W*in
   wire signed [9:0] m234_26;
   assign m234_26 =10'b0;

   // m234_27 = W*in
   wire signed [9:0] m234_27;
   assign m234_27 =10'b0;

   // m234_28 = W*in
   wire signed [9:0] m234_28;
   assign m234_28 =10'b0;

   // m234_29 = W*in
   wire signed [9:0] m234_29;
   assign m234_29 =10'b0;

   // m234_30 = W*in
   wire signed [9:0] m234_30;
   assign m234_30 =10'b0;

   // m234_31 = W*in
   wire signed [9:0] m234_31;
   assign m234_31 =10'b0;

   // m234_32 = W*in
   wire signed [9:0] m234_32;
   assign m234_32 =10'b0;

   // m234_33 = W*in
   wire signed [9:0] m234_33;
   assign m234_33 =10'b0;

   // m234_34 = W*in
   wire signed [9:0] m234_34;
   assign m234_34 =10'b0;

   // m234_35 = W*in
   wire signed [9:0] m234_35;
   assign m234_35 =10'b0;

   // m234_36 = W*in
   wire signed [9:0] m234_36;
   assign m234_36 =10'b0;

   // m234_37 = W*in
   wire signed [9:0] m234_37;
   assign m234_37 =10'b0;

   // m234_38 = W*in
   wire signed [9:0] m234_38;
   assign m234_38 =10'b0;

   // m234_39 = W*in
   wire signed [9:0] m234_39;
   assign m234_39 =10'b0;

   // m234_40 = W*in
   wire signed [9:0] m234_40;
   assign m234_40 =10'b0;

   // m234_41 = W*in
   wire signed [9:0] m234_41;
   assign m234_41 =10'b0;

   // m234_42 = W*in
   wire signed [9:0] m234_42;
   assign m234_42 =10'b0;

   // m234_43 = W*in
   wire signed [9:0] m234_43;
   assign m234_43 =10'b0;

   // m234_44 = W*in
   wire signed [9:0] m234_44;
   assign m234_44 =10'b0;

   // m234_45 = W*in
   wire signed [9:0] m234_45;
   assign m234_45 =10'b0;

   // m234_46 = W*in
   wire signed [9:0] m234_46;
   assign m234_46 =10'b0;

   // m234_47 = W*in
   wire signed [9:0] m234_47;
   assign m234_47 =10'b0;

   // m234_48 = W*in
   wire signed [9:0] m234_48;
   assign m234_48 =10'b0;

   // m234_49 = W*in
   wire signed [9:0] m234_49;
   assign m234_49 =10'b0;

   // m234_50 = W*in
   wire signed [9:0] m234_50;
   assign m234_50 =10'b0;

   // m234_51 = W*in
   wire signed [9:0] m234_51;
   assign m234_51 =10'b0;

   // m234_52 = W*in
   wire signed [9:0] m234_52;
   assign m234_52 =10'b0;

   // m234_53 = W*in
   wire signed [9:0] m234_53;
   assign m234_53 =10'b0;

   // m234_54 = W*in
   wire signed [9:0] m234_54;
   assign m234_54 =10'b0;

   // m234_55 = W*in
   wire signed [9:0] m234_55;
   assign m234_55 =10'b0;

   // m234_56 = W*in
   wire signed [9:0] m234_56;
   assign m234_56 =10'b0;

   // m234_57 = W*in
   wire signed [9:0] m234_57;
   assign m234_57 =10'b0;

   // m234_58 = W*in
   wire signed [9:0] m234_58;
   assign m234_58 =10'b0;

   // m234_59 = W*in
   wire signed [9:0] m234_59;
   assign m234_59 =10'b0;

   // m234_60 = W*in
   wire signed [9:0] m234_60;
   assign m234_60 =10'b0;

   // m234_61 = W*in
   wire signed [9:0] m234_61;
   assign m234_61 =10'b0;

   // m234_62 = W*in
   wire signed [9:0] m234_62;
   assign m234_62 =10'b0;

   // m234_63 = W*in
   wire signed [9:0] m234_63;
   assign m234_63 =10'b0;

   // m234_64 = W*in
   wire signed [9:0] m234_64;
   assign m234_64 =10'b0;

   // m234_65 = W*in
   wire signed [9:0] m234_65;
   assign m234_65 =10'b0;

   // m234_66 = W*in
   wire signed [9:0] m234_66;
   assign m234_66 =10'b0;

   // m234_67 = W*in
   wire signed [9:0] m234_67;
   assign m234_67 ={ {5{in234[5]}} , in234[5:1] };

   // m234_68 = W*in
   wire signed [9:0] m234_68;
   assign m234_68 =10'b0;

   // m234_69 = W*in
   wire signed [9:0] m234_69;
   assign m234_69 ={ {5{in234[5]}} , in234[5:1] };

   // m234_70 = W*in
   wire signed [9:0] m234_70;
   assign m234_70 =10'b0;

   // m234_71 = W*in
   wire signed [9:0] m234_71;
   assign m234_71 =10'b0;

   // m234_72 = W*in
   wire signed [9:0] m234_72;
   assign m234_72 =10'b0;

   // m234_73 = W*in
   wire signed [9:0] m234_73;
   assign m234_73 =10'b0;

   // m234_74 = W*in
   wire signed [9:0] m234_74;
   assign m234_74 =10'b0;

   // m234_75 = W*in
   wire signed [9:0] m234_75;
   assign m234_75 =10'b0;

   // m234_76 = W*in
   wire signed [9:0] m234_76;
   assign m234_76 =10'b0;

   // m234_77 = W*in
   wire signed [9:0] m234_77;
   assign m234_77 =10'b0;

   // m234_78 = W*in
   wire signed [9:0] m234_78;
   assign m234_78 =10'b0;

   // m234_79 = W*in
   wire signed [9:0] m234_79;
   assign m234_79 =10'b0;

   // m234_80 = W*in
   wire signed [9:0] m234_80;
   assign m234_80 =10'b0;

   // m234_81 = W*in
   wire signed [9:0] m234_81;
   assign m234_81 =10'b0;

   // m234_82 = W*in
   wire signed [9:0] m234_82;
   assign m234_82 =10'b0;

   // m234_83 = W*in
   wire signed [9:0] m234_83;
   assign m234_83 =10'b0;

   // m234_84 = W*in
   wire signed [9:0] m234_84;
   assign m234_84 =10'b0;

   // m234_85 = W*in
   wire signed [9:0] m234_85;
   assign m234_85 ={ {5{in234[5]}} , in234[5:1] };

   // m234_86 = W*in
   wire signed [9:0] m234_86;
   assign m234_86 =10'b0;

   // m234_87 = W*in
   wire signed [9:0] m234_87;
   assign m234_87 =10'b0;

   // m234_88 = W*in
   wire signed [9:0] m234_88;
   assign m234_88 =10'b0;

   // m234_89 = W*in
   wire signed [9:0] m234_89;
   assign m234_89 =10'b0;

   // m234_90 = W*in
   wire signed [9:0] m234_90;
   assign m234_90 =10'b0;

   // m234_91 = W*in
   wire signed [9:0] m234_91;
   assign m234_91 =10'b0;

   // m234_92 = W*in
   wire signed [9:0] m234_92;
   assign m234_92 =10'b0;

   // m234_93 = W*in
   wire signed [9:0] m234_93;
   assign m234_93 =10'b0;

   // m234_94 = W*in
   wire signed [9:0] m234_94;
   assign m234_94 =10'b0;

   // m234_95 = W*in
   wire signed [9:0] m234_95;
   assign m234_95 =10'b0;

   // m234_96 = W*in
   wire signed [9:0] m234_96;
   assign m234_96 =10'b0;

   // m234_97 = W*in
   wire signed [9:0] m234_97;
   assign m234_97 =10'b0;

   // m234_98 = W*in
   wire signed [9:0] m234_98;
   assign m234_98 =10'b0;

   // m234_99 = W*in
   wire signed [9:0] m234_99;
   assign m234_99 =10'b0;

   // m234_100 = W*in
   wire signed [9:0] m234_100;
   assign m234_100 =10'b0;

   // m234_101 = W*in
   wire signed [9:0] m234_101;
   assign m234_101 =10'b0;

   // m234_102 = W*in
   wire signed [9:0] m234_102;
   assign m234_102 =10'b0;

   // m234_103 = W*in
   wire signed [9:0] m234_103;
   assign m234_103 =10'b0;

   // m234_104 = W*in
   wire signed [9:0] m234_104;
   assign m234_104 =10'b0;

   // m234_105 = W*in
   wire signed [9:0] m234_105;
   assign m234_105 =10'b0;

   // m234_106 = W*in
   wire signed [9:0] m234_106;
   assign m234_106 =10'b0;

   // m234_107 = W*in
   wire signed [9:0] m234_107;
   assign m234_107 =10'b0;

   // m234_108 = W*in
   wire signed [9:0] m234_108;
   assign m234_108 =10'b0;

   // m234_109 = W*in
   wire signed [9:0] m234_109;
   assign m234_109 =10'b0;

   // m234_110 = W*in
   wire signed [9:0] m234_110;
   assign m234_110 =10'b0;

   // m234_111 = W*in
   wire signed [9:0] m234_111;
   assign m234_111 =10'b0;

   // m234_112 = W*in
   wire signed [9:0] m234_112;
   assign m234_112 =10'b0;

   // m234_113 = W*in
   wire signed [9:0] m234_113;
   assign m234_113 =10'b0;

   // m234_114 = W*in
   wire signed [9:0] m234_114;
   assign m234_114 =10'b0;

   // m234_115 = W*in
   wire signed [9:0] m234_115;
   assign m234_115 =10'b0;

   // m234_116 = W*in
   wire signed [9:0] m234_116;
   assign m234_116 =10'b0;

   // m234_117 = W*in
   wire signed [9:0] m234_117;
   assign m234_117 =10'b0;

   // m235_1 = W*in
   wire signed [9:0] m235_1;
   assign m235_1 =10'b0;

   // m235_2 = W*in
   wire signed [9:0] m235_2;
   assign m235_2 =10'b0;

   // m235_3 = W*in
   wire signed [9:0] m235_3;
   assign m235_3 =10'b0;

   // m235_4 = W*in
   wire signed [9:0] m235_4;
   assign m235_4 =10'b0;

   // m235_5 = W*in
   wire signed [9:0] m235_5;
   assign m235_5 ={ {4{in235[5]}} , in235[5:0] };

   // m235_6 = W*in
   wire signed [9:0] m235_6;
   assign m235_6 =10'b0;

   // m235_7 = W*in
   wire signed [9:0] m235_7;
   assign m235_7 =10'b0;

   // m235_8 = W*in
   wire signed [9:0] m235_8;
   assign m235_8 =10'b0;

   // m235_9 = W*in
   wire signed [9:0] m235_9;
   assign m235_9 =10'b0;

   // m235_10 = W*in
   wire signed [9:0] m235_10;
   assign m235_10 =10'b0;

   // m235_11 = W*in
   wire signed [9:0] m235_11;
   assign m235_11 =10'b0;

   // m235_12 = W*in
   wire signed [9:0] m235_12;
   assign m235_12 =10'b0;

   // m235_13 = W*in
   wire signed [9:0] m235_13;
   assign m235_13 =10'b0;

   // m235_14 = W*in
   wire signed [9:0] m235_14;
   assign m235_14 =10'b0;

   // m235_15 = W*in
   wire signed [9:0] m235_15;
   assign m235_15 =10'b0;

   // m235_16 = W*in
   wire signed [9:0] m235_16;
   assign m235_16 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_17 = W*in
   wire signed [9:0] m235_17;
   assign m235_17 =10'b0;

   // m235_18 = W*in
   wire signed [9:0] m235_18;
   assign m235_18 =10'b0;

   // m235_19 = W*in
   wire signed [9:0] m235_19;
   assign m235_19 =10'b0;

   // m235_20 = W*in
   wire signed [9:0] m235_20;
   assign m235_20 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_21 = W*in
   wire signed [9:0] m235_21;
   assign m235_21 ={ {5{in235[5]}} , in235[5:1] };

   // m235_22 = W*in
   wire signed [9:0] m235_22;
   assign m235_22 =10'b0;

   // m235_23 = W*in
   wire signed [9:0] m235_23;
   assign m235_23 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_24 = W*in
   wire signed [9:0] m235_24;
   assign m235_24 =10'b0;

   // m235_25 = W*in
   wire signed [9:0] m235_25;
   assign m235_25 =10'b0;

   // m235_26 = W*in
   wire signed [9:0] m235_26;
   assign m235_26 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_27 = W*in
   wire signed [9:0] m235_27;
   assign m235_27 =10'b0;

   // m235_28 = W*in
   wire signed [9:0] m235_28;
   assign m235_28 =10'b0;

   // m235_29 = W*in
   wire signed [9:0] m235_29;
   assign m235_29 =10'b0;

   // m235_30 = W*in
   wire signed [9:0] m235_30;
   assign m235_30 =10'b0;

   // m235_31 = W*in
   wire signed [9:0] m235_31;
   assign m235_31 =10'b0;

   // m235_32 = W*in
   wire signed [9:0] m235_32;
   assign m235_32 ={ {4{in235[5]}} , in235[5:0] };

   // m235_33 = W*in
   wire signed [9:0] m235_33;
   assign m235_33 =10'b0;

   // m235_34 = W*in
   wire signed [9:0] m235_34;
   assign m235_34 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_35 = W*in
   wire signed [9:0] m235_35;
   assign m235_35 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_36 = W*in
   wire signed [9:0] m235_36;
   assign m235_36 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_37 = W*in
   wire signed [9:0] m235_37;
   assign m235_37 =10'b0;

   // m235_38 = W*in
   wire signed [9:0] m235_38;
   assign m235_38 =10'b0;

   // m235_39 = W*in
   wire signed [9:0] m235_39;
   assign m235_39 =10'b0;

   // m235_40 = W*in
   wire signed [9:0] m235_40;
   assign m235_40 =10'b0;

   // m235_41 = W*in
   wire signed [9:0] m235_41;
   assign m235_41 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_42 = W*in
   wire signed [9:0] m235_42;
   assign m235_42 =10'b0;

   // m235_43 = W*in
   wire signed [9:0] m235_43;
   assign m235_43 =10'b0;

   // m235_44 = W*in
   wire signed [9:0] m235_44;
   assign m235_44 =10'b0;

   // m235_45 = W*in
   wire signed [9:0] m235_45;
   assign m235_45 =10'b0;

   // m235_46 = W*in
   wire signed [9:0] m235_46;
   assign m235_46 =10'b0;

   // m235_47 = W*in
   wire signed [9:0] m235_47;
   assign m235_47 =10'b0;

   // m235_48 = W*in
   wire signed [9:0] m235_48;
   assign m235_48 =10'b0;

   // m235_49 = W*in
   wire signed [9:0] m235_49;
   assign m235_49 ={ {4{in235[5]}} , in235[5:0] };

   // m235_50 = W*in
   wire signed [9:0] m235_50;
   assign m235_50 =10'b0;

   // m235_51 = W*in
   wire signed [9:0] m235_51;
   assign m235_51 =10'b0;

   // m235_52 = W*in
   wire signed [9:0] m235_52;
   assign m235_52 =10'b0;

   // m235_53 = W*in
   wire signed [9:0] m235_53;
   assign m235_53 ={ {4{in235[5]}} , in235[5:0] };

   // m235_54 = W*in
   wire signed [9:0] m235_54;
   assign m235_54 ={ {4{in235[5]}} , in235[5:0] };

   // m235_55 = W*in
   wire signed [9:0] m235_55;
   assign m235_55 =10'b0;

   // m235_56 = W*in
   wire signed [9:0] m235_56;
   assign m235_56 =10'b0;

   // m235_57 = W*in
   wire signed [9:0] m235_57;
   assign m235_57 =10'b0;

   // m235_58 = W*in
   wire signed [9:0] m235_58;
   assign m235_58 =10'b0;

   // m235_59 = W*in
   wire signed [9:0] m235_59;
   assign m235_59 =10'b0;

   // m235_60 = W*in
   wire signed [9:0] m235_60;
   assign m235_60 =10'b0;

   // m235_61 = W*in
   wire signed [9:0] m235_61;
   assign m235_61 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_62 = W*in
   wire signed [9:0] m235_62;
   assign m235_62 =10'b0;

   // m235_63 = W*in
   wire signed [9:0] m235_63;
   assign m235_63 =10'b0;

   // m235_64 = W*in
   wire signed [9:0] m235_64;
   assign m235_64 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_65 = W*in
   wire signed [9:0] m235_65;
   assign m235_65 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_66 = W*in
   wire signed [9:0] m235_66;
   assign m235_66 ={ {5{in235[5]}} , in235[5:1] };

   // m235_67 = W*in
   wire signed [9:0] m235_67;
   assign m235_67 =10'b0;

   // m235_68 = W*in
   wire signed [9:0] m235_68;
   assign m235_68 =10'b0;

   // m235_69 = W*in
   wire signed [9:0] m235_69;
   assign m235_69 =10'b0;

   // m235_70 = W*in
   wire signed [9:0] m235_70;
   assign m235_70 =10'b0;

   // m235_71 = W*in
   wire signed [9:0] m235_71;
   assign m235_71 =10'b0;

   // m235_72 = W*in
   wire signed [9:0] m235_72;
   assign m235_72 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_73 = W*in
   wire signed [9:0] m235_73;
   assign m235_73 =10'b0;

   // m235_74 = W*in
   wire signed [9:0] m235_74;
   assign m235_74 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_75 = W*in
   wire signed [9:0] m235_75;
   assign m235_75 ={ {5{neg235[5]}} , neg235[5:1] };

   // m235_76 = W*in
   wire signed [9:0] m235_76;
   assign m235_76 =10'b0;

   // m235_77 = W*in
   wire signed [9:0] m235_77;
   assign m235_77 =10'b0;

   // m235_78 = W*in
   wire signed [9:0] m235_78;
   assign m235_78 =10'b0;

   // m235_79 = W*in
   wire signed [9:0] m235_79;
   assign m235_79 =10'b0;

   // m235_80 = W*in
   wire signed [9:0] m235_80;
   assign m235_80 ={ {4{in235[5]}} , in235[5:0] };

   // m235_81 = W*in
   wire signed [9:0] m235_81;
   assign m235_81 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_82 = W*in
   wire signed [9:0] m235_82;
   assign m235_82 =10'b0;

   // m235_83 = W*in
   wire signed [9:0] m235_83;
   assign m235_83 =10'b0;

   // m235_84 = W*in
   wire signed [9:0] m235_84;
   assign m235_84 =10'b0;

   // m235_85 = W*in
   wire signed [9:0] m235_85;
   assign m235_85 ={ {5{in235[5]}} , in235[5:1] };

   // m235_86 = W*in
   wire signed [9:0] m235_86;
   assign m235_86 =10'b0;

   // m235_87 = W*in
   wire signed [9:0] m235_87;
   assign m235_87 =10'b0;

   // m235_88 = W*in
   wire signed [9:0] m235_88;
   assign m235_88 =10'b0;

   // m235_89 = W*in
   wire signed [9:0] m235_89;
   assign m235_89 =10'b0;

   // m235_90 = W*in
   wire signed [9:0] m235_90;
   assign m235_90 =10'b0;

   // m235_91 = W*in
   wire signed [9:0] m235_91;
   assign m235_91 =10'b0;

   // m235_92 = W*in
   wire signed [9:0] m235_92;
   assign m235_92 =10'b0;

   // m235_93 = W*in
   wire signed [9:0] m235_93;
   assign m235_93 =10'b0;

   // m235_94 = W*in
   wire signed [9:0] m235_94;
   assign m235_94 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_95 = W*in
   wire signed [9:0] m235_95;
   assign m235_95 ={ {4{in235[5]}} , in235[5:0] };

   // m235_96 = W*in
   wire signed [9:0] m235_96;
   assign m235_96 =10'b0;

   // m235_97 = W*in
   wire signed [9:0] m235_97;
   assign m235_97 =10'b0;

   // m235_98 = W*in
   wire signed [9:0] m235_98;
   assign m235_98 =10'b0;

   // m235_99 = W*in
   wire signed [9:0] m235_99;
   assign m235_99 =10'b0;

   // m235_100 = W*in
   wire signed [9:0] m235_100;
   assign m235_100 =10'b0;

   // m235_101 = W*in
   wire signed [9:0] m235_101;
   assign m235_101 =10'b0;

   // m235_102 = W*in
   wire signed [9:0] m235_102;
   assign m235_102 =10'b0;

   // m235_103 = W*in
   wire signed [9:0] m235_103;
   assign m235_103 =10'b0;

   // m235_104 = W*in
   wire signed [9:0] m235_104;
   assign m235_104 =10'b0;

   // m235_105 = W*in
   wire signed [9:0] m235_105;
   assign m235_105 =10'b0;

   // m235_106 = W*in
   wire signed [9:0] m235_106;
   assign m235_106 =10'b0;

   // m235_107 = W*in
   wire signed [9:0] m235_107;
   assign m235_107 =10'b0;

   // m235_108 = W*in
   wire signed [9:0] m235_108;
   assign m235_108 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_109 = W*in
   wire signed [9:0] m235_109;
   assign m235_109 ={ {4{neg235[5]}} , neg235[5:0] };

   // m235_110 = W*in
   wire signed [9:0] m235_110;
   assign m235_110 =10'b0;

   // m235_111 = W*in
   wire signed [9:0] m235_111;
   assign m235_111 =10'b0;

   // m235_112 = W*in
   wire signed [9:0] m235_112;
   assign m235_112 =10'b0;

   // m235_113 = W*in
   wire signed [9:0] m235_113;
   assign m235_113 =10'b0;

   // m235_114 = W*in
   wire signed [9:0] m235_114;
   assign m235_114 =10'b0;

   // m235_115 = W*in
   wire signed [9:0] m235_115;
   assign m235_115 =10'b0;

   // m235_116 = W*in
   wire signed [9:0] m235_116;
   assign m235_116 =10'b0;

   // m235_117 = W*in
   wire signed [9:0] m235_117;
   assign m235_117 =10'b0;

   // m236_1 = W*in
   wire signed [9:0] m236_1;
   assign m236_1 =10'b0;

   // m236_2 = W*in
   wire signed [9:0] m236_2;
   assign m236_2 =10'b0;

   // m236_3 = W*in
   wire signed [9:0] m236_3;
   assign m236_3 =10'b0;

   // m236_4 = W*in
   wire signed [9:0] m236_4;
   assign m236_4 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_5 = W*in
   wire signed [9:0] m236_5;
   assign m236_5 ={ {4{in236[5]}} , in236[5:0] };

   // m236_6 = W*in
   wire signed [9:0] m236_6;
   assign m236_6 ={ {4{in236[5]}} , in236[5:0] };

   // m236_7 = W*in
   wire signed [9:0] m236_7;
   assign m236_7 =10'b0;

   // m236_8 = W*in
   wire signed [9:0] m236_8;
   assign m236_8 ={ {4{in236[5]}} , in236[5:0] };

   // m236_9 = W*in
   wire signed [9:0] m236_9;
   assign m236_9 =10'b0;

   // m236_10 = W*in
   wire signed [9:0] m236_10;
   assign m236_10 =10'b0;

   // m236_11 = W*in
   wire signed [9:0] m236_11;
   assign m236_11 ={ {4{in236[5]}} , in236[5:0] };

   // m236_12 = W*in
   wire signed [9:0] m236_12;
   assign m236_12 =10'b0;

   // m236_13 = W*in
   wire signed [9:0] m236_13;
   assign m236_13 =10'b0;

   // m236_14 = W*in
   wire signed [9:0] m236_14;
   assign m236_14 =10'b0;

   // m236_15 = W*in
   wire signed [9:0] m236_15;
   assign m236_15 ={ {4{in236[5]}} , in236[5:0] };

   // m236_16 = W*in
   wire signed [9:0] m236_16;
   assign m236_16 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_17 = W*in
   wire signed [9:0] m236_17;
   assign m236_17 ={ {5{in236[5]}} , in236[5:1] };

   // m236_18 = W*in
   wire signed [9:0] m236_18;
   assign m236_18 =10'b0;

   // m236_19 = W*in
   wire signed [9:0] m236_19;
   assign m236_19 ={ {4{in236[5]}} , in236[5:0] };

   // m236_20 = W*in
   wire signed [9:0] m236_20;
   assign m236_20 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_21 = W*in
   wire signed [9:0] m236_21;
   assign m236_21 =10'b0;

   // m236_22 = W*in
   wire signed [9:0] m236_22;
   assign m236_22 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_23 = W*in
   wire signed [9:0] m236_23;
   assign m236_23 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_24 = W*in
   wire signed [9:0] m236_24;
   assign m236_24 =10'b0;

   // m236_25 = W*in
   wire signed [9:0] m236_25;
   assign m236_25 =10'b0;

   // m236_26 = W*in
   wire signed [9:0] m236_26;
   assign m236_26 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_27 = W*in
   wire signed [9:0] m236_27;
   assign m236_27 =10'b0;

   // m236_28 = W*in
   wire signed [9:0] m236_28;
   assign m236_28 =10'b0;

   // m236_29 = W*in
   wire signed [9:0] m236_29;
   assign m236_29 ={ {4{in236[5]}} , in236[5:0] };

   // m236_30 = W*in
   wire signed [9:0] m236_30;
   assign m236_30 =10'b0;

   // m236_31 = W*in
   wire signed [9:0] m236_31;
   assign m236_31 ={ {5{in236[5]}} , in236[5:1] };

   // m236_32 = W*in
   wire signed [9:0] m236_32;
   assign m236_32 ={ {5{in236[5]}} , in236[5:1] };

   // m236_33 = W*in
   wire signed [9:0] m236_33;
   assign m236_33 =10'b0;

   // m236_34 = W*in
   wire signed [9:0] m236_34;
   assign m236_34 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_35 = W*in
   wire signed [9:0] m236_35;
   assign m236_35 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_36 = W*in
   wire signed [9:0] m236_36;
   assign m236_36 =10'b0;

   // m236_37 = W*in
   wire signed [9:0] m236_37;
   assign m236_37 =10'b0;

   // m236_38 = W*in
   wire signed [9:0] m236_38;
   assign m236_38 ={ {4{in236[5]}} , in236[5:0] };

   // m236_39 = W*in
   wire signed [9:0] m236_39;
   assign m236_39 =10'b0;

   // m236_40 = W*in
   wire signed [9:0] m236_40;
   assign m236_40 =10'b0;

   // m236_41 = W*in
   wire signed [9:0] m236_41;
   assign m236_41 =10'b0;

   // m236_42 = W*in
   wire signed [9:0] m236_42;
   assign m236_42 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_43 = W*in
   wire signed [9:0] m236_43;
   assign m236_43 =10'b0;

   // m236_44 = W*in
   wire signed [9:0] m236_44;
   assign m236_44 ={ {4{in236[5]}} , in236[5:0] };

   // m236_45 = W*in
   wire signed [9:0] m236_45;
   assign m236_45 =10'b0;

   // m236_46 = W*in
   wire signed [9:0] m236_46;
   assign m236_46 =10'b0;

   // m236_47 = W*in
   wire signed [9:0] m236_47;
   assign m236_47 =10'b0;

   // m236_48 = W*in
   wire signed [9:0] m236_48;
   assign m236_48 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_49 = W*in
   wire signed [9:0] m236_49;
   assign m236_49 ={ {4{in236[5]}} , in236[5:0] };

   // m236_50 = W*in
   wire signed [9:0] m236_50;
   assign m236_50 =10'b0;

   // m236_51 = W*in
   wire signed [9:0] m236_51;
   assign m236_51 =10'b0;

   // m236_52 = W*in
   wire signed [9:0] m236_52;
   assign m236_52 =10'b0;

   // m236_53 = W*in
   wire signed [9:0] m236_53;
   assign m236_53 ={ {4{in236[5]}} , in236[5:0] };

   // m236_54 = W*in
   wire signed [9:0] m236_54;
   assign m236_54 =10'b0;

   // m236_55 = W*in
   wire signed [9:0] m236_55;
   assign m236_55 =10'b0;

   // m236_56 = W*in
   wire signed [9:0] m236_56;
   assign m236_56 =10'b0;

   // m236_57 = W*in
   wire signed [9:0] m236_57;
   assign m236_57 =10'b0;

   // m236_58 = W*in
   wire signed [9:0] m236_58;
   assign m236_58 =10'b0;

   // m236_59 = W*in
   wire signed [9:0] m236_59;
   assign m236_59 =10'b0;

   // m236_60 = W*in
   wire signed [9:0] m236_60;
   assign m236_60 =10'b0;

   // m236_61 = W*in
   wire signed [9:0] m236_61;
   assign m236_61 =10'b0;

   // m236_62 = W*in
   wire signed [9:0] m236_62;
   assign m236_62 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_63 = W*in
   wire signed [9:0] m236_63;
   assign m236_63 =10'b0;

   // m236_64 = W*in
   wire signed [9:0] m236_64;
   assign m236_64 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_65 = W*in
   wire signed [9:0] m236_65;
   assign m236_65 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_66 = W*in
   wire signed [9:0] m236_66;
   assign m236_66 ={ {4{in236[5]}} , in236[5:0] };

   // m236_67 = W*in
   wire signed [9:0] m236_67;
   assign m236_67 ={ {3{in236[5]}} , in236 , {1{1'b0}} };

   // m236_68 = W*in
   wire signed [9:0] m236_68;
   assign m236_68 ={ {4{in236[5]}} , in236[5:0] };

   // m236_69 = W*in
   wire signed [9:0] m236_69;
   assign m236_69 =10'b0;

   // m236_70 = W*in
   wire signed [9:0] m236_70;
   assign m236_70 =10'b0;

   // m236_71 = W*in
   wire signed [9:0] m236_71;
   assign m236_71 =10'b0;

   // m236_72 = W*in
   wire signed [9:0] m236_72;
   assign m236_72 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_73 = W*in
   wire signed [9:0] m236_73;
   assign m236_73 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_74 = W*in
   wire signed [9:0] m236_74;
   assign m236_74 =10'b0;

   // m236_75 = W*in
   wire signed [9:0] m236_75;
   assign m236_75 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_76 = W*in
   wire signed [9:0] m236_76;
   assign m236_76 =10'b0;

   // m236_77 = W*in
   wire signed [9:0] m236_77;
   assign m236_77 =10'b0;

   // m236_78 = W*in
   wire signed [9:0] m236_78;
   assign m236_78 =10'b0;

   // m236_79 = W*in
   wire signed [9:0] m236_79;
   assign m236_79 =10'b0;

   // m236_80 = W*in
   wire signed [9:0] m236_80;
   assign m236_80 ={ {4{in236[5]}} , in236[5:0] };

   // m236_81 = W*in
   wire signed [9:0] m236_81;
   assign m236_81 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_82 = W*in
   wire signed [9:0] m236_82;
   assign m236_82 =10'b0;

   // m236_83 = W*in
   wire signed [9:0] m236_83;
   assign m236_83 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_84 = W*in
   wire signed [9:0] m236_84;
   assign m236_84 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_85 = W*in
   wire signed [9:0] m236_85;
   assign m236_85 =10'b0;

   // m236_86 = W*in
   wire signed [9:0] m236_86;
   assign m236_86 =10'b0;

   // m236_87 = W*in
   wire signed [9:0] m236_87;
   assign m236_87 =10'b0;

   // m236_88 = W*in
   wire signed [9:0] m236_88;
   assign m236_88 =10'b0;

   // m236_89 = W*in
   wire signed [9:0] m236_89;
   assign m236_89 =10'b0;

   // m236_90 = W*in
   wire signed [9:0] m236_90;
   assign m236_90 =10'b0;

   // m236_91 = W*in
   wire signed [9:0] m236_91;
   assign m236_91 ={ {4{in236[5]}} , in236[5:0] };

   // m236_92 = W*in
   wire signed [9:0] m236_92;
   assign m236_92 =10'b0;

   // m236_93 = W*in
   wire signed [9:0] m236_93;
   assign m236_93 ={ {4{in236[5]}} , in236[5:0] };

   // m236_94 = W*in
   wire signed [9:0] m236_94;
   assign m236_94 =10'b0;

   // m236_95 = W*in
   wire signed [9:0] m236_95;
   assign m236_95 =10'b0;

   // m236_96 = W*in
   wire signed [9:0] m236_96;
   assign m236_96 =10'b0;

   // m236_97 = W*in
   wire signed [9:0] m236_97;
   assign m236_97 ={ {4{in236[5]}} , in236[5:0] };

   // m236_98 = W*in
   wire signed [9:0] m236_98;
   assign m236_98 =10'b0;

   // m236_99 = W*in
   wire signed [9:0] m236_99;
   assign m236_99 =10'b0;

   // m236_100 = W*in
   wire signed [9:0] m236_100;
   assign m236_100 =10'b0;

   // m236_101 = W*in
   wire signed [9:0] m236_101;
   assign m236_101 =10'b0;

   // m236_102 = W*in
   wire signed [9:0] m236_102;
   assign m236_102 =10'b0;

   // m236_103 = W*in
   wire signed [9:0] m236_103;
   assign m236_103 =10'b0;

   // m236_104 = W*in
   wire signed [9:0] m236_104;
   assign m236_104 =10'b0;

   // m236_105 = W*in
   wire signed [9:0] m236_105;
   assign m236_105 =10'b0;

   // m236_106 = W*in
   wire signed [9:0] m236_106;
   assign m236_106 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_107 = W*in
   wire signed [9:0] m236_107;
   assign m236_107 =10'b0;

   // m236_108 = W*in
   wire signed [9:0] m236_108;
   assign m236_108 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_109 = W*in
   wire signed [9:0] m236_109;
   assign m236_109 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_110 = W*in
   wire signed [9:0] m236_110;
   assign m236_110 =10'b0;

   // m236_111 = W*in
   wire signed [9:0] m236_111;
   assign m236_111 ={ {4{neg236[5]}} , neg236[5:0] };

   // m236_112 = W*in
   wire signed [9:0] m236_112;
   assign m236_112 =10'b0;

   // m236_113 = W*in
   wire signed [9:0] m236_113;
   assign m236_113 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_114 = W*in
   wire signed [9:0] m236_114;
   assign m236_114 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_115 = W*in
   wire signed [9:0] m236_115;
   assign m236_115 ={ {5{neg236[5]}} , neg236[5:1] };

   // m236_116 = W*in
   wire signed [9:0] m236_116;
   assign m236_116 =10'b0;

   // m236_117 = W*in
   wire signed [9:0] m236_117;
   assign m236_117 =10'b0;

   // m237_1 = W*in
   wire signed [9:0] m237_1;
   assign m237_1 =10'b0;

   // m237_2 = W*in
   wire signed [9:0] m237_2;
   assign m237_2 =10'b0;

   // m237_3 = W*in
   wire signed [9:0] m237_3;
   assign m237_3 =10'b0;

   // m237_4 = W*in
   wire signed [9:0] m237_4;
   assign m237_4 =10'b0;

   // m237_5 = W*in
   wire signed [9:0] m237_5;
   assign m237_5 =10'b0;

   // m237_6 = W*in
   wire signed [9:0] m237_6;
   assign m237_6 ={ {4{in237[5]}} , in237[5:0] };

   // m237_7 = W*in
   wire signed [9:0] m237_7;
   assign m237_7 =10'b0;

   // m237_8 = W*in
   wire signed [9:0] m237_8;
   assign m237_8 =10'b0;

   // m237_9 = W*in
   wire signed [9:0] m237_9;
   assign m237_9 =10'b0;

   // m237_10 = W*in
   wire signed [9:0] m237_10;
   assign m237_10 =10'b0;

   // m237_11 = W*in
   wire signed [9:0] m237_11;
   assign m237_11 =10'b0;

   // m237_12 = W*in
   wire signed [9:0] m237_12;
   assign m237_12 =10'b0;

   // m237_13 = W*in
   wire signed [9:0] m237_13;
   assign m237_13 =10'b0;

   // m237_14 = W*in
   wire signed [9:0] m237_14;
   assign m237_14 =10'b0;

   // m237_15 = W*in
   wire signed [9:0] m237_15;
   assign m237_15 ={ {4{in237[5]}} , in237[5:0] };

   // m237_16 = W*in
   wire signed [9:0] m237_16;
   assign m237_16 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_17 = W*in
   wire signed [9:0] m237_17;
   assign m237_17 =10'b0;

   // m237_18 = W*in
   wire signed [9:0] m237_18;
   assign m237_18 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_19 = W*in
   wire signed [9:0] m237_19;
   assign m237_19 ={ {4{in237[5]}} , in237[5:0] };

   // m237_20 = W*in
   wire signed [9:0] m237_20;
   assign m237_20 =10'b0;

   // m237_21 = W*in
   wire signed [9:0] m237_21;
   assign m237_21 =10'b0;

   // m237_22 = W*in
   wire signed [9:0] m237_22;
   assign m237_22 =10'b0;

   // m237_23 = W*in
   wire signed [9:0] m237_23;
   assign m237_23 ={ {5{neg237[5]}} , neg237[5:1] };

   // m237_24 = W*in
   wire signed [9:0] m237_24;
   assign m237_24 =10'b0;

   // m237_25 = W*in
   wire signed [9:0] m237_25;
   assign m237_25 =10'b0;

   // m237_26 = W*in
   wire signed [9:0] m237_26;
   assign m237_26 =10'b0;

   // m237_27 = W*in
   wire signed [9:0] m237_27;
   assign m237_27 =10'b0;

   // m237_28 = W*in
   wire signed [9:0] m237_28;
   assign m237_28 ={ {5{in237[5]}} , in237[5:1] };

   // m237_29 = W*in
   wire signed [9:0] m237_29;
   assign m237_29 =10'b0;

   // m237_30 = W*in
   wire signed [9:0] m237_30;
   assign m237_30 =10'b0;

   // m237_31 = W*in
   wire signed [9:0] m237_31;
   assign m237_31 =10'b0;

   // m237_32 = W*in
   wire signed [9:0] m237_32;
   assign m237_32 =10'b0;

   // m237_33 = W*in
   wire signed [9:0] m237_33;
   assign m237_33 =10'b0;

   // m237_34 = W*in
   wire signed [9:0] m237_34;
   assign m237_34 =10'b0;

   // m237_35 = W*in
   wire signed [9:0] m237_35;
   assign m237_35 ={ {5{neg237[5]}} , neg237[5:1] };

   // m237_36 = W*in
   wire signed [9:0] m237_36;
   assign m237_36 =10'b0;

   // m237_37 = W*in
   wire signed [9:0] m237_37;
   assign m237_37 =10'b0;

   // m237_38 = W*in
   wire signed [9:0] m237_38;
   assign m237_38 ={ {4{in237[5]}} , in237[5:0] };

   // m237_39 = W*in
   wire signed [9:0] m237_39;
   assign m237_39 =10'b0;

   // m237_40 = W*in
   wire signed [9:0] m237_40;
   assign m237_40 =10'b0;

   // m237_41 = W*in
   wire signed [9:0] m237_41;
   assign m237_41 =10'b0;

   // m237_42 = W*in
   wire signed [9:0] m237_42;
   assign m237_42 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_43 = W*in
   wire signed [9:0] m237_43;
   assign m237_43 =10'b0;

   // m237_44 = W*in
   wire signed [9:0] m237_44;
   assign m237_44 ={ {4{in237[5]}} , in237[5:0] };

   // m237_45 = W*in
   wire signed [9:0] m237_45;
   assign m237_45 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_46 = W*in
   wire signed [9:0] m237_46;
   assign m237_46 =10'b0;

   // m237_47 = W*in
   wire signed [9:0] m237_47;
   assign m237_47 =10'b0;

   // m237_48 = W*in
   wire signed [9:0] m237_48;
   assign m237_48 =10'b0;

   // m237_49 = W*in
   wire signed [9:0] m237_49;
   assign m237_49 =10'b0;

   // m237_50 = W*in
   wire signed [9:0] m237_50;
   assign m237_50 =10'b0;

   // m237_51 = W*in
   wire signed [9:0] m237_51;
   assign m237_51 =10'b0;

   // m237_52 = W*in
   wire signed [9:0] m237_52;
   assign m237_52 =10'b0;

   // m237_53 = W*in
   wire signed [9:0] m237_53;
   assign m237_53 ={ {4{in237[5]}} , in237[5:0] };

   // m237_54 = W*in
   wire signed [9:0] m237_54;
   assign m237_54 ={ {4{in237[5]}} , in237[5:0] };

   // m237_55 = W*in
   wire signed [9:0] m237_55;
   assign m237_55 =10'b0;

   // m237_56 = W*in
   wire signed [9:0] m237_56;
   assign m237_56 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_57 = W*in
   wire signed [9:0] m237_57;
   assign m237_57 =10'b0;

   // m237_58 = W*in
   wire signed [9:0] m237_58;
   assign m237_58 =10'b0;

   // m237_59 = W*in
   wire signed [9:0] m237_59;
   assign m237_59 =10'b0;

   // m237_60 = W*in
   wire signed [9:0] m237_60;
   assign m237_60 =10'b0;

   // m237_61 = W*in
   wire signed [9:0] m237_61;
   assign m237_61 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_62 = W*in
   wire signed [9:0] m237_62;
   assign m237_62 =10'b0;

   // m237_63 = W*in
   wire signed [9:0] m237_63;
   assign m237_63 =10'b0;

   // m237_64 = W*in
   wire signed [9:0] m237_64;
   assign m237_64 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_65 = W*in
   wire signed [9:0] m237_65;
   assign m237_65 =10'b0;

   // m237_66 = W*in
   wire signed [9:0] m237_66;
   assign m237_66 =10'b0;

   // m237_67 = W*in
   wire signed [9:0] m237_67;
   assign m237_67 ={ {4{in237[5]}} , in237[5:0] };

   // m237_68 = W*in
   wire signed [9:0] m237_68;
   assign m237_68 =10'b0;

   // m237_69 = W*in
   wire signed [9:0] m237_69;
   assign m237_69 =10'b0;

   // m237_70 = W*in
   wire signed [9:0] m237_70;
   assign m237_70 ={ {5{in237[5]}} , in237[5:1] };

   // m237_71 = W*in
   wire signed [9:0] m237_71;
   assign m237_71 ={ {5{in237[5]}} , in237[5:1] };

   // m237_72 = W*in
   wire signed [9:0] m237_72;
   assign m237_72 =10'b0;

   // m237_73 = W*in
   wire signed [9:0] m237_73;
   assign m237_73 =10'b0;

   // m237_74 = W*in
   wire signed [9:0] m237_74;
   assign m237_74 =10'b0;

   // m237_75 = W*in
   wire signed [9:0] m237_75;
   assign m237_75 =10'b0;

   // m237_76 = W*in
   wire signed [9:0] m237_76;
   assign m237_76 =10'b0;

   // m237_77 = W*in
   wire signed [9:0] m237_77;
   assign m237_77 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_78 = W*in
   wire signed [9:0] m237_78;
   assign m237_78 =10'b0;

   // m237_79 = W*in
   wire signed [9:0] m237_79;
   assign m237_79 =10'b0;

   // m237_80 = W*in
   wire signed [9:0] m237_80;
   assign m237_80 =10'b0;

   // m237_81 = W*in
   wire signed [9:0] m237_81;
   assign m237_81 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_82 = W*in
   wire signed [9:0] m237_82;
   assign m237_82 =10'b0;

   // m237_83 = W*in
   wire signed [9:0] m237_83;
   assign m237_83 ={ {5{neg237[5]}} , neg237[5:1] };

   // m237_84 = W*in
   wire signed [9:0] m237_84;
   assign m237_84 =10'b0;

   // m237_85 = W*in
   wire signed [9:0] m237_85;
   assign m237_85 =10'b0;

   // m237_86 = W*in
   wire signed [9:0] m237_86;
   assign m237_86 =10'b0;

   // m237_87 = W*in
   wire signed [9:0] m237_87;
   assign m237_87 =10'b0;

   // m237_88 = W*in
   wire signed [9:0] m237_88;
   assign m237_88 =10'b0;

   // m237_89 = W*in
   wire signed [9:0] m237_89;
   assign m237_89 =10'b0;

   // m237_90 = W*in
   wire signed [9:0] m237_90;
   assign m237_90 =10'b0;

   // m237_91 = W*in
   wire signed [9:0] m237_91;
   assign m237_91 =10'b0;

   // m237_92 = W*in
   wire signed [9:0] m237_92;
   assign m237_92 =10'b0;

   // m237_93 = W*in
   wire signed [9:0] m237_93;
   assign m237_93 =10'b0;

   // m237_94 = W*in
   wire signed [9:0] m237_94;
   assign m237_94 =10'b0;

   // m237_95 = W*in
   wire signed [9:0] m237_95;
   assign m237_95 =10'b0;

   // m237_96 = W*in
   wire signed [9:0] m237_96;
   assign m237_96 =10'b0;

   // m237_97 = W*in
   wire signed [9:0] m237_97;
   assign m237_97 ={ {4{in237[5]}} , in237[5:0] };

   // m237_98 = W*in
   wire signed [9:0] m237_98;
   assign m237_98 =10'b0;

   // m237_99 = W*in
   wire signed [9:0] m237_99;
   assign m237_99 =10'b0;

   // m237_100 = W*in
   wire signed [9:0] m237_100;
   assign m237_100 =10'b0;

   // m237_101 = W*in
   wire signed [9:0] m237_101;
   assign m237_101 ={ {5{in237[5]}} , in237[5:1] };

   // m237_102 = W*in
   wire signed [9:0] m237_102;
   assign m237_102 =10'b0;

   // m237_103 = W*in
   wire signed [9:0] m237_103;
   assign m237_103 =10'b0;

   // m237_104 = W*in
   wire signed [9:0] m237_104;
   assign m237_104 =10'b0;

   // m237_105 = W*in
   wire signed [9:0] m237_105;
   assign m237_105 =10'b0;

   // m237_106 = W*in
   wire signed [9:0] m237_106;
   assign m237_106 =10'b0;

   // m237_107 = W*in
   wire signed [9:0] m237_107;
   assign m237_107 =10'b0;

   // m237_108 = W*in
   wire signed [9:0] m237_108;
   assign m237_108 =10'b0;

   // m237_109 = W*in
   wire signed [9:0] m237_109;
   assign m237_109 ={ {4{neg237[5]}} , neg237[5:0] };

   // m237_110 = W*in
   wire signed [9:0] m237_110;
   assign m237_110 =10'b0;

   // m237_111 = W*in
   wire signed [9:0] m237_111;
   assign m237_111 =10'b0;

   // m237_112 = W*in
   wire signed [9:0] m237_112;
   assign m237_112 =10'b0;

   // m237_113 = W*in
   wire signed [9:0] m237_113;
   assign m237_113 =10'b0;

   // m237_114 = W*in
   wire signed [9:0] m237_114;
   assign m237_114 ={ {5{neg237[5]}} , neg237[5:1] };

   // m237_115 = W*in
   wire signed [9:0] m237_115;
   assign m237_115 ={ {5{neg237[5]}} , neg237[5:1] };

   // m237_116 = W*in
   wire signed [9:0] m237_116;
   assign m237_116 =10'b0;

   // m237_117 = W*in
   wire signed [9:0] m237_117;
   assign m237_117 =10'b0;

   // m238_1 = W*in
   wire signed [9:0] m238_1;
   assign m238_1 =10'b0;

   // m238_2 = W*in
   wire signed [9:0] m238_2;
   assign m238_2 =10'b0;

   // m238_3 = W*in
   wire signed [9:0] m238_3;
   assign m238_3 =10'b0;

   // m238_4 = W*in
   wire signed [9:0] m238_4;
   assign m238_4 =10'b0;

   // m238_5 = W*in
   wire signed [9:0] m238_5;
   assign m238_5 =10'b0;

   // m238_6 = W*in
   wire signed [9:0] m238_6;
   assign m238_6 =10'b0;

   // m238_7 = W*in
   wire signed [9:0] m238_7;
   assign m238_7 =10'b0;

   // m238_8 = W*in
   wire signed [9:0] m238_8;
   assign m238_8 =10'b0;

   // m238_9 = W*in
   wire signed [9:0] m238_9;
   assign m238_9 =10'b0;

   // m238_10 = W*in
   wire signed [9:0] m238_10;
   assign m238_10 =10'b0;

   // m238_11 = W*in
   wire signed [9:0] m238_11;
   assign m238_11 =10'b0;

   // m238_12 = W*in
   wire signed [9:0] m238_12;
   assign m238_12 =10'b0;

   // m238_13 = W*in
   wire signed [9:0] m238_13;
   assign m238_13 =10'b0;

   // m238_14 = W*in
   wire signed [9:0] m238_14;
   assign m238_14 =10'b0;

   // m238_15 = W*in
   wire signed [9:0] m238_15;
   assign m238_15 =10'b0;

   // m238_16 = W*in
   wire signed [9:0] m238_16;
   assign m238_16 =10'b0;

   // m238_17 = W*in
   wire signed [9:0] m238_17;
   assign m238_17 =10'b0;

   // m238_18 = W*in
   wire signed [9:0] m238_18;
   assign m238_18 =10'b0;

   // m238_19 = W*in
   wire signed [9:0] m238_19;
   assign m238_19 =10'b0;

   // m238_20 = W*in
   wire signed [9:0] m238_20;
   assign m238_20 =10'b0;

   // m238_21 = W*in
   wire signed [9:0] m238_21;
   assign m238_21 =10'b0;

   // m238_22 = W*in
   wire signed [9:0] m238_22;
   assign m238_22 =10'b0;

   // m238_23 = W*in
   wire signed [9:0] m238_23;
   assign m238_23 =10'b0;

   // m238_24 = W*in
   wire signed [9:0] m238_24;
   assign m238_24 =10'b0;

   // m238_25 = W*in
   wire signed [9:0] m238_25;
   assign m238_25 =10'b0;

   // m238_26 = W*in
   wire signed [9:0] m238_26;
   assign m238_26 =10'b0;

   // m238_27 = W*in
   wire signed [9:0] m238_27;
   assign m238_27 =10'b0;

   // m238_28 = W*in
   wire signed [9:0] m238_28;
   assign m238_28 =10'b0;

   // m238_29 = W*in
   wire signed [9:0] m238_29;
   assign m238_29 =10'b0;

   // m238_30 = W*in
   wire signed [9:0] m238_30;
   assign m238_30 =10'b0;

   // m238_31 = W*in
   wire signed [9:0] m238_31;
   assign m238_31 =10'b0;

   // m238_32 = W*in
   wire signed [9:0] m238_32;
   assign m238_32 =10'b0;

   // m238_33 = W*in
   wire signed [9:0] m238_33;
   assign m238_33 =10'b0;

   // m238_34 = W*in
   wire signed [9:0] m238_34;
   assign m238_34 =10'b0;

   // m238_35 = W*in
   wire signed [9:0] m238_35;
   assign m238_35 =10'b0;

   // m238_36 = W*in
   wire signed [9:0] m238_36;
   assign m238_36 =10'b0;

   // m238_37 = W*in
   wire signed [9:0] m238_37;
   assign m238_37 =10'b0;

   // m238_38 = W*in
   wire signed [9:0] m238_38;
   assign m238_38 =10'b0;

   // m238_39 = W*in
   wire signed [9:0] m238_39;
   assign m238_39 =10'b0;

   // m238_40 = W*in
   wire signed [9:0] m238_40;
   assign m238_40 =10'b0;

   // m238_41 = W*in
   wire signed [9:0] m238_41;
   assign m238_41 =10'b0;

   // m238_42 = W*in
   wire signed [9:0] m238_42;
   assign m238_42 =10'b0;

   // m238_43 = W*in
   wire signed [9:0] m238_43;
   assign m238_43 =10'b0;

   // m238_44 = W*in
   wire signed [9:0] m238_44;
   assign m238_44 =10'b0;

   // m238_45 = W*in
   wire signed [9:0] m238_45;
   assign m238_45 =10'b0;

   // m238_46 = W*in
   wire signed [9:0] m238_46;
   assign m238_46 =10'b0;

   // m238_47 = W*in
   wire signed [9:0] m238_47;
   assign m238_47 =10'b0;

   // m238_48 = W*in
   wire signed [9:0] m238_48;
   assign m238_48 =10'b0;

   // m238_49 = W*in
   wire signed [9:0] m238_49;
   assign m238_49 =10'b0;

   // m238_50 = W*in
   wire signed [9:0] m238_50;
   assign m238_50 =10'b0;

   // m238_51 = W*in
   wire signed [9:0] m238_51;
   assign m238_51 =10'b0;

   // m238_52 = W*in
   wire signed [9:0] m238_52;
   assign m238_52 =10'b0;

   // m238_53 = W*in
   wire signed [9:0] m238_53;
   assign m238_53 =10'b0;

   // m238_54 = W*in
   wire signed [9:0] m238_54;
   assign m238_54 =10'b0;

   // m238_55 = W*in
   wire signed [9:0] m238_55;
   assign m238_55 =10'b0;

   // m238_56 = W*in
   wire signed [9:0] m238_56;
   assign m238_56 =10'b0;

   // m238_57 = W*in
   wire signed [9:0] m238_57;
   assign m238_57 =10'b0;

   // m238_58 = W*in
   wire signed [9:0] m238_58;
   assign m238_58 =10'b0;

   // m238_59 = W*in
   wire signed [9:0] m238_59;
   assign m238_59 =10'b0;

   // m238_60 = W*in
   wire signed [9:0] m238_60;
   assign m238_60 =10'b0;

   // m238_61 = W*in
   wire signed [9:0] m238_61;
   assign m238_61 =10'b0;

   // m238_62 = W*in
   wire signed [9:0] m238_62;
   assign m238_62 =10'b0;

   // m238_63 = W*in
   wire signed [9:0] m238_63;
   assign m238_63 =10'b0;

   // m238_64 = W*in
   wire signed [9:0] m238_64;
   assign m238_64 ={ {5{in238[5]}} , in238[5:1] };

   // m238_65 = W*in
   wire signed [9:0] m238_65;
   assign m238_65 =10'b0;

   // m238_66 = W*in
   wire signed [9:0] m238_66;
   assign m238_66 =10'b0;

   // m238_67 = W*in
   wire signed [9:0] m238_67;
   assign m238_67 =10'b0;

   // m238_68 = W*in
   wire signed [9:0] m238_68;
   assign m238_68 =10'b0;

   // m238_69 = W*in
   wire signed [9:0] m238_69;
   assign m238_69 =10'b0;

   // m238_70 = W*in
   wire signed [9:0] m238_70;
   assign m238_70 =10'b0;

   // m238_71 = W*in
   wire signed [9:0] m238_71;
   assign m238_71 =10'b0;

   // m238_72 = W*in
   wire signed [9:0] m238_72;
   assign m238_72 =10'b0;

   // m238_73 = W*in
   wire signed [9:0] m238_73;
   assign m238_73 =10'b0;

   // m238_74 = W*in
   wire signed [9:0] m238_74;
   assign m238_74 =10'b0;

   // m238_75 = W*in
   wire signed [9:0] m238_75;
   assign m238_75 =10'b0;

   // m238_76 = W*in
   wire signed [9:0] m238_76;
   assign m238_76 =10'b0;

   // m238_77 = W*in
   wire signed [9:0] m238_77;
   assign m238_77 =10'b0;

   // m238_78 = W*in
   wire signed [9:0] m238_78;
   assign m238_78 =10'b0;

   // m238_79 = W*in
   wire signed [9:0] m238_79;
   assign m238_79 =10'b0;

   // m238_80 = W*in
   wire signed [9:0] m238_80;
   assign m238_80 =10'b0;

   // m238_81 = W*in
   wire signed [9:0] m238_81;
   assign m238_81 =10'b0;

   // m238_82 = W*in
   wire signed [9:0] m238_82;
   assign m238_82 =10'b0;

   // m238_83 = W*in
   wire signed [9:0] m238_83;
   assign m238_83 =10'b0;

   // m238_84 = W*in
   wire signed [9:0] m238_84;
   assign m238_84 =10'b0;

   // m238_85 = W*in
   wire signed [9:0] m238_85;
   assign m238_85 =10'b0;

   // m238_86 = W*in
   wire signed [9:0] m238_86;
   assign m238_86 =10'b0;

   // m238_87 = W*in
   wire signed [9:0] m238_87;
   assign m238_87 =10'b0;

   // m238_88 = W*in
   wire signed [9:0] m238_88;
   assign m238_88 =10'b0;

   // m238_89 = W*in
   wire signed [9:0] m238_89;
   assign m238_89 =10'b0;

   // m238_90 = W*in
   wire signed [9:0] m238_90;
   assign m238_90 =10'b0;

   // m238_91 = W*in
   wire signed [9:0] m238_91;
   assign m238_91 =10'b0;

   // m238_92 = W*in
   wire signed [9:0] m238_92;
   assign m238_92 =10'b0;

   // m238_93 = W*in
   wire signed [9:0] m238_93;
   assign m238_93 =10'b0;

   // m238_94 = W*in
   wire signed [9:0] m238_94;
   assign m238_94 =10'b0;

   // m238_95 = W*in
   wire signed [9:0] m238_95;
   assign m238_95 =10'b0;

   // m238_96 = W*in
   wire signed [9:0] m238_96;
   assign m238_96 =10'b0;

   // m238_97 = W*in
   wire signed [9:0] m238_97;
   assign m238_97 =10'b0;

   // m238_98 = W*in
   wire signed [9:0] m238_98;
   assign m238_98 =10'b0;

   // m238_99 = W*in
   wire signed [9:0] m238_99;
   assign m238_99 =10'b0;

   // m238_100 = W*in
   wire signed [9:0] m238_100;
   assign m238_100 =10'b0;

   // m238_101 = W*in
   wire signed [9:0] m238_101;
   assign m238_101 =10'b0;

   // m238_102 = W*in
   wire signed [9:0] m238_102;
   assign m238_102 =10'b0;

   // m238_103 = W*in
   wire signed [9:0] m238_103;
   assign m238_103 =10'b0;

   // m238_104 = W*in
   wire signed [9:0] m238_104;
   assign m238_104 =10'b0;

   // m238_105 = W*in
   wire signed [9:0] m238_105;
   assign m238_105 =10'b0;

   // m238_106 = W*in
   wire signed [9:0] m238_106;
   assign m238_106 =10'b0;

   // m238_107 = W*in
   wire signed [9:0] m238_107;
   assign m238_107 =10'b0;

   // m238_108 = W*in
   wire signed [9:0] m238_108;
   assign m238_108 =10'b0;

   // m238_109 = W*in
   wire signed [9:0] m238_109;
   assign m238_109 =10'b0;

   // m238_110 = W*in
   wire signed [9:0] m238_110;
   assign m238_110 =10'b0;

   // m238_111 = W*in
   wire signed [9:0] m238_111;
   assign m238_111 =10'b0;

   // m238_112 = W*in
   wire signed [9:0] m238_112;
   assign m238_112 =10'b0;

   // m238_113 = W*in
   wire signed [9:0] m238_113;
   assign m238_113 =10'b0;

   // m238_114 = W*in
   wire signed [9:0] m238_114;
   assign m238_114 =10'b0;

   // m238_115 = W*in
   wire signed [9:0] m238_115;
   assign m238_115 =10'b0;

   // m238_116 = W*in
   wire signed [9:0] m238_116;
   assign m238_116 =10'b0;

   // m238_117 = W*in
   wire signed [9:0] m238_117;
   assign m238_117 =10'b0;

   // m239_1 = W*in
   wire signed [9:0] m239_1;
   assign m239_1 =10'b0;

   // m239_2 = W*in
   wire signed [9:0] m239_2;
   assign m239_2 =10'b0;

   // m239_3 = W*in
   wire signed [9:0] m239_3;
   assign m239_3 =10'b0;

   // m239_4 = W*in
   wire signed [9:0] m239_4;
   assign m239_4 =10'b0;

   // m239_5 = W*in
   wire signed [9:0] m239_5;
   assign m239_5 ={ {4{in239[5]}} , in239[5:0] };

   // m239_6 = W*in
   wire signed [9:0] m239_6;
   assign m239_6 =10'b0;

   // m239_7 = W*in
   wire signed [9:0] m239_7;
   assign m239_7 =10'b0;

   // m239_8 = W*in
   wire signed [9:0] m239_8;
   assign m239_8 =10'b0;

   // m239_9 = W*in
   wire signed [9:0] m239_9;
   assign m239_9 =10'b0;

   // m239_10 = W*in
   wire signed [9:0] m239_10;
   assign m239_10 =10'b0;

   // m239_11 = W*in
   wire signed [9:0] m239_11;
   assign m239_11 =10'b0;

   // m239_12 = W*in
   wire signed [9:0] m239_12;
   assign m239_12 =10'b0;

   // m239_13 = W*in
   wire signed [9:0] m239_13;
   assign m239_13 =10'b0;

   // m239_14 = W*in
   wire signed [9:0] m239_14;
   assign m239_14 =10'b0;

   // m239_15 = W*in
   wire signed [9:0] m239_15;
   assign m239_15 =10'b0;

   // m239_16 = W*in
   wire signed [9:0] m239_16;
   assign m239_16 =10'b0;

   // m239_17 = W*in
   wire signed [9:0] m239_17;
   assign m239_17 =10'b0;

   // m239_18 = W*in
   wire signed [9:0] m239_18;
   assign m239_18 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_19 = W*in
   wire signed [9:0] m239_19;
   assign m239_19 ={ {5{in239[5]}} , in239[5:1] };

   // m239_20 = W*in
   wire signed [9:0] m239_20;
   assign m239_20 =10'b0;

   // m239_21 = W*in
   wire signed [9:0] m239_21;
   assign m239_21 =10'b0;

   // m239_22 = W*in
   wire signed [9:0] m239_22;
   assign m239_22 =10'b0;

   // m239_23 = W*in
   wire signed [9:0] m239_23;
   assign m239_23 =10'b0;

   // m239_24 = W*in
   wire signed [9:0] m239_24;
   assign m239_24 =10'b0;

   // m239_25 = W*in
   wire signed [9:0] m239_25;
   assign m239_25 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_26 = W*in
   wire signed [9:0] m239_26;
   assign m239_26 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_27 = W*in
   wire signed [9:0] m239_27;
   assign m239_27 =10'b0;

   // m239_28 = W*in
   wire signed [9:0] m239_28;
   assign m239_28 =10'b0;

   // m239_29 = W*in
   wire signed [9:0] m239_29;
   assign m239_29 =10'b0;

   // m239_30 = W*in
   wire signed [9:0] m239_30;
   assign m239_30 =10'b0;

   // m239_31 = W*in
   wire signed [9:0] m239_31;
   assign m239_31 =10'b0;

   // m239_32 = W*in
   wire signed [9:0] m239_32;
   assign m239_32 =10'b0;

   // m239_33 = W*in
   wire signed [9:0] m239_33;
   assign m239_33 =10'b0;

   // m239_34 = W*in
   wire signed [9:0] m239_34;
   assign m239_34 =10'b0;

   // m239_35 = W*in
   wire signed [9:0] m239_35;
   assign m239_35 =10'b0;

   // m239_36 = W*in
   wire signed [9:0] m239_36;
   assign m239_36 =10'b0;

   // m239_37 = W*in
   wire signed [9:0] m239_37;
   assign m239_37 =10'b0;

   // m239_38 = W*in
   wire signed [9:0] m239_38;
   assign m239_38 =10'b0;

   // m239_39 = W*in
   wire signed [9:0] m239_39;
   assign m239_39 =10'b0;

   // m239_40 = W*in
   wire signed [9:0] m239_40;
   assign m239_40 =10'b0;

   // m239_41 = W*in
   wire signed [9:0] m239_41;
   assign m239_41 =10'b0;

   // m239_42 = W*in
   wire signed [9:0] m239_42;
   assign m239_42 =10'b0;

   // m239_43 = W*in
   wire signed [9:0] m239_43;
   assign m239_43 ={ {4{neg239[5]}} , neg239[5:0] };

   // m239_44 = W*in
   wire signed [9:0] m239_44;
   assign m239_44 =10'b0;

   // m239_45 = W*in
   wire signed [9:0] m239_45;
   assign m239_45 =10'b0;

   // m239_46 = W*in
   wire signed [9:0] m239_46;
   assign m239_46 =10'b0;

   // m239_47 = W*in
   wire signed [9:0] m239_47;
   assign m239_47 =10'b0;

   // m239_48 = W*in
   wire signed [9:0] m239_48;
   assign m239_48 =10'b0;

   // m239_49 = W*in
   wire signed [9:0] m239_49;
   assign m239_49 =10'b0;

   // m239_50 = W*in
   wire signed [9:0] m239_50;
   assign m239_50 =10'b0;

   // m239_51 = W*in
   wire signed [9:0] m239_51;
   assign m239_51 =10'b0;

   // m239_52 = W*in
   wire signed [9:0] m239_52;
   assign m239_52 =10'b0;

   // m239_53 = W*in
   wire signed [9:0] m239_53;
   assign m239_53 =10'b0;

   // m239_54 = W*in
   wire signed [9:0] m239_54;
   assign m239_54 =10'b0;

   // m239_55 = W*in
   wire signed [9:0] m239_55;
   assign m239_55 =10'b0;

   // m239_56 = W*in
   wire signed [9:0] m239_56;
   assign m239_56 =10'b0;

   // m239_57 = W*in
   wire signed [9:0] m239_57;
   assign m239_57 =10'b0;

   // m239_58 = W*in
   wire signed [9:0] m239_58;
   assign m239_58 =10'b0;

   // m239_59 = W*in
   wire signed [9:0] m239_59;
   assign m239_59 =10'b0;

   // m239_60 = W*in
   wire signed [9:0] m239_60;
   assign m239_60 =10'b0;

   // m239_61 = W*in
   wire signed [9:0] m239_61;
   assign m239_61 =10'b0;

   // m239_62 = W*in
   wire signed [9:0] m239_62;
   assign m239_62 =10'b0;

   // m239_63 = W*in
   wire signed [9:0] m239_63;
   assign m239_63 =10'b0;

   // m239_64 = W*in
   wire signed [9:0] m239_64;
   assign m239_64 =10'b0;

   // m239_65 = W*in
   wire signed [9:0] m239_65;
   assign m239_65 ={ {5{in239[5]}} , in239[5:1] };

   // m239_66 = W*in
   wire signed [9:0] m239_66;
   assign m239_66 =10'b0;

   // m239_67 = W*in
   wire signed [9:0] m239_67;
   assign m239_67 ={ {4{in239[5]}} , in239[5:0] };

   // m239_68 = W*in
   wire signed [9:0] m239_68;
   assign m239_68 =10'b0;

   // m239_69 = W*in
   wire signed [9:0] m239_69;
   assign m239_69 =10'b0;

   // m239_70 = W*in
   wire signed [9:0] m239_70;
   assign m239_70 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_71 = W*in
   wire signed [9:0] m239_71;
   assign m239_71 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_72 = W*in
   wire signed [9:0] m239_72;
   assign m239_72 ={ {4{neg239[5]}} , neg239[5:0] };

   // m239_73 = W*in
   wire signed [9:0] m239_73;
   assign m239_73 ={ {5{in239[5]}} , in239[5:1] };

   // m239_74 = W*in
   wire signed [9:0] m239_74;
   assign m239_74 =10'b0;

   // m239_75 = W*in
   wire signed [9:0] m239_75;
   assign m239_75 =10'b0;

   // m239_76 = W*in
   wire signed [9:0] m239_76;
   assign m239_76 =10'b0;

   // m239_77 = W*in
   wire signed [9:0] m239_77;
   assign m239_77 =10'b0;

   // m239_78 = W*in
   wire signed [9:0] m239_78;
   assign m239_78 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_79 = W*in
   wire signed [9:0] m239_79;
   assign m239_79 =10'b0;

   // m239_80 = W*in
   wire signed [9:0] m239_80;
   assign m239_80 =10'b0;

   // m239_81 = W*in
   wire signed [9:0] m239_81;
   assign m239_81 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_82 = W*in
   wire signed [9:0] m239_82;
   assign m239_82 =10'b0;

   // m239_83 = W*in
   wire signed [9:0] m239_83;
   assign m239_83 =10'b0;

   // m239_84 = W*in
   wire signed [9:0] m239_84;
   assign m239_84 =10'b0;

   // m239_85 = W*in
   wire signed [9:0] m239_85;
   assign m239_85 =10'b0;

   // m239_86 = W*in
   wire signed [9:0] m239_86;
   assign m239_86 =10'b0;

   // m239_87 = W*in
   wire signed [9:0] m239_87;
   assign m239_87 =10'b0;

   // m239_88 = W*in
   wire signed [9:0] m239_88;
   assign m239_88 =10'b0;

   // m239_89 = W*in
   wire signed [9:0] m239_89;
   assign m239_89 =10'b0;

   // m239_90 = W*in
   wire signed [9:0] m239_90;
   assign m239_90 =10'b0;

   // m239_91 = W*in
   wire signed [9:0] m239_91;
   assign m239_91 =10'b0;

   // m239_92 = W*in
   wire signed [9:0] m239_92;
   assign m239_92 =10'b0;

   // m239_93 = W*in
   wire signed [9:0] m239_93;
   assign m239_93 =10'b0;

   // m239_94 = W*in
   wire signed [9:0] m239_94;
   assign m239_94 =10'b0;

   // m239_95 = W*in
   wire signed [9:0] m239_95;
   assign m239_95 =10'b0;

   // m239_96 = W*in
   wire signed [9:0] m239_96;
   assign m239_96 =10'b0;

   // m239_97 = W*in
   wire signed [9:0] m239_97;
   assign m239_97 =10'b0;

   // m239_98 = W*in
   wire signed [9:0] m239_98;
   assign m239_98 =10'b0;

   // m239_99 = W*in
   wire signed [9:0] m239_99;
   assign m239_99 ={ {4{neg239[5]}} , neg239[5:0] };

   // m239_100 = W*in
   wire signed [9:0] m239_100;
   assign m239_100 =10'b0;

   // m239_101 = W*in
   wire signed [9:0] m239_101;
   assign m239_101 =10'b0;

   // m239_102 = W*in
   wire signed [9:0] m239_102;
   assign m239_102 =10'b0;

   // m239_103 = W*in
   wire signed [9:0] m239_103;
   assign m239_103 ={ {4{neg239[5]}} , neg239[5:0] };

   // m239_104 = W*in
   wire signed [9:0] m239_104;
   assign m239_104 =10'b0;

   // m239_105 = W*in
   wire signed [9:0] m239_105;
   assign m239_105 ={ {5{in239[5]}} , in239[5:1] };

   // m239_106 = W*in
   wire signed [9:0] m239_106;
   assign m239_106 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_107 = W*in
   wire signed [9:0] m239_107;
   assign m239_107 =10'b0;

   // m239_108 = W*in
   wire signed [9:0] m239_108;
   assign m239_108 ={ {5{neg239[5]}} , neg239[5:1] };

   // m239_109 = W*in
   wire signed [9:0] m239_109;
   assign m239_109 =10'b0;

   // m239_110 = W*in
   wire signed [9:0] m239_110;
   assign m239_110 =10'b0;

   // m239_111 = W*in
   wire signed [9:0] m239_111;
   assign m239_111 =10'b0;

   // m239_112 = W*in
   wire signed [9:0] m239_112;
   assign m239_112 =10'b0;

   // m239_113 = W*in
   wire signed [9:0] m239_113;
   assign m239_113 =10'b0;

   // m239_114 = W*in
   wire signed [9:0] m239_114;
   assign m239_114 =10'b0;

   // m239_115 = W*in
   wire signed [9:0] m239_115;
   assign m239_115 =10'b0;

   // m239_116 = W*in
   wire signed [9:0] m239_116;
   assign m239_116 =10'b0;

   // m239_117 = W*in
   wire signed [9:0] m239_117;
   assign m239_117 =10'b0;

   // m240_1 = W*in
   wire signed [9:0] m240_1;
   assign m240_1 =10'b0;

   // m240_2 = W*in
   wire signed [9:0] m240_2;
   assign m240_2 =10'b0;

   // m240_3 = W*in
   wire signed [9:0] m240_3;
   assign m240_3 =10'b0;

   // m240_4 = W*in
   wire signed [9:0] m240_4;
   assign m240_4 =10'b0;

   // m240_5 = W*in
   wire signed [9:0] m240_5;
   assign m240_5 =10'b0;

   // m240_6 = W*in
   wire signed [9:0] m240_6;
   assign m240_6 =10'b0;

   // m240_7 = W*in
   wire signed [9:0] m240_7;
   assign m240_7 =10'b0;

   // m240_8 = W*in
   wire signed [9:0] m240_8;
   assign m240_8 =10'b0;

   // m240_9 = W*in
   wire signed [9:0] m240_9;
   assign m240_9 =10'b0;

   // m240_10 = W*in
   wire signed [9:0] m240_10;
   assign m240_10 =10'b0;

   // m240_11 = W*in
   wire signed [9:0] m240_11;
   assign m240_11 =10'b0;

   // m240_12 = W*in
   wire signed [9:0] m240_12;
   assign m240_12 =10'b0;

   // m240_13 = W*in
   wire signed [9:0] m240_13;
   assign m240_13 =10'b0;

   // m240_14 = W*in
   wire signed [9:0] m240_14;
   assign m240_14 =10'b0;

   // m240_15 = W*in
   wire signed [9:0] m240_15;
   assign m240_15 =10'b0;

   // m240_16 = W*in
   wire signed [9:0] m240_16;
   assign m240_16 =10'b0;

   // m240_17 = W*in
   wire signed [9:0] m240_17;
   assign m240_17 ={ {5{in240[5]}} , in240[5:1] };

   // m240_18 = W*in
   wire signed [9:0] m240_18;
   assign m240_18 =10'b0;

   // m240_19 = W*in
   wire signed [9:0] m240_19;
   assign m240_19 ={ {5{in240[5]}} , in240[5:1] };

   // m240_20 = W*in
   wire signed [9:0] m240_20;
   assign m240_20 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_21 = W*in
   wire signed [9:0] m240_21;
   assign m240_21 =10'b0;

   // m240_22 = W*in
   wire signed [9:0] m240_22;
   assign m240_22 =10'b0;

   // m240_23 = W*in
   wire signed [9:0] m240_23;
   assign m240_23 =10'b0;

   // m240_24 = W*in
   wire signed [9:0] m240_24;
   assign m240_24 =10'b0;

   // m240_25 = W*in
   wire signed [9:0] m240_25;
   assign m240_25 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_26 = W*in
   wire signed [9:0] m240_26;
   assign m240_26 =10'b0;

   // m240_27 = W*in
   wire signed [9:0] m240_27;
   assign m240_27 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_28 = W*in
   wire signed [9:0] m240_28;
   assign m240_28 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_29 = W*in
   wire signed [9:0] m240_29;
   assign m240_29 =10'b0;

   // m240_30 = W*in
   wire signed [9:0] m240_30;
   assign m240_30 =10'b0;

   // m240_31 = W*in
   wire signed [9:0] m240_31;
   assign m240_31 =10'b0;

   // m240_32 = W*in
   wire signed [9:0] m240_32;
   assign m240_32 =10'b0;

   // m240_33 = W*in
   wire signed [9:0] m240_33;
   assign m240_33 =10'b0;

   // m240_34 = W*in
   wire signed [9:0] m240_34;
   assign m240_34 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_35 = W*in
   wire signed [9:0] m240_35;
   assign m240_35 =10'b0;

   // m240_36 = W*in
   wire signed [9:0] m240_36;
   assign m240_36 =10'b0;

   // m240_37 = W*in
   wire signed [9:0] m240_37;
   assign m240_37 =10'b0;

   // m240_38 = W*in
   wire signed [9:0] m240_38;
   assign m240_38 =10'b0;

   // m240_39 = W*in
   wire signed [9:0] m240_39;
   assign m240_39 =10'b0;

   // m240_40 = W*in
   wire signed [9:0] m240_40;
   assign m240_40 =10'b0;

   // m240_41 = W*in
   wire signed [9:0] m240_41;
   assign m240_41 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_42 = W*in
   wire signed [9:0] m240_42;
   assign m240_42 =10'b0;

   // m240_43 = W*in
   wire signed [9:0] m240_43;
   assign m240_43 =10'b0;

   // m240_44 = W*in
   wire signed [9:0] m240_44;
   assign m240_44 =10'b0;

   // m240_45 = W*in
   wire signed [9:0] m240_45;
   assign m240_45 =10'b0;

   // m240_46 = W*in
   wire signed [9:0] m240_46;
   assign m240_46 =10'b0;

   // m240_47 = W*in
   wire signed [9:0] m240_47;
   assign m240_47 =10'b0;

   // m240_48 = W*in
   wire signed [9:0] m240_48;
   assign m240_48 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_49 = W*in
   wire signed [9:0] m240_49;
   assign m240_49 =10'b0;

   // m240_50 = W*in
   wire signed [9:0] m240_50;
   assign m240_50 =10'b0;

   // m240_51 = W*in
   wire signed [9:0] m240_51;
   assign m240_51 =10'b0;

   // m240_52 = W*in
   wire signed [9:0] m240_52;
   assign m240_52 =10'b0;

   // m240_53 = W*in
   wire signed [9:0] m240_53;
   assign m240_53 =10'b0;

   // m240_54 = W*in
   wire signed [9:0] m240_54;
   assign m240_54 =10'b0;

   // m240_55 = W*in
   wire signed [9:0] m240_55;
   assign m240_55 =10'b0;

   // m240_56 = W*in
   wire signed [9:0] m240_56;
   assign m240_56 =10'b0;

   // m240_57 = W*in
   wire signed [9:0] m240_57;
   assign m240_57 =10'b0;

   // m240_58 = W*in
   wire signed [9:0] m240_58;
   assign m240_58 =10'b0;

   // m240_59 = W*in
   wire signed [9:0] m240_59;
   assign m240_59 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_60 = W*in
   wire signed [9:0] m240_60;
   assign m240_60 =10'b0;

   // m240_61 = W*in
   wire signed [9:0] m240_61;
   assign m240_61 =10'b0;

   // m240_62 = W*in
   wire signed [9:0] m240_62;
   assign m240_62 =10'b0;

   // m240_63 = W*in
   wire signed [9:0] m240_63;
   assign m240_63 =10'b0;

   // m240_64 = W*in
   wire signed [9:0] m240_64;
   assign m240_64 =10'b0;

   // m240_65 = W*in
   wire signed [9:0] m240_65;
   assign m240_65 =10'b0;

   // m240_66 = W*in
   wire signed [9:0] m240_66;
   assign m240_66 =10'b0;

   // m240_67 = W*in
   wire signed [9:0] m240_67;
   assign m240_67 =10'b0;

   // m240_68 = W*in
   wire signed [9:0] m240_68;
   assign m240_68 =10'b0;

   // m240_69 = W*in
   wire signed [9:0] m240_69;
   assign m240_69 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_70 = W*in
   wire signed [9:0] m240_70;
   assign m240_70 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_71 = W*in
   wire signed [9:0] m240_71;
   assign m240_71 =10'b0;

   // m240_72 = W*in
   wire signed [9:0] m240_72;
   assign m240_72 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_73 = W*in
   wire signed [9:0] m240_73;
   assign m240_73 =10'b0;

   // m240_74 = W*in
   wire signed [9:0] m240_74;
   assign m240_74 =10'b0;

   // m240_75 = W*in
   wire signed [9:0] m240_75;
   assign m240_75 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_76 = W*in
   wire signed [9:0] m240_76;
   assign m240_76 =10'b0;

   // m240_77 = W*in
   wire signed [9:0] m240_77;
   assign m240_77 ={ {4{in240[5]}} , in240[5:0] };

   // m240_78 = W*in
   wire signed [9:0] m240_78;
   assign m240_78 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_79 = W*in
   wire signed [9:0] m240_79;
   assign m240_79 =10'b0;

   // m240_80 = W*in
   wire signed [9:0] m240_80;
   assign m240_80 =10'b0;

   // m240_81 = W*in
   wire signed [9:0] m240_81;
   assign m240_81 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_82 = W*in
   wire signed [9:0] m240_82;
   assign m240_82 =10'b0;

   // m240_83 = W*in
   wire signed [9:0] m240_83;
   assign m240_83 ={ {5{in240[5]}} , in240[5:1] };

   // m240_84 = W*in
   wire signed [9:0] m240_84;
   assign m240_84 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_85 = W*in
   wire signed [9:0] m240_85;
   assign m240_85 =10'b0;

   // m240_86 = W*in
   wire signed [9:0] m240_86;
   assign m240_86 =10'b0;

   // m240_87 = W*in
   wire signed [9:0] m240_87;
   assign m240_87 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_88 = W*in
   wire signed [9:0] m240_88;
   assign m240_88 =10'b0;

   // m240_89 = W*in
   wire signed [9:0] m240_89;
   assign m240_89 =10'b0;

   // m240_90 = W*in
   wire signed [9:0] m240_90;
   assign m240_90 =10'b0;

   // m240_91 = W*in
   wire signed [9:0] m240_91;
   assign m240_91 =10'b0;

   // m240_92 = W*in
   wire signed [9:0] m240_92;
   assign m240_92 =10'b0;

   // m240_93 = W*in
   wire signed [9:0] m240_93;
   assign m240_93 =10'b0;

   // m240_94 = W*in
   wire signed [9:0] m240_94;
   assign m240_94 =10'b0;

   // m240_95 = W*in
   wire signed [9:0] m240_95;
   assign m240_95 ={ {5{in240[5]}} , in240[5:1] };

   // m240_96 = W*in
   wire signed [9:0] m240_96;
   assign m240_96 =10'b0;

   // m240_97 = W*in
   wire signed [9:0] m240_97;
   assign m240_97 =10'b0;

   // m240_98 = W*in
   wire signed [9:0] m240_98;
   assign m240_98 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_99 = W*in
   wire signed [9:0] m240_99;
   assign m240_99 =10'b0;

   // m240_100 = W*in
   wire signed [9:0] m240_100;
   assign m240_100 =10'b0;

   // m240_101 = W*in
   wire signed [9:0] m240_101;
   assign m240_101 =10'b0;

   // m240_102 = W*in
   wire signed [9:0] m240_102;
   assign m240_102 =10'b0;

   // m240_103 = W*in
   wire signed [9:0] m240_103;
   assign m240_103 =10'b0;

   // m240_104 = W*in
   wire signed [9:0] m240_104;
   assign m240_104 =10'b0;

   // m240_105 = W*in
   wire signed [9:0] m240_105;
   assign m240_105 =10'b0;

   // m240_106 = W*in
   wire signed [9:0] m240_106;
   assign m240_106 ={ {5{neg240[5]}} , neg240[5:1] };

   // m240_107 = W*in
   wire signed [9:0] m240_107;
   assign m240_107 ={ {4{in240[5]}} , in240[5:0] };

   // m240_108 = W*in
   wire signed [9:0] m240_108;
   assign m240_108 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_109 = W*in
   wire signed [9:0] m240_109;
   assign m240_109 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_110 = W*in
   wire signed [9:0] m240_110;
   assign m240_110 =10'b0;

   // m240_111 = W*in
   wire signed [9:0] m240_111;
   assign m240_111 ={ {4{neg240[5]}} , neg240[5:0] };

   // m240_112 = W*in
   wire signed [9:0] m240_112;
   assign m240_112 =10'b0;

   // m240_113 = W*in
   wire signed [9:0] m240_113;
   assign m240_113 =10'b0;

   // m240_114 = W*in
   wire signed [9:0] m240_114;
   assign m240_114 =10'b0;

   // m240_115 = W*in
   wire signed [9:0] m240_115;
   assign m240_115 =10'b0;

   // m240_116 = W*in
   wire signed [9:0] m240_116;
   assign m240_116 =10'b0;

   // m240_117 = W*in
   wire signed [9:0] m240_117;
   assign m240_117 =10'b0;

   // m241_1 = W*in
   wire signed [9:0] m241_1;
   assign m241_1 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_2 = W*in
   wire signed [9:0] m241_2;
   assign m241_2 ={ {4{in241[5]}} , in241[5:0] };

   // m241_3 = W*in
   wire signed [9:0] m241_3;
   assign m241_3 ={ {4{in241[5]}} , in241[5:0] };

   // m241_4 = W*in
   wire signed [9:0] m241_4;
   assign m241_4 =10'b0;

   // m241_5 = W*in
   wire signed [9:0] m241_5;
   assign m241_5 =10'b0;

   // m241_6 = W*in
   wire signed [9:0] m241_6;
   assign m241_6 ={ {5{in241[5]}} , in241[5:1] };

   // m241_7 = W*in
   wire signed [9:0] m241_7;
   assign m241_7 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_8 = W*in
   wire signed [9:0] m241_8;
   assign m241_8 ={ {3{in241[5]}} , in241 , {1{1'b0}} };

   // m241_9 = W*in
   wire signed [9:0] m241_9;
   assign m241_9 =10'b0;

   // m241_10 = W*in
   wire signed [9:0] m241_10;
   assign m241_10 =10'b0;

   // m241_11 = W*in
   wire signed [9:0] m241_11;
   assign m241_11 =10'b0;

   // m241_12 = W*in
   wire signed [9:0] m241_12;
   assign m241_12 ={ {4{in241[5]}} , in241[5:0] };

   // m241_13 = W*in
   wire signed [9:0] m241_13;
   assign m241_13 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_14 = W*in
   wire signed [9:0] m241_14;
   assign m241_14 =10'b0;

   // m241_15 = W*in
   wire signed [9:0] m241_15;
   assign m241_15 =10'b0;

   // m241_16 = W*in
   wire signed [9:0] m241_16;
   assign m241_16 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_17 = W*in
   wire signed [9:0] m241_17;
   assign m241_17 ={ {4{in241[5]}} , in241[5:0] };

   // m241_18 = W*in
   wire signed [9:0] m241_18;
   assign m241_18 =10'b0;

   // m241_19 = W*in
   wire signed [9:0] m241_19;
   assign m241_19 ={ {4{in241[5]}} , in241[5:0] };

   // m241_20 = W*in
   wire signed [9:0] m241_20;
   assign m241_20 ={ {5{neg241[5]}} , neg241[5:1] };

   // m241_21 = W*in
   wire signed [9:0] m241_21;
   assign m241_21 =10'b0;

   // m241_22 = W*in
   wire signed [9:0] m241_22;
   assign m241_22 =10'b0;

   // m241_23 = W*in
   wire signed [9:0] m241_23;
   assign m241_23 =10'b0;

   // m241_24 = W*in
   wire signed [9:0] m241_24;
   assign m241_24 =10'b0;

   // m241_25 = W*in
   wire signed [9:0] m241_25;
   assign m241_25 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_26 = W*in
   wire signed [9:0] m241_26;
   assign m241_26 =10'b0;

   // m241_27 = W*in
   wire signed [9:0] m241_27;
   assign m241_27 ={ {5{in241[5]}} , in241[5:1] };

   // m241_28 = W*in
   wire signed [9:0] m241_28;
   assign m241_28 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_29 = W*in
   wire signed [9:0] m241_29;
   assign m241_29 =10'b0;

   // m241_30 = W*in
   wire signed [9:0] m241_30;
   assign m241_30 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_31 = W*in
   wire signed [9:0] m241_31;
   assign m241_31 ={ {4{in241[5]}} , in241[5:0] };

   // m241_32 = W*in
   wire signed [9:0] m241_32;
   assign m241_32 =10'b0;

   // m241_33 = W*in
   wire signed [9:0] m241_33;
   assign m241_33 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_34 = W*in
   wire signed [9:0] m241_34;
   assign m241_34 ={ {4{in241[5]}} , in241[5:0] };

   // m241_35 = W*in
   wire signed [9:0] m241_35;
   assign m241_35 =10'b0;

   // m241_36 = W*in
   wire signed [9:0] m241_36;
   assign m241_36 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_37 = W*in
   wire signed [9:0] m241_37;
   assign m241_37 ={ {4{in241[5]}} , in241[5:0] };

   // m241_38 = W*in
   wire signed [9:0] m241_38;
   assign m241_38 ={ {4{in241[5]}} , in241[5:0] };

   // m241_39 = W*in
   wire signed [9:0] m241_39;
   assign m241_39 =10'b0;

   // m241_40 = W*in
   wire signed [9:0] m241_40;
   assign m241_40 =10'b0;

   // m241_41 = W*in
   wire signed [9:0] m241_41;
   assign m241_41 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_42 = W*in
   wire signed [9:0] m241_42;
   assign m241_42 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_43 = W*in
   wire signed [9:0] m241_43;
   assign m241_43 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_44 = W*in
   wire signed [9:0] m241_44;
   assign m241_44 =10'b0;

   // m241_45 = W*in
   wire signed [9:0] m241_45;
   assign m241_45 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_46 = W*in
   wire signed [9:0] m241_46;
   assign m241_46 =10'b0;

   // m241_47 = W*in
   wire signed [9:0] m241_47;
   assign m241_47 =10'b0;

   // m241_48 = W*in
   wire signed [9:0] m241_48;
   assign m241_48 =10'b0;

   // m241_49 = W*in
   wire signed [9:0] m241_49;
   assign m241_49 =10'b0;

   // m241_50 = W*in
   wire signed [9:0] m241_50;
   assign m241_50 ={ {4{in241[5]}} , in241[5:0] };

   // m241_51 = W*in
   wire signed [9:0] m241_51;
   assign m241_51 =10'b0;

   // m241_52 = W*in
   wire signed [9:0] m241_52;
   assign m241_52 ={ {3{in241[5]}} , in241 , {1{1'b0}} };

   // m241_53 = W*in
   wire signed [9:0] m241_53;
   assign m241_53 ={ {4{in241[5]}} , in241[5:0] };

   // m241_54 = W*in
   wire signed [9:0] m241_54;
   assign m241_54 =10'b0;

   // m241_55 = W*in
   wire signed [9:0] m241_55;
   assign m241_55 =10'b0;

   // m241_56 = W*in
   wire signed [9:0] m241_56;
   assign m241_56 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_57 = W*in
   wire signed [9:0] m241_57;
   assign m241_57 =10'b0;

   // m241_58 = W*in
   wire signed [9:0] m241_58;
   assign m241_58 ={ {5{in241[5]}} , in241[5:1] };

   // m241_59 = W*in
   wire signed [9:0] m241_59;
   assign m241_59 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_60 = W*in
   wire signed [9:0] m241_60;
   assign m241_60 =10'b0;

   // m241_61 = W*in
   wire signed [9:0] m241_61;
   assign m241_61 =10'b0;

   // m241_62 = W*in
   wire signed [9:0] m241_62;
   assign m241_62 =10'b0;

   // m241_63 = W*in
   wire signed [9:0] m241_63;
   assign m241_63 ={ {4{in241[5]}} , in241[5:0] };

   // m241_64 = W*in
   wire signed [9:0] m241_64;
   assign m241_64 =10'b0;

   // m241_65 = W*in
   wire signed [9:0] m241_65;
   assign m241_65 =10'b0;

   // m241_66 = W*in
   wire signed [9:0] m241_66;
   assign m241_66 =10'b0;

   // m241_67 = W*in
   wire signed [9:0] m241_67;
   assign m241_67 ={ {4{in241[5]}} , in241[5:0] };

   // m241_68 = W*in
   wire signed [9:0] m241_68;
   assign m241_68 =10'b0;

   // m241_69 = W*in
   wire signed [9:0] m241_69;
   assign m241_69 =10'b0;

   // m241_70 = W*in
   wire signed [9:0] m241_70;
   assign m241_70 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_71 = W*in
   wire signed [9:0] m241_71;
   assign m241_71 =10'b0;

   // m241_72 = W*in
   wire signed [9:0] m241_72;
   assign m241_72 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_73 = W*in
   wire signed [9:0] m241_73;
   assign m241_73 ={ {5{in241[5]}} , in241[5:1] };

   // m241_74 = W*in
   wire signed [9:0] m241_74;
   assign m241_74 =10'b0;

   // m241_75 = W*in
   wire signed [9:0] m241_75;
   assign m241_75 ={ {5{neg241[5]}} , neg241[5:1] };

   // m241_76 = W*in
   wire signed [9:0] m241_76;
   assign m241_76 =10'b0;

   // m241_77 = W*in
   wire signed [9:0] m241_77;
   assign m241_77 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_78 = W*in
   wire signed [9:0] m241_78;
   assign m241_78 =10'b0;

   // m241_79 = W*in
   wire signed [9:0] m241_79;
   assign m241_79 =10'b0;

   // m241_80 = W*in
   wire signed [9:0] m241_80;
   assign m241_80 ={ {4{in241[5]}} , in241[5:0] };

   // m241_81 = W*in
   wire signed [9:0] m241_81;
   assign m241_81 =10'b0;

   // m241_82 = W*in
   wire signed [9:0] m241_82;
   assign m241_82 ={ {3{in241[5]}} , in241 , {1{1'b0}} };

   // m241_83 = W*in
   wire signed [9:0] m241_83;
   assign m241_83 ={ {5{neg241[5]}} , neg241[5:1] };

   // m241_84 = W*in
   wire signed [9:0] m241_84;
   assign m241_84 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_85 = W*in
   wire signed [9:0] m241_85;
   assign m241_85 =10'b0;

   // m241_86 = W*in
   wire signed [9:0] m241_86;
   assign m241_86 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_87 = W*in
   wire signed [9:0] m241_87;
   assign m241_87 =10'b0;

   // m241_88 = W*in
   wire signed [9:0] m241_88;
   assign m241_88 ={ {4{in241[5]}} , in241[5:0] };

   // m241_89 = W*in
   wire signed [9:0] m241_89;
   assign m241_89 =10'b0;

   // m241_90 = W*in
   wire signed [9:0] m241_90;
   assign m241_90 =10'b0;

   // m241_91 = W*in
   wire signed [9:0] m241_91;
   assign m241_91 =10'b0;

   // m241_92 = W*in
   wire signed [9:0] m241_92;
   assign m241_92 =10'b0;

   // m241_93 = W*in
   wire signed [9:0] m241_93;
   assign m241_93 =10'b0;

   // m241_94 = W*in
   wire signed [9:0] m241_94;
   assign m241_94 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_95 = W*in
   wire signed [9:0] m241_95;
   assign m241_95 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_96 = W*in
   wire signed [9:0] m241_96;
   assign m241_96 =10'b0;

   // m241_97 = W*in
   wire signed [9:0] m241_97;
   assign m241_97 =10'b0;

   // m241_98 = W*in
   wire signed [9:0] m241_98;
   assign m241_98 =10'b0;

   // m241_99 = W*in
   wire signed [9:0] m241_99;
   assign m241_99 =10'b0;

   // m241_100 = W*in
   wire signed [9:0] m241_100;
   assign m241_100 =10'b0;

   // m241_101 = W*in
   wire signed [9:0] m241_101;
   assign m241_101 =10'b0;

   // m241_102 = W*in
   wire signed [9:0] m241_102;
   assign m241_102 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_103 = W*in
   wire signed [9:0] m241_103;
   assign m241_103 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_104 = W*in
   wire signed [9:0] m241_104;
   assign m241_104 =10'b0;

   // m241_105 = W*in
   wire signed [9:0] m241_105;
   assign m241_105 ={ {4{in241[5]}} , in241[5:0] };

   // m241_106 = W*in
   wire signed [9:0] m241_106;
   assign m241_106 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_107 = W*in
   wire signed [9:0] m241_107;
   assign m241_107 =10'b0;

   // m241_108 = W*in
   wire signed [9:0] m241_108;
   assign m241_108 ={ {5{neg241[5]}} , neg241[5:1] };

   // m241_109 = W*in
   wire signed [9:0] m241_109;
   assign m241_109 =10'b0;

   // m241_110 = W*in
   wire signed [9:0] m241_110;
   assign m241_110 =10'b0;

   // m241_111 = W*in
   wire signed [9:0] m241_111;
   assign m241_111 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_112 = W*in
   wire signed [9:0] m241_112;
   assign m241_112 =10'b0;

   // m241_113 = W*in
   wire signed [9:0] m241_113;
   assign m241_113 =10'b0;

   // m241_114 = W*in
   wire signed [9:0] m241_114;
   assign m241_114 =10'b0;

   // m241_115 = W*in
   wire signed [9:0] m241_115;
   assign m241_115 ={ {5{neg241[5]}} , neg241[5:1] };

   // m241_116 = W*in
   wire signed [9:0] m241_116;
   assign m241_116 ={ {4{neg241[5]}} , neg241[5:0] };

   // m241_117 = W*in
   wire signed [9:0] m241_117;
   assign m241_117 =10'b0;

   // m242_1 = W*in
   wire signed [9:0] m242_1;
   assign m242_1 =10'b0;

   // m242_2 = W*in
   wire signed [9:0] m242_2;
   assign m242_2 =10'b0;

   // m242_3 = W*in
   wire signed [9:0] m242_3;
   assign m242_3 ={ {4{in242[5]}} , in242[5:0] };

   // m242_4 = W*in
   wire signed [9:0] m242_4;
   assign m242_4 =10'b0;

   // m242_5 = W*in
   wire signed [9:0] m242_5;
   assign m242_5 =10'b0;

   // m242_6 = W*in
   wire signed [9:0] m242_6;
   assign m242_6 =10'b0;

   // m242_7 = W*in
   wire signed [9:0] m242_7;
   assign m242_7 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_8 = W*in
   wire signed [9:0] m242_8;
   assign m242_8 ={ {4{in242[5]}} , in242[5:0] };

   // m242_9 = W*in
   wire signed [9:0] m242_9;
   assign m242_9 =10'b0;

   // m242_10 = W*in
   wire signed [9:0] m242_10;
   assign m242_10 =10'b0;

   // m242_11 = W*in
   wire signed [9:0] m242_11;
   assign m242_11 =10'b0;

   // m242_12 = W*in
   wire signed [9:0] m242_12;
   assign m242_12 ={ {4{in242[5]}} , in242[5:0] };

   // m242_13 = W*in
   wire signed [9:0] m242_13;
   assign m242_13 =10'b0;

   // m242_14 = W*in
   wire signed [9:0] m242_14;
   assign m242_14 ={ {4{in242[5]}} , in242[5:0] };

   // m242_15 = W*in
   wire signed [9:0] m242_15;
   assign m242_15 =10'b0;

   // m242_16 = W*in
   wire signed [9:0] m242_16;
   assign m242_16 =10'b0;

   // m242_17 = W*in
   wire signed [9:0] m242_17;
   assign m242_17 ={ {5{in242[5]}} , in242[5:1] };

   // m242_18 = W*in
   wire signed [9:0] m242_18;
   assign m242_18 =10'b0;

   // m242_19 = W*in
   wire signed [9:0] m242_19;
   assign m242_19 ={ {4{in242[5]}} , in242[5:0] };

   // m242_20 = W*in
   wire signed [9:0] m242_20;
   assign m242_20 =10'b0;

   // m242_21 = W*in
   wire signed [9:0] m242_21;
   assign m242_21 =10'b0;

   // m242_22 = W*in
   wire signed [9:0] m242_22;
   assign m242_22 =10'b0;

   // m242_23 = W*in
   wire signed [9:0] m242_23;
   assign m242_23 ={ {4{in242[5]}} , in242[5:0] };

   // m242_24 = W*in
   wire signed [9:0] m242_24;
   assign m242_24 =10'b0;

   // m242_25 = W*in
   wire signed [9:0] m242_25;
   assign m242_25 ={ {5{neg242[5]}} , neg242[5:1] };

   // m242_26 = W*in
   wire signed [9:0] m242_26;
   assign m242_26 =10'b0;

   // m242_27 = W*in
   wire signed [9:0] m242_27;
   assign m242_27 ={ {4{in242[5]}} , in242[5:0] };

   // m242_28 = W*in
   wire signed [9:0] m242_28;
   assign m242_28 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_29 = W*in
   wire signed [9:0] m242_29;
   assign m242_29 =10'b0;

   // m242_30 = W*in
   wire signed [9:0] m242_30;
   assign m242_30 =10'b0;

   // m242_31 = W*in
   wire signed [9:0] m242_31;
   assign m242_31 ={ {4{in242[5]}} , in242[5:0] };

   // m242_32 = W*in
   wire signed [9:0] m242_32;
   assign m242_32 =10'b0;

   // m242_33 = W*in
   wire signed [9:0] m242_33;
   assign m242_33 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_34 = W*in
   wire signed [9:0] m242_34;
   assign m242_34 =10'b0;

   // m242_35 = W*in
   wire signed [9:0] m242_35;
   assign m242_35 =10'b0;

   // m242_36 = W*in
   wire signed [9:0] m242_36;
   assign m242_36 =10'b0;

   // m242_37 = W*in
   wire signed [9:0] m242_37;
   assign m242_37 =10'b0;

   // m242_38 = W*in
   wire signed [9:0] m242_38;
   assign m242_38 =10'b0;

   // m242_39 = W*in
   wire signed [9:0] m242_39;
   assign m242_39 =10'b0;

   // m242_40 = W*in
   wire signed [9:0] m242_40;
   assign m242_40 =10'b0;

   // m242_41 = W*in
   wire signed [9:0] m242_41;
   assign m242_41 =10'b0;

   // m242_42 = W*in
   wire signed [9:0] m242_42;
   assign m242_42 =10'b0;

   // m242_43 = W*in
   wire signed [9:0] m242_43;
   assign m242_43 =10'b0;

   // m242_44 = W*in
   wire signed [9:0] m242_44;
   assign m242_44 =10'b0;

   // m242_45 = W*in
   wire signed [9:0] m242_45;
   assign m242_45 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_46 = W*in
   wire signed [9:0] m242_46;
   assign m242_46 =10'b0;

   // m242_47 = W*in
   wire signed [9:0] m242_47;
   assign m242_47 =10'b0;

   // m242_48 = W*in
   wire signed [9:0] m242_48;
   assign m242_48 =10'b0;

   // m242_49 = W*in
   wire signed [9:0] m242_49;
   assign m242_49 =10'b0;

   // m242_50 = W*in
   wire signed [9:0] m242_50;
   assign m242_50 =10'b0;

   // m242_51 = W*in
   wire signed [9:0] m242_51;
   assign m242_51 =10'b0;

   // m242_52 = W*in
   wire signed [9:0] m242_52;
   assign m242_52 ={ {4{in242[5]}} , in242[5:0] };

   // m242_53 = W*in
   wire signed [9:0] m242_53;
   assign m242_53 =10'b0;

   // m242_54 = W*in
   wire signed [9:0] m242_54;
   assign m242_54 =10'b0;

   // m242_55 = W*in
   wire signed [9:0] m242_55;
   assign m242_55 =10'b0;

   // m242_56 = W*in
   wire signed [9:0] m242_56;
   assign m242_56 =10'b0;

   // m242_57 = W*in
   wire signed [9:0] m242_57;
   assign m242_57 =10'b0;

   // m242_58 = W*in
   wire signed [9:0] m242_58;
   assign m242_58 =10'b0;

   // m242_59 = W*in
   wire signed [9:0] m242_59;
   assign m242_59 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_60 = W*in
   wire signed [9:0] m242_60;
   assign m242_60 =10'b0;

   // m242_61 = W*in
   wire signed [9:0] m242_61;
   assign m242_61 =10'b0;

   // m242_62 = W*in
   wire signed [9:0] m242_62;
   assign m242_62 =10'b0;

   // m242_63 = W*in
   wire signed [9:0] m242_63;
   assign m242_63 =10'b0;

   // m242_64 = W*in
   wire signed [9:0] m242_64;
   assign m242_64 =10'b0;

   // m242_65 = W*in
   wire signed [9:0] m242_65;
   assign m242_65 ={ {5{in242[5]}} , in242[5:1] };

   // m242_66 = W*in
   wire signed [9:0] m242_66;
   assign m242_66 =10'b0;

   // m242_67 = W*in
   wire signed [9:0] m242_67;
   assign m242_67 =10'b0;

   // m242_68 = W*in
   wire signed [9:0] m242_68;
   assign m242_68 =10'b0;

   // m242_69 = W*in
   wire signed [9:0] m242_69;
   assign m242_69 =10'b0;

   // m242_70 = W*in
   wire signed [9:0] m242_70;
   assign m242_70 ={ {4{in242[5]}} , in242[5:0] };

   // m242_71 = W*in
   wire signed [9:0] m242_71;
   assign m242_71 =10'b0;

   // m242_72 = W*in
   wire signed [9:0] m242_72;
   assign m242_72 =10'b0;

   // m242_73 = W*in
   wire signed [9:0] m242_73;
   assign m242_73 =10'b0;

   // m242_74 = W*in
   wire signed [9:0] m242_74;
   assign m242_74 =10'b0;

   // m242_75 = W*in
   wire signed [9:0] m242_75;
   assign m242_75 =10'b0;

   // m242_76 = W*in
   wire signed [9:0] m242_76;
   assign m242_76 ={ {4{in242[5]}} , in242[5:0] };

   // m242_77 = W*in
   wire signed [9:0] m242_77;
   assign m242_77 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_78 = W*in
   wire signed [9:0] m242_78;
   assign m242_78 =10'b0;

   // m242_79 = W*in
   wire signed [9:0] m242_79;
   assign m242_79 =10'b0;

   // m242_80 = W*in
   wire signed [9:0] m242_80;
   assign m242_80 =10'b0;

   // m242_81 = W*in
   wire signed [9:0] m242_81;
   assign m242_81 ={ {5{in242[5]}} , in242[5:1] };

   // m242_82 = W*in
   wire signed [9:0] m242_82;
   assign m242_82 =10'b0;

   // m242_83 = W*in
   wire signed [9:0] m242_83;
   assign m242_83 ={ {5{neg242[5]}} , neg242[5:1] };

   // m242_84 = W*in
   wire signed [9:0] m242_84;
   assign m242_84 =10'b0;

   // m242_85 = W*in
   wire signed [9:0] m242_85;
   assign m242_85 =10'b0;

   // m242_86 = W*in
   wire signed [9:0] m242_86;
   assign m242_86 =10'b0;

   // m242_87 = W*in
   wire signed [9:0] m242_87;
   assign m242_87 =10'b0;

   // m242_88 = W*in
   wire signed [9:0] m242_88;
   assign m242_88 =10'b0;

   // m242_89 = W*in
   wire signed [9:0] m242_89;
   assign m242_89 =10'b0;

   // m242_90 = W*in
   wire signed [9:0] m242_90;
   assign m242_90 =10'b0;

   // m242_91 = W*in
   wire signed [9:0] m242_91;
   assign m242_91 =10'b0;

   // m242_92 = W*in
   wire signed [9:0] m242_92;
   assign m242_92 =10'b0;

   // m242_93 = W*in
   wire signed [9:0] m242_93;
   assign m242_93 =10'b0;

   // m242_94 = W*in
   wire signed [9:0] m242_94;
   assign m242_94 =10'b0;

   // m242_95 = W*in
   wire signed [9:0] m242_95;
   assign m242_95 =10'b0;

   // m242_96 = W*in
   wire signed [9:0] m242_96;
   assign m242_96 =10'b0;

   // m242_97 = W*in
   wire signed [9:0] m242_97;
   assign m242_97 =10'b0;

   // m242_98 = W*in
   wire signed [9:0] m242_98;
   assign m242_98 ={ {4{in242[5]}} , in242[5:0] };

   // m242_99 = W*in
   wire signed [9:0] m242_99;
   assign m242_99 =10'b0;

   // m242_100 = W*in
   wire signed [9:0] m242_100;
   assign m242_100 =10'b0;

   // m242_101 = W*in
   wire signed [9:0] m242_101;
   assign m242_101 =10'b0;

   // m242_102 = W*in
   wire signed [9:0] m242_102;
   assign m242_102 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_103 = W*in
   wire signed [9:0] m242_103;
   assign m242_103 =10'b0;

   // m242_104 = W*in
   wire signed [9:0] m242_104;
   assign m242_104 =10'b0;

   // m242_105 = W*in
   wire signed [9:0] m242_105;
   assign m242_105 ={ {4{in242[5]}} , in242[5:0] };

   // m242_106 = W*in
   wire signed [9:0] m242_106;
   assign m242_106 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_107 = W*in
   wire signed [9:0] m242_107;
   assign m242_107 =10'b0;

   // m242_108 = W*in
   wire signed [9:0] m242_108;
   assign m242_108 =10'b0;

   // m242_109 = W*in
   wire signed [9:0] m242_109;
   assign m242_109 =10'b0;

   // m242_110 = W*in
   wire signed [9:0] m242_110;
   assign m242_110 =10'b0;

   // m242_111 = W*in
   wire signed [9:0] m242_111;
   assign m242_111 ={ {4{neg242[5]}} , neg242[5:0] };

   // m242_112 = W*in
   wire signed [9:0] m242_112;
   assign m242_112 =10'b0;

   // m242_113 = W*in
   wire signed [9:0] m242_113;
   assign m242_113 =10'b0;

   // m242_114 = W*in
   wire signed [9:0] m242_114;
   assign m242_114 =10'b0;

   // m242_115 = W*in
   wire signed [9:0] m242_115;
   assign m242_115 ={ {5{neg242[5]}} , neg242[5:1] };

   // m242_116 = W*in
   wire signed [9:0] m242_116;
   assign m242_116 =10'b0;

   // m242_117 = W*in
   wire signed [9:0] m242_117;
   assign m242_117 =10'b0;

   // m243_1 = W*in
   wire signed [9:0] m243_1;
   assign m243_1 =10'b0;

   // m243_2 = W*in
   wire signed [9:0] m243_2;
   assign m243_2 =10'b0;

   // m243_3 = W*in
   wire signed [9:0] m243_3;
   assign m243_3 =10'b0;

   // m243_4 = W*in
   wire signed [9:0] m243_4;
   assign m243_4 =10'b0;

   // m243_5 = W*in
   wire signed [9:0] m243_5;
   assign m243_5 =10'b0;

   // m243_6 = W*in
   wire signed [9:0] m243_6;
   assign m243_6 =10'b0;

   // m243_7 = W*in
   wire signed [9:0] m243_7;
   assign m243_7 =10'b0;

   // m243_8 = W*in
   wire signed [9:0] m243_8;
   assign m243_8 =10'b0;

   // m243_9 = W*in
   wire signed [9:0] m243_9;
   assign m243_9 =10'b0;

   // m243_10 = W*in
   wire signed [9:0] m243_10;
   assign m243_10 =10'b0;

   // m243_11 = W*in
   wire signed [9:0] m243_11;
   assign m243_11 =10'b0;

   // m243_12 = W*in
   wire signed [9:0] m243_12;
   assign m243_12 =10'b0;

   // m243_13 = W*in
   wire signed [9:0] m243_13;
   assign m243_13 ={ {4{in243[5]}} , in243[5:0] };

   // m243_14 = W*in
   wire signed [9:0] m243_14;
   assign m243_14 =10'b0;

   // m243_15 = W*in
   wire signed [9:0] m243_15;
   assign m243_15 =10'b0;

   // m243_16 = W*in
   wire signed [9:0] m243_16;
   assign m243_16 ={ {5{neg243[5]}} , neg243[5:1] };

   // m243_17 = W*in
   wire signed [9:0] m243_17;
   assign m243_17 =10'b0;

   // m243_18 = W*in
   wire signed [9:0] m243_18;
   assign m243_18 =10'b0;

   // m243_19 = W*in
   wire signed [9:0] m243_19;
   assign m243_19 ={ {4{neg243[5]}} , neg243[5:0] };

   // m243_20 = W*in
   wire signed [9:0] m243_20;
   assign m243_20 =10'b0;

   // m243_21 = W*in
   wire signed [9:0] m243_21;
   assign m243_21 =10'b0;

   // m243_22 = W*in
   wire signed [9:0] m243_22;
   assign m243_22 =10'b0;

   // m243_23 = W*in
   wire signed [9:0] m243_23;
   assign m243_23 ={ {4{in243[5]}} , in243[5:0] };

   // m243_24 = W*in
   wire signed [9:0] m243_24;
   assign m243_24 =10'b0;

   // m243_25 = W*in
   wire signed [9:0] m243_25;
   assign m243_25 ={ {5{neg243[5]}} , neg243[5:1] };

   // m243_26 = W*in
   wire signed [9:0] m243_26;
   assign m243_26 =10'b0;

   // m243_27 = W*in
   wire signed [9:0] m243_27;
   assign m243_27 ={ {5{in243[5]}} , in243[5:1] };

   // m243_28 = W*in
   wire signed [9:0] m243_28;
   assign m243_28 ={ {5{neg243[5]}} , neg243[5:1] };

   // m243_29 = W*in
   wire signed [9:0] m243_29;
   assign m243_29 =10'b0;

   // m243_30 = W*in
   wire signed [9:0] m243_30;
   assign m243_30 =10'b0;

   // m243_31 = W*in
   wire signed [9:0] m243_31;
   assign m243_31 =10'b0;

   // m243_32 = W*in
   wire signed [9:0] m243_32;
   assign m243_32 =10'b0;

   // m243_33 = W*in
   wire signed [9:0] m243_33;
   assign m243_33 =10'b0;

   // m243_34 = W*in
   wire signed [9:0] m243_34;
   assign m243_34 =10'b0;

   // m243_35 = W*in
   wire signed [9:0] m243_35;
   assign m243_35 =10'b0;

   // m243_36 = W*in
   wire signed [9:0] m243_36;
   assign m243_36 =10'b0;

   // m243_37 = W*in
   wire signed [9:0] m243_37;
   assign m243_37 =10'b0;

   // m243_38 = W*in
   wire signed [9:0] m243_38;
   assign m243_38 =10'b0;

   // m243_39 = W*in
   wire signed [9:0] m243_39;
   assign m243_39 =10'b0;

   // m243_40 = W*in
   wire signed [9:0] m243_40;
   assign m243_40 =10'b0;

   // m243_41 = W*in
   wire signed [9:0] m243_41;
   assign m243_41 ={ {4{in243[5]}} , in243[5:0] };

   // m243_42 = W*in
   wire signed [9:0] m243_42;
   assign m243_42 =10'b0;

   // m243_43 = W*in
   wire signed [9:0] m243_43;
   assign m243_43 =10'b0;

   // m243_44 = W*in
   wire signed [9:0] m243_44;
   assign m243_44 ={ {4{neg243[5]}} , neg243[5:0] };

   // m243_45 = W*in
   wire signed [9:0] m243_45;
   assign m243_45 =10'b0;

   // m243_46 = W*in
   wire signed [9:0] m243_46;
   assign m243_46 =10'b0;

   // m243_47 = W*in
   wire signed [9:0] m243_47;
   assign m243_47 =10'b0;

   // m243_48 = W*in
   wire signed [9:0] m243_48;
   assign m243_48 =10'b0;

   // m243_49 = W*in
   wire signed [9:0] m243_49;
   assign m243_49 =10'b0;

   // m243_50 = W*in
   wire signed [9:0] m243_50;
   assign m243_50 =10'b0;

   // m243_51 = W*in
   wire signed [9:0] m243_51;
   assign m243_51 =10'b0;

   // m243_52 = W*in
   wire signed [9:0] m243_52;
   assign m243_52 =10'b0;

   // m243_53 = W*in
   wire signed [9:0] m243_53;
   assign m243_53 =10'b0;

   // m243_54 = W*in
   wire signed [9:0] m243_54;
   assign m243_54 ={ {4{neg243[5]}} , neg243[5:0] };

   // m243_55 = W*in
   wire signed [9:0] m243_55;
   assign m243_55 =10'b0;

   // m243_56 = W*in
   wire signed [9:0] m243_56;
   assign m243_56 =10'b0;

   // m243_57 = W*in
   wire signed [9:0] m243_57;
   assign m243_57 =10'b0;

   // m243_58 = W*in
   wire signed [9:0] m243_58;
   assign m243_58 =10'b0;

   // m243_59 = W*in
   wire signed [9:0] m243_59;
   assign m243_59 =10'b0;

   // m243_60 = W*in
   wire signed [9:0] m243_60;
   assign m243_60 =10'b0;

   // m243_61 = W*in
   wire signed [9:0] m243_61;
   assign m243_61 =10'b0;

   // m243_62 = W*in
   wire signed [9:0] m243_62;
   assign m243_62 =10'b0;

   // m243_63 = W*in
   wire signed [9:0] m243_63;
   assign m243_63 =10'b0;

   // m243_64 = W*in
   wire signed [9:0] m243_64;
   assign m243_64 ={ {5{in243[5]}} , in243[5:1] };

   // m243_65 = W*in
   wire signed [9:0] m243_65;
   assign m243_65 =10'b0;

   // m243_66 = W*in
   wire signed [9:0] m243_66;
   assign m243_66 =10'b0;

   // m243_67 = W*in
   wire signed [9:0] m243_67;
   assign m243_67 ={ {4{neg243[5]}} , neg243[5:0] };

   // m243_68 = W*in
   wire signed [9:0] m243_68;
   assign m243_68 =10'b0;

   // m243_69 = W*in
   wire signed [9:0] m243_69;
   assign m243_69 ={ {5{in243[5]}} , in243[5:1] };

   // m243_70 = W*in
   wire signed [9:0] m243_70;
   assign m243_70 ={ {5{in243[5]}} , in243[5:1] };

   // m243_71 = W*in
   wire signed [9:0] m243_71;
   assign m243_71 =10'b0;

   // m243_72 = W*in
   wire signed [9:0] m243_72;
   assign m243_72 =10'b0;

   // m243_73 = W*in
   wire signed [9:0] m243_73;
   assign m243_73 =10'b0;

   // m243_74 = W*in
   wire signed [9:0] m243_74;
   assign m243_74 =10'b0;

   // m243_75 = W*in
   wire signed [9:0] m243_75;
   assign m243_75 ={ {5{neg243[5]}} , neg243[5:1] };

   // m243_76 = W*in
   wire signed [9:0] m243_76;
   assign m243_76 =10'b0;

   // m243_77 = W*in
   wire signed [9:0] m243_77;
   assign m243_77 =10'b0;

   // m243_78 = W*in
   wire signed [9:0] m243_78;
   assign m243_78 =10'b0;

   // m243_79 = W*in
   wire signed [9:0] m243_79;
   assign m243_79 =10'b0;

   // m243_80 = W*in
   wire signed [9:0] m243_80;
   assign m243_80 =10'b0;

   // m243_81 = W*in
   wire signed [9:0] m243_81;
   assign m243_81 =10'b0;

   // m243_82 = W*in
   wire signed [9:0] m243_82;
   assign m243_82 =10'b0;

   // m243_83 = W*in
   wire signed [9:0] m243_83;
   assign m243_83 =10'b0;

   // m243_84 = W*in
   wire signed [9:0] m243_84;
   assign m243_84 =10'b0;

   // m243_85 = W*in
   wire signed [9:0] m243_85;
   assign m243_85 =10'b0;

   // m243_86 = W*in
   wire signed [9:0] m243_86;
   assign m243_86 =10'b0;

   // m243_87 = W*in
   wire signed [9:0] m243_87;
   assign m243_87 =10'b0;

   // m243_88 = W*in
   wire signed [9:0] m243_88;
   assign m243_88 =10'b0;

   // m243_89 = W*in
   wire signed [9:0] m243_89;
   assign m243_89 =10'b0;

   // m243_90 = W*in
   wire signed [9:0] m243_90;
   assign m243_90 =10'b0;

   // m243_91 = W*in
   wire signed [9:0] m243_91;
   assign m243_91 ={ {4{neg243[5]}} , neg243[5:0] };

   // m243_92 = W*in
   wire signed [9:0] m243_92;
   assign m243_92 =10'b0;

   // m243_93 = W*in
   wire signed [9:0] m243_93;
   assign m243_93 =10'b0;

   // m243_94 = W*in
   wire signed [9:0] m243_94;
   assign m243_94 =10'b0;

   // m243_95 = W*in
   wire signed [9:0] m243_95;
   assign m243_95 =10'b0;

   // m243_96 = W*in
   wire signed [9:0] m243_96;
   assign m243_96 ={ {4{in243[5]}} , in243[5:0] };

   // m243_97 = W*in
   wire signed [9:0] m243_97;
   assign m243_97 ={ {4{neg243[5]}} , neg243[5:0] };

   // m243_98 = W*in
   wire signed [9:0] m243_98;
   assign m243_98 =10'b0;

   // m243_99 = W*in
   wire signed [9:0] m243_99;
   assign m243_99 =10'b0;

   // m243_100 = W*in
   wire signed [9:0] m243_100;
   assign m243_100 =10'b0;

   // m243_101 = W*in
   wire signed [9:0] m243_101;
   assign m243_101 =10'b0;

   // m243_102 = W*in
   wire signed [9:0] m243_102;
   assign m243_102 =10'b0;

   // m243_103 = W*in
   wire signed [9:0] m243_103;
   assign m243_103 =10'b0;

   // m243_104 = W*in
   wire signed [9:0] m243_104;
   assign m243_104 =10'b0;

   // m243_105 = W*in
   wire signed [9:0] m243_105;
   assign m243_105 =10'b0;

   // m243_106 = W*in
   wire signed [9:0] m243_106;
   assign m243_106 =10'b0;

   // m243_107 = W*in
   wire signed [9:0] m243_107;
   assign m243_107 =10'b0;

   // m243_108 = W*in
   wire signed [9:0] m243_108;
   assign m243_108 ={ {4{in243[5]}} , in243[5:0] };

   // m243_109 = W*in
   wire signed [9:0] m243_109;
   assign m243_109 ={ {4{in243[5]}} , in243[5:0] };

   // m243_110 = W*in
   wire signed [9:0] m243_110;
   assign m243_110 =10'b0;

   // m243_111 = W*in
   wire signed [9:0] m243_111;
   assign m243_111 =10'b0;

   // m243_112 = W*in
   wire signed [9:0] m243_112;
   assign m243_112 =10'b0;

   // m243_113 = W*in
   wire signed [9:0] m243_113;
   assign m243_113 =10'b0;

   // m243_114 = W*in
   wire signed [9:0] m243_114;
   assign m243_114 ={ {5{in243[5]}} , in243[5:1] };

   // m243_115 = W*in
   wire signed [9:0] m243_115;
   assign m243_115 =10'b0;

   // m243_116 = W*in
   wire signed [9:0] m243_116;
   assign m243_116 ={ {4{in243[5]}} , in243[5:0] };

   // m243_117 = W*in
   wire signed [9:0] m243_117;
   assign m243_117 =10'b0;

   // m244_1 = W*in
   wire signed [9:0] m244_1;
   assign m244_1 =10'b0;

   // m244_2 = W*in
   wire signed [9:0] m244_2;
   assign m244_2 =10'b0;

   // m244_3 = W*in
   wire signed [9:0] m244_3;
   assign m244_3 =10'b0;

   // m244_4 = W*in
   wire signed [9:0] m244_4;
   assign m244_4 =10'b0;

   // m244_5 = W*in
   wire signed [9:0] m244_5;
   assign m244_5 =10'b0;

   // m244_6 = W*in
   wire signed [9:0] m244_6;
   assign m244_6 =10'b0;

   // m244_7 = W*in
   wire signed [9:0] m244_7;
   assign m244_7 =10'b0;

   // m244_8 = W*in
   wire signed [9:0] m244_8;
   assign m244_8 =10'b0;

   // m244_9 = W*in
   wire signed [9:0] m244_9;
   assign m244_9 =10'b0;

   // m244_10 = W*in
   wire signed [9:0] m244_10;
   assign m244_10 =10'b0;

   // m244_11 = W*in
   wire signed [9:0] m244_11;
   assign m244_11 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_12 = W*in
   wire signed [9:0] m244_12;
   assign m244_12 =10'b0;

   // m244_13 = W*in
   wire signed [9:0] m244_13;
   assign m244_13 =10'b0;

   // m244_14 = W*in
   wire signed [9:0] m244_14;
   assign m244_14 =10'b0;

   // m244_15 = W*in
   wire signed [9:0] m244_15;
   assign m244_15 =10'b0;

   // m244_16 = W*in
   wire signed [9:0] m244_16;
   assign m244_16 ={ {5{neg244[5]}} , neg244[5:1] };

   // m244_17 = W*in
   wire signed [9:0] m244_17;
   assign m244_17 =10'b0;

   // m244_18 = W*in
   wire signed [9:0] m244_18;
   assign m244_18 ={ {5{in244[5]}} , in244[5:1] };

   // m244_19 = W*in
   wire signed [9:0] m244_19;
   assign m244_19 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_20 = W*in
   wire signed [9:0] m244_20;
   assign m244_20 =10'b0;

   // m244_21 = W*in
   wire signed [9:0] m244_21;
   assign m244_21 =10'b0;

   // m244_22 = W*in
   wire signed [9:0] m244_22;
   assign m244_22 =10'b0;

   // m244_23 = W*in
   wire signed [9:0] m244_23;
   assign m244_23 =10'b0;

   // m244_24 = W*in
   wire signed [9:0] m244_24;
   assign m244_24 =10'b0;

   // m244_25 = W*in
   wire signed [9:0] m244_25;
   assign m244_25 =10'b0;

   // m244_26 = W*in
   wire signed [9:0] m244_26;
   assign m244_26 ={ {4{in244[5]}} , in244[5:0] };

   // m244_27 = W*in
   wire signed [9:0] m244_27;
   assign m244_27 =10'b0;

   // m244_28 = W*in
   wire signed [9:0] m244_28;
   assign m244_28 =10'b0;

   // m244_29 = W*in
   wire signed [9:0] m244_29;
   assign m244_29 =10'b0;

   // m244_30 = W*in
   wire signed [9:0] m244_30;
   assign m244_30 =10'b0;

   // m244_31 = W*in
   wire signed [9:0] m244_31;
   assign m244_31 =10'b0;

   // m244_32 = W*in
   wire signed [9:0] m244_32;
   assign m244_32 =10'b0;

   // m244_33 = W*in
   wire signed [9:0] m244_33;
   assign m244_33 =10'b0;

   // m244_34 = W*in
   wire signed [9:0] m244_34;
   assign m244_34 =10'b0;

   // m244_35 = W*in
   wire signed [9:0] m244_35;
   assign m244_35 =10'b0;

   // m244_36 = W*in
   wire signed [9:0] m244_36;
   assign m244_36 =10'b0;

   // m244_37 = W*in
   wire signed [9:0] m244_37;
   assign m244_37 =10'b0;

   // m244_38 = W*in
   wire signed [9:0] m244_38;
   assign m244_38 =10'b0;

   // m244_39 = W*in
   wire signed [9:0] m244_39;
   assign m244_39 =10'b0;

   // m244_40 = W*in
   wire signed [9:0] m244_40;
   assign m244_40 =10'b0;

   // m244_41 = W*in
   wire signed [9:0] m244_41;
   assign m244_41 =10'b0;

   // m244_42 = W*in
   wire signed [9:0] m244_42;
   assign m244_42 =10'b0;

   // m244_43 = W*in
   wire signed [9:0] m244_43;
   assign m244_43 =10'b0;

   // m244_44 = W*in
   wire signed [9:0] m244_44;
   assign m244_44 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_45 = W*in
   wire signed [9:0] m244_45;
   assign m244_45 =10'b0;

   // m244_46 = W*in
   wire signed [9:0] m244_46;
   assign m244_46 =10'b0;

   // m244_47 = W*in
   wire signed [9:0] m244_47;
   assign m244_47 =10'b0;

   // m244_48 = W*in
   wire signed [9:0] m244_48;
   assign m244_48 =10'b0;

   // m244_49 = W*in
   wire signed [9:0] m244_49;
   assign m244_49 =10'b0;

   // m244_50 = W*in
   wire signed [9:0] m244_50;
   assign m244_50 =10'b0;

   // m244_51 = W*in
   wire signed [9:0] m244_51;
   assign m244_51 =10'b0;

   // m244_52 = W*in
   wire signed [9:0] m244_52;
   assign m244_52 =10'b0;

   // m244_53 = W*in
   wire signed [9:0] m244_53;
   assign m244_53 =10'b0;

   // m244_54 = W*in
   wire signed [9:0] m244_54;
   assign m244_54 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_55 = W*in
   wire signed [9:0] m244_55;
   assign m244_55 =10'b0;

   // m244_56 = W*in
   wire signed [9:0] m244_56;
   assign m244_56 =10'b0;

   // m244_57 = W*in
   wire signed [9:0] m244_57;
   assign m244_57 =10'b0;

   // m244_58 = W*in
   wire signed [9:0] m244_58;
   assign m244_58 =10'b0;

   // m244_59 = W*in
   wire signed [9:0] m244_59;
   assign m244_59 =10'b0;

   // m244_60 = W*in
   wire signed [9:0] m244_60;
   assign m244_60 =10'b0;

   // m244_61 = W*in
   wire signed [9:0] m244_61;
   assign m244_61 =10'b0;

   // m244_62 = W*in
   wire signed [9:0] m244_62;
   assign m244_62 =10'b0;

   // m244_63 = W*in
   wire signed [9:0] m244_63;
   assign m244_63 =10'b0;

   // m244_64 = W*in
   wire signed [9:0] m244_64;
   assign m244_64 =10'b0;

   // m244_65 = W*in
   wire signed [9:0] m244_65;
   assign m244_65 =10'b0;

   // m244_66 = W*in
   wire signed [9:0] m244_66;
   assign m244_66 =10'b0;

   // m244_67 = W*in
   wire signed [9:0] m244_67;
   assign m244_67 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_68 = W*in
   wire signed [9:0] m244_68;
   assign m244_68 =10'b0;

   // m244_69 = W*in
   wire signed [9:0] m244_69;
   assign m244_69 ={ {5{neg244[5]}} , neg244[5:1] };

   // m244_70 = W*in
   wire signed [9:0] m244_70;
   assign m244_70 =10'b0;

   // m244_71 = W*in
   wire signed [9:0] m244_71;
   assign m244_71 =10'b0;

   // m244_72 = W*in
   wire signed [9:0] m244_72;
   assign m244_72 =10'b0;

   // m244_73 = W*in
   wire signed [9:0] m244_73;
   assign m244_73 ={ {5{in244[5]}} , in244[5:1] };

   // m244_74 = W*in
   wire signed [9:0] m244_74;
   assign m244_74 =10'b0;

   // m244_75 = W*in
   wire signed [9:0] m244_75;
   assign m244_75 =10'b0;

   // m244_76 = W*in
   wire signed [9:0] m244_76;
   assign m244_76 =10'b0;

   // m244_77 = W*in
   wire signed [9:0] m244_77;
   assign m244_77 =10'b0;

   // m244_78 = W*in
   wire signed [9:0] m244_78;
   assign m244_78 ={ {4{in244[5]}} , in244[5:0] };

   // m244_79 = W*in
   wire signed [9:0] m244_79;
   assign m244_79 =10'b0;

   // m244_80 = W*in
   wire signed [9:0] m244_80;
   assign m244_80 =10'b0;

   // m244_81 = W*in
   wire signed [9:0] m244_81;
   assign m244_81 =10'b0;

   // m244_82 = W*in
   wire signed [9:0] m244_82;
   assign m244_82 =10'b0;

   // m244_83 = W*in
   wire signed [9:0] m244_83;
   assign m244_83 ={ {5{neg244[5]}} , neg244[5:1] };

   // m244_84 = W*in
   wire signed [9:0] m244_84;
   assign m244_84 =10'b0;

   // m244_85 = W*in
   wire signed [9:0] m244_85;
   assign m244_85 ={ {5{neg244[5]}} , neg244[5:1] };

   // m244_86 = W*in
   wire signed [9:0] m244_86;
   assign m244_86 =10'b0;

   // m244_87 = W*in
   wire signed [9:0] m244_87;
   assign m244_87 =10'b0;

   // m244_88 = W*in
   wire signed [9:0] m244_88;
   assign m244_88 =10'b0;

   // m244_89 = W*in
   wire signed [9:0] m244_89;
   assign m244_89 =10'b0;

   // m244_90 = W*in
   wire signed [9:0] m244_90;
   assign m244_90 =10'b0;

   // m244_91 = W*in
   wire signed [9:0] m244_91;
   assign m244_91 =10'b0;

   // m244_92 = W*in
   wire signed [9:0] m244_92;
   assign m244_92 =10'b0;

   // m244_93 = W*in
   wire signed [9:0] m244_93;
   assign m244_93 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_94 = W*in
   wire signed [9:0] m244_94;
   assign m244_94 =10'b0;

   // m244_95 = W*in
   wire signed [9:0] m244_95;
   assign m244_95 ={ {4{neg244[5]}} , neg244[5:0] };

   // m244_96 = W*in
   wire signed [9:0] m244_96;
   assign m244_96 =10'b0;

   // m244_97 = W*in
   wire signed [9:0] m244_97;
   assign m244_97 =10'b0;

   // m244_98 = W*in
   wire signed [9:0] m244_98;
   assign m244_98 =10'b0;

   // m244_99 = W*in
   wire signed [9:0] m244_99;
   assign m244_99 =10'b0;

   // m244_100 = W*in
   wire signed [9:0] m244_100;
   assign m244_100 =10'b0;

   // m244_101 = W*in
   wire signed [9:0] m244_101;
   assign m244_101 =10'b0;

   // m244_102 = W*in
   wire signed [9:0] m244_102;
   assign m244_102 =10'b0;

   // m244_103 = W*in
   wire signed [9:0] m244_103;
   assign m244_103 =10'b0;

   // m244_104 = W*in
   wire signed [9:0] m244_104;
   assign m244_104 =10'b0;

   // m244_105 = W*in
   wire signed [9:0] m244_105;
   assign m244_105 =10'b0;

   // m244_106 = W*in
   wire signed [9:0] m244_106;
   assign m244_106 =10'b0;

   // m244_107 = W*in
   wire signed [9:0] m244_107;
   assign m244_107 =10'b0;

   // m244_108 = W*in
   wire signed [9:0] m244_108;
   assign m244_108 =10'b0;

   // m244_109 = W*in
   wire signed [9:0] m244_109;
   assign m244_109 =10'b0;

   // m244_110 = W*in
   wire signed [9:0] m244_110;
   assign m244_110 =10'b0;

   // m244_111 = W*in
   wire signed [9:0] m244_111;
   assign m244_111 =10'b0;

   // m244_112 = W*in
   wire signed [9:0] m244_112;
   assign m244_112 =10'b0;

   // m244_113 = W*in
   wire signed [9:0] m244_113;
   assign m244_113 =10'b0;

   // m244_114 = W*in
   wire signed [9:0] m244_114;
   assign m244_114 =10'b0;

   // m244_115 = W*in
   wire signed [9:0] m244_115;
   assign m244_115 =10'b0;

   // m244_116 = W*in
   wire signed [9:0] m244_116;
   assign m244_116 =10'b0;

   // m244_117 = W*in
   wire signed [9:0] m244_117;
   assign m244_117 =10'b0;

   // m245_1 = W*in
   wire signed [9:0] m245_1;
   assign m245_1 ={ {4{in245[5]}} , in245[5:0] };

   // m245_2 = W*in
   wire signed [9:0] m245_2;
   assign m245_2 =10'b0;

   // m245_3 = W*in
   wire signed [9:0] m245_3;
   assign m245_3 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_4 = W*in
   wire signed [9:0] m245_4;
   assign m245_4 =10'b0;

   // m245_5 = W*in
   wire signed [9:0] m245_5;
   assign m245_5 =10'b0;

   // m245_6 = W*in
   wire signed [9:0] m245_6;
   assign m245_6 =10'b0;

   // m245_7 = W*in
   wire signed [9:0] m245_7;
   assign m245_7 =10'b0;

   // m245_8 = W*in
   wire signed [9:0] m245_8;
   assign m245_8 =10'b0;

   // m245_9 = W*in
   wire signed [9:0] m245_9;
   assign m245_9 =10'b0;

   // m245_10 = W*in
   wire signed [9:0] m245_10;
   assign m245_10 =10'b0;

   // m245_11 = W*in
   wire signed [9:0] m245_11;
   assign m245_11 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_12 = W*in
   wire signed [9:0] m245_12;
   assign m245_12 =10'b0;

   // m245_13 = W*in
   wire signed [9:0] m245_13;
   assign m245_13 =10'b0;

   // m245_14 = W*in
   wire signed [9:0] m245_14;
   assign m245_14 ={ {4{in245[5]}} , in245[5:0] };

   // m245_15 = W*in
   wire signed [9:0] m245_15;
   assign m245_15 =10'b0;

   // m245_16 = W*in
   wire signed [9:0] m245_16;
   assign m245_16 ={ {5{neg245[5]}} , neg245[5:1] };

   // m245_17 = W*in
   wire signed [9:0] m245_17;
   assign m245_17 ={ {5{in245[5]}} , in245[5:1] };

   // m245_18 = W*in
   wire signed [9:0] m245_18;
   assign m245_18 ={ {3{in245[5]}} , in245 , {1{1'b0}} };

   // m245_19 = W*in
   wire signed [9:0] m245_19;
   assign m245_19 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_20 = W*in
   wire signed [9:0] m245_20;
   assign m245_20 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_21 = W*in
   wire signed [9:0] m245_21;
   assign m245_21 ={ {4{in245[5]}} , in245[5:0] };

   // m245_22 = W*in
   wire signed [9:0] m245_22;
   assign m245_22 =10'b0;

   // m245_23 = W*in
   wire signed [9:0] m245_23;
   assign m245_23 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_24 = W*in
   wire signed [9:0] m245_24;
   assign m245_24 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_25 = W*in
   wire signed [9:0] m245_25;
   assign m245_25 =10'b0;

   // m245_26 = W*in
   wire signed [9:0] m245_26;
   assign m245_26 ={ {3{in245[5]}} , in245 , {1{1'b0}} };

   // m245_27 = W*in
   wire signed [9:0] m245_27;
   assign m245_27 ={ {5{neg245[5]}} , neg245[5:1] };

   // m245_28 = W*in
   wire signed [9:0] m245_28;
   assign m245_28 =10'b0;

   // m245_29 = W*in
   wire signed [9:0] m245_29;
   assign m245_29 =10'b0;

   // m245_30 = W*in
   wire signed [9:0] m245_30;
   assign m245_30 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_31 = W*in
   wire signed [9:0] m245_31;
   assign m245_31 =10'b0;

   // m245_32 = W*in
   wire signed [9:0] m245_32;
   assign m245_32 =10'b0;

   // m245_33 = W*in
   wire signed [9:0] m245_33;
   assign m245_33 ={ {4{in245[5]}} , in245[5:0] };

   // m245_34 = W*in
   wire signed [9:0] m245_34;
   assign m245_34 =10'b0;

   // m245_35 = W*in
   wire signed [9:0] m245_35;
   assign m245_35 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_36 = W*in
   wire signed [9:0] m245_36;
   assign m245_36 ={ {4{in245[5]}} , in245[5:0] };

   // m245_37 = W*in
   wire signed [9:0] m245_37;
   assign m245_37 =10'b0;

   // m245_38 = W*in
   wire signed [9:0] m245_38;
   assign m245_38 ={ {4{in245[5]}} , in245[5:0] };

   // m245_39 = W*in
   wire signed [9:0] m245_39;
   assign m245_39 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_40 = W*in
   wire signed [9:0] m245_40;
   assign m245_40 =10'b0;

   // m245_41 = W*in
   wire signed [9:0] m245_41;
   assign m245_41 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_42 = W*in
   wire signed [9:0] m245_42;
   assign m245_42 =10'b0;

   // m245_43 = W*in
   wire signed [9:0] m245_43;
   assign m245_43 ={ {4{in245[5]}} , in245[5:0] };

   // m245_44 = W*in
   wire signed [9:0] m245_44;
   assign m245_44 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_45 = W*in
   wire signed [9:0] m245_45;
   assign m245_45 =10'b0;

   // m245_46 = W*in
   wire signed [9:0] m245_46;
   assign m245_46 =10'b0;

   // m245_47 = W*in
   wire signed [9:0] m245_47;
   assign m245_47 =10'b0;

   // m245_48 = W*in
   wire signed [9:0] m245_48;
   assign m245_48 ={ {4{in245[5]}} , in245[5:0] };

   // m245_49 = W*in
   wire signed [9:0] m245_49;
   assign m245_49 =10'b0;

   // m245_50 = W*in
   wire signed [9:0] m245_50;
   assign m245_50 =10'b0;

   // m245_51 = W*in
   wire signed [9:0] m245_51;
   assign m245_51 =10'b0;

   // m245_52 = W*in
   wire signed [9:0] m245_52;
   assign m245_52 =10'b0;

   // m245_53 = W*in
   wire signed [9:0] m245_53;
   assign m245_53 =10'b0;

   // m245_54 = W*in
   wire signed [9:0] m245_54;
   assign m245_54 =10'b0;

   // m245_55 = W*in
   wire signed [9:0] m245_55;
   assign m245_55 =10'b0;

   // m245_56 = W*in
   wire signed [9:0] m245_56;
   assign m245_56 =10'b0;

   // m245_57 = W*in
   wire signed [9:0] m245_57;
   assign m245_57 =10'b0;

   // m245_58 = W*in
   wire signed [9:0] m245_58;
   assign m245_58 ={ {5{neg245[5]}} , neg245[5:1] };

   // m245_59 = W*in
   wire signed [9:0] m245_59;
   assign m245_59 =10'b0;

   // m245_60 = W*in
   wire signed [9:0] m245_60;
   assign m245_60 =10'b0;

   // m245_61 = W*in
   wire signed [9:0] m245_61;
   assign m245_61 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_62 = W*in
   wire signed [9:0] m245_62;
   assign m245_62 =10'b0;

   // m245_63 = W*in
   wire signed [9:0] m245_63;
   assign m245_63 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_64 = W*in
   wire signed [9:0] m245_64;
   assign m245_64 ={ {4{in245[5]}} , in245[5:0] };

   // m245_65 = W*in
   wire signed [9:0] m245_65;
   assign m245_65 =10'b0;

   // m245_66 = W*in
   wire signed [9:0] m245_66;
   assign m245_66 =10'b0;

   // m245_67 = W*in
   wire signed [9:0] m245_67;
   assign m245_67 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_68 = W*in
   wire signed [9:0] m245_68;
   assign m245_68 ={ {4{in245[5]}} , in245[5:0] };

   // m245_69 = W*in
   wire signed [9:0] m245_69;
   assign m245_69 =10'b0;

   // m245_70 = W*in
   wire signed [9:0] m245_70;
   assign m245_70 =10'b0;

   // m245_71 = W*in
   wire signed [9:0] m245_71;
   assign m245_71 ={ {4{in245[5]}} , in245[5:0] };

   // m245_72 = W*in
   wire signed [9:0] m245_72;
   assign m245_72 ={ {4{in245[5]}} , in245[5:0] };

   // m245_73 = W*in
   wire signed [9:0] m245_73;
   assign m245_73 ={ {4{in245[5]}} , in245[5:0] };

   // m245_74 = W*in
   wire signed [9:0] m245_74;
   assign m245_74 =10'b0;

   // m245_75 = W*in
   wire signed [9:0] m245_75;
   assign m245_75 =10'b0;

   // m245_76 = W*in
   wire signed [9:0] m245_76;
   assign m245_76 =10'b0;

   // m245_77 = W*in
   wire signed [9:0] m245_77;
   assign m245_77 =10'b0;

   // m245_78 = W*in
   wire signed [9:0] m245_78;
   assign m245_78 ={ {4{in245[5]}} , in245[5:0] };

   // m245_79 = W*in
   wire signed [9:0] m245_79;
   assign m245_79 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_80 = W*in
   wire signed [9:0] m245_80;
   assign m245_80 =10'b0;

   // m245_81 = W*in
   wire signed [9:0] m245_81;
   assign m245_81 =10'b0;

   // m245_82 = W*in
   wire signed [9:0] m245_82;
   assign m245_82 =10'b0;

   // m245_83 = W*in
   wire signed [9:0] m245_83;
   assign m245_83 =10'b0;

   // m245_84 = W*in
   wire signed [9:0] m245_84;
   assign m245_84 ={ {4{in245[5]}} , in245[5:0] };

   // m245_85 = W*in
   wire signed [9:0] m245_85;
   assign m245_85 =10'b0;

   // m245_86 = W*in
   wire signed [9:0] m245_86;
   assign m245_86 ={ {4{in245[5]}} , in245[5:0] };

   // m245_87 = W*in
   wire signed [9:0] m245_87;
   assign m245_87 ={ {4{in245[5]}} , in245[5:0] };

   // m245_88 = W*in
   wire signed [9:0] m245_88;
   assign m245_88 =10'b0;

   // m245_89 = W*in
   wire signed [9:0] m245_89;
   assign m245_89 =10'b0;

   // m245_90 = W*in
   wire signed [9:0] m245_90;
   assign m245_90 ={ {4{in245[5]}} , in245[5:0] };

   // m245_91 = W*in
   wire signed [9:0] m245_91;
   assign m245_91 =10'b0;

   // m245_92 = W*in
   wire signed [9:0] m245_92;
   assign m245_92 =10'b0;

   // m245_93 = W*in
   wire signed [9:0] m245_93;
   assign m245_93 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_94 = W*in
   wire signed [9:0] m245_94;
   assign m245_94 =10'b0;

   // m245_95 = W*in
   wire signed [9:0] m245_95;
   assign m245_95 =10'b0;

   // m245_96 = W*in
   wire signed [9:0] m245_96;
   assign m245_96 =10'b0;

   // m245_97 = W*in
   wire signed [9:0] m245_97;
   assign m245_97 =10'b0;

   // m245_98 = W*in
   wire signed [9:0] m245_98;
   assign m245_98 =10'b0;

   // m245_99 = W*in
   wire signed [9:0] m245_99;
   assign m245_99 =10'b0;

   // m245_100 = W*in
   wire signed [9:0] m245_100;
   assign m245_100 =10'b0;

   // m245_101 = W*in
   wire signed [9:0] m245_101;
   assign m245_101 =10'b0;

   // m245_102 = W*in
   wire signed [9:0] m245_102;
   assign m245_102 =10'b0;

   // m245_103 = W*in
   wire signed [9:0] m245_103;
   assign m245_103 =10'b0;

   // m245_104 = W*in
   wire signed [9:0] m245_104;
   assign m245_104 =10'b0;

   // m245_105 = W*in
   wire signed [9:0] m245_105;
   assign m245_105 =10'b0;

   // m245_106 = W*in
   wire signed [9:0] m245_106;
   assign m245_106 ={ {5{neg245[5]}} , neg245[5:1] };

   // m245_107 = W*in
   wire signed [9:0] m245_107;
   assign m245_107 =10'b0;

   // m245_108 = W*in
   wire signed [9:0] m245_108;
   assign m245_108 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_109 = W*in
   wire signed [9:0] m245_109;
   assign m245_109 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_110 = W*in
   wire signed [9:0] m245_110;
   assign m245_110 =10'b0;

   // m245_111 = W*in
   wire signed [9:0] m245_111;
   assign m245_111 ={ {4{in245[5]}} , in245[5:0] };

   // m245_112 = W*in
   wire signed [9:0] m245_112;
   assign m245_112 =10'b0;

   // m245_113 = W*in
   wire signed [9:0] m245_113;
   assign m245_113 =10'b0;

   // m245_114 = W*in
   wire signed [9:0] m245_114;
   assign m245_114 ={ {5{neg245[5]}} , neg245[5:1] };

   // m245_115 = W*in
   wire signed [9:0] m245_115;
   assign m245_115 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_116 = W*in
   wire signed [9:0] m245_116;
   assign m245_116 ={ {4{neg245[5]}} , neg245[5:0] };

   // m245_117 = W*in
   wire signed [9:0] m245_117;
   assign m245_117 ={ {4{neg245[5]}} , neg245[5:0] };

   // m246_1 = W*in
   wire signed [9:0] m246_1;
   assign m246_1 =10'b0;

   // m246_2 = W*in
   wire signed [9:0] m246_2;
   assign m246_2 =10'b0;

   // m246_3 = W*in
   wire signed [9:0] m246_3;
   assign m246_3 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_4 = W*in
   wire signed [9:0] m246_4;
   assign m246_4 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_5 = W*in
   wire signed [9:0] m246_5;
   assign m246_5 =10'b0;

   // m246_6 = W*in
   wire signed [9:0] m246_6;
   assign m246_6 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_7 = W*in
   wire signed [9:0] m246_7;
   assign m246_7 ={ {4{in246[5]}} , in246[5:0] };

   // m246_8 = W*in
   wire signed [9:0] m246_8;
   assign m246_8 =10'b0;

   // m246_9 = W*in
   wire signed [9:0] m246_9;
   assign m246_9 =10'b0;

   // m246_10 = W*in
   wire signed [9:0] m246_10;
   assign m246_10 =10'b0;

   // m246_11 = W*in
   wire signed [9:0] m246_11;
   assign m246_11 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_12 = W*in
   wire signed [9:0] m246_12;
   assign m246_12 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_13 = W*in
   wire signed [9:0] m246_13;
   assign m246_13 =10'b0;

   // m246_14 = W*in
   wire signed [9:0] m246_14;
   assign m246_14 =10'b0;

   // m246_15 = W*in
   wire signed [9:0] m246_15;
   assign m246_15 =10'b0;

   // m246_16 = W*in
   wire signed [9:0] m246_16;
   assign m246_16 =10'b0;

   // m246_17 = W*in
   wire signed [9:0] m246_17;
   assign m246_17 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_18 = W*in
   wire signed [9:0] m246_18;
   assign m246_18 =10'b0;

   // m246_19 = W*in
   wire signed [9:0] m246_19;
   assign m246_19 =10'b0;

   // m246_20 = W*in
   wire signed [9:0] m246_20;
   assign m246_20 ={ {5{neg246[5]}} , neg246[5:1] };

   // m246_21 = W*in
   wire signed [9:0] m246_21;
   assign m246_21 ={ {5{in246[5]}} , in246[5:1] };

   // m246_22 = W*in
   wire signed [9:0] m246_22;
   assign m246_22 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_23 = W*in
   wire signed [9:0] m246_23;
   assign m246_23 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_24 = W*in
   wire signed [9:0] m246_24;
   assign m246_24 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_25 = W*in
   wire signed [9:0] m246_25;
   assign m246_25 ={ {4{in246[5]}} , in246[5:0] };

   // m246_26 = W*in
   wire signed [9:0] m246_26;
   assign m246_26 ={ {4{in246[5]}} , in246[5:0] };

   // m246_27 = W*in
   wire signed [9:0] m246_27;
   assign m246_27 =10'b0;

   // m246_28 = W*in
   wire signed [9:0] m246_28;
   assign m246_28 ={ {4{in246[5]}} , in246[5:0] };

   // m246_29 = W*in
   wire signed [9:0] m246_29;
   assign m246_29 ={ {4{in246[5]}} , in246[5:0] };

   // m246_30 = W*in
   wire signed [9:0] m246_30;
   assign m246_30 =10'b0;

   // m246_31 = W*in
   wire signed [9:0] m246_31;
   assign m246_31 =10'b0;

   // m246_32 = W*in
   wire signed [9:0] m246_32;
   assign m246_32 =10'b0;

   // m246_33 = W*in
   wire signed [9:0] m246_33;
   assign m246_33 ={ {4{in246[5]}} , in246[5:0] };

   // m246_34 = W*in
   wire signed [9:0] m246_34;
   assign m246_34 =10'b0;

   // m246_35 = W*in
   wire signed [9:0] m246_35;
   assign m246_35 =10'b0;

   // m246_36 = W*in
   wire signed [9:0] m246_36;
   assign m246_36 ={ {4{in246[5]}} , in246[5:0] };

   // m246_37 = W*in
   wire signed [9:0] m246_37;
   assign m246_37 =10'b0;

   // m246_38 = W*in
   wire signed [9:0] m246_38;
   assign m246_38 =10'b0;

   // m246_39 = W*in
   wire signed [9:0] m246_39;
   assign m246_39 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_40 = W*in
   wire signed [9:0] m246_40;
   assign m246_40 =10'b0;

   // m246_41 = W*in
   wire signed [9:0] m246_41;
   assign m246_41 =10'b0;

   // m246_42 = W*in
   wire signed [9:0] m246_42;
   assign m246_42 =10'b0;

   // m246_43 = W*in
   wire signed [9:0] m246_43;
   assign m246_43 ={ {4{in246[5]}} , in246[5:0] };

   // m246_44 = W*in
   wire signed [9:0] m246_44;
   assign m246_44 =10'b0;

   // m246_45 = W*in
   wire signed [9:0] m246_45;
   assign m246_45 =10'b0;

   // m246_46 = W*in
   wire signed [9:0] m246_46;
   assign m246_46 =10'b0;

   // m246_47 = W*in
   wire signed [9:0] m246_47;
   assign m246_47 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_48 = W*in
   wire signed [9:0] m246_48;
   assign m246_48 ={ {4{in246[5]}} , in246[5:0] };

   // m246_49 = W*in
   wire signed [9:0] m246_49;
   assign m246_49 =10'b0;

   // m246_50 = W*in
   wire signed [9:0] m246_50;
   assign m246_50 =10'b0;

   // m246_51 = W*in
   wire signed [9:0] m246_51;
   assign m246_51 ={ {5{neg246[5]}} , neg246[5:1] };

   // m246_52 = W*in
   wire signed [9:0] m246_52;
   assign m246_52 =10'b0;

   // m246_53 = W*in
   wire signed [9:0] m246_53;
   assign m246_53 =10'b0;

   // m246_54 = W*in
   wire signed [9:0] m246_54;
   assign m246_54 =10'b0;

   // m246_55 = W*in
   wire signed [9:0] m246_55;
   assign m246_55 ={ {4{in246[5]}} , in246[5:0] };

   // m246_56 = W*in
   wire signed [9:0] m246_56;
   assign m246_56 =10'b0;

   // m246_57 = W*in
   wire signed [9:0] m246_57;
   assign m246_57 =10'b0;

   // m246_58 = W*in
   wire signed [9:0] m246_58;
   assign m246_58 =10'b0;

   // m246_59 = W*in
   wire signed [9:0] m246_59;
   assign m246_59 ={ {4{in246[5]}} , in246[5:0] };

   // m246_60 = W*in
   wire signed [9:0] m246_60;
   assign m246_60 =10'b0;

   // m246_61 = W*in
   wire signed [9:0] m246_61;
   assign m246_61 =10'b0;

   // m246_62 = W*in
   wire signed [9:0] m246_62;
   assign m246_62 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_63 = W*in
   wire signed [9:0] m246_63;
   assign m246_63 =10'b0;

   // m246_64 = W*in
   wire signed [9:0] m246_64;
   assign m246_64 ={ {5{neg246[5]}} , neg246[5:1] };

   // m246_65 = W*in
   wire signed [9:0] m246_65;
   assign m246_65 =10'b0;

   // m246_66 = W*in
   wire signed [9:0] m246_66;
   assign m246_66 =10'b0;

   // m246_67 = W*in
   wire signed [9:0] m246_67;
   assign m246_67 =10'b0;

   // m246_68 = W*in
   wire signed [9:0] m246_68;
   assign m246_68 ={ {4{in246[5]}} , in246[5:0] };

   // m246_69 = W*in
   wire signed [9:0] m246_69;
   assign m246_69 ={ {4{in246[5]}} , in246[5:0] };

   // m246_70 = W*in
   wire signed [9:0] m246_70;
   assign m246_70 ={ {4{in246[5]}} , in246[5:0] };

   // m246_71 = W*in
   wire signed [9:0] m246_71;
   assign m246_71 =10'b0;

   // m246_72 = W*in
   wire signed [9:0] m246_72;
   assign m246_72 ={ {4{in246[5]}} , in246[5:0] };

   // m246_73 = W*in
   wire signed [9:0] m246_73;
   assign m246_73 =10'b0;

   // m246_74 = W*in
   wire signed [9:0] m246_74;
   assign m246_74 =10'b0;

   // m246_75 = W*in
   wire signed [9:0] m246_75;
   assign m246_75 =10'b0;

   // m246_76 = W*in
   wire signed [9:0] m246_76;
   assign m246_76 =10'b0;

   // m246_77 = W*in
   wire signed [9:0] m246_77;
   assign m246_77 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_78 = W*in
   wire signed [9:0] m246_78;
   assign m246_78 =10'b0;

   // m246_79 = W*in
   wire signed [9:0] m246_79;
   assign m246_79 =10'b0;

   // m246_80 = W*in
   wire signed [9:0] m246_80;
   assign m246_80 =10'b0;

   // m246_81 = W*in
   wire signed [9:0] m246_81;
   assign m246_81 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_82 = W*in
   wire signed [9:0] m246_82;
   assign m246_82 ={ {4{in246[5]}} , in246[5:0] };

   // m246_83 = W*in
   wire signed [9:0] m246_83;
   assign m246_83 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_84 = W*in
   wire signed [9:0] m246_84;
   assign m246_84 ={ {4{in246[5]}} , in246[5:0] };

   // m246_85 = W*in
   wire signed [9:0] m246_85;
   assign m246_85 =10'b0;

   // m246_86 = W*in
   wire signed [9:0] m246_86;
   assign m246_86 =10'b0;

   // m246_87 = W*in
   wire signed [9:0] m246_87;
   assign m246_87 =10'b0;

   // m246_88 = W*in
   wire signed [9:0] m246_88;
   assign m246_88 =10'b0;

   // m246_89 = W*in
   wire signed [9:0] m246_89;
   assign m246_89 ={ {4{in246[5]}} , in246[5:0] };

   // m246_90 = W*in
   wire signed [9:0] m246_90;
   assign m246_90 =10'b0;

   // m246_91 = W*in
   wire signed [9:0] m246_91;
   assign m246_91 =10'b0;

   // m246_92 = W*in
   wire signed [9:0] m246_92;
   assign m246_92 =10'b0;

   // m246_93 = W*in
   wire signed [9:0] m246_93;
   assign m246_93 ={ {4{in246[5]}} , in246[5:0] };

   // m246_94 = W*in
   wire signed [9:0] m246_94;
   assign m246_94 =10'b0;

   // m246_95 = W*in
   wire signed [9:0] m246_95;
   assign m246_95 =10'b0;

   // m246_96 = W*in
   wire signed [9:0] m246_96;
   assign m246_96 =10'b0;

   // m246_97 = W*in
   wire signed [9:0] m246_97;
   assign m246_97 =10'b0;

   // m246_98 = W*in
   wire signed [9:0] m246_98;
   assign m246_98 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_99 = W*in
   wire signed [9:0] m246_99;
   assign m246_99 =10'b0;

   // m246_100 = W*in
   wire signed [9:0] m246_100;
   assign m246_100 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_101 = W*in
   wire signed [9:0] m246_101;
   assign m246_101 =10'b0;

   // m246_102 = W*in
   wire signed [9:0] m246_102;
   assign m246_102 =10'b0;

   // m246_103 = W*in
   wire signed [9:0] m246_103;
   assign m246_103 =10'b0;

   // m246_104 = W*in
   wire signed [9:0] m246_104;
   assign m246_104 =10'b0;

   // m246_105 = W*in
   wire signed [9:0] m246_105;
   assign m246_105 =10'b0;

   // m246_106 = W*in
   wire signed [9:0] m246_106;
   assign m246_106 ={ {4{in246[5]}} , in246[5:0] };

   // m246_107 = W*in
   wire signed [9:0] m246_107;
   assign m246_107 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_108 = W*in
   wire signed [9:0] m246_108;
   assign m246_108 =10'b0;

   // m246_109 = W*in
   wire signed [9:0] m246_109;
   assign m246_109 =10'b0;

   // m246_110 = W*in
   wire signed [9:0] m246_110;
   assign m246_110 =10'b0;

   // m246_111 = W*in
   wire signed [9:0] m246_111;
   assign m246_111 ={ {4{in246[5]}} , in246[5:0] };

   // m246_112 = W*in
   wire signed [9:0] m246_112;
   assign m246_112 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_113 = W*in
   wire signed [9:0] m246_113;
   assign m246_113 =10'b0;

   // m246_114 = W*in
   wire signed [9:0] m246_114;
   assign m246_114 ={ {4{neg246[5]}} , neg246[5:0] };

   // m246_115 = W*in
   wire signed [9:0] m246_115;
   assign m246_115 =10'b0;

   // m246_116 = W*in
   wire signed [9:0] m246_116;
   assign m246_116 =10'b0;

   // m246_117 = W*in
   wire signed [9:0] m246_117;
   assign m246_117 ={ {5{neg246[5]}} , neg246[5:1] };

   // m247_1 = W*in
   wire signed [9:0] m247_1;
   assign m247_1 =10'b0;

   // m247_2 = W*in
   wire signed [9:0] m247_2;
   assign m247_2 =10'b0;

   // m247_3 = W*in
   wire signed [9:0] m247_3;
   assign m247_3 =10'b0;

   // m247_4 = W*in
   wire signed [9:0] m247_4;
   assign m247_4 =10'b0;

   // m247_5 = W*in
   wire signed [9:0] m247_5;
   assign m247_5 =10'b0;

   // m247_6 = W*in
   wire signed [9:0] m247_6;
   assign m247_6 =10'b0;

   // m247_7 = W*in
   wire signed [9:0] m247_7;
   assign m247_7 =10'b0;

   // m247_8 = W*in
   wire signed [9:0] m247_8;
   assign m247_8 ={ {4{in247[5]}} , in247[5:0] };

   // m247_9 = W*in
   wire signed [9:0] m247_9;
   assign m247_9 =10'b0;

   // m247_10 = W*in
   wire signed [9:0] m247_10;
   assign m247_10 =10'b0;

   // m247_11 = W*in
   wire signed [9:0] m247_11;
   assign m247_11 =10'b0;

   // m247_12 = W*in
   wire signed [9:0] m247_12;
   assign m247_12 =10'b0;

   // m247_13 = W*in
   wire signed [9:0] m247_13;
   assign m247_13 =10'b0;

   // m247_14 = W*in
   wire signed [9:0] m247_14;
   assign m247_14 =10'b0;

   // m247_15 = W*in
   wire signed [9:0] m247_15;
   assign m247_15 =10'b0;

   // m247_16 = W*in
   wire signed [9:0] m247_16;
   assign m247_16 =10'b0;

   // m247_17 = W*in
   wire signed [9:0] m247_17;
   assign m247_17 =10'b0;

   // m247_18 = W*in
   wire signed [9:0] m247_18;
   assign m247_18 =10'b0;

   // m247_19 = W*in
   wire signed [9:0] m247_19;
   assign m247_19 =10'b0;

   // m247_20 = W*in
   wire signed [9:0] m247_20;
   assign m247_20 =10'b0;

   // m247_21 = W*in
   wire signed [9:0] m247_21;
   assign m247_21 =10'b0;

   // m247_22 = W*in
   wire signed [9:0] m247_22;
   assign m247_22 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_23 = W*in
   wire signed [9:0] m247_23;
   assign m247_23 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_24 = W*in
   wire signed [9:0] m247_24;
   assign m247_24 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_25 = W*in
   wire signed [9:0] m247_25;
   assign m247_25 =10'b0;

   // m247_26 = W*in
   wire signed [9:0] m247_26;
   assign m247_26 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_27 = W*in
   wire signed [9:0] m247_27;
   assign m247_27 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_28 = W*in
   wire signed [9:0] m247_28;
   assign m247_28 ={ {5{in247[5]}} , in247[5:1] };

   // m247_29 = W*in
   wire signed [9:0] m247_29;
   assign m247_29 =10'b0;

   // m247_30 = W*in
   wire signed [9:0] m247_30;
   assign m247_30 ={ {4{in247[5]}} , in247[5:0] };

   // m247_31 = W*in
   wire signed [9:0] m247_31;
   assign m247_31 ={ {5{in247[5]}} , in247[5:1] };

   // m247_32 = W*in
   wire signed [9:0] m247_32;
   assign m247_32 =10'b0;

   // m247_33 = W*in
   wire signed [9:0] m247_33;
   assign m247_33 =10'b0;

   // m247_34 = W*in
   wire signed [9:0] m247_34;
   assign m247_34 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_35 = W*in
   wire signed [9:0] m247_35;
   assign m247_35 =10'b0;

   // m247_36 = W*in
   wire signed [9:0] m247_36;
   assign m247_36 ={ {5{in247[5]}} , in247[5:1] };

   // m247_37 = W*in
   wire signed [9:0] m247_37;
   assign m247_37 =10'b0;

   // m247_38 = W*in
   wire signed [9:0] m247_38;
   assign m247_38 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_39 = W*in
   wire signed [9:0] m247_39;
   assign m247_39 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_40 = W*in
   wire signed [9:0] m247_40;
   assign m247_40 =10'b0;

   // m247_41 = W*in
   wire signed [9:0] m247_41;
   assign m247_41 =10'b0;

   // m247_42 = W*in
   wire signed [9:0] m247_42;
   assign m247_42 ={ {4{in247[5]}} , in247[5:0] };

   // m247_43 = W*in
   wire signed [9:0] m247_43;
   assign m247_43 =10'b0;

   // m247_44 = W*in
   wire signed [9:0] m247_44;
   assign m247_44 =10'b0;

   // m247_45 = W*in
   wire signed [9:0] m247_45;
   assign m247_45 =10'b0;

   // m247_46 = W*in
   wire signed [9:0] m247_46;
   assign m247_46 =10'b0;

   // m247_47 = W*in
   wire signed [9:0] m247_47;
   assign m247_47 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_48 = W*in
   wire signed [9:0] m247_48;
   assign m247_48 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_49 = W*in
   wire signed [9:0] m247_49;
   assign m247_49 ={ {4{in247[5]}} , in247[5:0] };

   // m247_50 = W*in
   wire signed [9:0] m247_50;
   assign m247_50 =10'b0;

   // m247_51 = W*in
   wire signed [9:0] m247_51;
   assign m247_51 =10'b0;

   // m247_52 = W*in
   wire signed [9:0] m247_52;
   assign m247_52 =10'b0;

   // m247_53 = W*in
   wire signed [9:0] m247_53;
   assign m247_53 ={ {4{in247[5]}} , in247[5:0] };

   // m247_54 = W*in
   wire signed [9:0] m247_54;
   assign m247_54 =10'b0;

   // m247_55 = W*in
   wire signed [9:0] m247_55;
   assign m247_55 =10'b0;

   // m247_56 = W*in
   wire signed [9:0] m247_56;
   assign m247_56 =10'b0;

   // m247_57 = W*in
   wire signed [9:0] m247_57;
   assign m247_57 =10'b0;

   // m247_58 = W*in
   wire signed [9:0] m247_58;
   assign m247_58 =10'b0;

   // m247_59 = W*in
   wire signed [9:0] m247_59;
   assign m247_59 =10'b0;

   // m247_60 = W*in
   wire signed [9:0] m247_60;
   assign m247_60 =10'b0;

   // m247_61 = W*in
   wire signed [9:0] m247_61;
   assign m247_61 =10'b0;

   // m247_62 = W*in
   wire signed [9:0] m247_62;
   assign m247_62 =10'b0;

   // m247_63 = W*in
   wire signed [9:0] m247_63;
   assign m247_63 =10'b0;

   // m247_64 = W*in
   wire signed [9:0] m247_64;
   assign m247_64 =10'b0;

   // m247_65 = W*in
   wire signed [9:0] m247_65;
   assign m247_65 ={ {5{in247[5]}} , in247[5:1] };

   // m247_66 = W*in
   wire signed [9:0] m247_66;
   assign m247_66 ={ {5{in247[5]}} , in247[5:1] };

   // m247_67 = W*in
   wire signed [9:0] m247_67;
   assign m247_67 ={ {4{in247[5]}} , in247[5:0] };

   // m247_68 = W*in
   wire signed [9:0] m247_68;
   assign m247_68 ={ {4{in247[5]}} , in247[5:0] };

   // m247_69 = W*in
   wire signed [9:0] m247_69;
   assign m247_69 =10'b0;

   // m247_70 = W*in
   wire signed [9:0] m247_70;
   assign m247_70 =10'b0;

   // m247_71 = W*in
   wire signed [9:0] m247_71;
   assign m247_71 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_72 = W*in
   wire signed [9:0] m247_72;
   assign m247_72 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_73 = W*in
   wire signed [9:0] m247_73;
   assign m247_73 ={ {4{in247[5]}} , in247[5:0] };

   // m247_74 = W*in
   wire signed [9:0] m247_74;
   assign m247_74 =10'b0;

   // m247_75 = W*in
   wire signed [9:0] m247_75;
   assign m247_75 =10'b0;

   // m247_76 = W*in
   wire signed [9:0] m247_76;
   assign m247_76 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_77 = W*in
   wire signed [9:0] m247_77;
   assign m247_77 =10'b0;

   // m247_78 = W*in
   wire signed [9:0] m247_78;
   assign m247_78 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_79 = W*in
   wire signed [9:0] m247_79;
   assign m247_79 =10'b0;

   // m247_80 = W*in
   wire signed [9:0] m247_80;
   assign m247_80 ={ {4{in247[5]}} , in247[5:0] };

   // m247_81 = W*in
   wire signed [9:0] m247_81;
   assign m247_81 =10'b0;

   // m247_82 = W*in
   wire signed [9:0] m247_82;
   assign m247_82 =10'b0;

   // m247_83 = W*in
   wire signed [9:0] m247_83;
   assign m247_83 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_84 = W*in
   wire signed [9:0] m247_84;
   assign m247_84 =10'b0;

   // m247_85 = W*in
   wire signed [9:0] m247_85;
   assign m247_85 =10'b0;

   // m247_86 = W*in
   wire signed [9:0] m247_86;
   assign m247_86 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_87 = W*in
   wire signed [9:0] m247_87;
   assign m247_87 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_88 = W*in
   wire signed [9:0] m247_88;
   assign m247_88 =10'b0;

   // m247_89 = W*in
   wire signed [9:0] m247_89;
   assign m247_89 =10'b0;

   // m247_90 = W*in
   wire signed [9:0] m247_90;
   assign m247_90 =10'b0;

   // m247_91 = W*in
   wire signed [9:0] m247_91;
   assign m247_91 =10'b0;

   // m247_92 = W*in
   wire signed [9:0] m247_92;
   assign m247_92 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_93 = W*in
   wire signed [9:0] m247_93;
   assign m247_93 =10'b0;

   // m247_94 = W*in
   wire signed [9:0] m247_94;
   assign m247_94 =10'b0;

   // m247_95 = W*in
   wire signed [9:0] m247_95;
   assign m247_95 =10'b0;

   // m247_96 = W*in
   wire signed [9:0] m247_96;
   assign m247_96 =10'b0;

   // m247_97 = W*in
   wire signed [9:0] m247_97;
   assign m247_97 =10'b0;

   // m247_98 = W*in
   wire signed [9:0] m247_98;
   assign m247_98 =10'b0;

   // m247_99 = W*in
   wire signed [9:0] m247_99;
   assign m247_99 =10'b0;

   // m247_100 = W*in
   wire signed [9:0] m247_100;
   assign m247_100 ={ {4{in247[5]}} , in247[5:0] };

   // m247_101 = W*in
   wire signed [9:0] m247_101;
   assign m247_101 =10'b0;

   // m247_102 = W*in
   wire signed [9:0] m247_102;
   assign m247_102 ={ {4{in247[5]}} , in247[5:0] };

   // m247_103 = W*in
   wire signed [9:0] m247_103;
   assign m247_103 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_104 = W*in
   wire signed [9:0] m247_104;
   assign m247_104 =10'b0;

   // m247_105 = W*in
   wire signed [9:0] m247_105;
   assign m247_105 =10'b0;

   // m247_106 = W*in
   wire signed [9:0] m247_106;
   assign m247_106 ={ {4{in247[5]}} , in247[5:0] };

   // m247_107 = W*in
   wire signed [9:0] m247_107;
   assign m247_107 =10'b0;

   // m247_108 = W*in
   wire signed [9:0] m247_108;
   assign m247_108 =10'b0;

   // m247_109 = W*in
   wire signed [9:0] m247_109;
   assign m247_109 ={ {5{neg247[5]}} , neg247[5:1] };

   // m247_110 = W*in
   wire signed [9:0] m247_110;
   assign m247_110 =10'b0;

   // m247_111 = W*in
   wire signed [9:0] m247_111;
   assign m247_111 =10'b0;

   // m247_112 = W*in
   wire signed [9:0] m247_112;
   assign m247_112 =10'b0;

   // m247_113 = W*in
   wire signed [9:0] m247_113;
   assign m247_113 =10'b0;

   // m247_114 = W*in
   wire signed [9:0] m247_114;
   assign m247_114 ={ {4{neg247[5]}} , neg247[5:0] };

   // m247_115 = W*in
   wire signed [9:0] m247_115;
   assign m247_115 =10'b0;

   // m247_116 = W*in
   wire signed [9:0] m247_116;
   assign m247_116 =10'b0;

   // m247_117 = W*in
   wire signed [9:0] m247_117;
   assign m247_117 =10'b0;

   // m248_1 = W*in
   wire signed [9:0] m248_1;
   assign m248_1 =10'b0;

   // m248_2 = W*in
   wire signed [9:0] m248_2;
   assign m248_2 =10'b0;

   // m248_3 = W*in
   wire signed [9:0] m248_3;
   assign m248_3 =10'b0;

   // m248_4 = W*in
   wire signed [9:0] m248_4;
   assign m248_4 =10'b0;

   // m248_5 = W*in
   wire signed [9:0] m248_5;
   assign m248_5 =10'b0;

   // m248_6 = W*in
   wire signed [9:0] m248_6;
   assign m248_6 =10'b0;

   // m248_7 = W*in
   wire signed [9:0] m248_7;
   assign m248_7 =10'b0;

   // m248_8 = W*in
   wire signed [9:0] m248_8;
   assign m248_8 =10'b0;

   // m248_9 = W*in
   wire signed [9:0] m248_9;
   assign m248_9 =10'b0;

   // m248_10 = W*in
   wire signed [9:0] m248_10;
   assign m248_10 =10'b0;

   // m248_11 = W*in
   wire signed [9:0] m248_11;
   assign m248_11 =10'b0;

   // m248_12 = W*in
   wire signed [9:0] m248_12;
   assign m248_12 =10'b0;

   // m248_13 = W*in
   wire signed [9:0] m248_13;
   assign m248_13 =10'b0;

   // m248_14 = W*in
   wire signed [9:0] m248_14;
   assign m248_14 =10'b0;

   // m248_15 = W*in
   wire signed [9:0] m248_15;
   assign m248_15 =10'b0;

   // m248_16 = W*in
   wire signed [9:0] m248_16;
   assign m248_16 =10'b0;

   // m248_17 = W*in
   wire signed [9:0] m248_17;
   assign m248_17 =10'b0;

   // m248_18 = W*in
   wire signed [9:0] m248_18;
   assign m248_18 =10'b0;

   // m248_19 = W*in
   wire signed [9:0] m248_19;
   assign m248_19 =10'b0;

   // m248_20 = W*in
   wire signed [9:0] m248_20;
   assign m248_20 =10'b0;

   // m248_21 = W*in
   wire signed [9:0] m248_21;
   assign m248_21 =10'b0;

   // m248_22 = W*in
   wire signed [9:0] m248_22;
   assign m248_22 =10'b0;

   // m248_23 = W*in
   wire signed [9:0] m248_23;
   assign m248_23 ={ {5{in248[5]}} , in248[5:1] };

   // m248_24 = W*in
   wire signed [9:0] m248_24;
   assign m248_24 =10'b0;

   // m248_25 = W*in
   wire signed [9:0] m248_25;
   assign m248_25 ={ {5{in248[5]}} , in248[5:1] };

   // m248_26 = W*in
   wire signed [9:0] m248_26;
   assign m248_26 ={ {5{neg248[5]}} , neg248[5:1] };

   // m248_27 = W*in
   wire signed [9:0] m248_27;
   assign m248_27 =10'b0;

   // m248_28 = W*in
   wire signed [9:0] m248_28;
   assign m248_28 ={ {5{in248[5]}} , in248[5:1] };

   // m248_29 = W*in
   wire signed [9:0] m248_29;
   assign m248_29 =10'b0;

   // m248_30 = W*in
   wire signed [9:0] m248_30;
   assign m248_30 =10'b0;

   // m248_31 = W*in
   wire signed [9:0] m248_31;
   assign m248_31 =10'b0;

   // m248_32 = W*in
   wire signed [9:0] m248_32;
   assign m248_32 =10'b0;

   // m248_33 = W*in
   wire signed [9:0] m248_33;
   assign m248_33 =10'b0;

   // m248_34 = W*in
   wire signed [9:0] m248_34;
   assign m248_34 =10'b0;

   // m248_35 = W*in
   wire signed [9:0] m248_35;
   assign m248_35 =10'b0;

   // m248_36 = W*in
   wire signed [9:0] m248_36;
   assign m248_36 ={ {5{in248[5]}} , in248[5:1] };

   // m248_37 = W*in
   wire signed [9:0] m248_37;
   assign m248_37 =10'b0;

   // m248_38 = W*in
   wire signed [9:0] m248_38;
   assign m248_38 =10'b0;

   // m248_39 = W*in
   wire signed [9:0] m248_39;
   assign m248_39 =10'b0;

   // m248_40 = W*in
   wire signed [9:0] m248_40;
   assign m248_40 =10'b0;

   // m248_41 = W*in
   wire signed [9:0] m248_41;
   assign m248_41 =10'b0;

   // m248_42 = W*in
   wire signed [9:0] m248_42;
   assign m248_42 =10'b0;

   // m248_43 = W*in
   wire signed [9:0] m248_43;
   assign m248_43 =10'b0;

   // m248_44 = W*in
   wire signed [9:0] m248_44;
   assign m248_44 =10'b0;

   // m248_45 = W*in
   wire signed [9:0] m248_45;
   assign m248_45 =10'b0;

   // m248_46 = W*in
   wire signed [9:0] m248_46;
   assign m248_46 =10'b0;

   // m248_47 = W*in
   wire signed [9:0] m248_47;
   assign m248_47 =10'b0;

   // m248_48 = W*in
   wire signed [9:0] m248_48;
   assign m248_48 =10'b0;

   // m248_49 = W*in
   wire signed [9:0] m248_49;
   assign m248_49 =10'b0;

   // m248_50 = W*in
   wire signed [9:0] m248_50;
   assign m248_50 =10'b0;

   // m248_51 = W*in
   wire signed [9:0] m248_51;
   assign m248_51 =10'b0;

   // m248_52 = W*in
   wire signed [9:0] m248_52;
   assign m248_52 =10'b0;

   // m248_53 = W*in
   wire signed [9:0] m248_53;
   assign m248_53 =10'b0;

   // m248_54 = W*in
   wire signed [9:0] m248_54;
   assign m248_54 =10'b0;

   // m248_55 = W*in
   wire signed [9:0] m248_55;
   assign m248_55 =10'b0;

   // m248_56 = W*in
   wire signed [9:0] m248_56;
   assign m248_56 =10'b0;

   // m248_57 = W*in
   wire signed [9:0] m248_57;
   assign m248_57 =10'b0;

   // m248_58 = W*in
   wire signed [9:0] m248_58;
   assign m248_58 =10'b0;

   // m248_59 = W*in
   wire signed [9:0] m248_59;
   assign m248_59 =10'b0;

   // m248_60 = W*in
   wire signed [9:0] m248_60;
   assign m248_60 =10'b0;

   // m248_61 = W*in
   wire signed [9:0] m248_61;
   assign m248_61 =10'b0;

   // m248_62 = W*in
   wire signed [9:0] m248_62;
   assign m248_62 =10'b0;

   // m248_63 = W*in
   wire signed [9:0] m248_63;
   assign m248_63 =10'b0;

   // m248_64 = W*in
   wire signed [9:0] m248_64;
   assign m248_64 =10'b0;

   // m248_65 = W*in
   wire signed [9:0] m248_65;
   assign m248_65 =10'b0;

   // m248_66 = W*in
   wire signed [9:0] m248_66;
   assign m248_66 =10'b0;

   // m248_67 = W*in
   wire signed [9:0] m248_67;
   assign m248_67 =10'b0;

   // m248_68 = W*in
   wire signed [9:0] m248_68;
   assign m248_68 =10'b0;

   // m248_69 = W*in
   wire signed [9:0] m248_69;
   assign m248_69 =10'b0;

   // m248_70 = W*in
   wire signed [9:0] m248_70;
   assign m248_70 =10'b0;

   // m248_71 = W*in
   wire signed [9:0] m248_71;
   assign m248_71 =10'b0;

   // m248_72 = W*in
   wire signed [9:0] m248_72;
   assign m248_72 =10'b0;

   // m248_73 = W*in
   wire signed [9:0] m248_73;
   assign m248_73 ={ {5{in248[5]}} , in248[5:1] };

   // m248_74 = W*in
   wire signed [9:0] m248_74;
   assign m248_74 =10'b0;

   // m248_75 = W*in
   wire signed [9:0] m248_75;
   assign m248_75 =10'b0;

   // m248_76 = W*in
   wire signed [9:0] m248_76;
   assign m248_76 ={ {4{neg248[5]}} , neg248[5:0] };

   // m248_77 = W*in
   wire signed [9:0] m248_77;
   assign m248_77 =10'b0;

   // m248_78 = W*in
   wire signed [9:0] m248_78;
   assign m248_78 =10'b0;

   // m248_79 = W*in
   wire signed [9:0] m248_79;
   assign m248_79 =10'b0;

   // m248_80 = W*in
   wire signed [9:0] m248_80;
   assign m248_80 =10'b0;

   // m248_81 = W*in
   wire signed [9:0] m248_81;
   assign m248_81 =10'b0;

   // m248_82 = W*in
   wire signed [9:0] m248_82;
   assign m248_82 =10'b0;

   // m248_83 = W*in
   wire signed [9:0] m248_83;
   assign m248_83 =10'b0;

   // m248_84 = W*in
   wire signed [9:0] m248_84;
   assign m248_84 =10'b0;

   // m248_85 = W*in
   wire signed [9:0] m248_85;
   assign m248_85 =10'b0;

   // m248_86 = W*in
   wire signed [9:0] m248_86;
   assign m248_86 =10'b0;

   // m248_87 = W*in
   wire signed [9:0] m248_87;
   assign m248_87 =10'b0;

   // m248_88 = W*in
   wire signed [9:0] m248_88;
   assign m248_88 =10'b0;

   // m248_89 = W*in
   wire signed [9:0] m248_89;
   assign m248_89 =10'b0;

   // m248_90 = W*in
   wire signed [9:0] m248_90;
   assign m248_90 =10'b0;

   // m248_91 = W*in
   wire signed [9:0] m248_91;
   assign m248_91 =10'b0;

   // m248_92 = W*in
   wire signed [9:0] m248_92;
   assign m248_92 =10'b0;

   // m248_93 = W*in
   wire signed [9:0] m248_93;
   assign m248_93 =10'b0;

   // m248_94 = W*in
   wire signed [9:0] m248_94;
   assign m248_94 =10'b0;

   // m248_95 = W*in
   wire signed [9:0] m248_95;
   assign m248_95 =10'b0;

   // m248_96 = W*in
   wire signed [9:0] m248_96;
   assign m248_96 =10'b0;

   // m248_97 = W*in
   wire signed [9:0] m248_97;
   assign m248_97 =10'b0;

   // m248_98 = W*in
   wire signed [9:0] m248_98;
   assign m248_98 =10'b0;

   // m248_99 = W*in
   wire signed [9:0] m248_99;
   assign m248_99 =10'b0;

   // m248_100 = W*in
   wire signed [9:0] m248_100;
   assign m248_100 =10'b0;

   // m248_101 = W*in
   wire signed [9:0] m248_101;
   assign m248_101 =10'b0;

   // m248_102 = W*in
   wire signed [9:0] m248_102;
   assign m248_102 =10'b0;

   // m248_103 = W*in
   wire signed [9:0] m248_103;
   assign m248_103 =10'b0;

   // m248_104 = W*in
   wire signed [9:0] m248_104;
   assign m248_104 =10'b0;

   // m248_105 = W*in
   wire signed [9:0] m248_105;
   assign m248_105 =10'b0;

   // m248_106 = W*in
   wire signed [9:0] m248_106;
   assign m248_106 =10'b0;

   // m248_107 = W*in
   wire signed [9:0] m248_107;
   assign m248_107 =10'b0;

   // m248_108 = W*in
   wire signed [9:0] m248_108;
   assign m248_108 =10'b0;

   // m248_109 = W*in
   wire signed [9:0] m248_109;
   assign m248_109 ={ {5{in248[5]}} , in248[5:1] };

   // m248_110 = W*in
   wire signed [9:0] m248_110;
   assign m248_110 =10'b0;

   // m248_111 = W*in
   wire signed [9:0] m248_111;
   assign m248_111 =10'b0;

   // m248_112 = W*in
   wire signed [9:0] m248_112;
   assign m248_112 =10'b0;

   // m248_113 = W*in
   wire signed [9:0] m248_113;
   assign m248_113 =10'b0;

   // m248_114 = W*in
   wire signed [9:0] m248_114;
   assign m248_114 =10'b0;

   // m248_115 = W*in
   wire signed [9:0] m248_115;
   assign m248_115 =10'b0;

   // m248_116 = W*in
   wire signed [9:0] m248_116;
   assign m248_116 =10'b0;

   // m248_117 = W*in
   wire signed [9:0] m248_117;
   assign m248_117 =10'b0;

   // m249_1 = W*in
   wire signed [9:0] m249_1;
   assign m249_1 =10'b0;

   // m249_2 = W*in
   wire signed [9:0] m249_2;
   assign m249_2 =10'b0;

   // m249_3 = W*in
   wire signed [9:0] m249_3;
   assign m249_3 =10'b0;

   // m249_4 = W*in
   wire signed [9:0] m249_4;
   assign m249_4 =10'b0;

   // m249_5 = W*in
   wire signed [9:0] m249_5;
   assign m249_5 =10'b0;

   // m249_6 = W*in
   wire signed [9:0] m249_6;
   assign m249_6 =10'b0;

   // m249_7 = W*in
   wire signed [9:0] m249_7;
   assign m249_7 ={ {4{in249[5]}} , in249[5:0] };

   // m249_8 = W*in
   wire signed [9:0] m249_8;
   assign m249_8 =10'b0;

   // m249_9 = W*in
   wire signed [9:0] m249_9;
   assign m249_9 =10'b0;

   // m249_10 = W*in
   wire signed [9:0] m249_10;
   assign m249_10 =10'b0;

   // m249_11 = W*in
   wire signed [9:0] m249_11;
   assign m249_11 =10'b0;

   // m249_12 = W*in
   wire signed [9:0] m249_12;
   assign m249_12 =10'b0;

   // m249_13 = W*in
   wire signed [9:0] m249_13;
   assign m249_13 =10'b0;

   // m249_14 = W*in
   wire signed [9:0] m249_14;
   assign m249_14 =10'b0;

   // m249_15 = W*in
   wire signed [9:0] m249_15;
   assign m249_15 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_16 = W*in
   wire signed [9:0] m249_16;
   assign m249_16 =10'b0;

   // m249_17 = W*in
   wire signed [9:0] m249_17;
   assign m249_17 =10'b0;

   // m249_18 = W*in
   wire signed [9:0] m249_18;
   assign m249_18 ={ {5{in249[5]}} , in249[5:1] };

   // m249_19 = W*in
   wire signed [9:0] m249_19;
   assign m249_19 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_20 = W*in
   wire signed [9:0] m249_20;
   assign m249_20 =10'b0;

   // m249_21 = W*in
   wire signed [9:0] m249_21;
   assign m249_21 =10'b0;

   // m249_22 = W*in
   wire signed [9:0] m249_22;
   assign m249_22 =10'b0;

   // m249_23 = W*in
   wire signed [9:0] m249_23;
   assign m249_23 =10'b0;

   // m249_24 = W*in
   wire signed [9:0] m249_24;
   assign m249_24 =10'b0;

   // m249_25 = W*in
   wire signed [9:0] m249_25;
   assign m249_25 =10'b0;

   // m249_26 = W*in
   wire signed [9:0] m249_26;
   assign m249_26 ={ {4{in249[5]}} , in249[5:0] };

   // m249_27 = W*in
   wire signed [9:0] m249_27;
   assign m249_27 ={ {5{neg249[5]}} , neg249[5:1] };

   // m249_28 = W*in
   wire signed [9:0] m249_28;
   assign m249_28 =10'b0;

   // m249_29 = W*in
   wire signed [9:0] m249_29;
   assign m249_29 =10'b0;

   // m249_30 = W*in
   wire signed [9:0] m249_30;
   assign m249_30 =10'b0;

   // m249_31 = W*in
   wire signed [9:0] m249_31;
   assign m249_31 =10'b0;

   // m249_32 = W*in
   wire signed [9:0] m249_32;
   assign m249_32 =10'b0;

   // m249_33 = W*in
   wire signed [9:0] m249_33;
   assign m249_33 =10'b0;

   // m249_34 = W*in
   wire signed [9:0] m249_34;
   assign m249_34 ={ {5{in249[5]}} , in249[5:1] };

   // m249_35 = W*in
   wire signed [9:0] m249_35;
   assign m249_35 =10'b0;

   // m249_36 = W*in
   wire signed [9:0] m249_36;
   assign m249_36 =10'b0;

   // m249_37 = W*in
   wire signed [9:0] m249_37;
   assign m249_37 =10'b0;

   // m249_38 = W*in
   wire signed [9:0] m249_38;
   assign m249_38 =10'b0;

   // m249_39 = W*in
   wire signed [9:0] m249_39;
   assign m249_39 =10'b0;

   // m249_40 = W*in
   wire signed [9:0] m249_40;
   assign m249_40 =10'b0;

   // m249_41 = W*in
   wire signed [9:0] m249_41;
   assign m249_41 =10'b0;

   // m249_42 = W*in
   wire signed [9:0] m249_42;
   assign m249_42 =10'b0;

   // m249_43 = W*in
   wire signed [9:0] m249_43;
   assign m249_43 =10'b0;

   // m249_44 = W*in
   wire signed [9:0] m249_44;
   assign m249_44 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_45 = W*in
   wire signed [9:0] m249_45;
   assign m249_45 =10'b0;

   // m249_46 = W*in
   wire signed [9:0] m249_46;
   assign m249_46 =10'b0;

   // m249_47 = W*in
   wire signed [9:0] m249_47;
   assign m249_47 ={ {4{in249[5]}} , in249[5:0] };

   // m249_48 = W*in
   wire signed [9:0] m249_48;
   assign m249_48 =10'b0;

   // m249_49 = W*in
   wire signed [9:0] m249_49;
   assign m249_49 =10'b0;

   // m249_50 = W*in
   wire signed [9:0] m249_50;
   assign m249_50 =10'b0;

   // m249_51 = W*in
   wire signed [9:0] m249_51;
   assign m249_51 =10'b0;

   // m249_52 = W*in
   wire signed [9:0] m249_52;
   assign m249_52 =10'b0;

   // m249_53 = W*in
   wire signed [9:0] m249_53;
   assign m249_53 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_54 = W*in
   wire signed [9:0] m249_54;
   assign m249_54 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_55 = W*in
   wire signed [9:0] m249_55;
   assign m249_55 =10'b0;

   // m249_56 = W*in
   wire signed [9:0] m249_56;
   assign m249_56 =10'b0;

   // m249_57 = W*in
   wire signed [9:0] m249_57;
   assign m249_57 =10'b0;

   // m249_58 = W*in
   wire signed [9:0] m249_58;
   assign m249_58 =10'b0;

   // m249_59 = W*in
   wire signed [9:0] m249_59;
   assign m249_59 =10'b0;

   // m249_60 = W*in
   wire signed [9:0] m249_60;
   assign m249_60 =10'b0;

   // m249_61 = W*in
   wire signed [9:0] m249_61;
   assign m249_61 =10'b0;

   // m249_62 = W*in
   wire signed [9:0] m249_62;
   assign m249_62 =10'b0;

   // m249_63 = W*in
   wire signed [9:0] m249_63;
   assign m249_63 =10'b0;

   // m249_64 = W*in
   wire signed [9:0] m249_64;
   assign m249_64 ={ {5{in249[5]}} , in249[5:1] };

   // m249_65 = W*in
   wire signed [9:0] m249_65;
   assign m249_65 ={ {5{neg249[5]}} , neg249[5:1] };

   // m249_66 = W*in
   wire signed [9:0] m249_66;
   assign m249_66 =10'b0;

   // m249_67 = W*in
   wire signed [9:0] m249_67;
   assign m249_67 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_68 = W*in
   wire signed [9:0] m249_68;
   assign m249_68 =10'b0;

   // m249_69 = W*in
   wire signed [9:0] m249_69;
   assign m249_69 =10'b0;

   // m249_70 = W*in
   wire signed [9:0] m249_70;
   assign m249_70 =10'b0;

   // m249_71 = W*in
   wire signed [9:0] m249_71;
   assign m249_71 =10'b0;

   // m249_72 = W*in
   wire signed [9:0] m249_72;
   assign m249_72 ={ {5{in249[5]}} , in249[5:1] };

   // m249_73 = W*in
   wire signed [9:0] m249_73;
   assign m249_73 =10'b0;

   // m249_74 = W*in
   wire signed [9:0] m249_74;
   assign m249_74 =10'b0;

   // m249_75 = W*in
   wire signed [9:0] m249_75;
   assign m249_75 ={ {5{in249[5]}} , in249[5:1] };

   // m249_76 = W*in
   wire signed [9:0] m249_76;
   assign m249_76 =10'b0;

   // m249_77 = W*in
   wire signed [9:0] m249_77;
   assign m249_77 =10'b0;

   // m249_78 = W*in
   wire signed [9:0] m249_78;
   assign m249_78 ={ {4{in249[5]}} , in249[5:0] };

   // m249_79 = W*in
   wire signed [9:0] m249_79;
   assign m249_79 =10'b0;

   // m249_80 = W*in
   wire signed [9:0] m249_80;
   assign m249_80 =10'b0;

   // m249_81 = W*in
   wire signed [9:0] m249_81;
   assign m249_81 =10'b0;

   // m249_82 = W*in
   wire signed [9:0] m249_82;
   assign m249_82 =10'b0;

   // m249_83 = W*in
   wire signed [9:0] m249_83;
   assign m249_83 =10'b0;

   // m249_84 = W*in
   wire signed [9:0] m249_84;
   assign m249_84 =10'b0;

   // m249_85 = W*in
   wire signed [9:0] m249_85;
   assign m249_85 ={ {5{neg249[5]}} , neg249[5:1] };

   // m249_86 = W*in
   wire signed [9:0] m249_86;
   assign m249_86 =10'b0;

   // m249_87 = W*in
   wire signed [9:0] m249_87;
   assign m249_87 =10'b0;

   // m249_88 = W*in
   wire signed [9:0] m249_88;
   assign m249_88 =10'b0;

   // m249_89 = W*in
   wire signed [9:0] m249_89;
   assign m249_89 =10'b0;

   // m249_90 = W*in
   wire signed [9:0] m249_90;
   assign m249_90 =10'b0;

   // m249_91 = W*in
   wire signed [9:0] m249_91;
   assign m249_91 =10'b0;

   // m249_92 = W*in
   wire signed [9:0] m249_92;
   assign m249_92 =10'b0;

   // m249_93 = W*in
   wire signed [9:0] m249_93;
   assign m249_93 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_94 = W*in
   wire signed [9:0] m249_94;
   assign m249_94 =10'b0;

   // m249_95 = W*in
   wire signed [9:0] m249_95;
   assign m249_95 =10'b0;

   // m249_96 = W*in
   wire signed [9:0] m249_96;
   assign m249_96 =10'b0;

   // m249_97 = W*in
   wire signed [9:0] m249_97;
   assign m249_97 ={ {4{neg249[5]}} , neg249[5:0] };

   // m249_98 = W*in
   wire signed [9:0] m249_98;
   assign m249_98 =10'b0;

   // m249_99 = W*in
   wire signed [9:0] m249_99;
   assign m249_99 =10'b0;

   // m249_100 = W*in
   wire signed [9:0] m249_100;
   assign m249_100 =10'b0;

   // m249_101 = W*in
   wire signed [9:0] m249_101;
   assign m249_101 =10'b0;

   // m249_102 = W*in
   wire signed [9:0] m249_102;
   assign m249_102 =10'b0;

   // m249_103 = W*in
   wire signed [9:0] m249_103;
   assign m249_103 =10'b0;

   // m249_104 = W*in
   wire signed [9:0] m249_104;
   assign m249_104 =10'b0;

   // m249_105 = W*in
   wire signed [9:0] m249_105;
   assign m249_105 =10'b0;

   // m249_106 = W*in
   wire signed [9:0] m249_106;
   assign m249_106 =10'b0;

   // m249_107 = W*in
   wire signed [9:0] m249_107;
   assign m249_107 =10'b0;

   // m249_108 = W*in
   wire signed [9:0] m249_108;
   assign m249_108 =10'b0;

   // m249_109 = W*in
   wire signed [9:0] m249_109;
   assign m249_109 =10'b0;

   // m249_110 = W*in
   wire signed [9:0] m249_110;
   assign m249_110 =10'b0;

   // m249_111 = W*in
   wire signed [9:0] m249_111;
   assign m249_111 =10'b0;

   // m249_112 = W*in
   wire signed [9:0] m249_112;
   assign m249_112 =10'b0;

   // m249_113 = W*in
   wire signed [9:0] m249_113;
   assign m249_113 =10'b0;

   // m249_114 = W*in
   wire signed [9:0] m249_114;
   assign m249_114 =10'b0;

   // m249_115 = W*in
   wire signed [9:0] m249_115;
   assign m249_115 =10'b0;

   // m249_116 = W*in
   wire signed [9:0] m249_116;
   assign m249_116 =10'b0;

   // m249_117 = W*in
   wire signed [9:0] m249_117;
   assign m249_117 =10'b0;

   // m250_1 = W*in
   wire signed [9:0] m250_1;
   assign m250_1 =10'b0;

   // m250_2 = W*in
   wire signed [9:0] m250_2;
   assign m250_2 ={ {4{in250[5]}} , in250[5:0] };

   // m250_3 = W*in
   wire signed [9:0] m250_3;
   assign m250_3 =10'b0;

   // m250_4 = W*in
   wire signed [9:0] m250_4;
   assign m250_4 =10'b0;

   // m250_5 = W*in
   wire signed [9:0] m250_5;
   assign m250_5 =10'b0;

   // m250_6 = W*in
   wire signed [9:0] m250_6;
   assign m250_6 =10'b0;

   // m250_7 = W*in
   wire signed [9:0] m250_7;
   assign m250_7 =10'b0;

   // m250_8 = W*in
   wire signed [9:0] m250_8;
   assign m250_8 =10'b0;

   // m250_9 = W*in
   wire signed [9:0] m250_9;
   assign m250_9 =10'b0;

   // m250_10 = W*in
   wire signed [9:0] m250_10;
   assign m250_10 =10'b0;

   // m250_11 = W*in
   wire signed [9:0] m250_11;
   assign m250_11 =10'b0;

   // m250_12 = W*in
   wire signed [9:0] m250_12;
   assign m250_12 =10'b0;

   // m250_13 = W*in
   wire signed [9:0] m250_13;
   assign m250_13 =10'b0;

   // m250_14 = W*in
   wire signed [9:0] m250_14;
   assign m250_14 ={ {4{in250[5]}} , in250[5:0] };

   // m250_15 = W*in
   wire signed [9:0] m250_15;
   assign m250_15 ={ {4{in250[5]}} , in250[5:0] };

   // m250_16 = W*in
   wire signed [9:0] m250_16;
   assign m250_16 =10'b0;

   // m250_17 = W*in
   wire signed [9:0] m250_17;
   assign m250_17 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_18 = W*in
   wire signed [9:0] m250_18;
   assign m250_18 ={ {4{in250[5]}} , in250[5:0] };

   // m250_19 = W*in
   wire signed [9:0] m250_19;
   assign m250_19 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_20 = W*in
   wire signed [9:0] m250_20;
   assign m250_20 =10'b0;

   // m250_21 = W*in
   wire signed [9:0] m250_21;
   assign m250_21 =10'b0;

   // m250_22 = W*in
   wire signed [9:0] m250_22;
   assign m250_22 =10'b0;

   // m250_23 = W*in
   wire signed [9:0] m250_23;
   assign m250_23 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_24 = W*in
   wire signed [9:0] m250_24;
   assign m250_24 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_25 = W*in
   wire signed [9:0] m250_25;
   assign m250_25 =10'b0;

   // m250_26 = W*in
   wire signed [9:0] m250_26;
   assign m250_26 ={ {4{in250[5]}} , in250[5:0] };

   // m250_27 = W*in
   wire signed [9:0] m250_27;
   assign m250_27 ={ {5{neg250[5]}} , neg250[5:1] };

   // m250_28 = W*in
   wire signed [9:0] m250_28;
   assign m250_28 =10'b0;

   // m250_29 = W*in
   wire signed [9:0] m250_29;
   assign m250_29 =10'b0;

   // m250_30 = W*in
   wire signed [9:0] m250_30;
   assign m250_30 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_31 = W*in
   wire signed [9:0] m250_31;
   assign m250_31 ={ {5{neg250[5]}} , neg250[5:1] };

   // m250_32 = W*in
   wire signed [9:0] m250_32;
   assign m250_32 =10'b0;

   // m250_33 = W*in
   wire signed [9:0] m250_33;
   assign m250_33 =10'b0;

   // m250_34 = W*in
   wire signed [9:0] m250_34;
   assign m250_34 =10'b0;

   // m250_35 = W*in
   wire signed [9:0] m250_35;
   assign m250_35 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_36 = W*in
   wire signed [9:0] m250_36;
   assign m250_36 ={ {4{in250[5]}} , in250[5:0] };

   // m250_37 = W*in
   wire signed [9:0] m250_37;
   assign m250_37 =10'b0;

   // m250_38 = W*in
   wire signed [9:0] m250_38;
   assign m250_38 ={ {4{in250[5]}} , in250[5:0] };

   // m250_39 = W*in
   wire signed [9:0] m250_39;
   assign m250_39 =10'b0;

   // m250_40 = W*in
   wire signed [9:0] m250_40;
   assign m250_40 =10'b0;

   // m250_41 = W*in
   wire signed [9:0] m250_41;
   assign m250_41 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_42 = W*in
   wire signed [9:0] m250_42;
   assign m250_42 =10'b0;

   // m250_43 = W*in
   wire signed [9:0] m250_43;
   assign m250_43 ={ {4{in250[5]}} , in250[5:0] };

   // m250_44 = W*in
   wire signed [9:0] m250_44;
   assign m250_44 ={ {3{neg250[5]}} , neg250 , {1{1'b0}} };

   // m250_45 = W*in
   wire signed [9:0] m250_45;
   assign m250_45 ={ {4{in250[5]}} , in250[5:0] };

   // m250_46 = W*in
   wire signed [9:0] m250_46;
   assign m250_46 =10'b0;

   // m250_47 = W*in
   wire signed [9:0] m250_47;
   assign m250_47 ={ {4{in250[5]}} , in250[5:0] };

   // m250_48 = W*in
   wire signed [9:0] m250_48;
   assign m250_48 ={ {4{in250[5]}} , in250[5:0] };

   // m250_49 = W*in
   wire signed [9:0] m250_49;
   assign m250_49 =10'b0;

   // m250_50 = W*in
   wire signed [9:0] m250_50;
   assign m250_50 =10'b0;

   // m250_51 = W*in
   wire signed [9:0] m250_51;
   assign m250_51 =10'b0;

   // m250_52 = W*in
   wire signed [9:0] m250_52;
   assign m250_52 =10'b0;

   // m250_53 = W*in
   wire signed [9:0] m250_53;
   assign m250_53 =10'b0;

   // m250_54 = W*in
   wire signed [9:0] m250_54;
   assign m250_54 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_55 = W*in
   wire signed [9:0] m250_55;
   assign m250_55 =10'b0;

   // m250_56 = W*in
   wire signed [9:0] m250_56;
   assign m250_56 =10'b0;

   // m250_57 = W*in
   wire signed [9:0] m250_57;
   assign m250_57 =10'b0;

   // m250_58 = W*in
   wire signed [9:0] m250_58;
   assign m250_58 =10'b0;

   // m250_59 = W*in
   wire signed [9:0] m250_59;
   assign m250_59 =10'b0;

   // m250_60 = W*in
   wire signed [9:0] m250_60;
   assign m250_60 =10'b0;

   // m250_61 = W*in
   wire signed [9:0] m250_61;
   assign m250_61 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_62 = W*in
   wire signed [9:0] m250_62;
   assign m250_62 =10'b0;

   // m250_63 = W*in
   wire signed [9:0] m250_63;
   assign m250_63 =10'b0;

   // m250_64 = W*in
   wire signed [9:0] m250_64;
   assign m250_64 =10'b0;

   // m250_65 = W*in
   wire signed [9:0] m250_65;
   assign m250_65 ={ {5{neg250[5]}} , neg250[5:1] };

   // m250_66 = W*in
   wire signed [9:0] m250_66;
   assign m250_66 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_67 = W*in
   wire signed [9:0] m250_67;
   assign m250_67 =10'b0;

   // m250_68 = W*in
   wire signed [9:0] m250_68;
   assign m250_68 ={ {4{in250[5]}} , in250[5:0] };

   // m250_69 = W*in
   wire signed [9:0] m250_69;
   assign m250_69 ={ {4{in250[5]}} , in250[5:0] };

   // m250_70 = W*in
   wire signed [9:0] m250_70;
   assign m250_70 ={ {4{in250[5]}} , in250[5:0] };

   // m250_71 = W*in
   wire signed [9:0] m250_71;
   assign m250_71 ={ {5{in250[5]}} , in250[5:1] };

   // m250_72 = W*in
   wire signed [9:0] m250_72;
   assign m250_72 ={ {4{in250[5]}} , in250[5:0] };

   // m250_73 = W*in
   wire signed [9:0] m250_73;
   assign m250_73 =10'b0;

   // m250_74 = W*in
   wire signed [9:0] m250_74;
   assign m250_74 ={ {4{in250[5]}} , in250[5:0] };

   // m250_75 = W*in
   wire signed [9:0] m250_75;
   assign m250_75 =10'b0;

   // m250_76 = W*in
   wire signed [9:0] m250_76;
   assign m250_76 =10'b0;

   // m250_77 = W*in
   wire signed [9:0] m250_77;
   assign m250_77 =10'b0;

   // m250_78 = W*in
   wire signed [9:0] m250_78;
   assign m250_78 ={ {4{in250[5]}} , in250[5:0] };

   // m250_79 = W*in
   wire signed [9:0] m250_79;
   assign m250_79 =10'b0;

   // m250_80 = W*in
   wire signed [9:0] m250_80;
   assign m250_80 =10'b0;

   // m250_81 = W*in
   wire signed [9:0] m250_81;
   assign m250_81 =10'b0;

   // m250_82 = W*in
   wire signed [9:0] m250_82;
   assign m250_82 =10'b0;

   // m250_83 = W*in
   wire signed [9:0] m250_83;
   assign m250_83 =10'b0;

   // m250_84 = W*in
   wire signed [9:0] m250_84;
   assign m250_84 ={ {4{in250[5]}} , in250[5:0] };

   // m250_85 = W*in
   wire signed [9:0] m250_85;
   assign m250_85 =10'b0;

   // m250_86 = W*in
   wire signed [9:0] m250_86;
   assign m250_86 ={ {4{in250[5]}} , in250[5:0] };

   // m250_87 = W*in
   wire signed [9:0] m250_87;
   assign m250_87 ={ {4{in250[5]}} , in250[5:0] };

   // m250_88 = W*in
   wire signed [9:0] m250_88;
   assign m250_88 ={ {4{in250[5]}} , in250[5:0] };

   // m250_89 = W*in
   wire signed [9:0] m250_89;
   assign m250_89 =10'b0;

   // m250_90 = W*in
   wire signed [9:0] m250_90;
   assign m250_90 ={ {4{in250[5]}} , in250[5:0] };

   // m250_91 = W*in
   wire signed [9:0] m250_91;
   assign m250_91 =10'b0;

   // m250_92 = W*in
   wire signed [9:0] m250_92;
   assign m250_92 =10'b0;

   // m250_93 = W*in
   wire signed [9:0] m250_93;
   assign m250_93 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_94 = W*in
   wire signed [9:0] m250_94;
   assign m250_94 =10'b0;

   // m250_95 = W*in
   wire signed [9:0] m250_95;
   assign m250_95 =10'b0;

   // m250_96 = W*in
   wire signed [9:0] m250_96;
   assign m250_96 =10'b0;

   // m250_97 = W*in
   wire signed [9:0] m250_97;
   assign m250_97 =10'b0;

   // m250_98 = W*in
   wire signed [9:0] m250_98;
   assign m250_98 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_99 = W*in
   wire signed [9:0] m250_99;
   assign m250_99 ={ {4{in250[5]}} , in250[5:0] };

   // m250_100 = W*in
   wire signed [9:0] m250_100;
   assign m250_100 =10'b0;

   // m250_101 = W*in
   wire signed [9:0] m250_101;
   assign m250_101 =10'b0;

   // m250_102 = W*in
   wire signed [9:0] m250_102;
   assign m250_102 =10'b0;

   // m250_103 = W*in
   wire signed [9:0] m250_103;
   assign m250_103 =10'b0;

   // m250_104 = W*in
   wire signed [9:0] m250_104;
   assign m250_104 =10'b0;

   // m250_105 = W*in
   wire signed [9:0] m250_105;
   assign m250_105 =10'b0;

   // m250_106 = W*in
   wire signed [9:0] m250_106;
   assign m250_106 =10'b0;

   // m250_107 = W*in
   wire signed [9:0] m250_107;
   assign m250_107 =10'b0;

   // m250_108 = W*in
   wire signed [9:0] m250_108;
   assign m250_108 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_109 = W*in
   wire signed [9:0] m250_109;
   assign m250_109 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_110 = W*in
   wire signed [9:0] m250_110;
   assign m250_110 ={ {4{neg250[5]}} , neg250[5:0] };

   // m250_111 = W*in
   wire signed [9:0] m250_111;
   assign m250_111 ={ {4{in250[5]}} , in250[5:0] };

   // m250_112 = W*in
   wire signed [9:0] m250_112;
   assign m250_112 =10'b0;

   // m250_113 = W*in
   wire signed [9:0] m250_113;
   assign m250_113 =10'b0;

   // m250_114 = W*in
   wire signed [9:0] m250_114;
   assign m250_114 =10'b0;

   // m250_115 = W*in
   wire signed [9:0] m250_115;
   assign m250_115 ={ {5{neg250[5]}} , neg250[5:1] };

   // m250_116 = W*in
   wire signed [9:0] m250_116;
   assign m250_116 =10'b0;

   // m250_117 = W*in
   wire signed [9:0] m250_117;
   assign m250_117 ={ {4{neg250[5]}} , neg250[5:0] };

   // m251_1 = W*in
   wire signed [9:0] m251_1;
   assign m251_1 ={ {4{in251[5]}} , in251[5:0] };

   // m251_2 = W*in
   wire signed [9:0] m251_2;
   assign m251_2 =10'b0;

   // m251_3 = W*in
   wire signed [9:0] m251_3;
   assign m251_3 =10'b0;

   // m251_4 = W*in
   wire signed [9:0] m251_4;
   assign m251_4 =10'b0;

   // m251_5 = W*in
   wire signed [9:0] m251_5;
   assign m251_5 ={ {4{in251[5]}} , in251[5:0] };

   // m251_6 = W*in
   wire signed [9:0] m251_6;
   assign m251_6 =10'b0;

   // m251_7 = W*in
   wire signed [9:0] m251_7;
   assign m251_7 ={ {4{in251[5]}} , in251[5:0] };

   // m251_8 = W*in
   wire signed [9:0] m251_8;
   assign m251_8 =10'b0;

   // m251_9 = W*in
   wire signed [9:0] m251_9;
   assign m251_9 =10'b0;

   // m251_10 = W*in
   wire signed [9:0] m251_10;
   assign m251_10 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_11 = W*in
   wire signed [9:0] m251_11;
   assign m251_11 =10'b0;

   // m251_12 = W*in
   wire signed [9:0] m251_12;
   assign m251_12 =10'b0;

   // m251_13 = W*in
   wire signed [9:0] m251_13;
   assign m251_13 ={ {4{in251[5]}} , in251[5:0] };

   // m251_14 = W*in
   wire signed [9:0] m251_14;
   assign m251_14 =10'b0;

   // m251_15 = W*in
   wire signed [9:0] m251_15;
   assign m251_15 =10'b0;

   // m251_16 = W*in
   wire signed [9:0] m251_16;
   assign m251_16 ={ {4{in251[5]}} , in251[5:0] };

   // m251_17 = W*in
   wire signed [9:0] m251_17;
   assign m251_17 =10'b0;

   // m251_18 = W*in
   wire signed [9:0] m251_18;
   assign m251_18 ={ {5{neg251[5]}} , neg251[5:1] };

   // m251_19 = W*in
   wire signed [9:0] m251_19;
   assign m251_19 =10'b0;

   // m251_20 = W*in
   wire signed [9:0] m251_20;
   assign m251_20 =10'b0;

   // m251_21 = W*in
   wire signed [9:0] m251_21;
   assign m251_21 =10'b0;

   // m251_22 = W*in
   wire signed [9:0] m251_22;
   assign m251_22 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_23 = W*in
   wire signed [9:0] m251_23;
   assign m251_23 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_24 = W*in
   wire signed [9:0] m251_24;
   assign m251_24 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_25 = W*in
   wire signed [9:0] m251_25;
   assign m251_25 ={ {4{in251[5]}} , in251[5:0] };

   // m251_26 = W*in
   wire signed [9:0] m251_26;
   assign m251_26 =10'b0;

   // m251_27 = W*in
   wire signed [9:0] m251_27;
   assign m251_27 ={ {5{neg251[5]}} , neg251[5:1] };

   // m251_28 = W*in
   wire signed [9:0] m251_28;
   assign m251_28 ={ {4{in251[5]}} , in251[5:0] };

   // m251_29 = W*in
   wire signed [9:0] m251_29;
   assign m251_29 =10'b0;

   // m251_30 = W*in
   wire signed [9:0] m251_30;
   assign m251_30 =10'b0;

   // m251_31 = W*in
   wire signed [9:0] m251_31;
   assign m251_31 =10'b0;

   // m251_32 = W*in
   wire signed [9:0] m251_32;
   assign m251_32 =10'b0;

   // m251_33 = W*in
   wire signed [9:0] m251_33;
   assign m251_33 ={ {4{in251[5]}} , in251[5:0] };

   // m251_34 = W*in
   wire signed [9:0] m251_34;
   assign m251_34 =10'b0;

   // m251_35 = W*in
   wire signed [9:0] m251_35;
   assign m251_35 =10'b0;

   // m251_36 = W*in
   wire signed [9:0] m251_36;
   assign m251_36 ={ {4{in251[5]}} , in251[5:0] };

   // m251_37 = W*in
   wire signed [9:0] m251_37;
   assign m251_37 =10'b0;

   // m251_38 = W*in
   wire signed [9:0] m251_38;
   assign m251_38 =10'b0;

   // m251_39 = W*in
   wire signed [9:0] m251_39;
   assign m251_39 =10'b0;

   // m251_40 = W*in
   wire signed [9:0] m251_40;
   assign m251_40 =10'b0;

   // m251_41 = W*in
   wire signed [9:0] m251_41;
   assign m251_41 =10'b0;

   // m251_42 = W*in
   wire signed [9:0] m251_42;
   assign m251_42 =10'b0;

   // m251_43 = W*in
   wire signed [9:0] m251_43;
   assign m251_43 =10'b0;

   // m251_44 = W*in
   wire signed [9:0] m251_44;
   assign m251_44 =10'b0;

   // m251_45 = W*in
   wire signed [9:0] m251_45;
   assign m251_45 =10'b0;

   // m251_46 = W*in
   wire signed [9:0] m251_46;
   assign m251_46 =10'b0;

   // m251_47 = W*in
   wire signed [9:0] m251_47;
   assign m251_47 =10'b0;

   // m251_48 = W*in
   wire signed [9:0] m251_48;
   assign m251_48 ={ {4{in251[5]}} , in251[5:0] };

   // m251_49 = W*in
   wire signed [9:0] m251_49;
   assign m251_49 =10'b0;

   // m251_50 = W*in
   wire signed [9:0] m251_50;
   assign m251_50 =10'b0;

   // m251_51 = W*in
   wire signed [9:0] m251_51;
   assign m251_51 =10'b0;

   // m251_52 = W*in
   wire signed [9:0] m251_52;
   assign m251_52 =10'b0;

   // m251_53 = W*in
   wire signed [9:0] m251_53;
   assign m251_53 ={ {4{in251[5]}} , in251[5:0] };

   // m251_54 = W*in
   wire signed [9:0] m251_54;
   assign m251_54 ={ {4{in251[5]}} , in251[5:0] };

   // m251_55 = W*in
   wire signed [9:0] m251_55;
   assign m251_55 =10'b0;

   // m251_56 = W*in
   wire signed [9:0] m251_56;
   assign m251_56 =10'b0;

   // m251_57 = W*in
   wire signed [9:0] m251_57;
   assign m251_57 =10'b0;

   // m251_58 = W*in
   wire signed [9:0] m251_58;
   assign m251_58 =10'b0;

   // m251_59 = W*in
   wire signed [9:0] m251_59;
   assign m251_59 ={ {4{in251[5]}} , in251[5:0] };

   // m251_60 = W*in
   wire signed [9:0] m251_60;
   assign m251_60 =10'b0;

   // m251_61 = W*in
   wire signed [9:0] m251_61;
   assign m251_61 =10'b0;

   // m251_62 = W*in
   wire signed [9:0] m251_62;
   assign m251_62 =10'b0;

   // m251_63 = W*in
   wire signed [9:0] m251_63;
   assign m251_63 =10'b0;

   // m251_64 = W*in
   wire signed [9:0] m251_64;
   assign m251_64 =10'b0;

   // m251_65 = W*in
   wire signed [9:0] m251_65;
   assign m251_65 =10'b0;

   // m251_66 = W*in
   wire signed [9:0] m251_66;
   assign m251_66 =10'b0;

   // m251_67 = W*in
   wire signed [9:0] m251_67;
   assign m251_67 =10'b0;

   // m251_68 = W*in
   wire signed [9:0] m251_68;
   assign m251_68 =10'b0;

   // m251_69 = W*in
   wire signed [9:0] m251_69;
   assign m251_69 =10'b0;

   // m251_70 = W*in
   wire signed [9:0] m251_70;
   assign m251_70 =10'b0;

   // m251_71 = W*in
   wire signed [9:0] m251_71;
   assign m251_71 =10'b0;

   // m251_72 = W*in
   wire signed [9:0] m251_72;
   assign m251_72 ={ {5{in251[5]}} , in251[5:1] };

   // m251_73 = W*in
   wire signed [9:0] m251_73;
   assign m251_73 ={ {4{in251[5]}} , in251[5:0] };

   // m251_74 = W*in
   wire signed [9:0] m251_74;
   assign m251_74 =10'b0;

   // m251_75 = W*in
   wire signed [9:0] m251_75;
   assign m251_75 =10'b0;

   // m251_76 = W*in
   wire signed [9:0] m251_76;
   assign m251_76 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_77 = W*in
   wire signed [9:0] m251_77;
   assign m251_77 =10'b0;

   // m251_78 = W*in
   wire signed [9:0] m251_78;
   assign m251_78 =10'b0;

   // m251_79 = W*in
   wire signed [9:0] m251_79;
   assign m251_79 =10'b0;

   // m251_80 = W*in
   wire signed [9:0] m251_80;
   assign m251_80 =10'b0;

   // m251_81 = W*in
   wire signed [9:0] m251_81;
   assign m251_81 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_82 = W*in
   wire signed [9:0] m251_82;
   assign m251_82 =10'b0;

   // m251_83 = W*in
   wire signed [9:0] m251_83;
   assign m251_83 =10'b0;

   // m251_84 = W*in
   wire signed [9:0] m251_84;
   assign m251_84 =10'b0;

   // m251_85 = W*in
   wire signed [9:0] m251_85;
   assign m251_85 =10'b0;

   // m251_86 = W*in
   wire signed [9:0] m251_86;
   assign m251_86 =10'b0;

   // m251_87 = W*in
   wire signed [9:0] m251_87;
   assign m251_87 =10'b0;

   // m251_88 = W*in
   wire signed [9:0] m251_88;
   assign m251_88 =10'b0;

   // m251_89 = W*in
   wire signed [9:0] m251_89;
   assign m251_89 =10'b0;

   // m251_90 = W*in
   wire signed [9:0] m251_90;
   assign m251_90 =10'b0;

   // m251_91 = W*in
   wire signed [9:0] m251_91;
   assign m251_91 =10'b0;

   // m251_92 = W*in
   wire signed [9:0] m251_92;
   assign m251_92 =10'b0;

   // m251_93 = W*in
   wire signed [9:0] m251_93;
   assign m251_93 =10'b0;

   // m251_94 = W*in
   wire signed [9:0] m251_94;
   assign m251_94 ={ {4{neg251[5]}} , neg251[5:0] };

   // m251_95 = W*in
   wire signed [9:0] m251_95;
   assign m251_95 =10'b0;

   // m251_96 = W*in
   wire signed [9:0] m251_96;
   assign m251_96 =10'b0;

   // m251_97 = W*in
   wire signed [9:0] m251_97;
   assign m251_97 =10'b0;

   // m251_98 = W*in
   wire signed [9:0] m251_98;
   assign m251_98 =10'b0;

   // m251_99 = W*in
   wire signed [9:0] m251_99;
   assign m251_99 =10'b0;

   // m251_100 = W*in
   wire signed [9:0] m251_100;
   assign m251_100 =10'b0;

   // m251_101 = W*in
   wire signed [9:0] m251_101;
   assign m251_101 =10'b0;

   // m251_102 = W*in
   wire signed [9:0] m251_102;
   assign m251_102 ={ {4{in251[5]}} , in251[5:0] };

   // m251_103 = W*in
   wire signed [9:0] m251_103;
   assign m251_103 =10'b0;

   // m251_104 = W*in
   wire signed [9:0] m251_104;
   assign m251_104 =10'b0;

   // m251_105 = W*in
   wire signed [9:0] m251_105;
   assign m251_105 =10'b0;

   // m251_106 = W*in
   wire signed [9:0] m251_106;
   assign m251_106 ={ {4{in251[5]}} , in251[5:0] };

   // m251_107 = W*in
   wire signed [9:0] m251_107;
   assign m251_107 =10'b0;

   // m251_108 = W*in
   wire signed [9:0] m251_108;
   assign m251_108 =10'b0;

   // m251_109 = W*in
   wire signed [9:0] m251_109;
   assign m251_109 =10'b0;

   // m251_110 = W*in
   wire signed [9:0] m251_110;
   assign m251_110 =10'b0;

   // m251_111 = W*in
   wire signed [9:0] m251_111;
   assign m251_111 =10'b0;

   // m251_112 = W*in
   wire signed [9:0] m251_112;
   assign m251_112 =10'b0;

   // m251_113 = W*in
   wire signed [9:0] m251_113;
   assign m251_113 =10'b0;

   // m251_114 = W*in
   wire signed [9:0] m251_114;
   assign m251_114 ={ {5{neg251[5]}} , neg251[5:1] };

   // m251_115 = W*in
   wire signed [9:0] m251_115;
   assign m251_115 =10'b0;

   // m251_116 = W*in
   wire signed [9:0] m251_116;
   assign m251_116 =10'b0;

   // m251_117 = W*in
   wire signed [9:0] m251_117;
   assign m251_117 =10'b0;

   // m252_1 = W*in
   wire signed [9:0] m252_1;
   assign m252_1 =10'b0;

   // m252_2 = W*in
   wire signed [9:0] m252_2;
   assign m252_2 =10'b0;

   // m252_3 = W*in
   wire signed [9:0] m252_3;
   assign m252_3 =10'b0;

   // m252_4 = W*in
   wire signed [9:0] m252_4;
   assign m252_4 =10'b0;

   // m252_5 = W*in
   wire signed [9:0] m252_5;
   assign m252_5 =10'b0;

   // m252_6 = W*in
   wire signed [9:0] m252_6;
   assign m252_6 =10'b0;

   // m252_7 = W*in
   wire signed [9:0] m252_7;
   assign m252_7 =10'b0;

   // m252_8 = W*in
   wire signed [9:0] m252_8;
   assign m252_8 =10'b0;

   // m252_9 = W*in
   wire signed [9:0] m252_9;
   assign m252_9 =10'b0;

   // m252_10 = W*in
   wire signed [9:0] m252_10;
   assign m252_10 =10'b0;

   // m252_11 = W*in
   wire signed [9:0] m252_11;
   assign m252_11 =10'b0;

   // m252_12 = W*in
   wire signed [9:0] m252_12;
   assign m252_12 =10'b0;

   // m252_13 = W*in
   wire signed [9:0] m252_13;
   assign m252_13 =10'b0;

   // m252_14 = W*in
   wire signed [9:0] m252_14;
   assign m252_14 =10'b0;

   // m252_15 = W*in
   wire signed [9:0] m252_15;
   assign m252_15 =10'b0;

   // m252_16 = W*in
   wire signed [9:0] m252_16;
   assign m252_16 =10'b0;

   // m252_17 = W*in
   wire signed [9:0] m252_17;
   assign m252_17 =10'b0;

   // m252_18 = W*in
   wire signed [9:0] m252_18;
   assign m252_18 =10'b0;

   // m252_19 = W*in
   wire signed [9:0] m252_19;
   assign m252_19 =10'b0;

   // m252_20 = W*in
   wire signed [9:0] m252_20;
   assign m252_20 ={ {5{neg252[5]}} , neg252[5:1] };

   // m252_21 = W*in
   wire signed [9:0] m252_21;
   assign m252_21 =10'b0;

   // m252_22 = W*in
   wire signed [9:0] m252_22;
   assign m252_22 =10'b0;

   // m252_23 = W*in
   wire signed [9:0] m252_23;
   assign m252_23 =10'b0;

   // m252_24 = W*in
   wire signed [9:0] m252_24;
   assign m252_24 =10'b0;

   // m252_25 = W*in
   wire signed [9:0] m252_25;
   assign m252_25 =10'b0;

   // m252_26 = W*in
   wire signed [9:0] m252_26;
   assign m252_26 ={ {5{neg252[5]}} , neg252[5:1] };

   // m252_27 = W*in
   wire signed [9:0] m252_27;
   assign m252_27 =10'b0;

   // m252_28 = W*in
   wire signed [9:0] m252_28;
   assign m252_28 =10'b0;

   // m252_29 = W*in
   wire signed [9:0] m252_29;
   assign m252_29 ={ {4{neg252[5]}} , neg252[5:0] };

   // m252_30 = W*in
   wire signed [9:0] m252_30;
   assign m252_30 =10'b0;

   // m252_31 = W*in
   wire signed [9:0] m252_31;
   assign m252_31 =10'b0;

   // m252_32 = W*in
   wire signed [9:0] m252_32;
   assign m252_32 ={ {4{in252[5]}} , in252[5:0] };

   // m252_33 = W*in
   wire signed [9:0] m252_33;
   assign m252_33 =10'b0;

   // m252_34 = W*in
   wire signed [9:0] m252_34;
   assign m252_34 ={ {4{neg252[5]}} , neg252[5:0] };

   // m252_35 = W*in
   wire signed [9:0] m252_35;
   assign m252_35 =10'b0;

   // m252_36 = W*in
   wire signed [9:0] m252_36;
   assign m252_36 ={ {5{in252[5]}} , in252[5:1] };

   // m252_37 = W*in
   wire signed [9:0] m252_37;
   assign m252_37 ={ {4{in252[5]}} , in252[5:0] };

   // m252_38 = W*in
   wire signed [9:0] m252_38;
   assign m252_38 =10'b0;

   // m252_39 = W*in
   wire signed [9:0] m252_39;
   assign m252_39 =10'b0;

   // m252_40 = W*in
   wire signed [9:0] m252_40;
   assign m252_40 ={ {4{in252[5]}} , in252[5:0] };

   // m252_41 = W*in
   wire signed [9:0] m252_41;
   assign m252_41 =10'b0;

   // m252_42 = W*in
   wire signed [9:0] m252_42;
   assign m252_42 =10'b0;

   // m252_43 = W*in
   wire signed [9:0] m252_43;
   assign m252_43 =10'b0;

   // m252_44 = W*in
   wire signed [9:0] m252_44;
   assign m252_44 ={ {4{in252[5]}} , in252[5:0] };

   // m252_45 = W*in
   wire signed [9:0] m252_45;
   assign m252_45 =10'b0;

   // m252_46 = W*in
   wire signed [9:0] m252_46;
   assign m252_46 =10'b0;

   // m252_47 = W*in
   wire signed [9:0] m252_47;
   assign m252_47 =10'b0;

   // m252_48 = W*in
   wire signed [9:0] m252_48;
   assign m252_48 =10'b0;

   // m252_49 = W*in
   wire signed [9:0] m252_49;
   assign m252_49 =10'b0;

   // m252_50 = W*in
   wire signed [9:0] m252_50;
   assign m252_50 =10'b0;

   // m252_51 = W*in
   wire signed [9:0] m252_51;
   assign m252_51 =10'b0;

   // m252_52 = W*in
   wire signed [9:0] m252_52;
   assign m252_52 =10'b0;

   // m252_53 = W*in
   wire signed [9:0] m252_53;
   assign m252_53 =10'b0;

   // m252_54 = W*in
   wire signed [9:0] m252_54;
   assign m252_54 ={ {4{in252[5]}} , in252[5:0] };

   // m252_55 = W*in
   wire signed [9:0] m252_55;
   assign m252_55 =10'b0;

   // m252_56 = W*in
   wire signed [9:0] m252_56;
   assign m252_56 =10'b0;

   // m252_57 = W*in
   wire signed [9:0] m252_57;
   assign m252_57 =10'b0;

   // m252_58 = W*in
   wire signed [9:0] m252_58;
   assign m252_58 =10'b0;

   // m252_59 = W*in
   wire signed [9:0] m252_59;
   assign m252_59 =10'b0;

   // m252_60 = W*in
   wire signed [9:0] m252_60;
   assign m252_60 =10'b0;

   // m252_61 = W*in
   wire signed [9:0] m252_61;
   assign m252_61 =10'b0;

   // m252_62 = W*in
   wire signed [9:0] m252_62;
   assign m252_62 =10'b0;

   // m252_63 = W*in
   wire signed [9:0] m252_63;
   assign m252_63 =10'b0;

   // m252_64 = W*in
   wire signed [9:0] m252_64;
   assign m252_64 ={ {5{neg252[5]}} , neg252[5:1] };

   // m252_65 = W*in
   wire signed [9:0] m252_65;
   assign m252_65 =10'b0;

   // m252_66 = W*in
   wire signed [9:0] m252_66;
   assign m252_66 =10'b0;

   // m252_67 = W*in
   wire signed [9:0] m252_67;
   assign m252_67 =10'b0;

   // m252_68 = W*in
   wire signed [9:0] m252_68;
   assign m252_68 =10'b0;

   // m252_69 = W*in
   wire signed [9:0] m252_69;
   assign m252_69 =10'b0;

   // m252_70 = W*in
   wire signed [9:0] m252_70;
   assign m252_70 ={ {4{neg252[5]}} , neg252[5:0] };

   // m252_71 = W*in
   wire signed [9:0] m252_71;
   assign m252_71 =10'b0;

   // m252_72 = W*in
   wire signed [9:0] m252_72;
   assign m252_72 ={ {5{neg252[5]}} , neg252[5:1] };

   // m252_73 = W*in
   wire signed [9:0] m252_73;
   assign m252_73 =10'b0;

   // m252_74 = W*in
   wire signed [9:0] m252_74;
   assign m252_74 ={ {5{neg252[5]}} , neg252[5:1] };

   // m252_75 = W*in
   wire signed [9:0] m252_75;
   assign m252_75 =10'b0;

   // m252_76 = W*in
   wire signed [9:0] m252_76;
   assign m252_76 ={ {4{neg252[5]}} , neg252[5:0] };

   // m252_77 = W*in
   wire signed [9:0] m252_77;
   assign m252_77 =10'b0;

   // m252_78 = W*in
   wire signed [9:0] m252_78;
   assign m252_78 =10'b0;

   // m252_79 = W*in
   wire signed [9:0] m252_79;
   assign m252_79 =10'b0;

   // m252_80 = W*in
   wire signed [9:0] m252_80;
   assign m252_80 =10'b0;

   // m252_81 = W*in
   wire signed [9:0] m252_81;
   assign m252_81 =10'b0;

   // m252_82 = W*in
   wire signed [9:0] m252_82;
   assign m252_82 =10'b0;

   // m252_83 = W*in
   wire signed [9:0] m252_83;
   assign m252_83 =10'b0;

   // m252_84 = W*in
   wire signed [9:0] m252_84;
   assign m252_84 =10'b0;

   // m252_85 = W*in
   wire signed [9:0] m252_85;
   assign m252_85 ={ {5{in252[5]}} , in252[5:1] };

   // m252_86 = W*in
   wire signed [9:0] m252_86;
   assign m252_86 =10'b0;

   // m252_87 = W*in
   wire signed [9:0] m252_87;
   assign m252_87 =10'b0;

   // m252_88 = W*in
   wire signed [9:0] m252_88;
   assign m252_88 ={ {4{neg252[5]}} , neg252[5:0] };

   // m252_89 = W*in
   wire signed [9:0] m252_89;
   assign m252_89 =10'b0;

   // m252_90 = W*in
   wire signed [9:0] m252_90;
   assign m252_90 =10'b0;

   // m252_91 = W*in
   wire signed [9:0] m252_91;
   assign m252_91 =10'b0;

   // m252_92 = W*in
   wire signed [9:0] m252_92;
   assign m252_92 =10'b0;

   // m252_93 = W*in
   wire signed [9:0] m252_93;
   assign m252_93 =10'b0;

   // m252_94 = W*in
   wire signed [9:0] m252_94;
   assign m252_94 =10'b0;

   // m252_95 = W*in
   wire signed [9:0] m252_95;
   assign m252_95 =10'b0;

   // m252_96 = W*in
   wire signed [9:0] m252_96;
   assign m252_96 =10'b0;

   // m252_97 = W*in
   wire signed [9:0] m252_97;
   assign m252_97 =10'b0;

   // m252_98 = W*in
   wire signed [9:0] m252_98;
   assign m252_98 =10'b0;

   // m252_99 = W*in
   wire signed [9:0] m252_99;
   assign m252_99 =10'b0;

   // m252_100 = W*in
   wire signed [9:0] m252_100;
   assign m252_100 =10'b0;

   // m252_101 = W*in
   wire signed [9:0] m252_101;
   assign m252_101 =10'b0;

   // m252_102 = W*in
   wire signed [9:0] m252_102;
   assign m252_102 =10'b0;

   // m252_103 = W*in
   wire signed [9:0] m252_103;
   assign m252_103 =10'b0;

   // m252_104 = W*in
   wire signed [9:0] m252_104;
   assign m252_104 =10'b0;

   // m252_105 = W*in
   wire signed [9:0] m252_105;
   assign m252_105 =10'b0;

   // m252_106 = W*in
   wire signed [9:0] m252_106;
   assign m252_106 =10'b0;

   // m252_107 = W*in
   wire signed [9:0] m252_107;
   assign m252_107 =10'b0;

   // m252_108 = W*in
   wire signed [9:0] m252_108;
   assign m252_108 =10'b0;

   // m252_109 = W*in
   wire signed [9:0] m252_109;
   assign m252_109 =10'b0;

   // m252_110 = W*in
   wire signed [9:0] m252_110;
   assign m252_110 =10'b0;

   // m252_111 = W*in
   wire signed [9:0] m252_111;
   assign m252_111 =10'b0;

   // m252_112 = W*in
   wire signed [9:0] m252_112;
   assign m252_112 =10'b0;

   // m252_113 = W*in
   wire signed [9:0] m252_113;
   assign m252_113 =10'b0;

   // m252_114 = W*in
   wire signed [9:0] m252_114;
   assign m252_114 ={ {5{neg252[5]}} , neg252[5:1] };

   // m252_115 = W*in
   wire signed [9:0] m252_115;
   assign m252_115 =10'b0;

   // m252_116 = W*in
   wire signed [9:0] m252_116;
   assign m252_116 =10'b0;

   // m252_117 = W*in
   wire signed [9:0] m252_117;
   assign m252_117 ={ {4{in252[5]}} , in252[5:0] };

   // m253_1 = W*in
   wire signed [9:0] m253_1;
   assign m253_1 =10'b0;

   // m253_2 = W*in
   wire signed [9:0] m253_2;
   assign m253_2 =10'b0;

   // m253_3 = W*in
   wire signed [9:0] m253_3;
   assign m253_3 =10'b0;

   // m253_4 = W*in
   wire signed [9:0] m253_4;
   assign m253_4 =10'b0;

   // m253_5 = W*in
   wire signed [9:0] m253_5;
   assign m253_5 =10'b0;

   // m253_6 = W*in
   wire signed [9:0] m253_6;
   assign m253_6 =10'b0;

   // m253_7 = W*in
   wire signed [9:0] m253_7;
   assign m253_7 =10'b0;

   // m253_8 = W*in
   wire signed [9:0] m253_8;
   assign m253_8 =10'b0;

   // m253_9 = W*in
   wire signed [9:0] m253_9;
   assign m253_9 =10'b0;

   // m253_10 = W*in
   wire signed [9:0] m253_10;
   assign m253_10 =10'b0;

   // m253_11 = W*in
   wire signed [9:0] m253_11;
   assign m253_11 =10'b0;

   // m253_12 = W*in
   wire signed [9:0] m253_12;
   assign m253_12 =10'b0;

   // m253_13 = W*in
   wire signed [9:0] m253_13;
   assign m253_13 =10'b0;

   // m253_14 = W*in
   wire signed [9:0] m253_14;
   assign m253_14 =10'b0;

   // m253_15 = W*in
   wire signed [9:0] m253_15;
   assign m253_15 =10'b0;

   // m253_16 = W*in
   wire signed [9:0] m253_16;
   assign m253_16 =10'b0;

   // m253_17 = W*in
   wire signed [9:0] m253_17;
   assign m253_17 ={ {5{in253[5]}} , in253[5:1] };

   // m253_18 = W*in
   wire signed [9:0] m253_18;
   assign m253_18 ={ {5{in253[5]}} , in253[5:1] };

   // m253_19 = W*in
   wire signed [9:0] m253_19;
   assign m253_19 =10'b0;

   // m253_20 = W*in
   wire signed [9:0] m253_20;
   assign m253_20 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_21 = W*in
   wire signed [9:0] m253_21;
   assign m253_21 ={ {4{neg253[5]}} , neg253[5:0] };

   // m253_22 = W*in
   wire signed [9:0] m253_22;
   assign m253_22 =10'b0;

   // m253_23 = W*in
   wire signed [9:0] m253_23;
   assign m253_23 =10'b0;

   // m253_24 = W*in
   wire signed [9:0] m253_24;
   assign m253_24 =10'b0;

   // m253_25 = W*in
   wire signed [9:0] m253_25;
   assign m253_25 ={ {5{in253[5]}} , in253[5:1] };

   // m253_26 = W*in
   wire signed [9:0] m253_26;
   assign m253_26 =10'b0;

   // m253_27 = W*in
   wire signed [9:0] m253_27;
   assign m253_27 ={ {5{in253[5]}} , in253[5:1] };

   // m253_28 = W*in
   wire signed [9:0] m253_28;
   assign m253_28 ={ {4{in253[5]}} , in253[5:0] };

   // m253_29 = W*in
   wire signed [9:0] m253_29;
   assign m253_29 =10'b0;

   // m253_30 = W*in
   wire signed [9:0] m253_30;
   assign m253_30 =10'b0;

   // m253_31 = W*in
   wire signed [9:0] m253_31;
   assign m253_31 =10'b0;

   // m253_32 = W*in
   wire signed [9:0] m253_32;
   assign m253_32 =10'b0;

   // m253_33 = W*in
   wire signed [9:0] m253_33;
   assign m253_33 =10'b0;

   // m253_34 = W*in
   wire signed [9:0] m253_34;
   assign m253_34 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_35 = W*in
   wire signed [9:0] m253_35;
   assign m253_35 =10'b0;

   // m253_36 = W*in
   wire signed [9:0] m253_36;
   assign m253_36 ={ {5{in253[5]}} , in253[5:1] };

   // m253_37 = W*in
   wire signed [9:0] m253_37;
   assign m253_37 =10'b0;

   // m253_38 = W*in
   wire signed [9:0] m253_38;
   assign m253_38 =10'b0;

   // m253_39 = W*in
   wire signed [9:0] m253_39;
   assign m253_39 =10'b0;

   // m253_40 = W*in
   wire signed [9:0] m253_40;
   assign m253_40 =10'b0;

   // m253_41 = W*in
   wire signed [9:0] m253_41;
   assign m253_41 =10'b0;

   // m253_42 = W*in
   wire signed [9:0] m253_42;
   assign m253_42 =10'b0;

   // m253_43 = W*in
   wire signed [9:0] m253_43;
   assign m253_43 =10'b0;

   // m253_44 = W*in
   wire signed [9:0] m253_44;
   assign m253_44 =10'b0;

   // m253_45 = W*in
   wire signed [9:0] m253_45;
   assign m253_45 =10'b0;

   // m253_46 = W*in
   wire signed [9:0] m253_46;
   assign m253_46 =10'b0;

   // m253_47 = W*in
   wire signed [9:0] m253_47;
   assign m253_47 =10'b0;

   // m253_48 = W*in
   wire signed [9:0] m253_48;
   assign m253_48 =10'b0;

   // m253_49 = W*in
   wire signed [9:0] m253_49;
   assign m253_49 =10'b0;

   // m253_50 = W*in
   wire signed [9:0] m253_50;
   assign m253_50 =10'b0;

   // m253_51 = W*in
   wire signed [9:0] m253_51;
   assign m253_51 =10'b0;

   // m253_52 = W*in
   wire signed [9:0] m253_52;
   assign m253_52 =10'b0;

   // m253_53 = W*in
   wire signed [9:0] m253_53;
   assign m253_53 =10'b0;

   // m253_54 = W*in
   wire signed [9:0] m253_54;
   assign m253_54 =10'b0;

   // m253_55 = W*in
   wire signed [9:0] m253_55;
   assign m253_55 =10'b0;

   // m253_56 = W*in
   wire signed [9:0] m253_56;
   assign m253_56 =10'b0;

   // m253_57 = W*in
   wire signed [9:0] m253_57;
   assign m253_57 =10'b0;

   // m253_58 = W*in
   wire signed [9:0] m253_58;
   assign m253_58 =10'b0;

   // m253_59 = W*in
   wire signed [9:0] m253_59;
   assign m253_59 =10'b0;

   // m253_60 = W*in
   wire signed [9:0] m253_60;
   assign m253_60 =10'b0;

   // m253_61 = W*in
   wire signed [9:0] m253_61;
   assign m253_61 =10'b0;

   // m253_62 = W*in
   wire signed [9:0] m253_62;
   assign m253_62 =10'b0;

   // m253_63 = W*in
   wire signed [9:0] m253_63;
   assign m253_63 =10'b0;

   // m253_64 = W*in
   wire signed [9:0] m253_64;
   assign m253_64 =10'b0;

   // m253_65 = W*in
   wire signed [9:0] m253_65;
   assign m253_65 =10'b0;

   // m253_66 = W*in
   wire signed [9:0] m253_66;
   assign m253_66 ={ {5{in253[5]}} , in253[5:1] };

   // m253_67 = W*in
   wire signed [9:0] m253_67;
   assign m253_67 ={ {4{neg253[5]}} , neg253[5:0] };

   // m253_68 = W*in
   wire signed [9:0] m253_68;
   assign m253_68 =10'b0;

   // m253_69 = W*in
   wire signed [9:0] m253_69;
   assign m253_69 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_70 = W*in
   wire signed [9:0] m253_70;
   assign m253_70 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_71 = W*in
   wire signed [9:0] m253_71;
   assign m253_71 ={ {5{in253[5]}} , in253[5:1] };

   // m253_72 = W*in
   wire signed [9:0] m253_72;
   assign m253_72 =10'b0;

   // m253_73 = W*in
   wire signed [9:0] m253_73;
   assign m253_73 ={ {5{in253[5]}} , in253[5:1] };

   // m253_74 = W*in
   wire signed [9:0] m253_74;
   assign m253_74 =10'b0;

   // m253_75 = W*in
   wire signed [9:0] m253_75;
   assign m253_75 =10'b0;

   // m253_76 = W*in
   wire signed [9:0] m253_76;
   assign m253_76 =10'b0;

   // m253_77 = W*in
   wire signed [9:0] m253_77;
   assign m253_77 ={ {4{in253[5]}} , in253[5:0] };

   // m253_78 = W*in
   wire signed [9:0] m253_78;
   assign m253_78 =10'b0;

   // m253_79 = W*in
   wire signed [9:0] m253_79;
   assign m253_79 =10'b0;

   // m253_80 = W*in
   wire signed [9:0] m253_80;
   assign m253_80 =10'b0;

   // m253_81 = W*in
   wire signed [9:0] m253_81;
   assign m253_81 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_82 = W*in
   wire signed [9:0] m253_82;
   assign m253_82 ={ {4{neg253[5]}} , neg253[5:0] };

   // m253_83 = W*in
   wire signed [9:0] m253_83;
   assign m253_83 =10'b0;

   // m253_84 = W*in
   wire signed [9:0] m253_84;
   assign m253_84 =10'b0;

   // m253_85 = W*in
   wire signed [9:0] m253_85;
   assign m253_85 =10'b0;

   // m253_86 = W*in
   wire signed [9:0] m253_86;
   assign m253_86 =10'b0;

   // m253_87 = W*in
   wire signed [9:0] m253_87;
   assign m253_87 =10'b0;

   // m253_88 = W*in
   wire signed [9:0] m253_88;
   assign m253_88 ={ {4{neg253[5]}} , neg253[5:0] };

   // m253_89 = W*in
   wire signed [9:0] m253_89;
   assign m253_89 =10'b0;

   // m253_90 = W*in
   wire signed [9:0] m253_90;
   assign m253_90 =10'b0;

   // m253_91 = W*in
   wire signed [9:0] m253_91;
   assign m253_91 =10'b0;

   // m253_92 = W*in
   wire signed [9:0] m253_92;
   assign m253_92 =10'b0;

   // m253_93 = W*in
   wire signed [9:0] m253_93;
   assign m253_93 =10'b0;

   // m253_94 = W*in
   wire signed [9:0] m253_94;
   assign m253_94 =10'b0;

   // m253_95 = W*in
   wire signed [9:0] m253_95;
   assign m253_95 =10'b0;

   // m253_96 = W*in
   wire signed [9:0] m253_96;
   assign m253_96 =10'b0;

   // m253_97 = W*in
   wire signed [9:0] m253_97;
   assign m253_97 =10'b0;

   // m253_98 = W*in
   wire signed [9:0] m253_98;
   assign m253_98 =10'b0;

   // m253_99 = W*in
   wire signed [9:0] m253_99;
   assign m253_99 =10'b0;

   // m253_100 = W*in
   wire signed [9:0] m253_100;
   assign m253_100 =10'b0;

   // m253_101 = W*in
   wire signed [9:0] m253_101;
   assign m253_101 =10'b0;

   // m253_102 = W*in
   wire signed [9:0] m253_102;
   assign m253_102 =10'b0;

   // m253_103 = W*in
   wire signed [9:0] m253_103;
   assign m253_103 =10'b0;

   // m253_104 = W*in
   wire signed [9:0] m253_104;
   assign m253_104 =10'b0;

   // m253_105 = W*in
   wire signed [9:0] m253_105;
   assign m253_105 =10'b0;

   // m253_106 = W*in
   wire signed [9:0] m253_106;
   assign m253_106 =10'b0;

   // m253_107 = W*in
   wire signed [9:0] m253_107;
   assign m253_107 =10'b0;

   // m253_108 = W*in
   wire signed [9:0] m253_108;
   assign m253_108 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_109 = W*in
   wire signed [9:0] m253_109;
   assign m253_109 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_110 = W*in
   wire signed [9:0] m253_110;
   assign m253_110 =10'b0;

   // m253_111 = W*in
   wire signed [9:0] m253_111;
   assign m253_111 =10'b0;

   // m253_112 = W*in
   wire signed [9:0] m253_112;
   assign m253_112 =10'b0;

   // m253_113 = W*in
   wire signed [9:0] m253_113;
   assign m253_113 =10'b0;

   // m253_114 = W*in
   wire signed [9:0] m253_114;
   assign m253_114 ={ {5{neg253[5]}} , neg253[5:1] };

   // m253_115 = W*in
   wire signed [9:0] m253_115;
   assign m253_115 =10'b0;

   // m253_116 = W*in
   wire signed [9:0] m253_116;
   assign m253_116 =10'b0;

   // m253_117 = W*in
   wire signed [9:0] m253_117;
   assign m253_117 =10'b0;

   // m254_1 = W*in
   wire signed [9:0] m254_1;
   assign m254_1 =10'b0;

   // m254_2 = W*in
   wire signed [9:0] m254_2;
   assign m254_2 =10'b0;

   // m254_3 = W*in
   wire signed [9:0] m254_3;
   assign m254_3 =10'b0;

   // m254_4 = W*in
   wire signed [9:0] m254_4;
   assign m254_4 =10'b0;

   // m254_5 = W*in
   wire signed [9:0] m254_5;
   assign m254_5 =10'b0;

   // m254_6 = W*in
   wire signed [9:0] m254_6;
   assign m254_6 =10'b0;

   // m254_7 = W*in
   wire signed [9:0] m254_7;
   assign m254_7 =10'b0;

   // m254_8 = W*in
   wire signed [9:0] m254_8;
   assign m254_8 =10'b0;

   // m254_9 = W*in
   wire signed [9:0] m254_9;
   assign m254_9 =10'b0;

   // m254_10 = W*in
   wire signed [9:0] m254_10;
   assign m254_10 =10'b0;

   // m254_11 = W*in
   wire signed [9:0] m254_11;
   assign m254_11 =10'b0;

   // m254_12 = W*in
   wire signed [9:0] m254_12;
   assign m254_12 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_13 = W*in
   wire signed [9:0] m254_13;
   assign m254_13 =10'b0;

   // m254_14 = W*in
   wire signed [9:0] m254_14;
   assign m254_14 =10'b0;

   // m254_15 = W*in
   wire signed [9:0] m254_15;
   assign m254_15 =10'b0;

   // m254_16 = W*in
   wire signed [9:0] m254_16;
   assign m254_16 =10'b0;

   // m254_17 = W*in
   wire signed [9:0] m254_17;
   assign m254_17 =10'b0;

   // m254_18 = W*in
   wire signed [9:0] m254_18;
   assign m254_18 =10'b0;

   // m254_19 = W*in
   wire signed [9:0] m254_19;
   assign m254_19 =10'b0;

   // m254_20 = W*in
   wire signed [9:0] m254_20;
   assign m254_20 ={ {5{in254[5]}} , in254[5:1] };

   // m254_21 = W*in
   wire signed [9:0] m254_21;
   assign m254_21 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_22 = W*in
   wire signed [9:0] m254_22;
   assign m254_22 =10'b0;

   // m254_23 = W*in
   wire signed [9:0] m254_23;
   assign m254_23 =10'b0;

   // m254_24 = W*in
   wire signed [9:0] m254_24;
   assign m254_24 =10'b0;

   // m254_25 = W*in
   wire signed [9:0] m254_25;
   assign m254_25 =10'b0;

   // m254_26 = W*in
   wire signed [9:0] m254_26;
   assign m254_26 =10'b0;

   // m254_27 = W*in
   wire signed [9:0] m254_27;
   assign m254_27 =10'b0;

   // m254_28 = W*in
   wire signed [9:0] m254_28;
   assign m254_28 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_29 = W*in
   wire signed [9:0] m254_29;
   assign m254_29 =10'b0;

   // m254_30 = W*in
   wire signed [9:0] m254_30;
   assign m254_30 =10'b0;

   // m254_31 = W*in
   wire signed [9:0] m254_31;
   assign m254_31 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_32 = W*in
   wire signed [9:0] m254_32;
   assign m254_32 =10'b0;

   // m254_33 = W*in
   wire signed [9:0] m254_33;
   assign m254_33 =10'b0;

   // m254_34 = W*in
   wire signed [9:0] m254_34;
   assign m254_34 =10'b0;

   // m254_35 = W*in
   wire signed [9:0] m254_35;
   assign m254_35 =10'b0;

   // m254_36 = W*in
   wire signed [9:0] m254_36;
   assign m254_36 =10'b0;

   // m254_37 = W*in
   wire signed [9:0] m254_37;
   assign m254_37 =10'b0;

   // m254_38 = W*in
   wire signed [9:0] m254_38;
   assign m254_38 =10'b0;

   // m254_39 = W*in
   wire signed [9:0] m254_39;
   assign m254_39 =10'b0;

   // m254_40 = W*in
   wire signed [9:0] m254_40;
   assign m254_40 =10'b0;

   // m254_41 = W*in
   wire signed [9:0] m254_41;
   assign m254_41 =10'b0;

   // m254_42 = W*in
   wire signed [9:0] m254_42;
   assign m254_42 =10'b0;

   // m254_43 = W*in
   wire signed [9:0] m254_43;
   assign m254_43 =10'b0;

   // m254_44 = W*in
   wire signed [9:0] m254_44;
   assign m254_44 =10'b0;

   // m254_45 = W*in
   wire signed [9:0] m254_45;
   assign m254_45 ={ {4{in254[5]}} , in254[5:0] };

   // m254_46 = W*in
   wire signed [9:0] m254_46;
   assign m254_46 =10'b0;

   // m254_47 = W*in
   wire signed [9:0] m254_47;
   assign m254_47 ={ {4{in254[5]}} , in254[5:0] };

   // m254_48 = W*in
   wire signed [9:0] m254_48;
   assign m254_48 =10'b0;

   // m254_49 = W*in
   wire signed [9:0] m254_49;
   assign m254_49 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_50 = W*in
   wire signed [9:0] m254_50;
   assign m254_50 =10'b0;

   // m254_51 = W*in
   wire signed [9:0] m254_51;
   assign m254_51 ={ {4{in254[5]}} , in254[5:0] };

   // m254_52 = W*in
   wire signed [9:0] m254_52;
   assign m254_52 =10'b0;

   // m254_53 = W*in
   wire signed [9:0] m254_53;
   assign m254_53 =10'b0;

   // m254_54 = W*in
   wire signed [9:0] m254_54;
   assign m254_54 =10'b0;

   // m254_55 = W*in
   wire signed [9:0] m254_55;
   assign m254_55 =10'b0;

   // m254_56 = W*in
   wire signed [9:0] m254_56;
   assign m254_56 =10'b0;

   // m254_57 = W*in
   wire signed [9:0] m254_57;
   assign m254_57 =10'b0;

   // m254_58 = W*in
   wire signed [9:0] m254_58;
   assign m254_58 =10'b0;

   // m254_59 = W*in
   wire signed [9:0] m254_59;
   assign m254_59 =10'b0;

   // m254_60 = W*in
   wire signed [9:0] m254_60;
   assign m254_60 =10'b0;

   // m254_61 = W*in
   wire signed [9:0] m254_61;
   assign m254_61 =10'b0;

   // m254_62 = W*in
   wire signed [9:0] m254_62;
   assign m254_62 =10'b0;

   // m254_63 = W*in
   wire signed [9:0] m254_63;
   assign m254_63 =10'b0;

   // m254_64 = W*in
   wire signed [9:0] m254_64;
   assign m254_64 ={ {5{in254[5]}} , in254[5:1] };

   // m254_65 = W*in
   wire signed [9:0] m254_65;
   assign m254_65 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_66 = W*in
   wire signed [9:0] m254_66;
   assign m254_66 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_67 = W*in
   wire signed [9:0] m254_67;
   assign m254_67 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_68 = W*in
   wire signed [9:0] m254_68;
   assign m254_68 =10'b0;

   // m254_69 = W*in
   wire signed [9:0] m254_69;
   assign m254_69 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_70 = W*in
   wire signed [9:0] m254_70;
   assign m254_70 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_71 = W*in
   wire signed [9:0] m254_71;
   assign m254_71 =10'b0;

   // m254_72 = W*in
   wire signed [9:0] m254_72;
   assign m254_72 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_73 = W*in
   wire signed [9:0] m254_73;
   assign m254_73 =10'b0;

   // m254_74 = W*in
   wire signed [9:0] m254_74;
   assign m254_74 =10'b0;

   // m254_75 = W*in
   wire signed [9:0] m254_75;
   assign m254_75 =10'b0;

   // m254_76 = W*in
   wire signed [9:0] m254_76;
   assign m254_76 =10'b0;

   // m254_77 = W*in
   wire signed [9:0] m254_77;
   assign m254_77 =10'b0;

   // m254_78 = W*in
   wire signed [9:0] m254_78;
   assign m254_78 =10'b0;

   // m254_79 = W*in
   wire signed [9:0] m254_79;
   assign m254_79 =10'b0;

   // m254_80 = W*in
   wire signed [9:0] m254_80;
   assign m254_80 =10'b0;

   // m254_81 = W*in
   wire signed [9:0] m254_81;
   assign m254_81 ={ {5{in254[5]}} , in254[5:1] };

   // m254_82 = W*in
   wire signed [9:0] m254_82;
   assign m254_82 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_83 = W*in
   wire signed [9:0] m254_83;
   assign m254_83 ={ {5{in254[5]}} , in254[5:1] };

   // m254_84 = W*in
   wire signed [9:0] m254_84;
   assign m254_84 =10'b0;

   // m254_85 = W*in
   wire signed [9:0] m254_85;
   assign m254_85 =10'b0;

   // m254_86 = W*in
   wire signed [9:0] m254_86;
   assign m254_86 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_87 = W*in
   wire signed [9:0] m254_87;
   assign m254_87 =10'b0;

   // m254_88 = W*in
   wire signed [9:0] m254_88;
   assign m254_88 =10'b0;

   // m254_89 = W*in
   wire signed [9:0] m254_89;
   assign m254_89 =10'b0;

   // m254_90 = W*in
   wire signed [9:0] m254_90;
   assign m254_90 =10'b0;

   // m254_91 = W*in
   wire signed [9:0] m254_91;
   assign m254_91 =10'b0;

   // m254_92 = W*in
   wire signed [9:0] m254_92;
   assign m254_92 =10'b0;

   // m254_93 = W*in
   wire signed [9:0] m254_93;
   assign m254_93 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_94 = W*in
   wire signed [9:0] m254_94;
   assign m254_94 =10'b0;

   // m254_95 = W*in
   wire signed [9:0] m254_95;
   assign m254_95 =10'b0;

   // m254_96 = W*in
   wire signed [9:0] m254_96;
   assign m254_96 =10'b0;

   // m254_97 = W*in
   wire signed [9:0] m254_97;
   assign m254_97 =10'b0;

   // m254_98 = W*in
   wire signed [9:0] m254_98;
   assign m254_98 =10'b0;

   // m254_99 = W*in
   wire signed [9:0] m254_99;
   assign m254_99 =10'b0;

   // m254_100 = W*in
   wire signed [9:0] m254_100;
   assign m254_100 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_101 = W*in
   wire signed [9:0] m254_101;
   assign m254_101 =10'b0;

   // m254_102 = W*in
   wire signed [9:0] m254_102;
   assign m254_102 =10'b0;

   // m254_103 = W*in
   wire signed [9:0] m254_103;
   assign m254_103 =10'b0;

   // m254_104 = W*in
   wire signed [9:0] m254_104;
   assign m254_104 ={ {4{neg254[5]}} , neg254[5:0] };

   // m254_105 = W*in
   wire signed [9:0] m254_105;
   assign m254_105 =10'b0;

   // m254_106 = W*in
   wire signed [9:0] m254_106;
   assign m254_106 =10'b0;

   // m254_107 = W*in
   wire signed [9:0] m254_107;
   assign m254_107 =10'b0;

   // m254_108 = W*in
   wire signed [9:0] m254_108;
   assign m254_108 ={ {5{neg254[5]}} , neg254[5:1] };

   // m254_109 = W*in
   wire signed [9:0] m254_109;
   assign m254_109 =10'b0;

   // m254_110 = W*in
   wire signed [9:0] m254_110;
   assign m254_110 =10'b0;

   // m254_111 = W*in
   wire signed [9:0] m254_111;
   assign m254_111 =10'b0;

   // m254_112 = W*in
   wire signed [9:0] m254_112;
   assign m254_112 =10'b0;

   // m254_113 = W*in
   wire signed [9:0] m254_113;
   assign m254_113 =10'b0;

   // m254_114 = W*in
   wire signed [9:0] m254_114;
   assign m254_114 =10'b0;

   // m254_115 = W*in
   wire signed [9:0] m254_115;
   assign m254_115 ={ {5{in254[5]}} , in254[5:1] };

   // m254_116 = W*in
   wire signed [9:0] m254_116;
   assign m254_116 =10'b0;

   // m254_117 = W*in
   wire signed [9:0] m254_117;
   assign m254_117 =10'b0;

   // m255_1 = W*in
   wire signed [9:0] m255_1;
   assign m255_1 =10'b0;

   // m255_2 = W*in
   wire signed [9:0] m255_2;
   assign m255_2 =10'b0;

   // m255_3 = W*in
   wire signed [9:0] m255_3;
   assign m255_3 =10'b0;

   // m255_4 = W*in
   wire signed [9:0] m255_4;
   assign m255_4 =10'b0;

   // m255_5 = W*in
   wire signed [9:0] m255_5;
   assign m255_5 =10'b0;

   // m255_6 = W*in
   wire signed [9:0] m255_6;
   assign m255_6 =10'b0;

   // m255_7 = W*in
   wire signed [9:0] m255_7;
   assign m255_7 =10'b0;

   // m255_8 = W*in
   wire signed [9:0] m255_8;
   assign m255_8 =10'b0;

   // m255_9 = W*in
   wire signed [9:0] m255_9;
   assign m255_9 =10'b0;

   // m255_10 = W*in
   wire signed [9:0] m255_10;
   assign m255_10 =10'b0;

   // m255_11 = W*in
   wire signed [9:0] m255_11;
   assign m255_11 =10'b0;

   // m255_12 = W*in
   wire signed [9:0] m255_12;
   assign m255_12 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_13 = W*in
   wire signed [9:0] m255_13;
   assign m255_13 =10'b0;

   // m255_14 = W*in
   wire signed [9:0] m255_14;
   assign m255_14 =10'b0;

   // m255_15 = W*in
   wire signed [9:0] m255_15;
   assign m255_15 =10'b0;

   // m255_16 = W*in
   wire signed [9:0] m255_16;
   assign m255_16 =10'b0;

   // m255_17 = W*in
   wire signed [9:0] m255_17;
   assign m255_17 =10'b0;

   // m255_18 = W*in
   wire signed [9:0] m255_18;
   assign m255_18 =10'b0;

   // m255_19 = W*in
   wire signed [9:0] m255_19;
   assign m255_19 =10'b0;

   // m255_20 = W*in
   wire signed [9:0] m255_20;
   assign m255_20 =10'b0;

   // m255_21 = W*in
   wire signed [9:0] m255_21;
   assign m255_21 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_22 = W*in
   wire signed [9:0] m255_22;
   assign m255_22 =10'b0;

   // m255_23 = W*in
   wire signed [9:0] m255_23;
   assign m255_23 =10'b0;

   // m255_24 = W*in
   wire signed [9:0] m255_24;
   assign m255_24 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_25 = W*in
   wire signed [9:0] m255_25;
   assign m255_25 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_26 = W*in
   wire signed [9:0] m255_26;
   assign m255_26 =10'b0;

   // m255_27 = W*in
   wire signed [9:0] m255_27;
   assign m255_27 =10'b0;

   // m255_28 = W*in
   wire signed [9:0] m255_28;
   assign m255_28 =10'b0;

   // m255_29 = W*in
   wire signed [9:0] m255_29;
   assign m255_29 =10'b0;

   // m255_30 = W*in
   wire signed [9:0] m255_30;
   assign m255_30 =10'b0;

   // m255_31 = W*in
   wire signed [9:0] m255_31;
   assign m255_31 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_32 = W*in
   wire signed [9:0] m255_32;
   assign m255_32 =10'b0;

   // m255_33 = W*in
   wire signed [9:0] m255_33;
   assign m255_33 =10'b0;

   // m255_34 = W*in
   wire signed [9:0] m255_34;
   assign m255_34 =10'b0;

   // m255_35 = W*in
   wire signed [9:0] m255_35;
   assign m255_35 =10'b0;

   // m255_36 = W*in
   wire signed [9:0] m255_36;
   assign m255_36 =10'b0;

   // m255_37 = W*in
   wire signed [9:0] m255_37;
   assign m255_37 =10'b0;

   // m255_38 = W*in
   wire signed [9:0] m255_38;
   assign m255_38 =10'b0;

   // m255_39 = W*in
   wire signed [9:0] m255_39;
   assign m255_39 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_40 = W*in
   wire signed [9:0] m255_40;
   assign m255_40 =10'b0;

   // m255_41 = W*in
   wire signed [9:0] m255_41;
   assign m255_41 =10'b0;

   // m255_42 = W*in
   wire signed [9:0] m255_42;
   assign m255_42 =10'b0;

   // m255_43 = W*in
   wire signed [9:0] m255_43;
   assign m255_43 =10'b0;

   // m255_44 = W*in
   wire signed [9:0] m255_44;
   assign m255_44 =10'b0;

   // m255_45 = W*in
   wire signed [9:0] m255_45;
   assign m255_45 =10'b0;

   // m255_46 = W*in
   wire signed [9:0] m255_46;
   assign m255_46 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_47 = W*in
   wire signed [9:0] m255_47;
   assign m255_47 =10'b0;

   // m255_48 = W*in
   wire signed [9:0] m255_48;
   assign m255_48 =10'b0;

   // m255_49 = W*in
   wire signed [9:0] m255_49;
   assign m255_49 =10'b0;

   // m255_50 = W*in
   wire signed [9:0] m255_50;
   assign m255_50 =10'b0;

   // m255_51 = W*in
   wire signed [9:0] m255_51;
   assign m255_51 ={ {4{in255[5]}} , in255[5:0] };

   // m255_52 = W*in
   wire signed [9:0] m255_52;
   assign m255_52 =10'b0;

   // m255_53 = W*in
   wire signed [9:0] m255_53;
   assign m255_53 =10'b0;

   // m255_54 = W*in
   wire signed [9:0] m255_54;
   assign m255_54 =10'b0;

   // m255_55 = W*in
   wire signed [9:0] m255_55;
   assign m255_55 =10'b0;

   // m255_56 = W*in
   wire signed [9:0] m255_56;
   assign m255_56 =10'b0;

   // m255_57 = W*in
   wire signed [9:0] m255_57;
   assign m255_57 =10'b0;

   // m255_58 = W*in
   wire signed [9:0] m255_58;
   assign m255_58 =10'b0;

   // m255_59 = W*in
   wire signed [9:0] m255_59;
   assign m255_59 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_60 = W*in
   wire signed [9:0] m255_60;
   assign m255_60 =10'b0;

   // m255_61 = W*in
   wire signed [9:0] m255_61;
   assign m255_61 =10'b0;

   // m255_62 = W*in
   wire signed [9:0] m255_62;
   assign m255_62 =10'b0;

   // m255_63 = W*in
   wire signed [9:0] m255_63;
   assign m255_63 =10'b0;

   // m255_64 = W*in
   wire signed [9:0] m255_64;
   assign m255_64 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_65 = W*in
   wire signed [9:0] m255_65;
   assign m255_65 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_66 = W*in
   wire signed [9:0] m255_66;
   assign m255_66 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_67 = W*in
   wire signed [9:0] m255_67;
   assign m255_67 =10'b0;

   // m255_68 = W*in
   wire signed [9:0] m255_68;
   assign m255_68 =10'b0;

   // m255_69 = W*in
   wire signed [9:0] m255_69;
   assign m255_69 =10'b0;

   // m255_70 = W*in
   wire signed [9:0] m255_70;
   assign m255_70 =10'b0;

   // m255_71 = W*in
   wire signed [9:0] m255_71;
   assign m255_71 =10'b0;

   // m255_72 = W*in
   wire signed [9:0] m255_72;
   assign m255_72 =10'b0;

   // m255_73 = W*in
   wire signed [9:0] m255_73;
   assign m255_73 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_74 = W*in
   wire signed [9:0] m255_74;
   assign m255_74 =10'b0;

   // m255_75 = W*in
   wire signed [9:0] m255_75;
   assign m255_75 =10'b0;

   // m255_76 = W*in
   wire signed [9:0] m255_76;
   assign m255_76 =10'b0;

   // m255_77 = W*in
   wire signed [9:0] m255_77;
   assign m255_77 =10'b0;

   // m255_78 = W*in
   wire signed [9:0] m255_78;
   assign m255_78 ={ {5{in255[5]}} , in255[5:1] };

   // m255_79 = W*in
   wire signed [9:0] m255_79;
   assign m255_79 =10'b0;

   // m255_80 = W*in
   wire signed [9:0] m255_80;
   assign m255_80 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_81 = W*in
   wire signed [9:0] m255_81;
   assign m255_81 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_82 = W*in
   wire signed [9:0] m255_82;
   assign m255_82 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_83 = W*in
   wire signed [9:0] m255_83;
   assign m255_83 ={ {5{in255[5]}} , in255[5:1] };

   // m255_84 = W*in
   wire signed [9:0] m255_84;
   assign m255_84 =10'b0;

   // m255_85 = W*in
   wire signed [9:0] m255_85;
   assign m255_85 =10'b0;

   // m255_86 = W*in
   wire signed [9:0] m255_86;
   assign m255_86 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_87 = W*in
   wire signed [9:0] m255_87;
   assign m255_87 =10'b0;

   // m255_88 = W*in
   wire signed [9:0] m255_88;
   assign m255_88 =10'b0;

   // m255_89 = W*in
   wire signed [9:0] m255_89;
   assign m255_89 =10'b0;

   // m255_90 = W*in
   wire signed [9:0] m255_90;
   assign m255_90 =10'b0;

   // m255_91 = W*in
   wire signed [9:0] m255_91;
   assign m255_91 ={ {4{neg255[5]}} , neg255[5:0] };

   // m255_92 = W*in
   wire signed [9:0] m255_92;
   assign m255_92 =10'b0;

   // m255_93 = W*in
   wire signed [9:0] m255_93;
   assign m255_93 =10'b0;

   // m255_94 = W*in
   wire signed [9:0] m255_94;
   assign m255_94 ={ {5{neg255[5]}} , neg255[5:1] };

   // m255_95 = W*in
   wire signed [9:0] m255_95;
   assign m255_95 =10'b0;

   // m255_96 = W*in
   wire signed [9:0] m255_96;
   assign m255_96 =10'b0;

   // m255_97 = W*in
   wire signed [9:0] m255_97;
   assign m255_97 =10'b0;

   // m255_98 = W*in
   wire signed [9:0] m255_98;
   assign m255_98 =10'b0;

   // m255_99 = W*in
   wire signed [9:0] m255_99;
   assign m255_99 =10'b0;

   // m255_100 = W*in
   wire signed [9:0] m255_100;
   assign m255_100 =10'b0;

   // m255_101 = W*in
   wire signed [9:0] m255_101;
   assign m255_101 =10'b0;

   // m255_102 = W*in
   wire signed [9:0] m255_102;
   assign m255_102 =10'b0;

   // m255_103 = W*in
   wire signed [9:0] m255_103;
   assign m255_103 =10'b0;

   // m255_104 = W*in
   wire signed [9:0] m255_104;
   assign m255_104 =10'b0;

   // m255_105 = W*in
   wire signed [9:0] m255_105;
   assign m255_105 =10'b0;

   // m255_106 = W*in
   wire signed [9:0] m255_106;
   assign m255_106 =10'b0;

   // m255_107 = W*in
   wire signed [9:0] m255_107;
   assign m255_107 =10'b0;

   // m255_108 = W*in
   wire signed [9:0] m255_108;
   assign m255_108 =10'b0;

   // m255_109 = W*in
   wire signed [9:0] m255_109;
   assign m255_109 =10'b0;

   // m255_110 = W*in
   wire signed [9:0] m255_110;
   assign m255_110 =10'b0;

   // m255_111 = W*in
   wire signed [9:0] m255_111;
   assign m255_111 =10'b0;

   // m255_112 = W*in
   wire signed [9:0] m255_112;
   assign m255_112 =10'b0;

   // m255_113 = W*in
   wire signed [9:0] m255_113;
   assign m255_113 =10'b0;

   // m255_114 = W*in
   wire signed [9:0] m255_114;
   assign m255_114 =10'b0;

   // m255_115 = W*in
   wire signed [9:0] m255_115;
   assign m255_115 =10'b0;

   // m255_116 = W*in
   wire signed [9:0] m255_116;
   assign m255_116 =10'b0;

   // m255_117 = W*in
   wire signed [9:0] m255_117;
   assign m255_117 ={ {4{neg255[5]}} , neg255[5:0] };

   // m256_1 = W*in
   wire signed [9:0] m256_1;
   assign m256_1 =10'b0;

   // m256_2 = W*in
   wire signed [9:0] m256_2;
   assign m256_2 =10'b0;

   // m256_3 = W*in
   wire signed [9:0] m256_3;
   assign m256_3 =10'b0;

   // m256_4 = W*in
   wire signed [9:0] m256_4;
   assign m256_4 =10'b0;

   // m256_5 = W*in
   wire signed [9:0] m256_5;
   assign m256_5 =10'b0;

   // m256_6 = W*in
   wire signed [9:0] m256_6;
   assign m256_6 =10'b0;

   // m256_7 = W*in
   wire signed [9:0] m256_7;
   assign m256_7 =10'b0;

   // m256_8 = W*in
   wire signed [9:0] m256_8;
   assign m256_8 =10'b0;

   // m256_9 = W*in
   wire signed [9:0] m256_9;
   assign m256_9 =10'b0;

   // m256_10 = W*in
   wire signed [9:0] m256_10;
   assign m256_10 =10'b0;

   // m256_11 = W*in
   wire signed [9:0] m256_11;
   assign m256_11 =10'b0;

   // m256_12 = W*in
   wire signed [9:0] m256_12;
   assign m256_12 =10'b0;

   // m256_13 = W*in
   wire signed [9:0] m256_13;
   assign m256_13 =10'b0;

   // m256_14 = W*in
   wire signed [9:0] m256_14;
   assign m256_14 =10'b0;

   // m256_15 = W*in
   wire signed [9:0] m256_15;
   assign m256_15 =10'b0;

   // m256_16 = W*in
   wire signed [9:0] m256_16;
   assign m256_16 =10'b0;

   // m256_17 = W*in
   wire signed [9:0] m256_17;
   assign m256_17 ={ {5{in256[5]}} , in256[5:1] };

   // m256_18 = W*in
   wire signed [9:0] m256_18;
   assign m256_18 ={ {4{neg256[5]}} , neg256[5:0] };

   // m256_19 = W*in
   wire signed [9:0] m256_19;
   assign m256_19 =10'b0;

   // m256_20 = W*in
   wire signed [9:0] m256_20;
   assign m256_20 =10'b0;

   // m256_21 = W*in
   wire signed [9:0] m256_21;
   assign m256_21 =10'b0;

   // m256_22 = W*in
   wire signed [9:0] m256_22;
   assign m256_22 =10'b0;

   // m256_23 = W*in
   wire signed [9:0] m256_23;
   assign m256_23 =10'b0;

   // m256_24 = W*in
   wire signed [9:0] m256_24;
   assign m256_24 =10'b0;

   // m256_25 = W*in
   wire signed [9:0] m256_25;
   assign m256_25 =10'b0;

   // m256_26 = W*in
   wire signed [9:0] m256_26;
   assign m256_26 =10'b0;

   // m256_27 = W*in
   wire signed [9:0] m256_27;
   assign m256_27 ={ {5{in256[5]}} , in256[5:1] };

   // m256_28 = W*in
   wire signed [9:0] m256_28;
   assign m256_28 =10'b0;

   // m256_29 = W*in
   wire signed [9:0] m256_29;
   assign m256_29 =10'b0;

   // m256_30 = W*in
   wire signed [9:0] m256_30;
   assign m256_30 =10'b0;

   // m256_31 = W*in
   wire signed [9:0] m256_31;
   assign m256_31 =10'b0;

   // m256_32 = W*in
   wire signed [9:0] m256_32;
   assign m256_32 =10'b0;

   // m256_33 = W*in
   wire signed [9:0] m256_33;
   assign m256_33 =10'b0;

   // m256_34 = W*in
   wire signed [9:0] m256_34;
   assign m256_34 ={ {5{in256[5]}} , in256[5:1] };

   // m256_35 = W*in
   wire signed [9:0] m256_35;
   assign m256_35 =10'b0;

   // m256_36 = W*in
   wire signed [9:0] m256_36;
   assign m256_36 ={ {5{neg256[5]}} , neg256[5:1] };

   // m256_37 = W*in
   wire signed [9:0] m256_37;
   assign m256_37 =10'b0;

   // m256_38 = W*in
   wire signed [9:0] m256_38;
   assign m256_38 =10'b0;

   // m256_39 = W*in
   wire signed [9:0] m256_39;
   assign m256_39 =10'b0;

   // m256_40 = W*in
   wire signed [9:0] m256_40;
   assign m256_40 =10'b0;

   // m256_41 = W*in
   wire signed [9:0] m256_41;
   assign m256_41 =10'b0;

   // m256_42 = W*in
   wire signed [9:0] m256_42;
   assign m256_42 ={ {4{neg256[5]}} , neg256[5:0] };

   // m256_43 = W*in
   wire signed [9:0] m256_43;
   assign m256_43 =10'b0;

   // m256_44 = W*in
   wire signed [9:0] m256_44;
   assign m256_44 =10'b0;

   // m256_45 = W*in
   wire signed [9:0] m256_45;
   assign m256_45 =10'b0;

   // m256_46 = W*in
   wire signed [9:0] m256_46;
   assign m256_46 =10'b0;

   // m256_47 = W*in
   wire signed [9:0] m256_47;
   assign m256_47 =10'b0;

   // m256_48 = W*in
   wire signed [9:0] m256_48;
   assign m256_48 =10'b0;

   // m256_49 = W*in
   wire signed [9:0] m256_49;
   assign m256_49 =10'b0;

   // m256_50 = W*in
   wire signed [9:0] m256_50;
   assign m256_50 =10'b0;

   // m256_51 = W*in
   wire signed [9:0] m256_51;
   assign m256_51 =10'b0;

   // m256_52 = W*in
   wire signed [9:0] m256_52;
   assign m256_52 =10'b0;

   // m256_53 = W*in
   wire signed [9:0] m256_53;
   assign m256_53 =10'b0;

   // m256_54 = W*in
   wire signed [9:0] m256_54;
   assign m256_54 ={ {4{in256[5]}} , in256[5:0] };

   // m256_55 = W*in
   wire signed [9:0] m256_55;
   assign m256_55 =10'b0;

   // m256_56 = W*in
   wire signed [9:0] m256_56;
   assign m256_56 =10'b0;

   // m256_57 = W*in
   wire signed [9:0] m256_57;
   assign m256_57 =10'b0;

   // m256_58 = W*in
   wire signed [9:0] m256_58;
   assign m256_58 =10'b0;

   // m256_59 = W*in
   wire signed [9:0] m256_59;
   assign m256_59 =10'b0;

   // m256_60 = W*in
   wire signed [9:0] m256_60;
   assign m256_60 =10'b0;

   // m256_61 = W*in
   wire signed [9:0] m256_61;
   assign m256_61 =10'b0;

   // m256_62 = W*in
   wire signed [9:0] m256_62;
   assign m256_62 =10'b0;

   // m256_63 = W*in
   wire signed [9:0] m256_63;
   assign m256_63 =10'b0;

   // m256_64 = W*in
   wire signed [9:0] m256_64;
   assign m256_64 =10'b0;

   // m256_65 = W*in
   wire signed [9:0] m256_65;
   assign m256_65 ={ {5{neg256[5]}} , neg256[5:1] };

   // m256_66 = W*in
   wire signed [9:0] m256_66;
   assign m256_66 ={ {5{neg256[5]}} , neg256[5:1] };

   // m256_67 = W*in
   wire signed [9:0] m256_67;
   assign m256_67 =10'b0;

   // m256_68 = W*in
   wire signed [9:0] m256_68;
   assign m256_68 =10'b0;

   // m256_69 = W*in
   wire signed [9:0] m256_69;
   assign m256_69 =10'b0;

   // m256_70 = W*in
   wire signed [9:0] m256_70;
   assign m256_70 =10'b0;

   // m256_71 = W*in
   wire signed [9:0] m256_71;
   assign m256_71 =10'b0;

   // m256_72 = W*in
   wire signed [9:0] m256_72;
   assign m256_72 =10'b0;

   // m256_73 = W*in
   wire signed [9:0] m256_73;
   assign m256_73 ={ {5{neg256[5]}} , neg256[5:1] };

   // m256_74 = W*in
   wire signed [9:0] m256_74;
   assign m256_74 =10'b0;

   // m256_75 = W*in
   wire signed [9:0] m256_75;
   assign m256_75 =10'b0;

   // m256_76 = W*in
   wire signed [9:0] m256_76;
   assign m256_76 =10'b0;

   // m256_77 = W*in
   wire signed [9:0] m256_77;
   assign m256_77 ={ {4{in256[5]}} , in256[5:0] };

   // m256_78 = W*in
   wire signed [9:0] m256_78;
   assign m256_78 =10'b0;

   // m256_79 = W*in
   wire signed [9:0] m256_79;
   assign m256_79 =10'b0;

   // m256_80 = W*in
   wire signed [9:0] m256_80;
   assign m256_80 =10'b0;

   // m256_81 = W*in
   wire signed [9:0] m256_81;
   assign m256_81 ={ {5{neg256[5]}} , neg256[5:1] };

   // m256_82 = W*in
   wire signed [9:0] m256_82;
   assign m256_82 =10'b0;

   // m256_83 = W*in
   wire signed [9:0] m256_83;
   assign m256_83 =10'b0;

   // m256_84 = W*in
   wire signed [9:0] m256_84;
   assign m256_84 =10'b0;

   // m256_85 = W*in
   wire signed [9:0] m256_85;
   assign m256_85 =10'b0;

   // m256_86 = W*in
   wire signed [9:0] m256_86;
   assign m256_86 =10'b0;

   // m256_87 = W*in
   wire signed [9:0] m256_87;
   assign m256_87 =10'b0;

   // m256_88 = W*in
   wire signed [9:0] m256_88;
   assign m256_88 =10'b0;

   // m256_89 = W*in
   wire signed [9:0] m256_89;
   assign m256_89 =10'b0;

   // m256_90 = W*in
   wire signed [9:0] m256_90;
   assign m256_90 ={ {4{in256[5]}} , in256[5:0] };

   // m256_91 = W*in
   wire signed [9:0] m256_91;
   assign m256_91 ={ {4{neg256[5]}} , neg256[5:0] };

   // m256_92 = W*in
   wire signed [9:0] m256_92;
   assign m256_92 =10'b0;

   // m256_93 = W*in
   wire signed [9:0] m256_93;
   assign m256_93 =10'b0;

   // m256_94 = W*in
   wire signed [9:0] m256_94;
   assign m256_94 =10'b0;

   // m256_95 = W*in
   wire signed [9:0] m256_95;
   assign m256_95 =10'b0;

   // m256_96 = W*in
   wire signed [9:0] m256_96;
   assign m256_96 =10'b0;

   // m256_97 = W*in
   wire signed [9:0] m256_97;
   assign m256_97 =10'b0;

   // m256_98 = W*in
   wire signed [9:0] m256_98;
   assign m256_98 =10'b0;

   // m256_99 = W*in
   wire signed [9:0] m256_99;
   assign m256_99 =10'b0;

   // m256_100 = W*in
   wire signed [9:0] m256_100;
   assign m256_100 =10'b0;

   // m256_101 = W*in
   wire signed [9:0] m256_101;
   assign m256_101 =10'b0;

   // m256_102 = W*in
   wire signed [9:0] m256_102;
   assign m256_102 =10'b0;

   // m256_103 = W*in
   wire signed [9:0] m256_103;
   assign m256_103 =10'b0;

   // m256_104 = W*in
   wire signed [9:0] m256_104;
   assign m256_104 =10'b0;

   // m256_105 = W*in
   wire signed [9:0] m256_105;
   assign m256_105 =10'b0;

   // m256_106 = W*in
   wire signed [9:0] m256_106;
   assign m256_106 =10'b0;

   // m256_107 = W*in
   wire signed [9:0] m256_107;
   assign m256_107 ={ {4{in256[5]}} , in256[5:0] };

   // m256_108 = W*in
   wire signed [9:0] m256_108;
   assign m256_108 =10'b0;

   // m256_109 = W*in
   wire signed [9:0] m256_109;
   assign m256_109 =10'b0;

   // m256_110 = W*in
   wire signed [9:0] m256_110;
   assign m256_110 =10'b0;

   // m256_111 = W*in
   wire signed [9:0] m256_111;
   assign m256_111 =10'b0;

   // m256_112 = W*in
   wire signed [9:0] m256_112;
   assign m256_112 =10'b0;

   // m256_113 = W*in
   wire signed [9:0] m256_113;
   assign m256_113 ={ {4{in256[5]}} , in256[5:0] };

   // m256_114 = W*in
   wire signed [9:0] m256_114;
   assign m256_114 =10'b0;

   // m256_115 = W*in
   wire signed [9:0] m256_115;
   assign m256_115 =10'b0;

   // m256_116 = W*in
   wire signed [9:0] m256_116;
   assign m256_116 =10'b0;

   // m256_117 = W*in
   wire signed [9:0] m256_117;
   assign m256_117 =10'b0;

   // m257_1 = W*in
   wire signed [9:0] m257_1;
   assign m257_1 =10'b0;

   // m257_2 = W*in
   wire signed [9:0] m257_2;
   assign m257_2 =10'b0;

   // m257_3 = W*in
   wire signed [9:0] m257_3;
   assign m257_3 ={ {4{in257[5]}} , in257[5:0] };

   // m257_4 = W*in
   wire signed [9:0] m257_4;
   assign m257_4 =10'b0;

   // m257_5 = W*in
   wire signed [9:0] m257_5;
   assign m257_5 =10'b0;

   // m257_6 = W*in
   wire signed [9:0] m257_6;
   assign m257_6 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_7 = W*in
   wire signed [9:0] m257_7;
   assign m257_7 =10'b0;

   // m257_8 = W*in
   wire signed [9:0] m257_8;
   assign m257_8 =10'b0;

   // m257_9 = W*in
   wire signed [9:0] m257_9;
   assign m257_9 =10'b0;

   // m257_10 = W*in
   wire signed [9:0] m257_10;
   assign m257_10 =10'b0;

   // m257_11 = W*in
   wire signed [9:0] m257_11;
   assign m257_11 =10'b0;

   // m257_12 = W*in
   wire signed [9:0] m257_12;
   assign m257_12 =10'b0;

   // m257_13 = W*in
   wire signed [9:0] m257_13;
   assign m257_13 =10'b0;

   // m257_14 = W*in
   wire signed [9:0] m257_14;
   assign m257_14 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_15 = W*in
   wire signed [9:0] m257_15;
   assign m257_15 =10'b0;

   // m257_16 = W*in
   wire signed [9:0] m257_16;
   assign m257_16 ={ {5{in257[5]}} , in257[5:1] };

   // m257_17 = W*in
   wire signed [9:0] m257_17;
   assign m257_17 ={ {4{in257[5]}} , in257[5:0] };

   // m257_18 = W*in
   wire signed [9:0] m257_18;
   assign m257_18 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_19 = W*in
   wire signed [9:0] m257_19;
   assign m257_19 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_20 = W*in
   wire signed [9:0] m257_20;
   assign m257_20 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_21 = W*in
   wire signed [9:0] m257_21;
   assign m257_21 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_22 = W*in
   wire signed [9:0] m257_22;
   assign m257_22 =10'b0;

   // m257_23 = W*in
   wire signed [9:0] m257_23;
   assign m257_23 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_24 = W*in
   wire signed [9:0] m257_24;
   assign m257_24 =10'b0;

   // m257_25 = W*in
   wire signed [9:0] m257_25;
   assign m257_25 =10'b0;

   // m257_26 = W*in
   wire signed [9:0] m257_26;
   assign m257_26 =10'b0;

   // m257_27 = W*in
   wire signed [9:0] m257_27;
   assign m257_27 ={ {4{in257[5]}} , in257[5:0] };

   // m257_28 = W*in
   wire signed [9:0] m257_28;
   assign m257_28 =10'b0;

   // m257_29 = W*in
   wire signed [9:0] m257_29;
   assign m257_29 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_30 = W*in
   wire signed [9:0] m257_30;
   assign m257_30 =10'b0;

   // m257_31 = W*in
   wire signed [9:0] m257_31;
   assign m257_31 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_32 = W*in
   wire signed [9:0] m257_32;
   assign m257_32 =10'b0;

   // m257_33 = W*in
   wire signed [9:0] m257_33;
   assign m257_33 =10'b0;

   // m257_34 = W*in
   wire signed [9:0] m257_34;
   assign m257_34 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_35 = W*in
   wire signed [9:0] m257_35;
   assign m257_35 =10'b0;

   // m257_36 = W*in
   wire signed [9:0] m257_36;
   assign m257_36 =10'b0;

   // m257_37 = W*in
   wire signed [9:0] m257_37;
   assign m257_37 =10'b0;

   // m257_38 = W*in
   wire signed [9:0] m257_38;
   assign m257_38 =10'b0;

   // m257_39 = W*in
   wire signed [9:0] m257_39;
   assign m257_39 =10'b0;

   // m257_40 = W*in
   wire signed [9:0] m257_40;
   assign m257_40 =10'b0;

   // m257_41 = W*in
   wire signed [9:0] m257_41;
   assign m257_41 =10'b0;

   // m257_42 = W*in
   wire signed [9:0] m257_42;
   assign m257_42 =10'b0;

   // m257_43 = W*in
   wire signed [9:0] m257_43;
   assign m257_43 =10'b0;

   // m257_44 = W*in
   wire signed [9:0] m257_44;
   assign m257_44 =10'b0;

   // m257_45 = W*in
   wire signed [9:0] m257_45;
   assign m257_45 ={ {4{in257[5]}} , in257[5:0] };

   // m257_46 = W*in
   wire signed [9:0] m257_46;
   assign m257_46 =10'b0;

   // m257_47 = W*in
   wire signed [9:0] m257_47;
   assign m257_47 =10'b0;

   // m257_48 = W*in
   wire signed [9:0] m257_48;
   assign m257_48 =10'b0;

   // m257_49 = W*in
   wire signed [9:0] m257_49;
   assign m257_49 =10'b0;

   // m257_50 = W*in
   wire signed [9:0] m257_50;
   assign m257_50 =10'b0;

   // m257_51 = W*in
   wire signed [9:0] m257_51;
   assign m257_51 ={ {4{in257[5]}} , in257[5:0] };

   // m257_52 = W*in
   wire signed [9:0] m257_52;
   assign m257_52 =10'b0;

   // m257_53 = W*in
   wire signed [9:0] m257_53;
   assign m257_53 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_54 = W*in
   wire signed [9:0] m257_54;
   assign m257_54 ={ {4{in257[5]}} , in257[5:0] };

   // m257_55 = W*in
   wire signed [9:0] m257_55;
   assign m257_55 =10'b0;

   // m257_56 = W*in
   wire signed [9:0] m257_56;
   assign m257_56 ={ {4{in257[5]}} , in257[5:0] };

   // m257_57 = W*in
   wire signed [9:0] m257_57;
   assign m257_57 =10'b0;

   // m257_58 = W*in
   wire signed [9:0] m257_58;
   assign m257_58 =10'b0;

   // m257_59 = W*in
   wire signed [9:0] m257_59;
   assign m257_59 ={ {4{in257[5]}} , in257[5:0] };

   // m257_60 = W*in
   wire signed [9:0] m257_60;
   assign m257_60 =10'b0;

   // m257_61 = W*in
   wire signed [9:0] m257_61;
   assign m257_61 ={ {5{in257[5]}} , in257[5:1] };

   // m257_62 = W*in
   wire signed [9:0] m257_62;
   assign m257_62 =10'b0;

   // m257_63 = W*in
   wire signed [9:0] m257_63;
   assign m257_63 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_64 = W*in
   wire signed [9:0] m257_64;
   assign m257_64 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_65 = W*in
   wire signed [9:0] m257_65;
   assign m257_65 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_66 = W*in
   wire signed [9:0] m257_66;
   assign m257_66 =10'b0;

   // m257_67 = W*in
   wire signed [9:0] m257_67;
   assign m257_67 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_68 = W*in
   wire signed [9:0] m257_68;
   assign m257_68 =10'b0;

   // m257_69 = W*in
   wire signed [9:0] m257_69;
   assign m257_69 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_70 = W*in
   wire signed [9:0] m257_70;
   assign m257_70 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_71 = W*in
   wire signed [9:0] m257_71;
   assign m257_71 =10'b0;

   // m257_72 = W*in
   wire signed [9:0] m257_72;
   assign m257_72 =10'b0;

   // m257_73 = W*in
   wire signed [9:0] m257_73;
   assign m257_73 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_74 = W*in
   wire signed [9:0] m257_74;
   assign m257_74 =10'b0;

   // m257_75 = W*in
   wire signed [9:0] m257_75;
   assign m257_75 =10'b0;

   // m257_76 = W*in
   wire signed [9:0] m257_76;
   assign m257_76 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_77 = W*in
   wire signed [9:0] m257_77;
   assign m257_77 ={ {4{in257[5]}} , in257[5:0] };

   // m257_78 = W*in
   wire signed [9:0] m257_78;
   assign m257_78 =10'b0;

   // m257_79 = W*in
   wire signed [9:0] m257_79;
   assign m257_79 =10'b0;

   // m257_80 = W*in
   wire signed [9:0] m257_80;
   assign m257_80 =10'b0;

   // m257_81 = W*in
   wire signed [9:0] m257_81;
   assign m257_81 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_82 = W*in
   wire signed [9:0] m257_82;
   assign m257_82 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_83 = W*in
   wire signed [9:0] m257_83;
   assign m257_83 ={ {4{in257[5]}} , in257[5:0] };

   // m257_84 = W*in
   wire signed [9:0] m257_84;
   assign m257_84 =10'b0;

   // m257_85 = W*in
   wire signed [9:0] m257_85;
   assign m257_85 =10'b0;

   // m257_86 = W*in
   wire signed [9:0] m257_86;
   assign m257_86 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_87 = W*in
   wire signed [9:0] m257_87;
   assign m257_87 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_88 = W*in
   wire signed [9:0] m257_88;
   assign m257_88 =10'b0;

   // m257_89 = W*in
   wire signed [9:0] m257_89;
   assign m257_89 =10'b0;

   // m257_90 = W*in
   wire signed [9:0] m257_90;
   assign m257_90 =10'b0;

   // m257_91 = W*in
   wire signed [9:0] m257_91;
   assign m257_91 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_92 = W*in
   wire signed [9:0] m257_92;
   assign m257_92 =10'b0;

   // m257_93 = W*in
   wire signed [9:0] m257_93;
   assign m257_93 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_94 = W*in
   wire signed [9:0] m257_94;
   assign m257_94 ={ {4{neg257[5]}} , neg257[5:0] };

   // m257_95 = W*in
   wire signed [9:0] m257_95;
   assign m257_95 ={ {4{in257[5]}} , in257[5:0] };

   // m257_96 = W*in
   wire signed [9:0] m257_96;
   assign m257_96 =10'b0;

   // m257_97 = W*in
   wire signed [9:0] m257_97;
   assign m257_97 =10'b0;

   // m257_98 = W*in
   wire signed [9:0] m257_98;
   assign m257_98 =10'b0;

   // m257_99 = W*in
   wire signed [9:0] m257_99;
   assign m257_99 ={ {3{neg257[5]}} , neg257 , {1{1'b0}} };

   // m257_100 = W*in
   wire signed [9:0] m257_100;
   assign m257_100 =10'b0;

   // m257_101 = W*in
   wire signed [9:0] m257_101;
   assign m257_101 =10'b0;

   // m257_102 = W*in
   wire signed [9:0] m257_102;
   assign m257_102 =10'b0;

   // m257_103 = W*in
   wire signed [9:0] m257_103;
   assign m257_103 ={ {4{in257[5]}} , in257[5:0] };

   // m257_104 = W*in
   wire signed [9:0] m257_104;
   assign m257_104 ={ {4{in257[5]}} , in257[5:0] };

   // m257_105 = W*in
   wire signed [9:0] m257_105;
   assign m257_105 =10'b0;

   // m257_106 = W*in
   wire signed [9:0] m257_106;
   assign m257_106 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_107 = W*in
   wire signed [9:0] m257_107;
   assign m257_107 ={ {4{in257[5]}} , in257[5:0] };

   // m257_108 = W*in
   wire signed [9:0] m257_108;
   assign m257_108 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_109 = W*in
   wire signed [9:0] m257_109;
   assign m257_109 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_110 = W*in
   wire signed [9:0] m257_110;
   assign m257_110 =10'b0;

   // m257_111 = W*in
   wire signed [9:0] m257_111;
   assign m257_111 =10'b0;

   // m257_112 = W*in
   wire signed [9:0] m257_112;
   assign m257_112 =10'b0;

   // m257_113 = W*in
   wire signed [9:0] m257_113;
   assign m257_113 =10'b0;

   // m257_114 = W*in
   wire signed [9:0] m257_114;
   assign m257_114 ={ {5{neg257[5]}} , neg257[5:1] };

   // m257_115 = W*in
   wire signed [9:0] m257_115;
   assign m257_115 =10'b0;

   // m257_116 = W*in
   wire signed [9:0] m257_116;
   assign m257_116 =10'b0;

   // m257_117 = W*in
   wire signed [9:0] m257_117;
   assign m257_117 =10'b0;

   // m258_1 = W*in
   wire signed [9:0] m258_1;
   assign m258_1 =10'b0;

   // m258_2 = W*in
   wire signed [9:0] m258_2;
   assign m258_2 =10'b0;

   // m258_3 = W*in
   wire signed [9:0] m258_3;
   assign m258_3 =10'b0;

   // m258_4 = W*in
   wire signed [9:0] m258_4;
   assign m258_4 =10'b0;

   // m258_5 = W*in
   wire signed [9:0] m258_5;
   assign m258_5 =10'b0;

   // m258_6 = W*in
   wire signed [9:0] m258_6;
   assign m258_6 =10'b0;

   // m258_7 = W*in
   wire signed [9:0] m258_7;
   assign m258_7 =10'b0;

   // m258_8 = W*in
   wire signed [9:0] m258_8;
   assign m258_8 =10'b0;

   // m258_9 = W*in
   wire signed [9:0] m258_9;
   assign m258_9 =10'b0;

   // m258_10 = W*in
   wire signed [9:0] m258_10;
   assign m258_10 =10'b0;

   // m258_11 = W*in
   wire signed [9:0] m258_11;
   assign m258_11 =10'b0;

   // m258_12 = W*in
   wire signed [9:0] m258_12;
   assign m258_12 =10'b0;

   // m258_13 = W*in
   wire signed [9:0] m258_13;
   assign m258_13 =10'b0;

   // m258_14 = W*in
   wire signed [9:0] m258_14;
   assign m258_14 =10'b0;

   // m258_15 = W*in
   wire signed [9:0] m258_15;
   assign m258_15 =10'b0;

   // m258_16 = W*in
   wire signed [9:0] m258_16;
   assign m258_16 =10'b0;

   // m258_17 = W*in
   wire signed [9:0] m258_17;
   assign m258_17 ={ {5{in258[5]}} , in258[5:1] };

   // m258_18 = W*in
   wire signed [9:0] m258_18;
   assign m258_18 =10'b0;

   // m258_19 = W*in
   wire signed [9:0] m258_19;
   assign m258_19 =10'b0;

   // m258_20 = W*in
   wire signed [9:0] m258_20;
   assign m258_20 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_21 = W*in
   wire signed [9:0] m258_21;
   assign m258_21 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_22 = W*in
   wire signed [9:0] m258_22;
   assign m258_22 =10'b0;

   // m258_23 = W*in
   wire signed [9:0] m258_23;
   assign m258_23 =10'b0;

   // m258_24 = W*in
   wire signed [9:0] m258_24;
   assign m258_24 =10'b0;

   // m258_25 = W*in
   wire signed [9:0] m258_25;
   assign m258_25 ={ {5{in258[5]}} , in258[5:1] };

   // m258_26 = W*in
   wire signed [9:0] m258_26;
   assign m258_26 =10'b0;

   // m258_27 = W*in
   wire signed [9:0] m258_27;
   assign m258_27 ={ {5{in258[5]}} , in258[5:1] };

   // m258_28 = W*in
   wire signed [9:0] m258_28;
   assign m258_28 ={ {4{in258[5]}} , in258[5:0] };

   // m258_29 = W*in
   wire signed [9:0] m258_29;
   assign m258_29 =10'b0;

   // m258_30 = W*in
   wire signed [9:0] m258_30;
   assign m258_30 =10'b0;

   // m258_31 = W*in
   wire signed [9:0] m258_31;
   assign m258_31 =10'b0;

   // m258_32 = W*in
   wire signed [9:0] m258_32;
   assign m258_32 =10'b0;

   // m258_33 = W*in
   wire signed [9:0] m258_33;
   assign m258_33 =10'b0;

   // m258_34 = W*in
   wire signed [9:0] m258_34;
   assign m258_34 =10'b0;

   // m258_35 = W*in
   wire signed [9:0] m258_35;
   assign m258_35 =10'b0;

   // m258_36 = W*in
   wire signed [9:0] m258_36;
   assign m258_36 =10'b0;

   // m258_37 = W*in
   wire signed [9:0] m258_37;
   assign m258_37 =10'b0;

   // m258_38 = W*in
   wire signed [9:0] m258_38;
   assign m258_38 =10'b0;

   // m258_39 = W*in
   wire signed [9:0] m258_39;
   assign m258_39 =10'b0;

   // m258_40 = W*in
   wire signed [9:0] m258_40;
   assign m258_40 =10'b0;

   // m258_41 = W*in
   wire signed [9:0] m258_41;
   assign m258_41 =10'b0;

   // m258_42 = W*in
   wire signed [9:0] m258_42;
   assign m258_42 =10'b0;

   // m258_43 = W*in
   wire signed [9:0] m258_43;
   assign m258_43 ={ {4{in258[5]}} , in258[5:0] };

   // m258_44 = W*in
   wire signed [9:0] m258_44;
   assign m258_44 =10'b0;

   // m258_45 = W*in
   wire signed [9:0] m258_45;
   assign m258_45 =10'b0;

   // m258_46 = W*in
   wire signed [9:0] m258_46;
   assign m258_46 ={ {4{in258[5]}} , in258[5:0] };

   // m258_47 = W*in
   wire signed [9:0] m258_47;
   assign m258_47 =10'b0;

   // m258_48 = W*in
   wire signed [9:0] m258_48;
   assign m258_48 =10'b0;

   // m258_49 = W*in
   wire signed [9:0] m258_49;
   assign m258_49 =10'b0;

   // m258_50 = W*in
   wire signed [9:0] m258_50;
   assign m258_50 =10'b0;

   // m258_51 = W*in
   wire signed [9:0] m258_51;
   assign m258_51 =10'b0;

   // m258_52 = W*in
   wire signed [9:0] m258_52;
   assign m258_52 =10'b0;

   // m258_53 = W*in
   wire signed [9:0] m258_53;
   assign m258_53 =10'b0;

   // m258_54 = W*in
   wire signed [9:0] m258_54;
   assign m258_54 =10'b0;

   // m258_55 = W*in
   wire signed [9:0] m258_55;
   assign m258_55 =10'b0;

   // m258_56 = W*in
   wire signed [9:0] m258_56;
   assign m258_56 =10'b0;

   // m258_57 = W*in
   wire signed [9:0] m258_57;
   assign m258_57 =10'b0;

   // m258_58 = W*in
   wire signed [9:0] m258_58;
   assign m258_58 =10'b0;

   // m258_59 = W*in
   wire signed [9:0] m258_59;
   assign m258_59 ={ {4{in258[5]}} , in258[5:0] };

   // m258_60 = W*in
   wire signed [9:0] m258_60;
   assign m258_60 =10'b0;

   // m258_61 = W*in
   wire signed [9:0] m258_61;
   assign m258_61 =10'b0;

   // m258_62 = W*in
   wire signed [9:0] m258_62;
   assign m258_62 =10'b0;

   // m258_63 = W*in
   wire signed [9:0] m258_63;
   assign m258_63 =10'b0;

   // m258_64 = W*in
   wire signed [9:0] m258_64;
   assign m258_64 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_65 = W*in
   wire signed [9:0] m258_65;
   assign m258_65 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_66 = W*in
   wire signed [9:0] m258_66;
   assign m258_66 =10'b0;

   // m258_67 = W*in
   wire signed [9:0] m258_67;
   assign m258_67 ={ {4{neg258[5]}} , neg258[5:0] };

   // m258_68 = W*in
   wire signed [9:0] m258_68;
   assign m258_68 =10'b0;

   // m258_69 = W*in
   wire signed [9:0] m258_69;
   assign m258_69 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_70 = W*in
   wire signed [9:0] m258_70;
   assign m258_70 =10'b0;

   // m258_71 = W*in
   wire signed [9:0] m258_71;
   assign m258_71 ={ {4{in258[5]}} , in258[5:0] };

   // m258_72 = W*in
   wire signed [9:0] m258_72;
   assign m258_72 ={ {5{in258[5]}} , in258[5:1] };

   // m258_73 = W*in
   wire signed [9:0] m258_73;
   assign m258_73 =10'b0;

   // m258_74 = W*in
   wire signed [9:0] m258_74;
   assign m258_74 =10'b0;

   // m258_75 = W*in
   wire signed [9:0] m258_75;
   assign m258_75 =10'b0;

   // m258_76 = W*in
   wire signed [9:0] m258_76;
   assign m258_76 =10'b0;

   // m258_77 = W*in
   wire signed [9:0] m258_77;
   assign m258_77 ={ {4{in258[5]}} , in258[5:0] };

   // m258_78 = W*in
   wire signed [9:0] m258_78;
   assign m258_78 =10'b0;

   // m258_79 = W*in
   wire signed [9:0] m258_79;
   assign m258_79 =10'b0;

   // m258_80 = W*in
   wire signed [9:0] m258_80;
   assign m258_80 =10'b0;

   // m258_81 = W*in
   wire signed [9:0] m258_81;
   assign m258_81 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_82 = W*in
   wire signed [9:0] m258_82;
   assign m258_82 =10'b0;

   // m258_83 = W*in
   wire signed [9:0] m258_83;
   assign m258_83 ={ {5{in258[5]}} , in258[5:1] };

   // m258_84 = W*in
   wire signed [9:0] m258_84;
   assign m258_84 =10'b0;

   // m258_85 = W*in
   wire signed [9:0] m258_85;
   assign m258_85 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_86 = W*in
   wire signed [9:0] m258_86;
   assign m258_86 =10'b0;

   // m258_87 = W*in
   wire signed [9:0] m258_87;
   assign m258_87 =10'b0;

   // m258_88 = W*in
   wire signed [9:0] m258_88;
   assign m258_88 =10'b0;

   // m258_89 = W*in
   wire signed [9:0] m258_89;
   assign m258_89 =10'b0;

   // m258_90 = W*in
   wire signed [9:0] m258_90;
   assign m258_90 =10'b0;

   // m258_91 = W*in
   wire signed [9:0] m258_91;
   assign m258_91 =10'b0;

   // m258_92 = W*in
   wire signed [9:0] m258_92;
   assign m258_92 =10'b0;

   // m258_93 = W*in
   wire signed [9:0] m258_93;
   assign m258_93 ={ {4{neg258[5]}} , neg258[5:0] };

   // m258_94 = W*in
   wire signed [9:0] m258_94;
   assign m258_94 =10'b0;

   // m258_95 = W*in
   wire signed [9:0] m258_95;
   assign m258_95 =10'b0;

   // m258_96 = W*in
   wire signed [9:0] m258_96;
   assign m258_96 =10'b0;

   // m258_97 = W*in
   wire signed [9:0] m258_97;
   assign m258_97 =10'b0;

   // m258_98 = W*in
   wire signed [9:0] m258_98;
   assign m258_98 =10'b0;

   // m258_99 = W*in
   wire signed [9:0] m258_99;
   assign m258_99 =10'b0;

   // m258_100 = W*in
   wire signed [9:0] m258_100;
   assign m258_100 =10'b0;

   // m258_101 = W*in
   wire signed [9:0] m258_101;
   assign m258_101 =10'b0;

   // m258_102 = W*in
   wire signed [9:0] m258_102;
   assign m258_102 =10'b0;

   // m258_103 = W*in
   wire signed [9:0] m258_103;
   assign m258_103 ={ {4{in258[5]}} , in258[5:0] };

   // m258_104 = W*in
   wire signed [9:0] m258_104;
   assign m258_104 ={ {4{in258[5]}} , in258[5:0] };

   // m258_105 = W*in
   wire signed [9:0] m258_105;
   assign m258_105 =10'b0;

   // m258_106 = W*in
   wire signed [9:0] m258_106;
   assign m258_106 =10'b0;

   // m258_107 = W*in
   wire signed [9:0] m258_107;
   assign m258_107 =10'b0;

   // m258_108 = W*in
   wire signed [9:0] m258_108;
   assign m258_108 =10'b0;

   // m258_109 = W*in
   wire signed [9:0] m258_109;
   assign m258_109 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_110 = W*in
   wire signed [9:0] m258_110;
   assign m258_110 =10'b0;

   // m258_111 = W*in
   wire signed [9:0] m258_111;
   assign m258_111 =10'b0;

   // m258_112 = W*in
   wire signed [9:0] m258_112;
   assign m258_112 =10'b0;

   // m258_113 = W*in
   wire signed [9:0] m258_113;
   assign m258_113 =10'b0;

   // m258_114 = W*in
   wire signed [9:0] m258_114;
   assign m258_114 ={ {5{neg258[5]}} , neg258[5:1] };

   // m258_115 = W*in
   wire signed [9:0] m258_115;
   assign m258_115 =10'b0;

   // m258_116 = W*in
   wire signed [9:0] m258_116;
   assign m258_116 =10'b0;

   // m258_117 = W*in
   wire signed [9:0] m258_117;
   assign m258_117 =10'b0;

   // m259_1 = W*in
   wire signed [9:0] m259_1;
   assign m259_1 =10'b0;

   // m259_2 = W*in
   wire signed [9:0] m259_2;
   assign m259_2 =10'b0;

   // m259_3 = W*in
   wire signed [9:0] m259_3;
   assign m259_3 =10'b0;

   // m259_4 = W*in
   wire signed [9:0] m259_4;
   assign m259_4 =10'b0;

   // m259_5 = W*in
   wire signed [9:0] m259_5;
   assign m259_5 =10'b0;

   // m259_6 = W*in
   wire signed [9:0] m259_6;
   assign m259_6 =10'b0;

   // m259_7 = W*in
   wire signed [9:0] m259_7;
   assign m259_7 =10'b0;

   // m259_8 = W*in
   wire signed [9:0] m259_8;
   assign m259_8 =10'b0;

   // m259_9 = W*in
   wire signed [9:0] m259_9;
   assign m259_9 =10'b0;

   // m259_10 = W*in
   wire signed [9:0] m259_10;
   assign m259_10 =10'b0;

   // m259_11 = W*in
   wire signed [9:0] m259_11;
   assign m259_11 =10'b0;

   // m259_12 = W*in
   wire signed [9:0] m259_12;
   assign m259_12 =10'b0;

   // m259_13 = W*in
   wire signed [9:0] m259_13;
   assign m259_13 =10'b0;

   // m259_14 = W*in
   wire signed [9:0] m259_14;
   assign m259_14 =10'b0;

   // m259_15 = W*in
   wire signed [9:0] m259_15;
   assign m259_15 =10'b0;

   // m259_16 = W*in
   wire signed [9:0] m259_16;
   assign m259_16 =10'b0;

   // m259_17 = W*in
   wire signed [9:0] m259_17;
   assign m259_17 =10'b0;

   // m259_18 = W*in
   wire signed [9:0] m259_18;
   assign m259_18 =10'b0;

   // m259_19 = W*in
   wire signed [9:0] m259_19;
   assign m259_19 ={ {4{in259[5]}} , in259[5:0] };

   // m259_20 = W*in
   wire signed [9:0] m259_20;
   assign m259_20 =10'b0;

   // m259_21 = W*in
   wire signed [9:0] m259_21;
   assign m259_21 =10'b0;

   // m259_22 = W*in
   wire signed [9:0] m259_22;
   assign m259_22 =10'b0;

   // m259_23 = W*in
   wire signed [9:0] m259_23;
   assign m259_23 =10'b0;

   // m259_24 = W*in
   wire signed [9:0] m259_24;
   assign m259_24 =10'b0;

   // m259_25 = W*in
   wire signed [9:0] m259_25;
   assign m259_25 =10'b0;

   // m259_26 = W*in
   wire signed [9:0] m259_26;
   assign m259_26 =10'b0;

   // m259_27 = W*in
   wire signed [9:0] m259_27;
   assign m259_27 =10'b0;

   // m259_28 = W*in
   wire signed [9:0] m259_28;
   assign m259_28 =10'b0;

   // m259_29 = W*in
   wire signed [9:0] m259_29;
   assign m259_29 =10'b0;

   // m259_30 = W*in
   wire signed [9:0] m259_30;
   assign m259_30 =10'b0;

   // m259_31 = W*in
   wire signed [9:0] m259_31;
   assign m259_31 =10'b0;

   // m259_32 = W*in
   wire signed [9:0] m259_32;
   assign m259_32 =10'b0;

   // m259_33 = W*in
   wire signed [9:0] m259_33;
   assign m259_33 =10'b0;

   // m259_34 = W*in
   wire signed [9:0] m259_34;
   assign m259_34 ={ {5{neg259[5]}} , neg259[5:1] };

   // m259_35 = W*in
   wire signed [9:0] m259_35;
   assign m259_35 =10'b0;

   // m259_36 = W*in
   wire signed [9:0] m259_36;
   assign m259_36 =10'b0;

   // m259_37 = W*in
   wire signed [9:0] m259_37;
   assign m259_37 =10'b0;

   // m259_38 = W*in
   wire signed [9:0] m259_38;
   assign m259_38 =10'b0;

   // m259_39 = W*in
   wire signed [9:0] m259_39;
   assign m259_39 =10'b0;

   // m259_40 = W*in
   wire signed [9:0] m259_40;
   assign m259_40 =10'b0;

   // m259_41 = W*in
   wire signed [9:0] m259_41;
   assign m259_41 =10'b0;

   // m259_42 = W*in
   wire signed [9:0] m259_42;
   assign m259_42 =10'b0;

   // m259_43 = W*in
   wire signed [9:0] m259_43;
   assign m259_43 =10'b0;

   // m259_44 = W*in
   wire signed [9:0] m259_44;
   assign m259_44 ={ {4{in259[5]}} , in259[5:0] };

   // m259_45 = W*in
   wire signed [9:0] m259_45;
   assign m259_45 =10'b0;

   // m259_46 = W*in
   wire signed [9:0] m259_46;
   assign m259_46 =10'b0;

   // m259_47 = W*in
   wire signed [9:0] m259_47;
   assign m259_47 =10'b0;

   // m259_48 = W*in
   wire signed [9:0] m259_48;
   assign m259_48 =10'b0;

   // m259_49 = W*in
   wire signed [9:0] m259_49;
   assign m259_49 =10'b0;

   // m259_50 = W*in
   wire signed [9:0] m259_50;
   assign m259_50 =10'b0;

   // m259_51 = W*in
   wire signed [9:0] m259_51;
   assign m259_51 =10'b0;

   // m259_52 = W*in
   wire signed [9:0] m259_52;
   assign m259_52 =10'b0;

   // m259_53 = W*in
   wire signed [9:0] m259_53;
   assign m259_53 ={ {4{in259[5]}} , in259[5:0] };

   // m259_54 = W*in
   wire signed [9:0] m259_54;
   assign m259_54 =10'b0;

   // m259_55 = W*in
   wire signed [9:0] m259_55;
   assign m259_55 =10'b0;

   // m259_56 = W*in
   wire signed [9:0] m259_56;
   assign m259_56 =10'b0;

   // m259_57 = W*in
   wire signed [9:0] m259_57;
   assign m259_57 =10'b0;

   // m259_58 = W*in
   wire signed [9:0] m259_58;
   assign m259_58 =10'b0;

   // m259_59 = W*in
   wire signed [9:0] m259_59;
   assign m259_59 =10'b0;

   // m259_60 = W*in
   wire signed [9:0] m259_60;
   assign m259_60 =10'b0;

   // m259_61 = W*in
   wire signed [9:0] m259_61;
   assign m259_61 =10'b0;

   // m259_62 = W*in
   wire signed [9:0] m259_62;
   assign m259_62 =10'b0;

   // m259_63 = W*in
   wire signed [9:0] m259_63;
   assign m259_63 =10'b0;

   // m259_64 = W*in
   wire signed [9:0] m259_64;
   assign m259_64 =10'b0;

   // m259_65 = W*in
   wire signed [9:0] m259_65;
   assign m259_65 =10'b0;

   // m259_66 = W*in
   wire signed [9:0] m259_66;
   assign m259_66 =10'b0;

   // m259_67 = W*in
   wire signed [9:0] m259_67;
   assign m259_67 ={ {4{in259[5]}} , in259[5:0] };

   // m259_68 = W*in
   wire signed [9:0] m259_68;
   assign m259_68 =10'b0;

   // m259_69 = W*in
   wire signed [9:0] m259_69;
   assign m259_69 =10'b0;

   // m259_70 = W*in
   wire signed [9:0] m259_70;
   assign m259_70 ={ {5{neg259[5]}} , neg259[5:1] };

   // m259_71 = W*in
   wire signed [9:0] m259_71;
   assign m259_71 =10'b0;

   // m259_72 = W*in
   wire signed [9:0] m259_72;
   assign m259_72 =10'b0;

   // m259_73 = W*in
   wire signed [9:0] m259_73;
   assign m259_73 =10'b0;

   // m259_74 = W*in
   wire signed [9:0] m259_74;
   assign m259_74 =10'b0;

   // m259_75 = W*in
   wire signed [9:0] m259_75;
   assign m259_75 =10'b0;

   // m259_76 = W*in
   wire signed [9:0] m259_76;
   assign m259_76 =10'b0;

   // m259_77 = W*in
   wire signed [9:0] m259_77;
   assign m259_77 =10'b0;

   // m259_78 = W*in
   wire signed [9:0] m259_78;
   assign m259_78 =10'b0;

   // m259_79 = W*in
   wire signed [9:0] m259_79;
   assign m259_79 =10'b0;

   // m259_80 = W*in
   wire signed [9:0] m259_80;
   assign m259_80 =10'b0;

   // m259_81 = W*in
   wire signed [9:0] m259_81;
   assign m259_81 ={ {5{neg259[5]}} , neg259[5:1] };

   // m259_82 = W*in
   wire signed [9:0] m259_82;
   assign m259_82 =10'b0;

   // m259_83 = W*in
   wire signed [9:0] m259_83;
   assign m259_83 ={ {5{neg259[5]}} , neg259[5:1] };

   // m259_84 = W*in
   wire signed [9:0] m259_84;
   assign m259_84 =10'b0;

   // m259_85 = W*in
   wire signed [9:0] m259_85;
   assign m259_85 =10'b0;

   // m259_86 = W*in
   wire signed [9:0] m259_86;
   assign m259_86 =10'b0;

   // m259_87 = W*in
   wire signed [9:0] m259_87;
   assign m259_87 =10'b0;

   // m259_88 = W*in
   wire signed [9:0] m259_88;
   assign m259_88 =10'b0;

   // m259_89 = W*in
   wire signed [9:0] m259_89;
   assign m259_89 =10'b0;

   // m259_90 = W*in
   wire signed [9:0] m259_90;
   assign m259_90 =10'b0;

   // m259_91 = W*in
   wire signed [9:0] m259_91;
   assign m259_91 =10'b0;

   // m259_92 = W*in
   wire signed [9:0] m259_92;
   assign m259_92 =10'b0;

   // m259_93 = W*in
   wire signed [9:0] m259_93;
   assign m259_93 ={ {4{in259[5]}} , in259[5:0] };

   // m259_94 = W*in
   wire signed [9:0] m259_94;
   assign m259_94 =10'b0;

   // m259_95 = W*in
   wire signed [9:0] m259_95;
   assign m259_95 =10'b0;

   // m259_96 = W*in
   wire signed [9:0] m259_96;
   assign m259_96 =10'b0;

   // m259_97 = W*in
   wire signed [9:0] m259_97;
   assign m259_97 =10'b0;

   // m259_98 = W*in
   wire signed [9:0] m259_98;
   assign m259_98 =10'b0;

   // m259_99 = W*in
   wire signed [9:0] m259_99;
   assign m259_99 =10'b0;

   // m259_100 = W*in
   wire signed [9:0] m259_100;
   assign m259_100 =10'b0;

   // m259_101 = W*in
   wire signed [9:0] m259_101;
   assign m259_101 =10'b0;

   // m259_102 = W*in
   wire signed [9:0] m259_102;
   assign m259_102 =10'b0;

   // m259_103 = W*in
   wire signed [9:0] m259_103;
   assign m259_103 =10'b0;

   // m259_104 = W*in
   wire signed [9:0] m259_104;
   assign m259_104 =10'b0;

   // m259_105 = W*in
   wire signed [9:0] m259_105;
   assign m259_105 =10'b0;

   // m259_106 = W*in
   wire signed [9:0] m259_106;
   assign m259_106 =10'b0;

   // m259_107 = W*in
   wire signed [9:0] m259_107;
   assign m259_107 =10'b0;

   // m259_108 = W*in
   wire signed [9:0] m259_108;
   assign m259_108 ={ {5{neg259[5]}} , neg259[5:1] };

   // m259_109 = W*in
   wire signed [9:0] m259_109;
   assign m259_109 ={ {5{neg259[5]}} , neg259[5:1] };

   // m259_110 = W*in
   wire signed [9:0] m259_110;
   assign m259_110 =10'b0;

   // m259_111 = W*in
   wire signed [9:0] m259_111;
   assign m259_111 =10'b0;

   // m259_112 = W*in
   wire signed [9:0] m259_112;
   assign m259_112 =10'b0;

   // m259_113 = W*in
   wire signed [9:0] m259_113;
   assign m259_113 =10'b0;

   // m259_114 = W*in
   wire signed [9:0] m259_114;
   assign m259_114 =10'b0;

   // m259_115 = W*in
   wire signed [9:0] m259_115;
   assign m259_115 =10'b0;

   // m259_116 = W*in
   wire signed [9:0] m259_116;
   assign m259_116 =10'b0;

   // m259_117 = W*in
   wire signed [9:0] m259_117;
   assign m259_117 =10'b0;

   // m260_1 = W*in
   wire signed [9:0] m260_1;
   assign m260_1 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_2 = W*in
   wire signed [9:0] m260_2;
   assign m260_2 ={ {4{in260[5]}} , in260[5:0] };

   // m260_3 = W*in
   wire signed [9:0] m260_3;
   assign m260_3 =10'b0;

   // m260_4 = W*in
   wire signed [9:0] m260_4;
   assign m260_4 =10'b0;

   // m260_5 = W*in
   wire signed [9:0] m260_5;
   assign m260_5 ={ {4{in260[5]}} , in260[5:0] };

   // m260_6 = W*in
   wire signed [9:0] m260_6;
   assign m260_6 =10'b0;

   // m260_7 = W*in
   wire signed [9:0] m260_7;
   assign m260_7 =10'b0;

   // m260_8 = W*in
   wire signed [9:0] m260_8;
   assign m260_8 ={ {4{in260[5]}} , in260[5:0] };

   // m260_9 = W*in
   wire signed [9:0] m260_9;
   assign m260_9 =10'b0;

   // m260_10 = W*in
   wire signed [9:0] m260_10;
   assign m260_10 =10'b0;

   // m260_11 = W*in
   wire signed [9:0] m260_11;
   assign m260_11 =10'b0;

   // m260_12 = W*in
   wire signed [9:0] m260_12;
   assign m260_12 =10'b0;

   // m260_13 = W*in
   wire signed [9:0] m260_13;
   assign m260_13 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_14 = W*in
   wire signed [9:0] m260_14;
   assign m260_14 =10'b0;

   // m260_15 = W*in
   wire signed [9:0] m260_15;
   assign m260_15 =10'b0;

   // m260_16 = W*in
   wire signed [9:0] m260_16;
   assign m260_16 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_17 = W*in
   wire signed [9:0] m260_17;
   assign m260_17 =10'b0;

   // m260_18 = W*in
   wire signed [9:0] m260_18;
   assign m260_18 =10'b0;

   // m260_19 = W*in
   wire signed [9:0] m260_19;
   assign m260_19 ={ {4{in260[5]}} , in260[5:0] };

   // m260_20 = W*in
   wire signed [9:0] m260_20;
   assign m260_20 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_21 = W*in
   wire signed [9:0] m260_21;
   assign m260_21 =10'b0;

   // m260_22 = W*in
   wire signed [9:0] m260_22;
   assign m260_22 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_23 = W*in
   wire signed [9:0] m260_23;
   assign m260_23 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_24 = W*in
   wire signed [9:0] m260_24;
   assign m260_24 =10'b0;

   // m260_25 = W*in
   wire signed [9:0] m260_25;
   assign m260_25 =10'b0;

   // m260_26 = W*in
   wire signed [9:0] m260_26;
   assign m260_26 =10'b0;

   // m260_27 = W*in
   wire signed [9:0] m260_27;
   assign m260_27 =10'b0;

   // m260_28 = W*in
   wire signed [9:0] m260_28;
   assign m260_28 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_29 = W*in
   wire signed [9:0] m260_29;
   assign m260_29 =10'b0;

   // m260_30 = W*in
   wire signed [9:0] m260_30;
   assign m260_30 =10'b0;

   // m260_31 = W*in
   wire signed [9:0] m260_31;
   assign m260_31 =10'b0;

   // m260_32 = W*in
   wire signed [9:0] m260_32;
   assign m260_32 ={ {4{in260[5]}} , in260[5:0] };

   // m260_33 = W*in
   wire signed [9:0] m260_33;
   assign m260_33 =10'b0;

   // m260_34 = W*in
   wire signed [9:0] m260_34;
   assign m260_34 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_35 = W*in
   wire signed [9:0] m260_35;
   assign m260_35 =10'b0;

   // m260_36 = W*in
   wire signed [9:0] m260_36;
   assign m260_36 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_37 = W*in
   wire signed [9:0] m260_37;
   assign m260_37 =10'b0;

   // m260_38 = W*in
   wire signed [9:0] m260_38;
   assign m260_38 =10'b0;

   // m260_39 = W*in
   wire signed [9:0] m260_39;
   assign m260_39 =10'b0;

   // m260_40 = W*in
   wire signed [9:0] m260_40;
   assign m260_40 =10'b0;

   // m260_41 = W*in
   wire signed [9:0] m260_41;
   assign m260_41 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_42 = W*in
   wire signed [9:0] m260_42;
   assign m260_42 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_43 = W*in
   wire signed [9:0] m260_43;
   assign m260_43 =10'b0;

   // m260_44 = W*in
   wire signed [9:0] m260_44;
   assign m260_44 ={ {4{in260[5]}} , in260[5:0] };

   // m260_45 = W*in
   wire signed [9:0] m260_45;
   assign m260_45 =10'b0;

   // m260_46 = W*in
   wire signed [9:0] m260_46;
   assign m260_46 =10'b0;

   // m260_47 = W*in
   wire signed [9:0] m260_47;
   assign m260_47 =10'b0;

   // m260_48 = W*in
   wire signed [9:0] m260_48;
   assign m260_48 =10'b0;

   // m260_49 = W*in
   wire signed [9:0] m260_49;
   assign m260_49 =10'b0;

   // m260_50 = W*in
   wire signed [9:0] m260_50;
   assign m260_50 =10'b0;

   // m260_51 = W*in
   wire signed [9:0] m260_51;
   assign m260_51 =10'b0;

   // m260_52 = W*in
   wire signed [9:0] m260_52;
   assign m260_52 =10'b0;

   // m260_53 = W*in
   wire signed [9:0] m260_53;
   assign m260_53 ={ {4{in260[5]}} , in260[5:0] };

   // m260_54 = W*in
   wire signed [9:0] m260_54;
   assign m260_54 ={ {4{in260[5]}} , in260[5:0] };

   // m260_55 = W*in
   wire signed [9:0] m260_55;
   assign m260_55 =10'b0;

   // m260_56 = W*in
   wire signed [9:0] m260_56;
   assign m260_56 =10'b0;

   // m260_57 = W*in
   wire signed [9:0] m260_57;
   assign m260_57 =10'b0;

   // m260_58 = W*in
   wire signed [9:0] m260_58;
   assign m260_58 =10'b0;

   // m260_59 = W*in
   wire signed [9:0] m260_59;
   assign m260_59 =10'b0;

   // m260_60 = W*in
   wire signed [9:0] m260_60;
   assign m260_60 =10'b0;

   // m260_61 = W*in
   wire signed [9:0] m260_61;
   assign m260_61 =10'b0;

   // m260_62 = W*in
   wire signed [9:0] m260_62;
   assign m260_62 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_63 = W*in
   wire signed [9:0] m260_63;
   assign m260_63 =10'b0;

   // m260_64 = W*in
   wire signed [9:0] m260_64;
   assign m260_64 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_65 = W*in
   wire signed [9:0] m260_65;
   assign m260_65 =10'b0;

   // m260_66 = W*in
   wire signed [9:0] m260_66;
   assign m260_66 =10'b0;

   // m260_67 = W*in
   wire signed [9:0] m260_67;
   assign m260_67 ={ {4{in260[5]}} , in260[5:0] };

   // m260_68 = W*in
   wire signed [9:0] m260_68;
   assign m260_68 ={ {4{in260[5]}} , in260[5:0] };

   // m260_69 = W*in
   wire signed [9:0] m260_69;
   assign m260_69 =10'b0;

   // m260_70 = W*in
   wire signed [9:0] m260_70;
   assign m260_70 =10'b0;

   // m260_71 = W*in
   wire signed [9:0] m260_71;
   assign m260_71 =10'b0;

   // m260_72 = W*in
   wire signed [9:0] m260_72;
   assign m260_72 =10'b0;

   // m260_73 = W*in
   wire signed [9:0] m260_73;
   assign m260_73 =10'b0;

   // m260_74 = W*in
   wire signed [9:0] m260_74;
   assign m260_74 =10'b0;

   // m260_75 = W*in
   wire signed [9:0] m260_75;
   assign m260_75 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_76 = W*in
   wire signed [9:0] m260_76;
   assign m260_76 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_77 = W*in
   wire signed [9:0] m260_77;
   assign m260_77 =10'b0;

   // m260_78 = W*in
   wire signed [9:0] m260_78;
   assign m260_78 =10'b0;

   // m260_79 = W*in
   wire signed [9:0] m260_79;
   assign m260_79 =10'b0;

   // m260_80 = W*in
   wire signed [9:0] m260_80;
   assign m260_80 ={ {4{in260[5]}} , in260[5:0] };

   // m260_81 = W*in
   wire signed [9:0] m260_81;
   assign m260_81 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_82 = W*in
   wire signed [9:0] m260_82;
   assign m260_82 =10'b0;

   // m260_83 = W*in
   wire signed [9:0] m260_83;
   assign m260_83 =10'b0;

   // m260_84 = W*in
   wire signed [9:0] m260_84;
   assign m260_84 =10'b0;

   // m260_85 = W*in
   wire signed [9:0] m260_85;
   assign m260_85 =10'b0;

   // m260_86 = W*in
   wire signed [9:0] m260_86;
   assign m260_86 =10'b0;

   // m260_87 = W*in
   wire signed [9:0] m260_87;
   assign m260_87 =10'b0;

   // m260_88 = W*in
   wire signed [9:0] m260_88;
   assign m260_88 =10'b0;

   // m260_89 = W*in
   wire signed [9:0] m260_89;
   assign m260_89 =10'b0;

   // m260_90 = W*in
   wire signed [9:0] m260_90;
   assign m260_90 =10'b0;

   // m260_91 = W*in
   wire signed [9:0] m260_91;
   assign m260_91 =10'b0;

   // m260_92 = W*in
   wire signed [9:0] m260_92;
   assign m260_92 =10'b0;

   // m260_93 = W*in
   wire signed [9:0] m260_93;
   assign m260_93 =10'b0;

   // m260_94 = W*in
   wire signed [9:0] m260_94;
   assign m260_94 =10'b0;

   // m260_95 = W*in
   wire signed [9:0] m260_95;
   assign m260_95 =10'b0;

   // m260_96 = W*in
   wire signed [9:0] m260_96;
   assign m260_96 =10'b0;

   // m260_97 = W*in
   wire signed [9:0] m260_97;
   assign m260_97 =10'b0;

   // m260_98 = W*in
   wire signed [9:0] m260_98;
   assign m260_98 =10'b0;

   // m260_99 = W*in
   wire signed [9:0] m260_99;
   assign m260_99 =10'b0;

   // m260_100 = W*in
   wire signed [9:0] m260_100;
   assign m260_100 =10'b0;

   // m260_101 = W*in
   wire signed [9:0] m260_101;
   assign m260_101 =10'b0;

   // m260_102 = W*in
   wire signed [9:0] m260_102;
   assign m260_102 =10'b0;

   // m260_103 = W*in
   wire signed [9:0] m260_103;
   assign m260_103 =10'b0;

   // m260_104 = W*in
   wire signed [9:0] m260_104;
   assign m260_104 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_105 = W*in
   wire signed [9:0] m260_105;
   assign m260_105 =10'b0;

   // m260_106 = W*in
   wire signed [9:0] m260_106;
   assign m260_106 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_107 = W*in
   wire signed [9:0] m260_107;
   assign m260_107 =10'b0;

   // m260_108 = W*in
   wire signed [9:0] m260_108;
   assign m260_108 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_109 = W*in
   wire signed [9:0] m260_109;
   assign m260_109 ={ {4{neg260[5]}} , neg260[5:0] };

   // m260_110 = W*in
   wire signed [9:0] m260_110;
   assign m260_110 =10'b0;

   // m260_111 = W*in
   wire signed [9:0] m260_111;
   assign m260_111 =10'b0;

   // m260_112 = W*in
   wire signed [9:0] m260_112;
   assign m260_112 =10'b0;

   // m260_113 = W*in
   wire signed [9:0] m260_113;
   assign m260_113 =10'b0;

   // m260_114 = W*in
   wire signed [9:0] m260_114;
   assign m260_114 ={ {5{neg260[5]}} , neg260[5:1] };

   // m260_115 = W*in
   wire signed [9:0] m260_115;
   assign m260_115 =10'b0;

   // m260_116 = W*in
   wire signed [9:0] m260_116;
   assign m260_116 =10'b0;

   // m260_117 = W*in
   wire signed [9:0] m260_117;
   assign m260_117 =10'b0;

   // m261_1 = W*in
   wire signed [9:0] m261_1;
   assign m261_1 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_2 = W*in
   wire signed [9:0] m261_2;
   assign m261_2 =10'b0;

   // m261_3 = W*in
   wire signed [9:0] m261_3;
   assign m261_3 =10'b0;

   // m261_4 = W*in
   wire signed [9:0] m261_4;
   assign m261_4 =10'b0;

   // m261_5 = W*in
   wire signed [9:0] m261_5;
   assign m261_5 ={ {4{in261[5]}} , in261[5:0] };

   // m261_6 = W*in
   wire signed [9:0] m261_6;
   assign m261_6 ={ {4{in261[5]}} , in261[5:0] };

   // m261_7 = W*in
   wire signed [9:0] m261_7;
   assign m261_7 =10'b0;

   // m261_8 = W*in
   wire signed [9:0] m261_8;
   assign m261_8 =10'b0;

   // m261_9 = W*in
   wire signed [9:0] m261_9;
   assign m261_9 =10'b0;

   // m261_10 = W*in
   wire signed [9:0] m261_10;
   assign m261_10 =10'b0;

   // m261_11 = W*in
   wire signed [9:0] m261_11;
   assign m261_11 =10'b0;

   // m261_12 = W*in
   wire signed [9:0] m261_12;
   assign m261_12 =10'b0;

   // m261_13 = W*in
   wire signed [9:0] m261_13;
   assign m261_13 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_14 = W*in
   wire signed [9:0] m261_14;
   assign m261_14 =10'b0;

   // m261_15 = W*in
   wire signed [9:0] m261_15;
   assign m261_15 =10'b0;

   // m261_16 = W*in
   wire signed [9:0] m261_16;
   assign m261_16 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_17 = W*in
   wire signed [9:0] m261_17;
   assign m261_17 =10'b0;

   // m261_18 = W*in
   wire signed [9:0] m261_18;
   assign m261_18 =10'b0;

   // m261_19 = W*in
   wire signed [9:0] m261_19;
   assign m261_19 ={ {4{in261[5]}} , in261[5:0] };

   // m261_20 = W*in
   wire signed [9:0] m261_20;
   assign m261_20 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_21 = W*in
   wire signed [9:0] m261_21;
   assign m261_21 ={ {4{in261[5]}} , in261[5:0] };

   // m261_22 = W*in
   wire signed [9:0] m261_22;
   assign m261_22 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_23 = W*in
   wire signed [9:0] m261_23;
   assign m261_23 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_24 = W*in
   wire signed [9:0] m261_24;
   assign m261_24 =10'b0;

   // m261_25 = W*in
   wire signed [9:0] m261_25;
   assign m261_25 =10'b0;

   // m261_26 = W*in
   wire signed [9:0] m261_26;
   assign m261_26 =10'b0;

   // m261_27 = W*in
   wire signed [9:0] m261_27;
   assign m261_27 =10'b0;

   // m261_28 = W*in
   wire signed [9:0] m261_28;
   assign m261_28 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_29 = W*in
   wire signed [9:0] m261_29;
   assign m261_29 =10'b0;

   // m261_30 = W*in
   wire signed [9:0] m261_30;
   assign m261_30 =10'b0;

   // m261_31 = W*in
   wire signed [9:0] m261_31;
   assign m261_31 ={ {5{in261[5]}} , in261[5:1] };

   // m261_32 = W*in
   wire signed [9:0] m261_32;
   assign m261_32 =10'b0;

   // m261_33 = W*in
   wire signed [9:0] m261_33;
   assign m261_33 =10'b0;

   // m261_34 = W*in
   wire signed [9:0] m261_34;
   assign m261_34 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_35 = W*in
   wire signed [9:0] m261_35;
   assign m261_35 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_36 = W*in
   wire signed [9:0] m261_36;
   assign m261_36 =10'b0;

   // m261_37 = W*in
   wire signed [9:0] m261_37;
   assign m261_37 =10'b0;

   // m261_38 = W*in
   wire signed [9:0] m261_38;
   assign m261_38 ={ {4{in261[5]}} , in261[5:0] };

   // m261_39 = W*in
   wire signed [9:0] m261_39;
   assign m261_39 =10'b0;

   // m261_40 = W*in
   wire signed [9:0] m261_40;
   assign m261_40 =10'b0;

   // m261_41 = W*in
   wire signed [9:0] m261_41;
   assign m261_41 =10'b0;

   // m261_42 = W*in
   wire signed [9:0] m261_42;
   assign m261_42 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_43 = W*in
   wire signed [9:0] m261_43;
   assign m261_43 =10'b0;

   // m261_44 = W*in
   wire signed [9:0] m261_44;
   assign m261_44 ={ {4{in261[5]}} , in261[5:0] };

   // m261_45 = W*in
   wire signed [9:0] m261_45;
   assign m261_45 =10'b0;

   // m261_46 = W*in
   wire signed [9:0] m261_46;
   assign m261_46 =10'b0;

   // m261_47 = W*in
   wire signed [9:0] m261_47;
   assign m261_47 =10'b0;

   // m261_48 = W*in
   wire signed [9:0] m261_48;
   assign m261_48 =10'b0;

   // m261_49 = W*in
   wire signed [9:0] m261_49;
   assign m261_49 =10'b0;

   // m261_50 = W*in
   wire signed [9:0] m261_50;
   assign m261_50 =10'b0;

   // m261_51 = W*in
   wire signed [9:0] m261_51;
   assign m261_51 =10'b0;

   // m261_52 = W*in
   wire signed [9:0] m261_52;
   assign m261_52 =10'b0;

   // m261_53 = W*in
   wire signed [9:0] m261_53;
   assign m261_53 ={ {4{in261[5]}} , in261[5:0] };

   // m261_54 = W*in
   wire signed [9:0] m261_54;
   assign m261_54 ={ {4{in261[5]}} , in261[5:0] };

   // m261_55 = W*in
   wire signed [9:0] m261_55;
   assign m261_55 =10'b0;

   // m261_56 = W*in
   wire signed [9:0] m261_56;
   assign m261_56 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_57 = W*in
   wire signed [9:0] m261_57;
   assign m261_57 =10'b0;

   // m261_58 = W*in
   wire signed [9:0] m261_58;
   assign m261_58 =10'b0;

   // m261_59 = W*in
   wire signed [9:0] m261_59;
   assign m261_59 =10'b0;

   // m261_60 = W*in
   wire signed [9:0] m261_60;
   assign m261_60 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_61 = W*in
   wire signed [9:0] m261_61;
   assign m261_61 =10'b0;

   // m261_62 = W*in
   wire signed [9:0] m261_62;
   assign m261_62 =10'b0;

   // m261_63 = W*in
   wire signed [9:0] m261_63;
   assign m261_63 ={ {4{in261[5]}} , in261[5:0] };

   // m261_64 = W*in
   wire signed [9:0] m261_64;
   assign m261_64 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_65 = W*in
   wire signed [9:0] m261_65;
   assign m261_65 =10'b0;

   // m261_66 = W*in
   wire signed [9:0] m261_66;
   assign m261_66 =10'b0;

   // m261_67 = W*in
   wire signed [9:0] m261_67;
   assign m261_67 =10'b0;

   // m261_68 = W*in
   wire signed [9:0] m261_68;
   assign m261_68 =10'b0;

   // m261_69 = W*in
   wire signed [9:0] m261_69;
   assign m261_69 ={ {4{in261[5]}} , in261[5:0] };

   // m261_70 = W*in
   wire signed [9:0] m261_70;
   assign m261_70 ={ {4{in261[5]}} , in261[5:0] };

   // m261_71 = W*in
   wire signed [9:0] m261_71;
   assign m261_71 =10'b0;

   // m261_72 = W*in
   wire signed [9:0] m261_72;
   assign m261_72 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_73 = W*in
   wire signed [9:0] m261_73;
   assign m261_73 =10'b0;

   // m261_74 = W*in
   wire signed [9:0] m261_74;
   assign m261_74 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_75 = W*in
   wire signed [9:0] m261_75;
   assign m261_75 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_76 = W*in
   wire signed [9:0] m261_76;
   assign m261_76 =10'b0;

   // m261_77 = W*in
   wire signed [9:0] m261_77;
   assign m261_77 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_78 = W*in
   wire signed [9:0] m261_78;
   assign m261_78 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_79 = W*in
   wire signed [9:0] m261_79;
   assign m261_79 ={ {4{in261[5]}} , in261[5:0] };

   // m261_80 = W*in
   wire signed [9:0] m261_80;
   assign m261_80 =10'b0;

   // m261_81 = W*in
   wire signed [9:0] m261_81;
   assign m261_81 ={ {4{neg261[5]}} , neg261[5:0] };

   // m261_82 = W*in
   wire signed [9:0] m261_82;
   assign m261_82 ={ {4{in261[5]}} , in261[5:0] };

   // m261_83 = W*in
   wire signed [9:0] m261_83;
   assign m261_83 =10'b0;

   // m261_84 = W*in
   wire signed [9:0] m261_84;
   assign m261_84 =10'b0;

   // m261_85 = W*in
   wire signed [9:0] m261_85;
   assign m261_85 ={ {4{in261[5]}} , in261[5:0] };

   // m261_86 = W*in
   wire signed [9:0] m261_86;
   assign m261_86 =10'b0;

   // m261_87 = W*in
   wire signed [9:0] m261_87;
   assign m261_87 =10'b0;

   // m261_88 = W*in
   wire signed [9:0] m261_88;
   assign m261_88 =10'b0;

   // m261_89 = W*in
   wire signed [9:0] m261_89;
   assign m261_89 =10'b0;

   // m261_90 = W*in
   wire signed [9:0] m261_90;
   assign m261_90 =10'b0;

   // m261_91 = W*in
   wire signed [9:0] m261_91;
   assign m261_91 =10'b0;

   // m261_92 = W*in
   wire signed [9:0] m261_92;
   assign m261_92 =10'b0;

   // m261_93 = W*in
   wire signed [9:0] m261_93;
   assign m261_93 ={ {4{in261[5]}} , in261[5:0] };

   // m261_94 = W*in
   wire signed [9:0] m261_94;
   assign m261_94 =10'b0;

   // m261_95 = W*in
   wire signed [9:0] m261_95;
   assign m261_95 =10'b0;

   // m261_96 = W*in
   wire signed [9:0] m261_96;
   assign m261_96 =10'b0;

   // m261_97 = W*in
   wire signed [9:0] m261_97;
   assign m261_97 =10'b0;

   // m261_98 = W*in
   wire signed [9:0] m261_98;
   assign m261_98 =10'b0;

   // m261_99 = W*in
   wire signed [9:0] m261_99;
   assign m261_99 =10'b0;

   // m261_100 = W*in
   wire signed [9:0] m261_100;
   assign m261_100 =10'b0;

   // m261_101 = W*in
   wire signed [9:0] m261_101;
   assign m261_101 =10'b0;

   // m261_102 = W*in
   wire signed [9:0] m261_102;
   assign m261_102 =10'b0;

   // m261_103 = W*in
   wire signed [9:0] m261_103;
   assign m261_103 =10'b0;

   // m261_104 = W*in
   wire signed [9:0] m261_104;
   assign m261_104 =10'b0;

   // m261_105 = W*in
   wire signed [9:0] m261_105;
   assign m261_105 =10'b0;

   // m261_106 = W*in
   wire signed [9:0] m261_106;
   assign m261_106 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_107 = W*in
   wire signed [9:0] m261_107;
   assign m261_107 =10'b0;

   // m261_108 = W*in
   wire signed [9:0] m261_108;
   assign m261_108 =10'b0;

   // m261_109 = W*in
   wire signed [9:0] m261_109;
   assign m261_109 =10'b0;

   // m261_110 = W*in
   wire signed [9:0] m261_110;
   assign m261_110 =10'b0;

   // m261_111 = W*in
   wire signed [9:0] m261_111;
   assign m261_111 =10'b0;

   // m261_112 = W*in
   wire signed [9:0] m261_112;
   assign m261_112 =10'b0;

   // m261_113 = W*in
   wire signed [9:0] m261_113;
   assign m261_113 =10'b0;

   // m261_114 = W*in
   wire signed [9:0] m261_114;
   assign m261_114 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_115 = W*in
   wire signed [9:0] m261_115;
   assign m261_115 ={ {5{neg261[5]}} , neg261[5:1] };

   // m261_116 = W*in
   wire signed [9:0] m261_116;
   assign m261_116 =10'b0;

   // m261_117 = W*in
   wire signed [9:0] m261_117;
   assign m261_117 ={ {4{neg261[5]}} , neg261[5:0] };

   // m262_1 = W*in
   wire signed [9:0] m262_1;
   assign m262_1 =10'b0;

   // m262_2 = W*in
   wire signed [9:0] m262_2;
   assign m262_2 =10'b0;

   // m262_3 = W*in
   wire signed [9:0] m262_3;
   assign m262_3 =10'b0;

   // m262_4 = W*in
   wire signed [9:0] m262_4;
   assign m262_4 =10'b0;

   // m262_5 = W*in
   wire signed [9:0] m262_5;
   assign m262_5 =10'b0;

   // m262_6 = W*in
   wire signed [9:0] m262_6;
   assign m262_6 ={ {4{neg262[5]}} , neg262[5:0] };

   // m262_7 = W*in
   wire signed [9:0] m262_7;
   assign m262_7 =10'b0;

   // m262_8 = W*in
   wire signed [9:0] m262_8;
   assign m262_8 =10'b0;

   // m262_9 = W*in
   wire signed [9:0] m262_9;
   assign m262_9 =10'b0;

   // m262_10 = W*in
   wire signed [9:0] m262_10;
   assign m262_10 =10'b0;

   // m262_11 = W*in
   wire signed [9:0] m262_11;
   assign m262_11 ={ {4{neg262[5]}} , neg262[5:0] };

   // m262_12 = W*in
   wire signed [9:0] m262_12;
   assign m262_12 =10'b0;

   // m262_13 = W*in
   wire signed [9:0] m262_13;
   assign m262_13 ={ {4{in262[5]}} , in262[5:0] };

   // m262_14 = W*in
   wire signed [9:0] m262_14;
   assign m262_14 =10'b0;

   // m262_15 = W*in
   wire signed [9:0] m262_15;
   assign m262_15 =10'b0;

   // m262_16 = W*in
   wire signed [9:0] m262_16;
   assign m262_16 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_17 = W*in
   wire signed [9:0] m262_17;
   assign m262_17 =10'b0;

   // m262_18 = W*in
   wire signed [9:0] m262_18;
   assign m262_18 =10'b0;

   // m262_19 = W*in
   wire signed [9:0] m262_19;
   assign m262_19 =10'b0;

   // m262_20 = W*in
   wire signed [9:0] m262_20;
   assign m262_20 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_21 = W*in
   wire signed [9:0] m262_21;
   assign m262_21 ={ {5{in262[5]}} , in262[5:1] };

   // m262_22 = W*in
   wire signed [9:0] m262_22;
   assign m262_22 =10'b0;

   // m262_23 = W*in
   wire signed [9:0] m262_23;
   assign m262_23 =10'b0;

   // m262_24 = W*in
   wire signed [9:0] m262_24;
   assign m262_24 =10'b0;

   // m262_25 = W*in
   wire signed [9:0] m262_25;
   assign m262_25 =10'b0;

   // m262_26 = W*in
   wire signed [9:0] m262_26;
   assign m262_26 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_27 = W*in
   wire signed [9:0] m262_27;
   assign m262_27 =10'b0;

   // m262_28 = W*in
   wire signed [9:0] m262_28;
   assign m262_28 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_29 = W*in
   wire signed [9:0] m262_29;
   assign m262_29 =10'b0;

   // m262_30 = W*in
   wire signed [9:0] m262_30;
   assign m262_30 =10'b0;

   // m262_31 = W*in
   wire signed [9:0] m262_31;
   assign m262_31 =10'b0;

   // m262_32 = W*in
   wire signed [9:0] m262_32;
   assign m262_32 =10'b0;

   // m262_33 = W*in
   wire signed [9:0] m262_33;
   assign m262_33 =10'b0;

   // m262_34 = W*in
   wire signed [9:0] m262_34;
   assign m262_34 =10'b0;

   // m262_35 = W*in
   wire signed [9:0] m262_35;
   assign m262_35 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_36 = W*in
   wire signed [9:0] m262_36;
   assign m262_36 =10'b0;

   // m262_37 = W*in
   wire signed [9:0] m262_37;
   assign m262_37 ={ {4{in262[5]}} , in262[5:0] };

   // m262_38 = W*in
   wire signed [9:0] m262_38;
   assign m262_38 =10'b0;

   // m262_39 = W*in
   wire signed [9:0] m262_39;
   assign m262_39 =10'b0;

   // m262_40 = W*in
   wire signed [9:0] m262_40;
   assign m262_40 =10'b0;

   // m262_41 = W*in
   wire signed [9:0] m262_41;
   assign m262_41 ={ {4{in262[5]}} , in262[5:0] };

   // m262_42 = W*in
   wire signed [9:0] m262_42;
   assign m262_42 =10'b0;

   // m262_43 = W*in
   wire signed [9:0] m262_43;
   assign m262_43 =10'b0;

   // m262_44 = W*in
   wire signed [9:0] m262_44;
   assign m262_44 =10'b0;

   // m262_45 = W*in
   wire signed [9:0] m262_45;
   assign m262_45 =10'b0;

   // m262_46 = W*in
   wire signed [9:0] m262_46;
   assign m262_46 =10'b0;

   // m262_47 = W*in
   wire signed [9:0] m262_47;
   assign m262_47 =10'b0;

   // m262_48 = W*in
   wire signed [9:0] m262_48;
   assign m262_48 =10'b0;

   // m262_49 = W*in
   wire signed [9:0] m262_49;
   assign m262_49 ={ {4{neg262[5]}} , neg262[5:0] };

   // m262_50 = W*in
   wire signed [9:0] m262_50;
   assign m262_50 =10'b0;

   // m262_51 = W*in
   wire signed [9:0] m262_51;
   assign m262_51 =10'b0;

   // m262_52 = W*in
   wire signed [9:0] m262_52;
   assign m262_52 =10'b0;

   // m262_53 = W*in
   wire signed [9:0] m262_53;
   assign m262_53 =10'b0;

   // m262_54 = W*in
   wire signed [9:0] m262_54;
   assign m262_54 ={ {4{neg262[5]}} , neg262[5:0] };

   // m262_55 = W*in
   wire signed [9:0] m262_55;
   assign m262_55 =10'b0;

   // m262_56 = W*in
   wire signed [9:0] m262_56;
   assign m262_56 =10'b0;

   // m262_57 = W*in
   wire signed [9:0] m262_57;
   assign m262_57 =10'b0;

   // m262_58 = W*in
   wire signed [9:0] m262_58;
   assign m262_58 =10'b0;

   // m262_59 = W*in
   wire signed [9:0] m262_59;
   assign m262_59 =10'b0;

   // m262_60 = W*in
   wire signed [9:0] m262_60;
   assign m262_60 =10'b0;

   // m262_61 = W*in
   wire signed [9:0] m262_61;
   assign m262_61 =10'b0;

   // m262_62 = W*in
   wire signed [9:0] m262_62;
   assign m262_62 =10'b0;

   // m262_63 = W*in
   wire signed [9:0] m262_63;
   assign m262_63 =10'b0;

   // m262_64 = W*in
   wire signed [9:0] m262_64;
   assign m262_64 ={ {4{neg262[5]}} , neg262[5:0] };

   // m262_65 = W*in
   wire signed [9:0] m262_65;
   assign m262_65 ={ {4{in262[5]}} , in262[5:0] };

   // m262_66 = W*in
   wire signed [9:0] m262_66;
   assign m262_66 ={ {4{in262[5]}} , in262[5:0] };

   // m262_67 = W*in
   wire signed [9:0] m262_67;
   assign m262_67 ={ {4{neg262[5]}} , neg262[5:0] };

   // m262_68 = W*in
   wire signed [9:0] m262_68;
   assign m262_68 =10'b0;

   // m262_69 = W*in
   wire signed [9:0] m262_69;
   assign m262_69 ={ {4{in262[5]}} , in262[5:0] };

   // m262_70 = W*in
   wire signed [9:0] m262_70;
   assign m262_70 ={ {4{in262[5]}} , in262[5:0] };

   // m262_71 = W*in
   wire signed [9:0] m262_71;
   assign m262_71 =10'b0;

   // m262_72 = W*in
   wire signed [9:0] m262_72;
   assign m262_72 =10'b0;

   // m262_73 = W*in
   wire signed [9:0] m262_73;
   assign m262_73 =10'b0;

   // m262_74 = W*in
   wire signed [9:0] m262_74;
   assign m262_74 =10'b0;

   // m262_75 = W*in
   wire signed [9:0] m262_75;
   assign m262_75 =10'b0;

   // m262_76 = W*in
   wire signed [9:0] m262_76;
   assign m262_76 =10'b0;

   // m262_77 = W*in
   wire signed [9:0] m262_77;
   assign m262_77 =10'b0;

   // m262_78 = W*in
   wire signed [9:0] m262_78;
   assign m262_78 =10'b0;

   // m262_79 = W*in
   wire signed [9:0] m262_79;
   assign m262_79 ={ {4{in262[5]}} , in262[5:0] };

   // m262_80 = W*in
   wire signed [9:0] m262_80;
   assign m262_80 =10'b0;

   // m262_81 = W*in
   wire signed [9:0] m262_81;
   assign m262_81 =10'b0;

   // m262_82 = W*in
   wire signed [9:0] m262_82;
   assign m262_82 ={ {4{in262[5]}} , in262[5:0] };

   // m262_83 = W*in
   wire signed [9:0] m262_83;
   assign m262_83 =10'b0;

   // m262_84 = W*in
   wire signed [9:0] m262_84;
   assign m262_84 =10'b0;

   // m262_85 = W*in
   wire signed [9:0] m262_85;
   assign m262_85 ={ {4{in262[5]}} , in262[5:0] };

   // m262_86 = W*in
   wire signed [9:0] m262_86;
   assign m262_86 =10'b0;

   // m262_87 = W*in
   wire signed [9:0] m262_87;
   assign m262_87 =10'b0;

   // m262_88 = W*in
   wire signed [9:0] m262_88;
   assign m262_88 =10'b0;

   // m262_89 = W*in
   wire signed [9:0] m262_89;
   assign m262_89 ={ {4{in262[5]}} , in262[5:0] };

   // m262_90 = W*in
   wire signed [9:0] m262_90;
   assign m262_90 =10'b0;

   // m262_91 = W*in
   wire signed [9:0] m262_91;
   assign m262_91 =10'b0;

   // m262_92 = W*in
   wire signed [9:0] m262_92;
   assign m262_92 =10'b0;

   // m262_93 = W*in
   wire signed [9:0] m262_93;
   assign m262_93 ={ {4{in262[5]}} , in262[5:0] };

   // m262_94 = W*in
   wire signed [9:0] m262_94;
   assign m262_94 =10'b0;

   // m262_95 = W*in
   wire signed [9:0] m262_95;
   assign m262_95 =10'b0;

   // m262_96 = W*in
   wire signed [9:0] m262_96;
   assign m262_96 ={ {4{in262[5]}} , in262[5:0] };

   // m262_97 = W*in
   wire signed [9:0] m262_97;
   assign m262_97 =10'b0;

   // m262_98 = W*in
   wire signed [9:0] m262_98;
   assign m262_98 =10'b0;

   // m262_99 = W*in
   wire signed [9:0] m262_99;
   assign m262_99 =10'b0;

   // m262_100 = W*in
   wire signed [9:0] m262_100;
   assign m262_100 =10'b0;

   // m262_101 = W*in
   wire signed [9:0] m262_101;
   assign m262_101 =10'b0;

   // m262_102 = W*in
   wire signed [9:0] m262_102;
   assign m262_102 =10'b0;

   // m262_103 = W*in
   wire signed [9:0] m262_103;
   assign m262_103 =10'b0;

   // m262_104 = W*in
   wire signed [9:0] m262_104;
   assign m262_104 =10'b0;

   // m262_105 = W*in
   wire signed [9:0] m262_105;
   assign m262_105 =10'b0;

   // m262_106 = W*in
   wire signed [9:0] m262_106;
   assign m262_106 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_107 = W*in
   wire signed [9:0] m262_107;
   assign m262_107 =10'b0;

   // m262_108 = W*in
   wire signed [9:0] m262_108;
   assign m262_108 ={ {4{in262[5]}} , in262[5:0] };

   // m262_109 = W*in
   wire signed [9:0] m262_109;
   assign m262_109 ={ {4{in262[5]}} , in262[5:0] };

   // m262_110 = W*in
   wire signed [9:0] m262_110;
   assign m262_110 =10'b0;

   // m262_111 = W*in
   wire signed [9:0] m262_111;
   assign m262_111 =10'b0;

   // m262_112 = W*in
   wire signed [9:0] m262_112;
   assign m262_112 =10'b0;

   // m262_113 = W*in
   wire signed [9:0] m262_113;
   assign m262_113 =10'b0;

   // m262_114 = W*in
   wire signed [9:0] m262_114;
   assign m262_114 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_115 = W*in
   wire signed [9:0] m262_115;
   assign m262_115 ={ {5{neg262[5]}} , neg262[5:1] };

   // m262_116 = W*in
   wire signed [9:0] m262_116;
   assign m262_116 ={ {4{in262[5]}} , in262[5:0] };

   // m262_117 = W*in
   wire signed [9:0] m262_117;
   assign m262_117 ={ {4{neg262[5]}} , neg262[5:0] };

   // m263_1 = W*in
   wire signed [9:0] m263_1;
   assign m263_1 =10'b0;

   // m263_2 = W*in
   wire signed [9:0] m263_2;
   assign m263_2 =10'b0;

   // m263_3 = W*in
   wire signed [9:0] m263_3;
   assign m263_3 =10'b0;

   // m263_4 = W*in
   wire signed [9:0] m263_4;
   assign m263_4 =10'b0;

   // m263_5 = W*in
   wire signed [9:0] m263_5;
   assign m263_5 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_6 = W*in
   wire signed [9:0] m263_6;
   assign m263_6 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_7 = W*in
   wire signed [9:0] m263_7;
   assign m263_7 =10'b0;

   // m263_8 = W*in
   wire signed [9:0] m263_8;
   assign m263_8 =10'b0;

   // m263_9 = W*in
   wire signed [9:0] m263_9;
   assign m263_9 =10'b0;

   // m263_10 = W*in
   wire signed [9:0] m263_10;
   assign m263_10 =10'b0;

   // m263_11 = W*in
   wire signed [9:0] m263_11;
   assign m263_11 =10'b0;

   // m263_12 = W*in
   wire signed [9:0] m263_12;
   assign m263_12 =10'b0;

   // m263_13 = W*in
   wire signed [9:0] m263_13;
   assign m263_13 ={ {4{in263[5]}} , in263[5:0] };

   // m263_14 = W*in
   wire signed [9:0] m263_14;
   assign m263_14 =10'b0;

   // m263_15 = W*in
   wire signed [9:0] m263_15;
   assign m263_15 =10'b0;

   // m263_16 = W*in
   wire signed [9:0] m263_16;
   assign m263_16 =10'b0;

   // m263_17 = W*in
   wire signed [9:0] m263_17;
   assign m263_17 =10'b0;

   // m263_18 = W*in
   wire signed [9:0] m263_18;
   assign m263_18 =10'b0;

   // m263_19 = W*in
   wire signed [9:0] m263_19;
   assign m263_19 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_20 = W*in
   wire signed [9:0] m263_20;
   assign m263_20 ={ {5{in263[5]}} , in263[5:1] };

   // m263_21 = W*in
   wire signed [9:0] m263_21;
   assign m263_21 =10'b0;

   // m263_22 = W*in
   wire signed [9:0] m263_22;
   assign m263_22 =10'b0;

   // m263_23 = W*in
   wire signed [9:0] m263_23;
   assign m263_23 =10'b0;

   // m263_24 = W*in
   wire signed [9:0] m263_24;
   assign m263_24 =10'b0;

   // m263_25 = W*in
   wire signed [9:0] m263_25;
   assign m263_25 =10'b0;

   // m263_26 = W*in
   wire signed [9:0] m263_26;
   assign m263_26 ={ {5{neg263[5]}} , neg263[5:1] };

   // m263_27 = W*in
   wire signed [9:0] m263_27;
   assign m263_27 =10'b0;

   // m263_28 = W*in
   wire signed [9:0] m263_28;
   assign m263_28 ={ {5{neg263[5]}} , neg263[5:1] };

   // m263_29 = W*in
   wire signed [9:0] m263_29;
   assign m263_29 =10'b0;

   // m263_30 = W*in
   wire signed [9:0] m263_30;
   assign m263_30 =10'b0;

   // m263_31 = W*in
   wire signed [9:0] m263_31;
   assign m263_31 =10'b0;

   // m263_32 = W*in
   wire signed [9:0] m263_32;
   assign m263_32 =10'b0;

   // m263_33 = W*in
   wire signed [9:0] m263_33;
   assign m263_33 =10'b0;

   // m263_34 = W*in
   wire signed [9:0] m263_34;
   assign m263_34 =10'b0;

   // m263_35 = W*in
   wire signed [9:0] m263_35;
   assign m263_35 =10'b0;

   // m263_36 = W*in
   wire signed [9:0] m263_36;
   assign m263_36 =10'b0;

   // m263_37 = W*in
   wire signed [9:0] m263_37;
   assign m263_37 =10'b0;

   // m263_38 = W*in
   wire signed [9:0] m263_38;
   assign m263_38 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_39 = W*in
   wire signed [9:0] m263_39;
   assign m263_39 =10'b0;

   // m263_40 = W*in
   wire signed [9:0] m263_40;
   assign m263_40 =10'b0;

   // m263_41 = W*in
   wire signed [9:0] m263_41;
   assign m263_41 ={ {4{in263[5]}} , in263[5:0] };

   // m263_42 = W*in
   wire signed [9:0] m263_42;
   assign m263_42 =10'b0;

   // m263_43 = W*in
   wire signed [9:0] m263_43;
   assign m263_43 =10'b0;

   // m263_44 = W*in
   wire signed [9:0] m263_44;
   assign m263_44 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_45 = W*in
   wire signed [9:0] m263_45;
   assign m263_45 =10'b0;

   // m263_46 = W*in
   wire signed [9:0] m263_46;
   assign m263_46 =10'b0;

   // m263_47 = W*in
   wire signed [9:0] m263_47;
   assign m263_47 =10'b0;

   // m263_48 = W*in
   wire signed [9:0] m263_48;
   assign m263_48 =10'b0;

   // m263_49 = W*in
   wire signed [9:0] m263_49;
   assign m263_49 =10'b0;

   // m263_50 = W*in
   wire signed [9:0] m263_50;
   assign m263_50 =10'b0;

   // m263_51 = W*in
   wire signed [9:0] m263_51;
   assign m263_51 =10'b0;

   // m263_52 = W*in
   wire signed [9:0] m263_52;
   assign m263_52 =10'b0;

   // m263_53 = W*in
   wire signed [9:0] m263_53;
   assign m263_53 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_54 = W*in
   wire signed [9:0] m263_54;
   assign m263_54 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_55 = W*in
   wire signed [9:0] m263_55;
   assign m263_55 =10'b0;

   // m263_56 = W*in
   wire signed [9:0] m263_56;
   assign m263_56 =10'b0;

   // m263_57 = W*in
   wire signed [9:0] m263_57;
   assign m263_57 =10'b0;

   // m263_58 = W*in
   wire signed [9:0] m263_58;
   assign m263_58 =10'b0;

   // m263_59 = W*in
   wire signed [9:0] m263_59;
   assign m263_59 =10'b0;

   // m263_60 = W*in
   wire signed [9:0] m263_60;
   assign m263_60 =10'b0;

   // m263_61 = W*in
   wire signed [9:0] m263_61;
   assign m263_61 =10'b0;

   // m263_62 = W*in
   wire signed [9:0] m263_62;
   assign m263_62 =10'b0;

   // m263_63 = W*in
   wire signed [9:0] m263_63;
   assign m263_63 =10'b0;

   // m263_64 = W*in
   wire signed [9:0] m263_64;
   assign m263_64 =10'b0;

   // m263_65 = W*in
   wire signed [9:0] m263_65;
   assign m263_65 ={ {5{in263[5]}} , in263[5:1] };

   // m263_66 = W*in
   wire signed [9:0] m263_66;
   assign m263_66 =10'b0;

   // m263_67 = W*in
   wire signed [9:0] m263_67;
   assign m263_67 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_68 = W*in
   wire signed [9:0] m263_68;
   assign m263_68 =10'b0;

   // m263_69 = W*in
   wire signed [9:0] m263_69;
   assign m263_69 ={ {5{in263[5]}} , in263[5:1] };

   // m263_70 = W*in
   wire signed [9:0] m263_70;
   assign m263_70 ={ {5{in263[5]}} , in263[5:1] };

   // m263_71 = W*in
   wire signed [9:0] m263_71;
   assign m263_71 ={ {5{neg263[5]}} , neg263[5:1] };

   // m263_72 = W*in
   wire signed [9:0] m263_72;
   assign m263_72 =10'b0;

   // m263_73 = W*in
   wire signed [9:0] m263_73;
   assign m263_73 =10'b0;

   // m263_74 = W*in
   wire signed [9:0] m263_74;
   assign m263_74 =10'b0;

   // m263_75 = W*in
   wire signed [9:0] m263_75;
   assign m263_75 =10'b0;

   // m263_76 = W*in
   wire signed [9:0] m263_76;
   assign m263_76 =10'b0;

   // m263_77 = W*in
   wire signed [9:0] m263_77;
   assign m263_77 =10'b0;

   // m263_78 = W*in
   wire signed [9:0] m263_78;
   assign m263_78 =10'b0;

   // m263_79 = W*in
   wire signed [9:0] m263_79;
   assign m263_79 =10'b0;

   // m263_80 = W*in
   wire signed [9:0] m263_80;
   assign m263_80 =10'b0;

   // m263_81 = W*in
   wire signed [9:0] m263_81;
   assign m263_81 =10'b0;

   // m263_82 = W*in
   wire signed [9:0] m263_82;
   assign m263_82 =10'b0;

   // m263_83 = W*in
   wire signed [9:0] m263_83;
   assign m263_83 =10'b0;

   // m263_84 = W*in
   wire signed [9:0] m263_84;
   assign m263_84 =10'b0;

   // m263_85 = W*in
   wire signed [9:0] m263_85;
   assign m263_85 =10'b0;

   // m263_86 = W*in
   wire signed [9:0] m263_86;
   assign m263_86 =10'b0;

   // m263_87 = W*in
   wire signed [9:0] m263_87;
   assign m263_87 =10'b0;

   // m263_88 = W*in
   wire signed [9:0] m263_88;
   assign m263_88 =10'b0;

   // m263_89 = W*in
   wire signed [9:0] m263_89;
   assign m263_89 ={ {4{in263[5]}} , in263[5:0] };

   // m263_90 = W*in
   wire signed [9:0] m263_90;
   assign m263_90 =10'b0;

   // m263_91 = W*in
   wire signed [9:0] m263_91;
   assign m263_91 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_92 = W*in
   wire signed [9:0] m263_92;
   assign m263_92 =10'b0;

   // m263_93 = W*in
   wire signed [9:0] m263_93;
   assign m263_93 =10'b0;

   // m263_94 = W*in
   wire signed [9:0] m263_94;
   assign m263_94 =10'b0;

   // m263_95 = W*in
   wire signed [9:0] m263_95;
   assign m263_95 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_96 = W*in
   wire signed [9:0] m263_96;
   assign m263_96 ={ {4{in263[5]}} , in263[5:0] };

   // m263_97 = W*in
   wire signed [9:0] m263_97;
   assign m263_97 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_98 = W*in
   wire signed [9:0] m263_98;
   assign m263_98 =10'b0;

   // m263_99 = W*in
   wire signed [9:0] m263_99;
   assign m263_99 =10'b0;

   // m263_100 = W*in
   wire signed [9:0] m263_100;
   assign m263_100 =10'b0;

   // m263_101 = W*in
   wire signed [9:0] m263_101;
   assign m263_101 =10'b0;

   // m263_102 = W*in
   wire signed [9:0] m263_102;
   assign m263_102 =10'b0;

   // m263_103 = W*in
   wire signed [9:0] m263_103;
   assign m263_103 =10'b0;

   // m263_104 = W*in
   wire signed [9:0] m263_104;
   assign m263_104 =10'b0;

   // m263_105 = W*in
   wire signed [9:0] m263_105;
   assign m263_105 =10'b0;

   // m263_106 = W*in
   wire signed [9:0] m263_106;
   assign m263_106 =10'b0;

   // m263_107 = W*in
   wire signed [9:0] m263_107;
   assign m263_107 =10'b0;

   // m263_108 = W*in
   wire signed [9:0] m263_108;
   assign m263_108 ={ {4{in263[5]}} , in263[5:0] };

   // m263_109 = W*in
   wire signed [9:0] m263_109;
   assign m263_109 ={ {4{in263[5]}} , in263[5:0] };

   // m263_110 = W*in
   wire signed [9:0] m263_110;
   assign m263_110 ={ {4{neg263[5]}} , neg263[5:0] };

   // m263_111 = W*in
   wire signed [9:0] m263_111;
   assign m263_111 =10'b0;

   // m263_112 = W*in
   wire signed [9:0] m263_112;
   assign m263_112 =10'b0;

   // m263_113 = W*in
   wire signed [9:0] m263_113;
   assign m263_113 =10'b0;

   // m263_114 = W*in
   wire signed [9:0] m263_114;
   assign m263_114 =10'b0;

   // m263_115 = W*in
   wire signed [9:0] m263_115;
   assign m263_115 ={ {5{in263[5]}} , in263[5:1] };

   // m263_116 = W*in
   wire signed [9:0] m263_116;
   assign m263_116 ={ {4{in263[5]}} , in263[5:0] };

   // m263_117 = W*in
   wire signed [9:0] m263_117;
   assign m263_117 =10'b0;

   // m264_1 = W*in
   wire signed [9:0] m264_1;
   assign m264_1 =10'b0;

   // m264_2 = W*in
   wire signed [9:0] m264_2;
   assign m264_2 =10'b0;

   // m264_3 = W*in
   wire signed [9:0] m264_3;
   assign m264_3 =10'b0;

   // m264_4 = W*in
   wire signed [9:0] m264_4;
   assign m264_4 =10'b0;

   // m264_5 = W*in
   wire signed [9:0] m264_5;
   assign m264_5 =10'b0;

   // m264_6 = W*in
   wire signed [9:0] m264_6;
   assign m264_6 =10'b0;

   // m264_7 = W*in
   wire signed [9:0] m264_7;
   assign m264_7 =10'b0;

   // m264_8 = W*in
   wire signed [9:0] m264_8;
   assign m264_8 =10'b0;

   // m264_9 = W*in
   wire signed [9:0] m264_9;
   assign m264_9 =10'b0;

   // m264_10 = W*in
   wire signed [9:0] m264_10;
   assign m264_10 =10'b0;

   // m264_11 = W*in
   wire signed [9:0] m264_11;
   assign m264_11 =10'b0;

   // m264_12 = W*in
   wire signed [9:0] m264_12;
   assign m264_12 =10'b0;

   // m264_13 = W*in
   wire signed [9:0] m264_13;
   assign m264_13 =10'b0;

   // m264_14 = W*in
   wire signed [9:0] m264_14;
   assign m264_14 =10'b0;

   // m264_15 = W*in
   wire signed [9:0] m264_15;
   assign m264_15 =10'b0;

   // m264_16 = W*in
   wire signed [9:0] m264_16;
   assign m264_16 =10'b0;

   // m264_17 = W*in
   wire signed [9:0] m264_17;
   assign m264_17 ={ {5{in264[5]}} , in264[5:1] };

   // m264_18 = W*in
   wire signed [9:0] m264_18;
   assign m264_18 ={ {5{neg264[5]}} , neg264[5:1] };

   // m264_19 = W*in
   wire signed [9:0] m264_19;
   assign m264_19 ={ {5{in264[5]}} , in264[5:1] };

   // m264_20 = W*in
   wire signed [9:0] m264_20;
   assign m264_20 =10'b0;

   // m264_21 = W*in
   wire signed [9:0] m264_21;
   assign m264_21 =10'b0;

   // m264_22 = W*in
   wire signed [9:0] m264_22;
   assign m264_22 =10'b0;

   // m264_23 = W*in
   wire signed [9:0] m264_23;
   assign m264_23 =10'b0;

   // m264_24 = W*in
   wire signed [9:0] m264_24;
   assign m264_24 =10'b0;

   // m264_25 = W*in
   wire signed [9:0] m264_25;
   assign m264_25 =10'b0;

   // m264_26 = W*in
   wire signed [9:0] m264_26;
   assign m264_26 ={ {5{neg264[5]}} , neg264[5:1] };

   // m264_27 = W*in
   wire signed [9:0] m264_27;
   assign m264_27 =10'b0;

   // m264_28 = W*in
   wire signed [9:0] m264_28;
   assign m264_28 =10'b0;

   // m264_29 = W*in
   wire signed [9:0] m264_29;
   assign m264_29 =10'b0;

   // m264_30 = W*in
   wire signed [9:0] m264_30;
   assign m264_30 =10'b0;

   // m264_31 = W*in
   wire signed [9:0] m264_31;
   assign m264_31 =10'b0;

   // m264_32 = W*in
   wire signed [9:0] m264_32;
   assign m264_32 =10'b0;

   // m264_33 = W*in
   wire signed [9:0] m264_33;
   assign m264_33 =10'b0;

   // m264_34 = W*in
   wire signed [9:0] m264_34;
   assign m264_34 ={ {4{neg264[5]}} , neg264[5:0] };

   // m264_35 = W*in
   wire signed [9:0] m264_35;
   assign m264_35 =10'b0;

   // m264_36 = W*in
   wire signed [9:0] m264_36;
   assign m264_36 =10'b0;

   // m264_37 = W*in
   wire signed [9:0] m264_37;
   assign m264_37 =10'b0;

   // m264_38 = W*in
   wire signed [9:0] m264_38;
   assign m264_38 =10'b0;

   // m264_39 = W*in
   wire signed [9:0] m264_39;
   assign m264_39 =10'b0;

   // m264_40 = W*in
   wire signed [9:0] m264_40;
   assign m264_40 =10'b0;

   // m264_41 = W*in
   wire signed [9:0] m264_41;
   assign m264_41 =10'b0;

   // m264_42 = W*in
   wire signed [9:0] m264_42;
   assign m264_42 =10'b0;

   // m264_43 = W*in
   wire signed [9:0] m264_43;
   assign m264_43 =10'b0;

   // m264_44 = W*in
   wire signed [9:0] m264_44;
   assign m264_44 =10'b0;

   // m264_45 = W*in
   wire signed [9:0] m264_45;
   assign m264_45 =10'b0;

   // m264_46 = W*in
   wire signed [9:0] m264_46;
   assign m264_46 =10'b0;

   // m264_47 = W*in
   wire signed [9:0] m264_47;
   assign m264_47 =10'b0;

   // m264_48 = W*in
   wire signed [9:0] m264_48;
   assign m264_48 =10'b0;

   // m264_49 = W*in
   wire signed [9:0] m264_49;
   assign m264_49 =10'b0;

   // m264_50 = W*in
   wire signed [9:0] m264_50;
   assign m264_50 =10'b0;

   // m264_51 = W*in
   wire signed [9:0] m264_51;
   assign m264_51 =10'b0;

   // m264_52 = W*in
   wire signed [9:0] m264_52;
   assign m264_52 =10'b0;

   // m264_53 = W*in
   wire signed [9:0] m264_53;
   assign m264_53 =10'b0;

   // m264_54 = W*in
   wire signed [9:0] m264_54;
   assign m264_54 =10'b0;

   // m264_55 = W*in
   wire signed [9:0] m264_55;
   assign m264_55 =10'b0;

   // m264_56 = W*in
   wire signed [9:0] m264_56;
   assign m264_56 =10'b0;

   // m264_57 = W*in
   wire signed [9:0] m264_57;
   assign m264_57 =10'b0;

   // m264_58 = W*in
   wire signed [9:0] m264_58;
   assign m264_58 =10'b0;

   // m264_59 = W*in
   wire signed [9:0] m264_59;
   assign m264_59 =10'b0;

   // m264_60 = W*in
   wire signed [9:0] m264_60;
   assign m264_60 =10'b0;

   // m264_61 = W*in
   wire signed [9:0] m264_61;
   assign m264_61 =10'b0;

   // m264_62 = W*in
   wire signed [9:0] m264_62;
   assign m264_62 =10'b0;

   // m264_63 = W*in
   wire signed [9:0] m264_63;
   assign m264_63 =10'b0;

   // m264_64 = W*in
   wire signed [9:0] m264_64;
   assign m264_64 ={ {5{neg264[5]}} , neg264[5:1] };

   // m264_65 = W*in
   wire signed [9:0] m264_65;
   assign m264_65 =10'b0;

   // m264_66 = W*in
   wire signed [9:0] m264_66;
   assign m264_66 ={ {5{in264[5]}} , in264[5:1] };

   // m264_67 = W*in
   wire signed [9:0] m264_67;
   assign m264_67 ={ {4{in264[5]}} , in264[5:0] };

   // m264_68 = W*in
   wire signed [9:0] m264_68;
   assign m264_68 =10'b0;

   // m264_69 = W*in
   wire signed [9:0] m264_69;
   assign m264_69 =10'b0;

   // m264_70 = W*in
   wire signed [9:0] m264_70;
   assign m264_70 =10'b0;

   // m264_71 = W*in
   wire signed [9:0] m264_71;
   assign m264_71 =10'b0;

   // m264_72 = W*in
   wire signed [9:0] m264_72;
   assign m264_72 =10'b0;

   // m264_73 = W*in
   wire signed [9:0] m264_73;
   assign m264_73 =10'b0;

   // m264_74 = W*in
   wire signed [9:0] m264_74;
   assign m264_74 =10'b0;

   // m264_75 = W*in
   wire signed [9:0] m264_75;
   assign m264_75 =10'b0;

   // m264_76 = W*in
   wire signed [9:0] m264_76;
   assign m264_76 =10'b0;

   // m264_77 = W*in
   wire signed [9:0] m264_77;
   assign m264_77 =10'b0;

   // m264_78 = W*in
   wire signed [9:0] m264_78;
   assign m264_78 ={ {5{neg264[5]}} , neg264[5:1] };

   // m264_79 = W*in
   wire signed [9:0] m264_79;
   assign m264_79 =10'b0;

   // m264_80 = W*in
   wire signed [9:0] m264_80;
   assign m264_80 =10'b0;

   // m264_81 = W*in
   wire signed [9:0] m264_81;
   assign m264_81 ={ {5{neg264[5]}} , neg264[5:1] };

   // m264_82 = W*in
   wire signed [9:0] m264_82;
   assign m264_82 =10'b0;

   // m264_83 = W*in
   wire signed [9:0] m264_83;
   assign m264_83 =10'b0;

   // m264_84 = W*in
   wire signed [9:0] m264_84;
   assign m264_84 =10'b0;

   // m264_85 = W*in
   wire signed [9:0] m264_85;
   assign m264_85 =10'b0;

   // m264_86 = W*in
   wire signed [9:0] m264_86;
   assign m264_86 =10'b0;

   // m264_87 = W*in
   wire signed [9:0] m264_87;
   assign m264_87 =10'b0;

   // m264_88 = W*in
   wire signed [9:0] m264_88;
   assign m264_88 =10'b0;

   // m264_89 = W*in
   wire signed [9:0] m264_89;
   assign m264_89 =10'b0;

   // m264_90 = W*in
   wire signed [9:0] m264_90;
   assign m264_90 =10'b0;

   // m264_91 = W*in
   wire signed [9:0] m264_91;
   assign m264_91 =10'b0;

   // m264_92 = W*in
   wire signed [9:0] m264_92;
   assign m264_92 =10'b0;

   // m264_93 = W*in
   wire signed [9:0] m264_93;
   assign m264_93 =10'b0;

   // m264_94 = W*in
   wire signed [9:0] m264_94;
   assign m264_94 =10'b0;

   // m264_95 = W*in
   wire signed [9:0] m264_95;
   assign m264_95 =10'b0;

   // m264_96 = W*in
   wire signed [9:0] m264_96;
   assign m264_96 =10'b0;

   // m264_97 = W*in
   wire signed [9:0] m264_97;
   assign m264_97 ={ {4{in264[5]}} , in264[5:0] };

   // m264_98 = W*in
   wire signed [9:0] m264_98;
   assign m264_98 =10'b0;

   // m264_99 = W*in
   wire signed [9:0] m264_99;
   assign m264_99 =10'b0;

   // m264_100 = W*in
   wire signed [9:0] m264_100;
   assign m264_100 =10'b0;

   // m264_101 = W*in
   wire signed [9:0] m264_101;
   assign m264_101 =10'b0;

   // m264_102 = W*in
   wire signed [9:0] m264_102;
   assign m264_102 =10'b0;

   // m264_103 = W*in
   wire signed [9:0] m264_103;
   assign m264_103 =10'b0;

   // m264_104 = W*in
   wire signed [9:0] m264_104;
   assign m264_104 =10'b0;

   // m264_105 = W*in
   wire signed [9:0] m264_105;
   assign m264_105 =10'b0;

   // m264_106 = W*in
   wire signed [9:0] m264_106;
   assign m264_106 =10'b0;

   // m264_107 = W*in
   wire signed [9:0] m264_107;
   assign m264_107 =10'b0;

   // m264_108 = W*in
   wire signed [9:0] m264_108;
   assign m264_108 =10'b0;

   // m264_109 = W*in
   wire signed [9:0] m264_109;
   assign m264_109 ={ {5{neg264[5]}} , neg264[5:1] };

   // m264_110 = W*in
   wire signed [9:0] m264_110;
   assign m264_110 =10'b0;

   // m264_111 = W*in
   wire signed [9:0] m264_111;
   assign m264_111 =10'b0;

   // m264_112 = W*in
   wire signed [9:0] m264_112;
   assign m264_112 =10'b0;

   // m264_113 = W*in
   wire signed [9:0] m264_113;
   assign m264_113 =10'b0;

   // m264_114 = W*in
   wire signed [9:0] m264_114;
   assign m264_114 =10'b0;

   // m264_115 = W*in
   wire signed [9:0] m264_115;
   assign m264_115 =10'b0;

   // m264_116 = W*in
   wire signed [9:0] m264_116;
   assign m264_116 =10'b0;

   // m264_117 = W*in
   wire signed [9:0] m264_117;
   assign m264_117 =10'b0;

   // m265_1 = W*in
   wire signed [9:0] m265_1;
   assign m265_1 =10'b0;

   // m265_2 = W*in
   wire signed [9:0] m265_2;
   assign m265_2 =10'b0;

   // m265_3 = W*in
   wire signed [9:0] m265_3;
   assign m265_3 =10'b0;

   // m265_4 = W*in
   wire signed [9:0] m265_4;
   assign m265_4 =10'b0;

   // m265_5 = W*in
   wire signed [9:0] m265_5;
   assign m265_5 =10'b0;

   // m265_6 = W*in
   wire signed [9:0] m265_6;
   assign m265_6 =10'b0;

   // m265_7 = W*in
   wire signed [9:0] m265_7;
   assign m265_7 =10'b0;

   // m265_8 = W*in
   wire signed [9:0] m265_8;
   assign m265_8 ={ {4{in265[5]}} , in265[5:0] };

   // m265_9 = W*in
   wire signed [9:0] m265_9;
   assign m265_9 =10'b0;

   // m265_10 = W*in
   wire signed [9:0] m265_10;
   assign m265_10 =10'b0;

   // m265_11 = W*in
   wire signed [9:0] m265_11;
   assign m265_11 =10'b0;

   // m265_12 = W*in
   wire signed [9:0] m265_12;
   assign m265_12 =10'b0;

   // m265_13 = W*in
   wire signed [9:0] m265_13;
   assign m265_13 =10'b0;

   // m265_14 = W*in
   wire signed [9:0] m265_14;
   assign m265_14 =10'b0;

   // m265_15 = W*in
   wire signed [9:0] m265_15;
   assign m265_15 =10'b0;

   // m265_16 = W*in
   wire signed [9:0] m265_16;
   assign m265_16 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_17 = W*in
   wire signed [9:0] m265_17;
   assign m265_17 ={ {3{in265[5]}} , in265 , {1{1'b0}} };

   // m265_18 = W*in
   wire signed [9:0] m265_18;
   assign m265_18 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_19 = W*in
   wire signed [9:0] m265_19;
   assign m265_19 ={ {4{in265[5]}} , in265[5:0] };

   // m265_20 = W*in
   wire signed [9:0] m265_20;
   assign m265_20 =10'b0;

   // m265_21 = W*in
   wire signed [9:0] m265_21;
   assign m265_21 =10'b0;

   // m265_22 = W*in
   wire signed [9:0] m265_22;
   assign m265_22 =10'b0;

   // m265_23 = W*in
   wire signed [9:0] m265_23;
   assign m265_23 =10'b0;

   // m265_24 = W*in
   wire signed [9:0] m265_24;
   assign m265_24 =10'b0;

   // m265_25 = W*in
   wire signed [9:0] m265_25;
   assign m265_25 =10'b0;

   // m265_26 = W*in
   wire signed [9:0] m265_26;
   assign m265_26 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_27 = W*in
   wire signed [9:0] m265_27;
   assign m265_27 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_28 = W*in
   wire signed [9:0] m265_28;
   assign m265_28 =10'b0;

   // m265_29 = W*in
   wire signed [9:0] m265_29;
   assign m265_29 =10'b0;

   // m265_30 = W*in
   wire signed [9:0] m265_30;
   assign m265_30 =10'b0;

   // m265_31 = W*in
   wire signed [9:0] m265_31;
   assign m265_31 =10'b0;

   // m265_32 = W*in
   wire signed [9:0] m265_32;
   assign m265_32 =10'b0;

   // m265_33 = W*in
   wire signed [9:0] m265_33;
   assign m265_33 =10'b0;

   // m265_34 = W*in
   wire signed [9:0] m265_34;
   assign m265_34 =10'b0;

   // m265_35 = W*in
   wire signed [9:0] m265_35;
   assign m265_35 =10'b0;

   // m265_36 = W*in
   wire signed [9:0] m265_36;
   assign m265_36 ={ {4{in265[5]}} , in265[5:0] };

   // m265_37 = W*in
   wire signed [9:0] m265_37;
   assign m265_37 =10'b0;

   // m265_38 = W*in
   wire signed [9:0] m265_38;
   assign m265_38 =10'b0;

   // m265_39 = W*in
   wire signed [9:0] m265_39;
   assign m265_39 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_40 = W*in
   wire signed [9:0] m265_40;
   assign m265_40 =10'b0;

   // m265_41 = W*in
   wire signed [9:0] m265_41;
   assign m265_41 =10'b0;

   // m265_42 = W*in
   wire signed [9:0] m265_42;
   assign m265_42 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_43 = W*in
   wire signed [9:0] m265_43;
   assign m265_43 =10'b0;

   // m265_44 = W*in
   wire signed [9:0] m265_44;
   assign m265_44 ={ {4{in265[5]}} , in265[5:0] };

   // m265_45 = W*in
   wire signed [9:0] m265_45;
   assign m265_45 =10'b0;

   // m265_46 = W*in
   wire signed [9:0] m265_46;
   assign m265_46 =10'b0;

   // m265_47 = W*in
   wire signed [9:0] m265_47;
   assign m265_47 =10'b0;

   // m265_48 = W*in
   wire signed [9:0] m265_48;
   assign m265_48 =10'b0;

   // m265_49 = W*in
   wire signed [9:0] m265_49;
   assign m265_49 ={ {4{in265[5]}} , in265[5:0] };

   // m265_50 = W*in
   wire signed [9:0] m265_50;
   assign m265_50 =10'b0;

   // m265_51 = W*in
   wire signed [9:0] m265_51;
   assign m265_51 ={ {4{in265[5]}} , in265[5:0] };

   // m265_52 = W*in
   wire signed [9:0] m265_52;
   assign m265_52 =10'b0;

   // m265_53 = W*in
   wire signed [9:0] m265_53;
   assign m265_53 ={ {3{in265[5]}} , in265 , {1{1'b0}} };

   // m265_54 = W*in
   wire signed [9:0] m265_54;
   assign m265_54 ={ {4{in265[5]}} , in265[5:0] };

   // m265_55 = W*in
   wire signed [9:0] m265_55;
   assign m265_55 =10'b0;

   // m265_56 = W*in
   wire signed [9:0] m265_56;
   assign m265_56 =10'b0;

   // m265_57 = W*in
   wire signed [9:0] m265_57;
   assign m265_57 =10'b0;

   // m265_58 = W*in
   wire signed [9:0] m265_58;
   assign m265_58 =10'b0;

   // m265_59 = W*in
   wire signed [9:0] m265_59;
   assign m265_59 =10'b0;

   // m265_60 = W*in
   wire signed [9:0] m265_60;
   assign m265_60 =10'b0;

   // m265_61 = W*in
   wire signed [9:0] m265_61;
   assign m265_61 =10'b0;

   // m265_62 = W*in
   wire signed [9:0] m265_62;
   assign m265_62 =10'b0;

   // m265_63 = W*in
   wire signed [9:0] m265_63;
   assign m265_63 =10'b0;

   // m265_64 = W*in
   wire signed [9:0] m265_64;
   assign m265_64 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_65 = W*in
   wire signed [9:0] m265_65;
   assign m265_65 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_66 = W*in
   wire signed [9:0] m265_66;
   assign m265_66 =10'b0;

   // m265_67 = W*in
   wire signed [9:0] m265_67;
   assign m265_67 ={ {4{in265[5]}} , in265[5:0] };

   // m265_68 = W*in
   wire signed [9:0] m265_68;
   assign m265_68 =10'b0;

   // m265_69 = W*in
   wire signed [9:0] m265_69;
   assign m265_69 =10'b0;

   // m265_70 = W*in
   wire signed [9:0] m265_70;
   assign m265_70 =10'b0;

   // m265_71 = W*in
   wire signed [9:0] m265_71;
   assign m265_71 =10'b0;

   // m265_72 = W*in
   wire signed [9:0] m265_72;
   assign m265_72 ={ {5{in265[5]}} , in265[5:1] };

   // m265_73 = W*in
   wire signed [9:0] m265_73;
   assign m265_73 =10'b0;

   // m265_74 = W*in
   wire signed [9:0] m265_74;
   assign m265_74 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_75 = W*in
   wire signed [9:0] m265_75;
   assign m265_75 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_76 = W*in
   wire signed [9:0] m265_76;
   assign m265_76 =10'b0;

   // m265_77 = W*in
   wire signed [9:0] m265_77;
   assign m265_77 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_78 = W*in
   wire signed [9:0] m265_78;
   assign m265_78 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_79 = W*in
   wire signed [9:0] m265_79;
   assign m265_79 =10'b0;

   // m265_80 = W*in
   wire signed [9:0] m265_80;
   assign m265_80 =10'b0;

   // m265_81 = W*in
   wire signed [9:0] m265_81;
   assign m265_81 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_82 = W*in
   wire signed [9:0] m265_82;
   assign m265_82 =10'b0;

   // m265_83 = W*in
   wire signed [9:0] m265_83;
   assign m265_83 =10'b0;

   // m265_84 = W*in
   wire signed [9:0] m265_84;
   assign m265_84 =10'b0;

   // m265_85 = W*in
   wire signed [9:0] m265_85;
   assign m265_85 =10'b0;

   // m265_86 = W*in
   wire signed [9:0] m265_86;
   assign m265_86 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_87 = W*in
   wire signed [9:0] m265_87;
   assign m265_87 =10'b0;

   // m265_88 = W*in
   wire signed [9:0] m265_88;
   assign m265_88 =10'b0;

   // m265_89 = W*in
   wire signed [9:0] m265_89;
   assign m265_89 =10'b0;

   // m265_90 = W*in
   wire signed [9:0] m265_90;
   assign m265_90 =10'b0;

   // m265_91 = W*in
   wire signed [9:0] m265_91;
   assign m265_91 =10'b0;

   // m265_92 = W*in
   wire signed [9:0] m265_92;
   assign m265_92 =10'b0;

   // m265_93 = W*in
   wire signed [9:0] m265_93;
   assign m265_93 =10'b0;

   // m265_94 = W*in
   wire signed [9:0] m265_94;
   assign m265_94 =10'b0;

   // m265_95 = W*in
   wire signed [9:0] m265_95;
   assign m265_95 ={ {5{in265[5]}} , in265[5:1] };

   // m265_96 = W*in
   wire signed [9:0] m265_96;
   assign m265_96 =10'b0;

   // m265_97 = W*in
   wire signed [9:0] m265_97;
   assign m265_97 =10'b0;

   // m265_98 = W*in
   wire signed [9:0] m265_98;
   assign m265_98 =10'b0;

   // m265_99 = W*in
   wire signed [9:0] m265_99;
   assign m265_99 =10'b0;

   // m265_100 = W*in
   wire signed [9:0] m265_100;
   assign m265_100 =10'b0;

   // m265_101 = W*in
   wire signed [9:0] m265_101;
   assign m265_101 =10'b0;

   // m265_102 = W*in
   wire signed [9:0] m265_102;
   assign m265_102 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_103 = W*in
   wire signed [9:0] m265_103;
   assign m265_103 =10'b0;

   // m265_104 = W*in
   wire signed [9:0] m265_104;
   assign m265_104 =10'b0;

   // m265_105 = W*in
   wire signed [9:0] m265_105;
   assign m265_105 =10'b0;

   // m265_106 = W*in
   wire signed [9:0] m265_106;
   assign m265_106 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_107 = W*in
   wire signed [9:0] m265_107;
   assign m265_107 ={ {4{in265[5]}} , in265[5:0] };

   // m265_108 = W*in
   wire signed [9:0] m265_108;
   assign m265_108 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_109 = W*in
   wire signed [9:0] m265_109;
   assign m265_109 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_110 = W*in
   wire signed [9:0] m265_110;
   assign m265_110 =10'b0;

   // m265_111 = W*in
   wire signed [9:0] m265_111;
   assign m265_111 =10'b0;

   // m265_112 = W*in
   wire signed [9:0] m265_112;
   assign m265_112 ={ {4{neg265[5]}} , neg265[5:0] };

   // m265_113 = W*in
   wire signed [9:0] m265_113;
   assign m265_113 =10'b0;

   // m265_114 = W*in
   wire signed [9:0] m265_114;
   assign m265_114 ={ {5{neg265[5]}} , neg265[5:1] };

   // m265_115 = W*in
   wire signed [9:0] m265_115;
   assign m265_115 =10'b0;

   // m265_116 = W*in
   wire signed [9:0] m265_116;
   assign m265_116 =10'b0;

   // m265_117 = W*in
   wire signed [9:0] m265_117;
   assign m265_117 =10'b0;

   // m266_1 = W*in
   wire signed [9:0] m266_1;
   assign m266_1 =10'b0;

   // m266_2 = W*in
   wire signed [9:0] m266_2;
   assign m266_2 =10'b0;

   // m266_3 = W*in
   wire signed [9:0] m266_3;
   assign m266_3 =10'b0;

   // m266_4 = W*in
   wire signed [9:0] m266_4;
   assign m266_4 =10'b0;

   // m266_5 = W*in
   wire signed [9:0] m266_5;
   assign m266_5 =10'b0;

   // m266_6 = W*in
   wire signed [9:0] m266_6;
   assign m266_6 =10'b0;

   // m266_7 = W*in
   wire signed [9:0] m266_7;
   assign m266_7 =10'b0;

   // m266_8 = W*in
   wire signed [9:0] m266_8;
   assign m266_8 =10'b0;

   // m266_9 = W*in
   wire signed [9:0] m266_9;
   assign m266_9 =10'b0;

   // m266_10 = W*in
   wire signed [9:0] m266_10;
   assign m266_10 =10'b0;

   // m266_11 = W*in
   wire signed [9:0] m266_11;
   assign m266_11 =10'b0;

   // m266_12 = W*in
   wire signed [9:0] m266_12;
   assign m266_12 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_13 = W*in
   wire signed [9:0] m266_13;
   assign m266_13 =10'b0;

   // m266_14 = W*in
   wire signed [9:0] m266_14;
   assign m266_14 =10'b0;

   // m266_15 = W*in
   wire signed [9:0] m266_15;
   assign m266_15 =10'b0;

   // m266_16 = W*in
   wire signed [9:0] m266_16;
   assign m266_16 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_17 = W*in
   wire signed [9:0] m266_17;
   assign m266_17 =10'b0;

   // m266_18 = W*in
   wire signed [9:0] m266_18;
   assign m266_18 ={ {5{neg266[5]}} , neg266[5:1] };

   // m266_19 = W*in
   wire signed [9:0] m266_19;
   assign m266_19 ={ {5{in266[5]}} , in266[5:1] };

   // m266_20 = W*in
   wire signed [9:0] m266_20;
   assign m266_20 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_21 = W*in
   wire signed [9:0] m266_21;
   assign m266_21 ={ {5{in266[5]}} , in266[5:1] };

   // m266_22 = W*in
   wire signed [9:0] m266_22;
   assign m266_22 =10'b0;

   // m266_23 = W*in
   wire signed [9:0] m266_23;
   assign m266_23 =10'b0;

   // m266_24 = W*in
   wire signed [9:0] m266_24;
   assign m266_24 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_25 = W*in
   wire signed [9:0] m266_25;
   assign m266_25 =10'b0;

   // m266_26 = W*in
   wire signed [9:0] m266_26;
   assign m266_26 =10'b0;

   // m266_27 = W*in
   wire signed [9:0] m266_27;
   assign m266_27 =10'b0;

   // m266_28 = W*in
   wire signed [9:0] m266_28;
   assign m266_28 =10'b0;

   // m266_29 = W*in
   wire signed [9:0] m266_29;
   assign m266_29 =10'b0;

   // m266_30 = W*in
   wire signed [9:0] m266_30;
   assign m266_30 =10'b0;

   // m266_31 = W*in
   wire signed [9:0] m266_31;
   assign m266_31 =10'b0;

   // m266_32 = W*in
   wire signed [9:0] m266_32;
   assign m266_32 =10'b0;

   // m266_33 = W*in
   wire signed [9:0] m266_33;
   assign m266_33 =10'b0;

   // m266_34 = W*in
   wire signed [9:0] m266_34;
   assign m266_34 =10'b0;

   // m266_35 = W*in
   wire signed [9:0] m266_35;
   assign m266_35 =10'b0;

   // m266_36 = W*in
   wire signed [9:0] m266_36;
   assign m266_36 ={ {5{in266[5]}} , in266[5:1] };

   // m266_37 = W*in
   wire signed [9:0] m266_37;
   assign m266_37 =10'b0;

   // m266_38 = W*in
   wire signed [9:0] m266_38;
   assign m266_38 =10'b0;

   // m266_39 = W*in
   wire signed [9:0] m266_39;
   assign m266_39 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_40 = W*in
   wire signed [9:0] m266_40;
   assign m266_40 =10'b0;

   // m266_41 = W*in
   wire signed [9:0] m266_41;
   assign m266_41 =10'b0;

   // m266_42 = W*in
   wire signed [9:0] m266_42;
   assign m266_42 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_43 = W*in
   wire signed [9:0] m266_43;
   assign m266_43 ={ {4{in266[5]}} , in266[5:0] };

   // m266_44 = W*in
   wire signed [9:0] m266_44;
   assign m266_44 ={ {4{in266[5]}} , in266[5:0] };

   // m266_45 = W*in
   wire signed [9:0] m266_45;
   assign m266_45 =10'b0;

   // m266_46 = W*in
   wire signed [9:0] m266_46;
   assign m266_46 =10'b0;

   // m266_47 = W*in
   wire signed [9:0] m266_47;
   assign m266_47 =10'b0;

   // m266_48 = W*in
   wire signed [9:0] m266_48;
   assign m266_48 =10'b0;

   // m266_49 = W*in
   wire signed [9:0] m266_49;
   assign m266_49 =10'b0;

   // m266_50 = W*in
   wire signed [9:0] m266_50;
   assign m266_50 ={ {4{in266[5]}} , in266[5:0] };

   // m266_51 = W*in
   wire signed [9:0] m266_51;
   assign m266_51 =10'b0;

   // m266_52 = W*in
   wire signed [9:0] m266_52;
   assign m266_52 =10'b0;

   // m266_53 = W*in
   wire signed [9:0] m266_53;
   assign m266_53 ={ {4{in266[5]}} , in266[5:0] };

   // m266_54 = W*in
   wire signed [9:0] m266_54;
   assign m266_54 ={ {4{in266[5]}} , in266[5:0] };

   // m266_55 = W*in
   wire signed [9:0] m266_55;
   assign m266_55 =10'b0;

   // m266_56 = W*in
   wire signed [9:0] m266_56;
   assign m266_56 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_57 = W*in
   wire signed [9:0] m266_57;
   assign m266_57 =10'b0;

   // m266_58 = W*in
   wire signed [9:0] m266_58;
   assign m266_58 =10'b0;

   // m266_59 = W*in
   wire signed [9:0] m266_59;
   assign m266_59 =10'b0;

   // m266_60 = W*in
   wire signed [9:0] m266_60;
   assign m266_60 =10'b0;

   // m266_61 = W*in
   wire signed [9:0] m266_61;
   assign m266_61 =10'b0;

   // m266_62 = W*in
   wire signed [9:0] m266_62;
   assign m266_62 =10'b0;

   // m266_63 = W*in
   wire signed [9:0] m266_63;
   assign m266_63 =10'b0;

   // m266_64 = W*in
   wire signed [9:0] m266_64;
   assign m266_64 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_65 = W*in
   wire signed [9:0] m266_65;
   assign m266_65 =10'b0;

   // m266_66 = W*in
   wire signed [9:0] m266_66;
   assign m266_66 =10'b0;

   // m266_67 = W*in
   wire signed [9:0] m266_67;
   assign m266_67 ={ {4{in266[5]}} , in266[5:0] };

   // m266_68 = W*in
   wire signed [9:0] m266_68;
   assign m266_68 =10'b0;

   // m266_69 = W*in
   wire signed [9:0] m266_69;
   assign m266_69 ={ {5{in266[5]}} , in266[5:1] };

   // m266_70 = W*in
   wire signed [9:0] m266_70;
   assign m266_70 =10'b0;

   // m266_71 = W*in
   wire signed [9:0] m266_71;
   assign m266_71 =10'b0;

   // m266_72 = W*in
   wire signed [9:0] m266_72;
   assign m266_72 ={ {4{in266[5]}} , in266[5:0] };

   // m266_73 = W*in
   wire signed [9:0] m266_73;
   assign m266_73 =10'b0;

   // m266_74 = W*in
   wire signed [9:0] m266_74;
   assign m266_74 =10'b0;

   // m266_75 = W*in
   wire signed [9:0] m266_75;
   assign m266_75 =10'b0;

   // m266_76 = W*in
   wire signed [9:0] m266_76;
   assign m266_76 =10'b0;

   // m266_77 = W*in
   wire signed [9:0] m266_77;
   assign m266_77 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_78 = W*in
   wire signed [9:0] m266_78;
   assign m266_78 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_79 = W*in
   wire signed [9:0] m266_79;
   assign m266_79 =10'b0;

   // m266_80 = W*in
   wire signed [9:0] m266_80;
   assign m266_80 =10'b0;

   // m266_81 = W*in
   wire signed [9:0] m266_81;
   assign m266_81 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_82 = W*in
   wire signed [9:0] m266_82;
   assign m266_82 =10'b0;

   // m266_83 = W*in
   wire signed [9:0] m266_83;
   assign m266_83 ={ {5{neg266[5]}} , neg266[5:1] };

   // m266_84 = W*in
   wire signed [9:0] m266_84;
   assign m266_84 ={ {4{in266[5]}} , in266[5:0] };

   // m266_85 = W*in
   wire signed [9:0] m266_85;
   assign m266_85 =10'b0;

   // m266_86 = W*in
   wire signed [9:0] m266_86;
   assign m266_86 =10'b0;

   // m266_87 = W*in
   wire signed [9:0] m266_87;
   assign m266_87 =10'b0;

   // m266_88 = W*in
   wire signed [9:0] m266_88;
   assign m266_88 =10'b0;

   // m266_89 = W*in
   wire signed [9:0] m266_89;
   assign m266_89 =10'b0;

   // m266_90 = W*in
   wire signed [9:0] m266_90;
   assign m266_90 =10'b0;

   // m266_91 = W*in
   wire signed [9:0] m266_91;
   assign m266_91 =10'b0;

   // m266_92 = W*in
   wire signed [9:0] m266_92;
   assign m266_92 =10'b0;

   // m266_93 = W*in
   wire signed [9:0] m266_93;
   assign m266_93 =10'b0;

   // m266_94 = W*in
   wire signed [9:0] m266_94;
   assign m266_94 =10'b0;

   // m266_95 = W*in
   wire signed [9:0] m266_95;
   assign m266_95 =10'b0;

   // m266_96 = W*in
   wire signed [9:0] m266_96;
   assign m266_96 =10'b0;

   // m266_97 = W*in
   wire signed [9:0] m266_97;
   assign m266_97 =10'b0;

   // m266_98 = W*in
   wire signed [9:0] m266_98;
   assign m266_98 =10'b0;

   // m266_99 = W*in
   wire signed [9:0] m266_99;
   assign m266_99 =10'b0;

   // m266_100 = W*in
   wire signed [9:0] m266_100;
   assign m266_100 =10'b0;

   // m266_101 = W*in
   wire signed [9:0] m266_101;
   assign m266_101 =10'b0;

   // m266_102 = W*in
   wire signed [9:0] m266_102;
   assign m266_102 =10'b0;

   // m266_103 = W*in
   wire signed [9:0] m266_103;
   assign m266_103 =10'b0;

   // m266_104 = W*in
   wire signed [9:0] m266_104;
   assign m266_104 =10'b0;

   // m266_105 = W*in
   wire signed [9:0] m266_105;
   assign m266_105 =10'b0;

   // m266_106 = W*in
   wire signed [9:0] m266_106;
   assign m266_106 ={ {5{neg266[5]}} , neg266[5:1] };

   // m266_107 = W*in
   wire signed [9:0] m266_107;
   assign m266_107 =10'b0;

   // m266_108 = W*in
   wire signed [9:0] m266_108;
   assign m266_108 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_109 = W*in
   wire signed [9:0] m266_109;
   assign m266_109 =10'b0;

   // m266_110 = W*in
   wire signed [9:0] m266_110;
   assign m266_110 =10'b0;

   // m266_111 = W*in
   wire signed [9:0] m266_111;
   assign m266_111 =10'b0;

   // m266_112 = W*in
   wire signed [9:0] m266_112;
   assign m266_112 =10'b0;

   // m266_113 = W*in
   wire signed [9:0] m266_113;
   assign m266_113 =10'b0;

   // m266_114 = W*in
   wire signed [9:0] m266_114;
   assign m266_114 =10'b0;

   // m266_115 = W*in
   wire signed [9:0] m266_115;
   assign m266_115 ={ {5{neg266[5]}} , neg266[5:1] };

   // m266_116 = W*in
   wire signed [9:0] m266_116;
   assign m266_116 ={ {4{neg266[5]}} , neg266[5:0] };

   // m266_117 = W*in
   wire signed [9:0] m266_117;
   assign m266_117 =10'b0;

   // m267_1 = W*in
   wire signed [9:0] m267_1;
   assign m267_1 =10'b0;

   // m267_2 = W*in
   wire signed [9:0] m267_2;
   assign m267_2 =10'b0;

   // m267_3 = W*in
   wire signed [9:0] m267_3;
   assign m267_3 =10'b0;

   // m267_4 = W*in
   wire signed [9:0] m267_4;
   assign m267_4 =10'b0;

   // m267_5 = W*in
   wire signed [9:0] m267_5;
   assign m267_5 =10'b0;

   // m267_6 = W*in
   wire signed [9:0] m267_6;
   assign m267_6 =10'b0;

   // m267_7 = W*in
   wire signed [9:0] m267_7;
   assign m267_7 =10'b0;

   // m267_8 = W*in
   wire signed [9:0] m267_8;
   assign m267_8 =10'b0;

   // m267_9 = W*in
   wire signed [9:0] m267_9;
   assign m267_9 =10'b0;

   // m267_10 = W*in
   wire signed [9:0] m267_10;
   assign m267_10 =10'b0;

   // m267_11 = W*in
   wire signed [9:0] m267_11;
   assign m267_11 =10'b0;

   // m267_12 = W*in
   wire signed [9:0] m267_12;
   assign m267_12 =10'b0;

   // m267_13 = W*in
   wire signed [9:0] m267_13;
   assign m267_13 =10'b0;

   // m267_14 = W*in
   wire signed [9:0] m267_14;
   assign m267_14 =10'b0;

   // m267_15 = W*in
   wire signed [9:0] m267_15;
   assign m267_15 =10'b0;

   // m267_16 = W*in
   wire signed [9:0] m267_16;
   assign m267_16 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_17 = W*in
   wire signed [9:0] m267_17;
   assign m267_17 =10'b0;

   // m267_18 = W*in
   wire signed [9:0] m267_18;
   assign m267_18 =10'b0;

   // m267_19 = W*in
   wire signed [9:0] m267_19;
   assign m267_19 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_20 = W*in
   wire signed [9:0] m267_20;
   assign m267_20 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_21 = W*in
   wire signed [9:0] m267_21;
   assign m267_21 ={ {5{in267[5]}} , in267[5:1] };

   // m267_22 = W*in
   wire signed [9:0] m267_22;
   assign m267_22 =10'b0;

   // m267_23 = W*in
   wire signed [9:0] m267_23;
   assign m267_23 =10'b0;

   // m267_24 = W*in
   wire signed [9:0] m267_24;
   assign m267_24 =10'b0;

   // m267_25 = W*in
   wire signed [9:0] m267_25;
   assign m267_25 ={ {4{neg267[5]}} , neg267[5:0] };

   // m267_26 = W*in
   wire signed [9:0] m267_26;
   assign m267_26 =10'b0;

   // m267_27 = W*in
   wire signed [9:0] m267_27;
   assign m267_27 =10'b0;

   // m267_28 = W*in
   wire signed [9:0] m267_28;
   assign m267_28 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_29 = W*in
   wire signed [9:0] m267_29;
   assign m267_29 =10'b0;

   // m267_30 = W*in
   wire signed [9:0] m267_30;
   assign m267_30 =10'b0;

   // m267_31 = W*in
   wire signed [9:0] m267_31;
   assign m267_31 =10'b0;

   // m267_32 = W*in
   wire signed [9:0] m267_32;
   assign m267_32 =10'b0;

   // m267_33 = W*in
   wire signed [9:0] m267_33;
   assign m267_33 =10'b0;

   // m267_34 = W*in
   wire signed [9:0] m267_34;
   assign m267_34 =10'b0;

   // m267_35 = W*in
   wire signed [9:0] m267_35;
   assign m267_35 =10'b0;

   // m267_36 = W*in
   wire signed [9:0] m267_36;
   assign m267_36 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_37 = W*in
   wire signed [9:0] m267_37;
   assign m267_37 =10'b0;

   // m267_38 = W*in
   wire signed [9:0] m267_38;
   assign m267_38 =10'b0;

   // m267_39 = W*in
   wire signed [9:0] m267_39;
   assign m267_39 =10'b0;

   // m267_40 = W*in
   wire signed [9:0] m267_40;
   assign m267_40 =10'b0;

   // m267_41 = W*in
   wire signed [9:0] m267_41;
   assign m267_41 =10'b0;

   // m267_42 = W*in
   wire signed [9:0] m267_42;
   assign m267_42 =10'b0;

   // m267_43 = W*in
   wire signed [9:0] m267_43;
   assign m267_43 =10'b0;

   // m267_44 = W*in
   wire signed [9:0] m267_44;
   assign m267_44 =10'b0;

   // m267_45 = W*in
   wire signed [9:0] m267_45;
   assign m267_45 =10'b0;

   // m267_46 = W*in
   wire signed [9:0] m267_46;
   assign m267_46 =10'b0;

   // m267_47 = W*in
   wire signed [9:0] m267_47;
   assign m267_47 =10'b0;

   // m267_48 = W*in
   wire signed [9:0] m267_48;
   assign m267_48 =10'b0;

   // m267_49 = W*in
   wire signed [9:0] m267_49;
   assign m267_49 =10'b0;

   // m267_50 = W*in
   wire signed [9:0] m267_50;
   assign m267_50 =10'b0;

   // m267_51 = W*in
   wire signed [9:0] m267_51;
   assign m267_51 =10'b0;

   // m267_52 = W*in
   wire signed [9:0] m267_52;
   assign m267_52 =10'b0;

   // m267_53 = W*in
   wire signed [9:0] m267_53;
   assign m267_53 =10'b0;

   // m267_54 = W*in
   wire signed [9:0] m267_54;
   assign m267_54 =10'b0;

   // m267_55 = W*in
   wire signed [9:0] m267_55;
   assign m267_55 =10'b0;

   // m267_56 = W*in
   wire signed [9:0] m267_56;
   assign m267_56 =10'b0;

   // m267_57 = W*in
   wire signed [9:0] m267_57;
   assign m267_57 =10'b0;

   // m267_58 = W*in
   wire signed [9:0] m267_58;
   assign m267_58 =10'b0;

   // m267_59 = W*in
   wire signed [9:0] m267_59;
   assign m267_59 =10'b0;

   // m267_60 = W*in
   wire signed [9:0] m267_60;
   assign m267_60 =10'b0;

   // m267_61 = W*in
   wire signed [9:0] m267_61;
   assign m267_61 =10'b0;

   // m267_62 = W*in
   wire signed [9:0] m267_62;
   assign m267_62 =10'b0;

   // m267_63 = W*in
   wire signed [9:0] m267_63;
   assign m267_63 =10'b0;

   // m267_64 = W*in
   wire signed [9:0] m267_64;
   assign m267_64 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_65 = W*in
   wire signed [9:0] m267_65;
   assign m267_65 ={ {5{in267[5]}} , in267[5:1] };

   // m267_66 = W*in
   wire signed [9:0] m267_66;
   assign m267_66 ={ {5{in267[5]}} , in267[5:1] };

   // m267_67 = W*in
   wire signed [9:0] m267_67;
   assign m267_67 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_68 = W*in
   wire signed [9:0] m267_68;
   assign m267_68 =10'b0;

   // m267_69 = W*in
   wire signed [9:0] m267_69;
   assign m267_69 ={ {5{in267[5]}} , in267[5:1] };

   // m267_70 = W*in
   wire signed [9:0] m267_70;
   assign m267_70 ={ {4{in267[5]}} , in267[5:0] };

   // m267_71 = W*in
   wire signed [9:0] m267_71;
   assign m267_71 =10'b0;

   // m267_72 = W*in
   wire signed [9:0] m267_72;
   assign m267_72 =10'b0;

   // m267_73 = W*in
   wire signed [9:0] m267_73;
   assign m267_73 =10'b0;

   // m267_74 = W*in
   wire signed [9:0] m267_74;
   assign m267_74 =10'b0;

   // m267_75 = W*in
   wire signed [9:0] m267_75;
   assign m267_75 =10'b0;

   // m267_76 = W*in
   wire signed [9:0] m267_76;
   assign m267_76 =10'b0;

   // m267_77 = W*in
   wire signed [9:0] m267_77;
   assign m267_77 =10'b0;

   // m267_78 = W*in
   wire signed [9:0] m267_78;
   assign m267_78 =10'b0;

   // m267_79 = W*in
   wire signed [9:0] m267_79;
   assign m267_79 =10'b0;

   // m267_80 = W*in
   wire signed [9:0] m267_80;
   assign m267_80 =10'b0;

   // m267_81 = W*in
   wire signed [9:0] m267_81;
   assign m267_81 =10'b0;

   // m267_82 = W*in
   wire signed [9:0] m267_82;
   assign m267_82 ={ {5{in267[5]}} , in267[5:1] };

   // m267_83 = W*in
   wire signed [9:0] m267_83;
   assign m267_83 =10'b0;

   // m267_84 = W*in
   wire signed [9:0] m267_84;
   assign m267_84 =10'b0;

   // m267_85 = W*in
   wire signed [9:0] m267_85;
   assign m267_85 =10'b0;

   // m267_86 = W*in
   wire signed [9:0] m267_86;
   assign m267_86 ={ {4{in267[5]}} , in267[5:0] };

   // m267_87 = W*in
   wire signed [9:0] m267_87;
   assign m267_87 =10'b0;

   // m267_88 = W*in
   wire signed [9:0] m267_88;
   assign m267_88 =10'b0;

   // m267_89 = W*in
   wire signed [9:0] m267_89;
   assign m267_89 =10'b0;

   // m267_90 = W*in
   wire signed [9:0] m267_90;
   assign m267_90 =10'b0;

   // m267_91 = W*in
   wire signed [9:0] m267_91;
   assign m267_91 =10'b0;

   // m267_92 = W*in
   wire signed [9:0] m267_92;
   assign m267_92 =10'b0;

   // m267_93 = W*in
   wire signed [9:0] m267_93;
   assign m267_93 =10'b0;

   // m267_94 = W*in
   wire signed [9:0] m267_94;
   assign m267_94 =10'b0;

   // m267_95 = W*in
   wire signed [9:0] m267_95;
   assign m267_95 =10'b0;

   // m267_96 = W*in
   wire signed [9:0] m267_96;
   assign m267_96 =10'b0;

   // m267_97 = W*in
   wire signed [9:0] m267_97;
   assign m267_97 =10'b0;

   // m267_98 = W*in
   wire signed [9:0] m267_98;
   assign m267_98 =10'b0;

   // m267_99 = W*in
   wire signed [9:0] m267_99;
   assign m267_99 =10'b0;

   // m267_100 = W*in
   wire signed [9:0] m267_100;
   assign m267_100 =10'b0;

   // m267_101 = W*in
   wire signed [9:0] m267_101;
   assign m267_101 =10'b0;

   // m267_102 = W*in
   wire signed [9:0] m267_102;
   assign m267_102 =10'b0;

   // m267_103 = W*in
   wire signed [9:0] m267_103;
   assign m267_103 =10'b0;

   // m267_104 = W*in
   wire signed [9:0] m267_104;
   assign m267_104 =10'b0;

   // m267_105 = W*in
   wire signed [9:0] m267_105;
   assign m267_105 =10'b0;

   // m267_106 = W*in
   wire signed [9:0] m267_106;
   assign m267_106 ={ {4{neg267[5]}} , neg267[5:0] };

   // m267_107 = W*in
   wire signed [9:0] m267_107;
   assign m267_107 =10'b0;

   // m267_108 = W*in
   wire signed [9:0] m267_108;
   assign m267_108 =10'b0;

   // m267_109 = W*in
   wire signed [9:0] m267_109;
   assign m267_109 =10'b0;

   // m267_110 = W*in
   wire signed [9:0] m267_110;
   assign m267_110 =10'b0;

   // m267_111 = W*in
   wire signed [9:0] m267_111;
   assign m267_111 =10'b0;

   // m267_112 = W*in
   wire signed [9:0] m267_112;
   assign m267_112 =10'b0;

   // m267_113 = W*in
   wire signed [9:0] m267_113;
   assign m267_113 =10'b0;

   // m267_114 = W*in
   wire signed [9:0] m267_114;
   assign m267_114 =10'b0;

   // m267_115 = W*in
   wire signed [9:0] m267_115;
   assign m267_115 ={ {5{neg267[5]}} , neg267[5:1] };

   // m267_116 = W*in
   wire signed [9:0] m267_116;
   assign m267_116 =10'b0;

   // m267_117 = W*in
   wire signed [9:0] m267_117;
   assign m267_117 =10'b0;

   // m268_1 = W*in
   wire signed [9:0] m268_1;
   assign m268_1 =10'b0;

   // m268_2 = W*in
   wire signed [9:0] m268_2;
   assign m268_2 =10'b0;

   // m268_3 = W*in
   wire signed [9:0] m268_3;
   assign m268_3 =10'b0;

   // m268_4 = W*in
   wire signed [9:0] m268_4;
   assign m268_4 =10'b0;

   // m268_5 = W*in
   wire signed [9:0] m268_5;
   assign m268_5 =10'b0;

   // m268_6 = W*in
   wire signed [9:0] m268_6;
   assign m268_6 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_7 = W*in
   wire signed [9:0] m268_7;
   assign m268_7 =10'b0;

   // m268_8 = W*in
   wire signed [9:0] m268_8;
   assign m268_8 =10'b0;

   // m268_9 = W*in
   wire signed [9:0] m268_9;
   assign m268_9 =10'b0;

   // m268_10 = W*in
   wire signed [9:0] m268_10;
   assign m268_10 =10'b0;

   // m268_11 = W*in
   wire signed [9:0] m268_11;
   assign m268_11 =10'b0;

   // m268_12 = W*in
   wire signed [9:0] m268_12;
   assign m268_12 =10'b0;

   // m268_13 = W*in
   wire signed [9:0] m268_13;
   assign m268_13 ={ {4{in268[5]}} , in268[5:0] };

   // m268_14 = W*in
   wire signed [9:0] m268_14;
   assign m268_14 =10'b0;

   // m268_15 = W*in
   wire signed [9:0] m268_15;
   assign m268_15 =10'b0;

   // m268_16 = W*in
   wire signed [9:0] m268_16;
   assign m268_16 =10'b0;

   // m268_17 = W*in
   wire signed [9:0] m268_17;
   assign m268_17 =10'b0;

   // m268_18 = W*in
   wire signed [9:0] m268_18;
   assign m268_18 =10'b0;

   // m268_19 = W*in
   wire signed [9:0] m268_19;
   assign m268_19 ={ {5{neg268[5]}} , neg268[5:1] };

   // m268_20 = W*in
   wire signed [9:0] m268_20;
   assign m268_20 ={ {5{neg268[5]}} , neg268[5:1] };

   // m268_21 = W*in
   wire signed [9:0] m268_21;
   assign m268_21 ={ {5{in268[5]}} , in268[5:1] };

   // m268_22 = W*in
   wire signed [9:0] m268_22;
   assign m268_22 =10'b0;

   // m268_23 = W*in
   wire signed [9:0] m268_23;
   assign m268_23 ={ {4{in268[5]}} , in268[5:0] };

   // m268_24 = W*in
   wire signed [9:0] m268_24;
   assign m268_24 =10'b0;

   // m268_25 = W*in
   wire signed [9:0] m268_25;
   assign m268_25 =10'b0;

   // m268_26 = W*in
   wire signed [9:0] m268_26;
   assign m268_26 =10'b0;

   // m268_27 = W*in
   wire signed [9:0] m268_27;
   assign m268_27 =10'b0;

   // m268_28 = W*in
   wire signed [9:0] m268_28;
   assign m268_28 =10'b0;

   // m268_29 = W*in
   wire signed [9:0] m268_29;
   assign m268_29 ={ {4{in268[5]}} , in268[5:0] };

   // m268_30 = W*in
   wire signed [9:0] m268_30;
   assign m268_30 =10'b0;

   // m268_31 = W*in
   wire signed [9:0] m268_31;
   assign m268_31 =10'b0;

   // m268_32 = W*in
   wire signed [9:0] m268_32;
   assign m268_32 =10'b0;

   // m268_33 = W*in
   wire signed [9:0] m268_33;
   assign m268_33 =10'b0;

   // m268_34 = W*in
   wire signed [9:0] m268_34;
   assign m268_34 =10'b0;

   // m268_35 = W*in
   wire signed [9:0] m268_35;
   assign m268_35 ={ {5{neg268[5]}} , neg268[5:1] };

   // m268_36 = W*in
   wire signed [9:0] m268_36;
   assign m268_36 =10'b0;

   // m268_37 = W*in
   wire signed [9:0] m268_37;
   assign m268_37 =10'b0;

   // m268_38 = W*in
   wire signed [9:0] m268_38;
   assign m268_38 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_39 = W*in
   wire signed [9:0] m268_39;
   assign m268_39 =10'b0;

   // m268_40 = W*in
   wire signed [9:0] m268_40;
   assign m268_40 =10'b0;

   // m268_41 = W*in
   wire signed [9:0] m268_41;
   assign m268_41 ={ {4{in268[5]}} , in268[5:0] };

   // m268_42 = W*in
   wire signed [9:0] m268_42;
   assign m268_42 =10'b0;

   // m268_43 = W*in
   wire signed [9:0] m268_43;
   assign m268_43 =10'b0;

   // m268_44 = W*in
   wire signed [9:0] m268_44;
   assign m268_44 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_45 = W*in
   wire signed [9:0] m268_45;
   assign m268_45 =10'b0;

   // m268_46 = W*in
   wire signed [9:0] m268_46;
   assign m268_46 =10'b0;

   // m268_47 = W*in
   wire signed [9:0] m268_47;
   assign m268_47 =10'b0;

   // m268_48 = W*in
   wire signed [9:0] m268_48;
   assign m268_48 =10'b0;

   // m268_49 = W*in
   wire signed [9:0] m268_49;
   assign m268_49 =10'b0;

   // m268_50 = W*in
   wire signed [9:0] m268_50;
   assign m268_50 =10'b0;

   // m268_51 = W*in
   wire signed [9:0] m268_51;
   assign m268_51 =10'b0;

   // m268_52 = W*in
   wire signed [9:0] m268_52;
   assign m268_52 =10'b0;

   // m268_53 = W*in
   wire signed [9:0] m268_53;
   assign m268_53 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_54 = W*in
   wire signed [9:0] m268_54;
   assign m268_54 =10'b0;

   // m268_55 = W*in
   wire signed [9:0] m268_55;
   assign m268_55 =10'b0;

   // m268_56 = W*in
   wire signed [9:0] m268_56;
   assign m268_56 =10'b0;

   // m268_57 = W*in
   wire signed [9:0] m268_57;
   assign m268_57 =10'b0;

   // m268_58 = W*in
   wire signed [9:0] m268_58;
   assign m268_58 =10'b0;

   // m268_59 = W*in
   wire signed [9:0] m268_59;
   assign m268_59 =10'b0;

   // m268_60 = W*in
   wire signed [9:0] m268_60;
   assign m268_60 =10'b0;

   // m268_61 = W*in
   wire signed [9:0] m268_61;
   assign m268_61 =10'b0;

   // m268_62 = W*in
   wire signed [9:0] m268_62;
   assign m268_62 =10'b0;

   // m268_63 = W*in
   wire signed [9:0] m268_63;
   assign m268_63 =10'b0;

   // m268_64 = W*in
   wire signed [9:0] m268_64;
   assign m268_64 ={ {5{neg268[5]}} , neg268[5:1] };

   // m268_65 = W*in
   wire signed [9:0] m268_65;
   assign m268_65 ={ {5{in268[5]}} , in268[5:1] };

   // m268_66 = W*in
   wire signed [9:0] m268_66;
   assign m268_66 ={ {5{in268[5]}} , in268[5:1] };

   // m268_67 = W*in
   wire signed [9:0] m268_67;
   assign m268_67 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_68 = W*in
   wire signed [9:0] m268_68;
   assign m268_68 =10'b0;

   // m268_69 = W*in
   wire signed [9:0] m268_69;
   assign m268_69 ={ {4{in268[5]}} , in268[5:0] };

   // m268_70 = W*in
   wire signed [9:0] m268_70;
   assign m268_70 ={ {4{in268[5]}} , in268[5:0] };

   // m268_71 = W*in
   wire signed [9:0] m268_71;
   assign m268_71 =10'b0;

   // m268_72 = W*in
   wire signed [9:0] m268_72;
   assign m268_72 =10'b0;

   // m268_73 = W*in
   wire signed [9:0] m268_73;
   assign m268_73 =10'b0;

   // m268_74 = W*in
   wire signed [9:0] m268_74;
   assign m268_74 =10'b0;

   // m268_75 = W*in
   wire signed [9:0] m268_75;
   assign m268_75 =10'b0;

   // m268_76 = W*in
   wire signed [9:0] m268_76;
   assign m268_76 =10'b0;

   // m268_77 = W*in
   wire signed [9:0] m268_77;
   assign m268_77 =10'b0;

   // m268_78 = W*in
   wire signed [9:0] m268_78;
   assign m268_78 =10'b0;

   // m268_79 = W*in
   wire signed [9:0] m268_79;
   assign m268_79 =10'b0;

   // m268_80 = W*in
   wire signed [9:0] m268_80;
   assign m268_80 =10'b0;

   // m268_81 = W*in
   wire signed [9:0] m268_81;
   assign m268_81 =10'b0;

   // m268_82 = W*in
   wire signed [9:0] m268_82;
   assign m268_82 =10'b0;

   // m268_83 = W*in
   wire signed [9:0] m268_83;
   assign m268_83 =10'b0;

   // m268_84 = W*in
   wire signed [9:0] m268_84;
   assign m268_84 =10'b0;

   // m268_85 = W*in
   wire signed [9:0] m268_85;
   assign m268_85 =10'b0;

   // m268_86 = W*in
   wire signed [9:0] m268_86;
   assign m268_86 ={ {4{in268[5]}} , in268[5:0] };

   // m268_87 = W*in
   wire signed [9:0] m268_87;
   assign m268_87 =10'b0;

   // m268_88 = W*in
   wire signed [9:0] m268_88;
   assign m268_88 =10'b0;

   // m268_89 = W*in
   wire signed [9:0] m268_89;
   assign m268_89 =10'b0;

   // m268_90 = W*in
   wire signed [9:0] m268_90;
   assign m268_90 =10'b0;

   // m268_91 = W*in
   wire signed [9:0] m268_91;
   assign m268_91 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_92 = W*in
   wire signed [9:0] m268_92;
   assign m268_92 =10'b0;

   // m268_93 = W*in
   wire signed [9:0] m268_93;
   assign m268_93 =10'b0;

   // m268_94 = W*in
   wire signed [9:0] m268_94;
   assign m268_94 =10'b0;

   // m268_95 = W*in
   wire signed [9:0] m268_95;
   assign m268_95 =10'b0;

   // m268_96 = W*in
   wire signed [9:0] m268_96;
   assign m268_96 ={ {4{in268[5]}} , in268[5:0] };

   // m268_97 = W*in
   wire signed [9:0] m268_97;
   assign m268_97 ={ {4{neg268[5]}} , neg268[5:0] };

   // m268_98 = W*in
   wire signed [9:0] m268_98;
   assign m268_98 =10'b0;

   // m268_99 = W*in
   wire signed [9:0] m268_99;
   assign m268_99 =10'b0;

   // m268_100 = W*in
   wire signed [9:0] m268_100;
   assign m268_100 =10'b0;

   // m268_101 = W*in
   wire signed [9:0] m268_101;
   assign m268_101 =10'b0;

   // m268_102 = W*in
   wire signed [9:0] m268_102;
   assign m268_102 =10'b0;

   // m268_103 = W*in
   wire signed [9:0] m268_103;
   assign m268_103 =10'b0;

   // m268_104 = W*in
   wire signed [9:0] m268_104;
   assign m268_104 =10'b0;

   // m268_105 = W*in
   wire signed [9:0] m268_105;
   assign m268_105 =10'b0;

   // m268_106 = W*in
   wire signed [9:0] m268_106;
   assign m268_106 ={ {5{neg268[5]}} , neg268[5:1] };

   // m268_107 = W*in
   wire signed [9:0] m268_107;
   assign m268_107 =10'b0;

   // m268_108 = W*in
   wire signed [9:0] m268_108;
   assign m268_108 ={ {4{in268[5]}} , in268[5:0] };

   // m268_109 = W*in
   wire signed [9:0] m268_109;
   assign m268_109 ={ {4{in268[5]}} , in268[5:0] };

   // m268_110 = W*in
   wire signed [9:0] m268_110;
   assign m268_110 =10'b0;

   // m268_111 = W*in
   wire signed [9:0] m268_111;
   assign m268_111 =10'b0;

   // m268_112 = W*in
   wire signed [9:0] m268_112;
   assign m268_112 =10'b0;

   // m268_113 = W*in
   wire signed [9:0] m268_113;
   assign m268_113 =10'b0;

   // m268_114 = W*in
   wire signed [9:0] m268_114;
   assign m268_114 =10'b0;

   // m268_115 = W*in
   wire signed [9:0] m268_115;
   assign m268_115 ={ {5{neg268[5]}} , neg268[5:1] };

   // m268_116 = W*in
   wire signed [9:0] m268_116;
   assign m268_116 ={ {4{in268[5]}} , in268[5:0] };

   // m268_117 = W*in
   wire signed [9:0] m268_117;
   assign m268_117 =10'b0;

   // m269_1 = W*in
   wire signed [9:0] m269_1;
   assign m269_1 =10'b0;

   // m269_2 = W*in
   wire signed [9:0] m269_2;
   assign m269_2 =10'b0;

   // m269_3 = W*in
   wire signed [9:0] m269_3;
   assign m269_3 =10'b0;

   // m269_4 = W*in
   wire signed [9:0] m269_4;
   assign m269_4 =10'b0;

   // m269_5 = W*in
   wire signed [9:0] m269_5;
   assign m269_5 =10'b0;

   // m269_6 = W*in
   wire signed [9:0] m269_6;
   assign m269_6 =10'b0;

   // m269_7 = W*in
   wire signed [9:0] m269_7;
   assign m269_7 ={ {4{in269[5]}} , in269[5:0] };

   // m269_8 = W*in
   wire signed [9:0] m269_8;
   assign m269_8 =10'b0;

   // m269_9 = W*in
   wire signed [9:0] m269_9;
   assign m269_9 =10'b0;

   // m269_10 = W*in
   wire signed [9:0] m269_10;
   assign m269_10 =10'b0;

   // m269_11 = W*in
   wire signed [9:0] m269_11;
   assign m269_11 =10'b0;

   // m269_12 = W*in
   wire signed [9:0] m269_12;
   assign m269_12 =10'b0;

   // m269_13 = W*in
   wire signed [9:0] m269_13;
   assign m269_13 =10'b0;

   // m269_14 = W*in
   wire signed [9:0] m269_14;
   assign m269_14 =10'b0;

   // m269_15 = W*in
   wire signed [9:0] m269_15;
   assign m269_15 =10'b0;

   // m269_16 = W*in
   wire signed [9:0] m269_16;
   assign m269_16 ={ {5{in269[5]}} , in269[5:1] };

   // m269_17 = W*in
   wire signed [9:0] m269_17;
   assign m269_17 =10'b0;

   // m269_18 = W*in
   wire signed [9:0] m269_18;
   assign m269_18 =10'b0;

   // m269_19 = W*in
   wire signed [9:0] m269_19;
   assign m269_19 =10'b0;

   // m269_20 = W*in
   wire signed [9:0] m269_20;
   assign m269_20 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_21 = W*in
   wire signed [9:0] m269_21;
   assign m269_21 ={ {5{in269[5]}} , in269[5:1] };

   // m269_22 = W*in
   wire signed [9:0] m269_22;
   assign m269_22 =10'b0;

   // m269_23 = W*in
   wire signed [9:0] m269_23;
   assign m269_23 =10'b0;

   // m269_24 = W*in
   wire signed [9:0] m269_24;
   assign m269_24 =10'b0;

   // m269_25 = W*in
   wire signed [9:0] m269_25;
   assign m269_25 =10'b0;

   // m269_26 = W*in
   wire signed [9:0] m269_26;
   assign m269_26 =10'b0;

   // m269_27 = W*in
   wire signed [9:0] m269_27;
   assign m269_27 =10'b0;

   // m269_28 = W*in
   wire signed [9:0] m269_28;
   assign m269_28 =10'b0;

   // m269_29 = W*in
   wire signed [9:0] m269_29;
   assign m269_29 =10'b0;

   // m269_30 = W*in
   wire signed [9:0] m269_30;
   assign m269_30 =10'b0;

   // m269_31 = W*in
   wire signed [9:0] m269_31;
   assign m269_31 =10'b0;

   // m269_32 = W*in
   wire signed [9:0] m269_32;
   assign m269_32 =10'b0;

   // m269_33 = W*in
   wire signed [9:0] m269_33;
   assign m269_33 ={ {4{in269[5]}} , in269[5:0] };

   // m269_34 = W*in
   wire signed [9:0] m269_34;
   assign m269_34 =10'b0;

   // m269_35 = W*in
   wire signed [9:0] m269_35;
   assign m269_35 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_36 = W*in
   wire signed [9:0] m269_36;
   assign m269_36 ={ {5{in269[5]}} , in269[5:1] };

   // m269_37 = W*in
   wire signed [9:0] m269_37;
   assign m269_37 =10'b0;

   // m269_38 = W*in
   wire signed [9:0] m269_38;
   assign m269_38 =10'b0;

   // m269_39 = W*in
   wire signed [9:0] m269_39;
   assign m269_39 =10'b0;

   // m269_40 = W*in
   wire signed [9:0] m269_40;
   assign m269_40 =10'b0;

   // m269_41 = W*in
   wire signed [9:0] m269_41;
   assign m269_41 =10'b0;

   // m269_42 = W*in
   wire signed [9:0] m269_42;
   assign m269_42 =10'b0;

   // m269_43 = W*in
   wire signed [9:0] m269_43;
   assign m269_43 =10'b0;

   // m269_44 = W*in
   wire signed [9:0] m269_44;
   assign m269_44 =10'b0;

   // m269_45 = W*in
   wire signed [9:0] m269_45;
   assign m269_45 =10'b0;

   // m269_46 = W*in
   wire signed [9:0] m269_46;
   assign m269_46 =10'b0;

   // m269_47 = W*in
   wire signed [9:0] m269_47;
   assign m269_47 =10'b0;

   // m269_48 = W*in
   wire signed [9:0] m269_48;
   assign m269_48 =10'b0;

   // m269_49 = W*in
   wire signed [9:0] m269_49;
   assign m269_49 =10'b0;

   // m269_50 = W*in
   wire signed [9:0] m269_50;
   assign m269_50 =10'b0;

   // m269_51 = W*in
   wire signed [9:0] m269_51;
   assign m269_51 =10'b0;

   // m269_52 = W*in
   wire signed [9:0] m269_52;
   assign m269_52 =10'b0;

   // m269_53 = W*in
   wire signed [9:0] m269_53;
   assign m269_53 =10'b0;

   // m269_54 = W*in
   wire signed [9:0] m269_54;
   assign m269_54 =10'b0;

   // m269_55 = W*in
   wire signed [9:0] m269_55;
   assign m269_55 =10'b0;

   // m269_56 = W*in
   wire signed [9:0] m269_56;
   assign m269_56 =10'b0;

   // m269_57 = W*in
   wire signed [9:0] m269_57;
   assign m269_57 =10'b0;

   // m269_58 = W*in
   wire signed [9:0] m269_58;
   assign m269_58 =10'b0;

   // m269_59 = W*in
   wire signed [9:0] m269_59;
   assign m269_59 =10'b0;

   // m269_60 = W*in
   wire signed [9:0] m269_60;
   assign m269_60 =10'b0;

   // m269_61 = W*in
   wire signed [9:0] m269_61;
   assign m269_61 =10'b0;

   // m269_62 = W*in
   wire signed [9:0] m269_62;
   assign m269_62 =10'b0;

   // m269_63 = W*in
   wire signed [9:0] m269_63;
   assign m269_63 =10'b0;

   // m269_64 = W*in
   wire signed [9:0] m269_64;
   assign m269_64 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_65 = W*in
   wire signed [9:0] m269_65;
   assign m269_65 =10'b0;

   // m269_66 = W*in
   wire signed [9:0] m269_66;
   assign m269_66 ={ {5{in269[5]}} , in269[5:1] };

   // m269_67 = W*in
   wire signed [9:0] m269_67;
   assign m269_67 =10'b0;

   // m269_68 = W*in
   wire signed [9:0] m269_68;
   assign m269_68 =10'b0;

   // m269_69 = W*in
   wire signed [9:0] m269_69;
   assign m269_69 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_70 = W*in
   wire signed [9:0] m269_70;
   assign m269_70 =10'b0;

   // m269_71 = W*in
   wire signed [9:0] m269_71;
   assign m269_71 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_72 = W*in
   wire signed [9:0] m269_72;
   assign m269_72 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_73 = W*in
   wire signed [9:0] m269_73;
   assign m269_73 ={ {5{in269[5]}} , in269[5:1] };

   // m269_74 = W*in
   wire signed [9:0] m269_74;
   assign m269_74 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_75 = W*in
   wire signed [9:0] m269_75;
   assign m269_75 =10'b0;

   // m269_76 = W*in
   wire signed [9:0] m269_76;
   assign m269_76 =10'b0;

   // m269_77 = W*in
   wire signed [9:0] m269_77;
   assign m269_77 =10'b0;

   // m269_78 = W*in
   wire signed [9:0] m269_78;
   assign m269_78 ={ {5{in269[5]}} , in269[5:1] };

   // m269_79 = W*in
   wire signed [9:0] m269_79;
   assign m269_79 =10'b0;

   // m269_80 = W*in
   wire signed [9:0] m269_80;
   assign m269_80 =10'b0;

   // m269_81 = W*in
   wire signed [9:0] m269_81;
   assign m269_81 =10'b0;

   // m269_82 = W*in
   wire signed [9:0] m269_82;
   assign m269_82 =10'b0;

   // m269_83 = W*in
   wire signed [9:0] m269_83;
   assign m269_83 =10'b0;

   // m269_84 = W*in
   wire signed [9:0] m269_84;
   assign m269_84 =10'b0;

   // m269_85 = W*in
   wire signed [9:0] m269_85;
   assign m269_85 =10'b0;

   // m269_86 = W*in
   wire signed [9:0] m269_86;
   assign m269_86 =10'b0;

   // m269_87 = W*in
   wire signed [9:0] m269_87;
   assign m269_87 =10'b0;

   // m269_88 = W*in
   wire signed [9:0] m269_88;
   assign m269_88 =10'b0;

   // m269_89 = W*in
   wire signed [9:0] m269_89;
   assign m269_89 =10'b0;

   // m269_90 = W*in
   wire signed [9:0] m269_90;
   assign m269_90 =10'b0;

   // m269_91 = W*in
   wire signed [9:0] m269_91;
   assign m269_91 =10'b0;

   // m269_92 = W*in
   wire signed [9:0] m269_92;
   assign m269_92 ={ {4{neg269[5]}} , neg269[5:0] };

   // m269_93 = W*in
   wire signed [9:0] m269_93;
   assign m269_93 =10'b0;

   // m269_94 = W*in
   wire signed [9:0] m269_94;
   assign m269_94 =10'b0;

   // m269_95 = W*in
   wire signed [9:0] m269_95;
   assign m269_95 =10'b0;

   // m269_96 = W*in
   wire signed [9:0] m269_96;
   assign m269_96 =10'b0;

   // m269_97 = W*in
   wire signed [9:0] m269_97;
   assign m269_97 =10'b0;

   // m269_98 = W*in
   wire signed [9:0] m269_98;
   assign m269_98 =10'b0;

   // m269_99 = W*in
   wire signed [9:0] m269_99;
   assign m269_99 =10'b0;

   // m269_100 = W*in
   wire signed [9:0] m269_100;
   assign m269_100 =10'b0;

   // m269_101 = W*in
   wire signed [9:0] m269_101;
   assign m269_101 =10'b0;

   // m269_102 = W*in
   wire signed [9:0] m269_102;
   assign m269_102 =10'b0;

   // m269_103 = W*in
   wire signed [9:0] m269_103;
   assign m269_103 =10'b0;

   // m269_104 = W*in
   wire signed [9:0] m269_104;
   assign m269_104 =10'b0;

   // m269_105 = W*in
   wire signed [9:0] m269_105;
   assign m269_105 =10'b0;

   // m269_106 = W*in
   wire signed [9:0] m269_106;
   assign m269_106 =10'b0;

   // m269_107 = W*in
   wire signed [9:0] m269_107;
   assign m269_107 =10'b0;

   // m269_108 = W*in
   wire signed [9:0] m269_108;
   assign m269_108 =10'b0;

   // m269_109 = W*in
   wire signed [9:0] m269_109;
   assign m269_109 =10'b0;

   // m269_110 = W*in
   wire signed [9:0] m269_110;
   assign m269_110 =10'b0;

   // m269_111 = W*in
   wire signed [9:0] m269_111;
   assign m269_111 =10'b0;

   // m269_112 = W*in
   wire signed [9:0] m269_112;
   assign m269_112 =10'b0;

   // m269_113 = W*in
   wire signed [9:0] m269_113;
   assign m269_113 =10'b0;

   // m269_114 = W*in
   wire signed [9:0] m269_114;
   assign m269_114 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_115 = W*in
   wire signed [9:0] m269_115;
   assign m269_115 ={ {5{neg269[5]}} , neg269[5:1] };

   // m269_116 = W*in
   wire signed [9:0] m269_116;
   assign m269_116 =10'b0;

   // m269_117 = W*in
   wire signed [9:0] m269_117;
   assign m269_117 =10'b0;

   // m270_1 = W*in
   wire signed [9:0] m270_1;
   assign m270_1 =10'b0;

   // m270_2 = W*in
   wire signed [9:0] m270_2;
   assign m270_2 =10'b0;

   // m270_3 = W*in
   wire signed [9:0] m270_3;
   assign m270_3 =10'b0;

   // m270_4 = W*in
   wire signed [9:0] m270_4;
   assign m270_4 =10'b0;

   // m270_5 = W*in
   wire signed [9:0] m270_5;
   assign m270_5 =10'b0;

   // m270_6 = W*in
   wire signed [9:0] m270_6;
   assign m270_6 =10'b0;

   // m270_7 = W*in
   wire signed [9:0] m270_7;
   assign m270_7 =10'b0;

   // m270_8 = W*in
   wire signed [9:0] m270_8;
   assign m270_8 =10'b0;

   // m270_9 = W*in
   wire signed [9:0] m270_9;
   assign m270_9 =10'b0;

   // m270_10 = W*in
   wire signed [9:0] m270_10;
   assign m270_10 ={ {4{in270[5]}} , in270[5:0] };

   // m270_11 = W*in
   wire signed [9:0] m270_11;
   assign m270_11 =10'b0;

   // m270_12 = W*in
   wire signed [9:0] m270_12;
   assign m270_12 =10'b0;

   // m270_13 = W*in
   wire signed [9:0] m270_13;
   assign m270_13 =10'b0;

   // m270_14 = W*in
   wire signed [9:0] m270_14;
   assign m270_14 =10'b0;

   // m270_15 = W*in
   wire signed [9:0] m270_15;
   assign m270_15 =10'b0;

   // m270_16 = W*in
   wire signed [9:0] m270_16;
   assign m270_16 =10'b0;

   // m270_17 = W*in
   wire signed [9:0] m270_17;
   assign m270_17 ={ {5{in270[5]}} , in270[5:1] };

   // m270_18 = W*in
   wire signed [9:0] m270_18;
   assign m270_18 =10'b0;

   // m270_19 = W*in
   wire signed [9:0] m270_19;
   assign m270_19 =10'b0;

   // m270_20 = W*in
   wire signed [9:0] m270_20;
   assign m270_20 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_21 = W*in
   wire signed [9:0] m270_21;
   assign m270_21 ={ {4{in270[5]}} , in270[5:0] };

   // m270_22 = W*in
   wire signed [9:0] m270_22;
   assign m270_22 =10'b0;

   // m270_23 = W*in
   wire signed [9:0] m270_23;
   assign m270_23 =10'b0;

   // m270_24 = W*in
   wire signed [9:0] m270_24;
   assign m270_24 =10'b0;

   // m270_25 = W*in
   wire signed [9:0] m270_25;
   assign m270_25 =10'b0;

   // m270_26 = W*in
   wire signed [9:0] m270_26;
   assign m270_26 ={ {4{in270[5]}} , in270[5:0] };

   // m270_27 = W*in
   wire signed [9:0] m270_27;
   assign m270_27 ={ {5{neg270[5]}} , neg270[5:1] };

   // m270_28 = W*in
   wire signed [9:0] m270_28;
   assign m270_28 =10'b0;

   // m270_29 = W*in
   wire signed [9:0] m270_29;
   assign m270_29 ={ {4{in270[5]}} , in270[5:0] };

   // m270_30 = W*in
   wire signed [9:0] m270_30;
   assign m270_30 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_31 = W*in
   wire signed [9:0] m270_31;
   assign m270_31 ={ {5{neg270[5]}} , neg270[5:1] };

   // m270_32 = W*in
   wire signed [9:0] m270_32;
   assign m270_32 =10'b0;

   // m270_33 = W*in
   wire signed [9:0] m270_33;
   assign m270_33 =10'b0;

   // m270_34 = W*in
   wire signed [9:0] m270_34;
   assign m270_34 ={ {5{neg270[5]}} , neg270[5:1] };

   // m270_35 = W*in
   wire signed [9:0] m270_35;
   assign m270_35 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_36 = W*in
   wire signed [9:0] m270_36;
   assign m270_36 =10'b0;

   // m270_37 = W*in
   wire signed [9:0] m270_37;
   assign m270_37 ={ {4{in270[5]}} , in270[5:0] };

   // m270_38 = W*in
   wire signed [9:0] m270_38;
   assign m270_38 =10'b0;

   // m270_39 = W*in
   wire signed [9:0] m270_39;
   assign m270_39 =10'b0;

   // m270_40 = W*in
   wire signed [9:0] m270_40;
   assign m270_40 =10'b0;

   // m270_41 = W*in
   wire signed [9:0] m270_41;
   assign m270_41 =10'b0;

   // m270_42 = W*in
   wire signed [9:0] m270_42;
   assign m270_42 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_43 = W*in
   wire signed [9:0] m270_43;
   assign m270_43 =10'b0;

   // m270_44 = W*in
   wire signed [9:0] m270_44;
   assign m270_44 =10'b0;

   // m270_45 = W*in
   wire signed [9:0] m270_45;
   assign m270_45 =10'b0;

   // m270_46 = W*in
   wire signed [9:0] m270_46;
   assign m270_46 =10'b0;

   // m270_47 = W*in
   wire signed [9:0] m270_47;
   assign m270_47 =10'b0;

   // m270_48 = W*in
   wire signed [9:0] m270_48;
   assign m270_48 =10'b0;

   // m270_49 = W*in
   wire signed [9:0] m270_49;
   assign m270_49 =10'b0;

   // m270_50 = W*in
   wire signed [9:0] m270_50;
   assign m270_50 =10'b0;

   // m270_51 = W*in
   wire signed [9:0] m270_51;
   assign m270_51 =10'b0;

   // m270_52 = W*in
   wire signed [9:0] m270_52;
   assign m270_52 =10'b0;

   // m270_53 = W*in
   wire signed [9:0] m270_53;
   assign m270_53 ={ {4{in270[5]}} , in270[5:0] };

   // m270_54 = W*in
   wire signed [9:0] m270_54;
   assign m270_54 =10'b0;

   // m270_55 = W*in
   wire signed [9:0] m270_55;
   assign m270_55 ={ {4{in270[5]}} , in270[5:0] };

   // m270_56 = W*in
   wire signed [9:0] m270_56;
   assign m270_56 =10'b0;

   // m270_57 = W*in
   wire signed [9:0] m270_57;
   assign m270_57 =10'b0;

   // m270_58 = W*in
   wire signed [9:0] m270_58;
   assign m270_58 =10'b0;

   // m270_59 = W*in
   wire signed [9:0] m270_59;
   assign m270_59 =10'b0;

   // m270_60 = W*in
   wire signed [9:0] m270_60;
   assign m270_60 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_61 = W*in
   wire signed [9:0] m270_61;
   assign m270_61 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_62 = W*in
   wire signed [9:0] m270_62;
   assign m270_62 =10'b0;

   // m270_63 = W*in
   wire signed [9:0] m270_63;
   assign m270_63 ={ {4{in270[5]}} , in270[5:0] };

   // m270_64 = W*in
   wire signed [9:0] m270_64;
   assign m270_64 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_65 = W*in
   wire signed [9:0] m270_65;
   assign m270_65 =10'b0;

   // m270_66 = W*in
   wire signed [9:0] m270_66;
   assign m270_66 =10'b0;

   // m270_67 = W*in
   wire signed [9:0] m270_67;
   assign m270_67 =10'b0;

   // m270_68 = W*in
   wire signed [9:0] m270_68;
   assign m270_68 =10'b0;

   // m270_69 = W*in
   wire signed [9:0] m270_69;
   assign m270_69 ={ {4{in270[5]}} , in270[5:0] };

   // m270_70 = W*in
   wire signed [9:0] m270_70;
   assign m270_70 ={ {4{in270[5]}} , in270[5:0] };

   // m270_71 = W*in
   wire signed [9:0] m270_71;
   assign m270_71 =10'b0;

   // m270_72 = W*in
   wire signed [9:0] m270_72;
   assign m270_72 =10'b0;

   // m270_73 = W*in
   wire signed [9:0] m270_73;
   assign m270_73 =10'b0;

   // m270_74 = W*in
   wire signed [9:0] m270_74;
   assign m270_74 =10'b0;

   // m270_75 = W*in
   wire signed [9:0] m270_75;
   assign m270_75 ={ {5{neg270[5]}} , neg270[5:1] };

   // m270_76 = W*in
   wire signed [9:0] m270_76;
   assign m270_76 =10'b0;

   // m270_77 = W*in
   wire signed [9:0] m270_77;
   assign m270_77 =10'b0;

   // m270_78 = W*in
   wire signed [9:0] m270_78;
   assign m270_78 ={ {4{in270[5]}} , in270[5:0] };

   // m270_79 = W*in
   wire signed [9:0] m270_79;
   assign m270_79 =10'b0;

   // m270_80 = W*in
   wire signed [9:0] m270_80;
   assign m270_80 =10'b0;

   // m270_81 = W*in
   wire signed [9:0] m270_81;
   assign m270_81 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_82 = W*in
   wire signed [9:0] m270_82;
   assign m270_82 ={ {3{in270[5]}} , in270 , {1{1'b0}} };

   // m270_83 = W*in
   wire signed [9:0] m270_83;
   assign m270_83 =10'b0;

   // m270_84 = W*in
   wire signed [9:0] m270_84;
   assign m270_84 =10'b0;

   // m270_85 = W*in
   wire signed [9:0] m270_85;
   assign m270_85 ={ {4{in270[5]}} , in270[5:0] };

   // m270_86 = W*in
   wire signed [9:0] m270_86;
   assign m270_86 ={ {4{in270[5]}} , in270[5:0] };

   // m270_87 = W*in
   wire signed [9:0] m270_87;
   assign m270_87 ={ {4{in270[5]}} , in270[5:0] };

   // m270_88 = W*in
   wire signed [9:0] m270_88;
   assign m270_88 =10'b0;

   // m270_89 = W*in
   wire signed [9:0] m270_89;
   assign m270_89 =10'b0;

   // m270_90 = W*in
   wire signed [9:0] m270_90;
   assign m270_90 =10'b0;

   // m270_91 = W*in
   wire signed [9:0] m270_91;
   assign m270_91 =10'b0;

   // m270_92 = W*in
   wire signed [9:0] m270_92;
   assign m270_92 =10'b0;

   // m270_93 = W*in
   wire signed [9:0] m270_93;
   assign m270_93 =10'b0;

   // m270_94 = W*in
   wire signed [9:0] m270_94;
   assign m270_94 =10'b0;

   // m270_95 = W*in
   wire signed [9:0] m270_95;
   assign m270_95 =10'b0;

   // m270_96 = W*in
   wire signed [9:0] m270_96;
   assign m270_96 =10'b0;

   // m270_97 = W*in
   wire signed [9:0] m270_97;
   assign m270_97 =10'b0;

   // m270_98 = W*in
   wire signed [9:0] m270_98;
   assign m270_98 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_99 = W*in
   wire signed [9:0] m270_99;
   assign m270_99 ={ {4{in270[5]}} , in270[5:0] };

   // m270_100 = W*in
   wire signed [9:0] m270_100;
   assign m270_100 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_101 = W*in
   wire signed [9:0] m270_101;
   assign m270_101 =10'b0;

   // m270_102 = W*in
   wire signed [9:0] m270_102;
   assign m270_102 =10'b0;

   // m270_103 = W*in
   wire signed [9:0] m270_103;
   assign m270_103 =10'b0;

   // m270_104 = W*in
   wire signed [9:0] m270_104;
   assign m270_104 =10'b0;

   // m270_105 = W*in
   wire signed [9:0] m270_105;
   assign m270_105 =10'b0;

   // m270_106 = W*in
   wire signed [9:0] m270_106;
   assign m270_106 =10'b0;

   // m270_107 = W*in
   wire signed [9:0] m270_107;
   assign m270_107 =10'b0;

   // m270_108 = W*in
   wire signed [9:0] m270_108;
   assign m270_108 =10'b0;

   // m270_109 = W*in
   wire signed [9:0] m270_109;
   assign m270_109 =10'b0;

   // m270_110 = W*in
   wire signed [9:0] m270_110;
   assign m270_110 =10'b0;

   // m270_111 = W*in
   wire signed [9:0] m270_111;
   assign m270_111 =10'b0;

   // m270_112 = W*in
   wire signed [9:0] m270_112;
   assign m270_112 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_113 = W*in
   wire signed [9:0] m270_113;
   assign m270_113 =10'b0;

   // m270_114 = W*in
   wire signed [9:0] m270_114;
   assign m270_114 ={ {5{neg270[5]}} , neg270[5:1] };

   // m270_115 = W*in
   wire signed [9:0] m270_115;
   assign m270_115 ={ {4{neg270[5]}} , neg270[5:0] };

   // m270_116 = W*in
   wire signed [9:0] m270_116;
   assign m270_116 =10'b0;

   // m270_117 = W*in
   wire signed [9:0] m270_117;
   assign m270_117 ={ {4{neg270[5]}} , neg270[5:0] };

   // m271_1 = W*in
   wire signed [9:0] m271_1;
   assign m271_1 =10'b0;

   // m271_2 = W*in
   wire signed [9:0] m271_2;
   assign m271_2 =10'b0;

   // m271_3 = W*in
   wire signed [9:0] m271_3;
   assign m271_3 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_4 = W*in
   wire signed [9:0] m271_4;
   assign m271_4 =10'b0;

   // m271_5 = W*in
   wire signed [9:0] m271_5;
   assign m271_5 ={ {4{in271[5]}} , in271[5:0] };

   // m271_6 = W*in
   wire signed [9:0] m271_6;
   assign m271_6 =10'b0;

   // m271_7 = W*in
   wire signed [9:0] m271_7;
   assign m271_7 =10'b0;

   // m271_8 = W*in
   wire signed [9:0] m271_8;
   assign m271_8 =10'b0;

   // m271_9 = W*in
   wire signed [9:0] m271_9;
   assign m271_9 =10'b0;

   // m271_10 = W*in
   wire signed [9:0] m271_10;
   assign m271_10 ={ {4{in271[5]}} , in271[5:0] };

   // m271_11 = W*in
   wire signed [9:0] m271_11;
   assign m271_11 =10'b0;

   // m271_12 = W*in
   wire signed [9:0] m271_12;
   assign m271_12 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_13 = W*in
   wire signed [9:0] m271_13;
   assign m271_13 =10'b0;

   // m271_14 = W*in
   wire signed [9:0] m271_14;
   assign m271_14 ={ {4{in271[5]}} , in271[5:0] };

   // m271_15 = W*in
   wire signed [9:0] m271_15;
   assign m271_15 =10'b0;

   // m271_16 = W*in
   wire signed [9:0] m271_16;
   assign m271_16 =10'b0;

   // m271_17 = W*in
   wire signed [9:0] m271_17;
   assign m271_17 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_18 = W*in
   wire signed [9:0] m271_18;
   assign m271_18 =10'b0;

   // m271_19 = W*in
   wire signed [9:0] m271_19;
   assign m271_19 ={ {4{in271[5]}} , in271[5:0] };

   // m271_20 = W*in
   wire signed [9:0] m271_20;
   assign m271_20 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_21 = W*in
   wire signed [9:0] m271_21;
   assign m271_21 ={ {5{in271[5]}} , in271[5:1] };

   // m271_22 = W*in
   wire signed [9:0] m271_22;
   assign m271_22 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_23 = W*in
   wire signed [9:0] m271_23;
   assign m271_23 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_24 = W*in
   wire signed [9:0] m271_24;
   assign m271_24 =10'b0;

   // m271_25 = W*in
   wire signed [9:0] m271_25;
   assign m271_25 =10'b0;

   // m271_26 = W*in
   wire signed [9:0] m271_26;
   assign m271_26 ={ {4{in271[5]}} , in271[5:0] };

   // m271_27 = W*in
   wire signed [9:0] m271_27;
   assign m271_27 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_28 = W*in
   wire signed [9:0] m271_28;
   assign m271_28 =10'b0;

   // m271_29 = W*in
   wire signed [9:0] m271_29;
   assign m271_29 =10'b0;

   // m271_30 = W*in
   wire signed [9:0] m271_30;
   assign m271_30 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_31 = W*in
   wire signed [9:0] m271_31;
   assign m271_31 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_32 = W*in
   wire signed [9:0] m271_32;
   assign m271_32 ={ {4{in271[5]}} , in271[5:0] };

   // m271_33 = W*in
   wire signed [9:0] m271_33;
   assign m271_33 =10'b0;

   // m271_34 = W*in
   wire signed [9:0] m271_34;
   assign m271_34 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_35 = W*in
   wire signed [9:0] m271_35;
   assign m271_35 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_36 = W*in
   wire signed [9:0] m271_36;
   assign m271_36 =10'b0;

   // m271_37 = W*in
   wire signed [9:0] m271_37;
   assign m271_37 =10'b0;

   // m271_38 = W*in
   wire signed [9:0] m271_38;
   assign m271_38 =10'b0;

   // m271_39 = W*in
   wire signed [9:0] m271_39;
   assign m271_39 =10'b0;

   // m271_40 = W*in
   wire signed [9:0] m271_40;
   assign m271_40 =10'b0;

   // m271_41 = W*in
   wire signed [9:0] m271_41;
   assign m271_41 =10'b0;

   // m271_42 = W*in
   wire signed [9:0] m271_42;
   assign m271_42 =10'b0;

   // m271_43 = W*in
   wire signed [9:0] m271_43;
   assign m271_43 =10'b0;

   // m271_44 = W*in
   wire signed [9:0] m271_44;
   assign m271_44 =10'b0;

   // m271_45 = W*in
   wire signed [9:0] m271_45;
   assign m271_45 =10'b0;

   // m271_46 = W*in
   wire signed [9:0] m271_46;
   assign m271_46 =10'b0;

   // m271_47 = W*in
   wire signed [9:0] m271_47;
   assign m271_47 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_48 = W*in
   wire signed [9:0] m271_48;
   assign m271_48 ={ {4{in271[5]}} , in271[5:0] };

   // m271_49 = W*in
   wire signed [9:0] m271_49;
   assign m271_49 =10'b0;

   // m271_50 = W*in
   wire signed [9:0] m271_50;
   assign m271_50 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_51 = W*in
   wire signed [9:0] m271_51;
   assign m271_51 =10'b0;

   // m271_52 = W*in
   wire signed [9:0] m271_52;
   assign m271_52 =10'b0;

   // m271_53 = W*in
   wire signed [9:0] m271_53;
   assign m271_53 ={ {4{in271[5]}} , in271[5:0] };

   // m271_54 = W*in
   wire signed [9:0] m271_54;
   assign m271_54 ={ {4{in271[5]}} , in271[5:0] };

   // m271_55 = W*in
   wire signed [9:0] m271_55;
   assign m271_55 ={ {4{in271[5]}} , in271[5:0] };

   // m271_56 = W*in
   wire signed [9:0] m271_56;
   assign m271_56 =10'b0;

   // m271_57 = W*in
   wire signed [9:0] m271_57;
   assign m271_57 =10'b0;

   // m271_58 = W*in
   wire signed [9:0] m271_58;
   assign m271_58 =10'b0;

   // m271_59 = W*in
   wire signed [9:0] m271_59;
   assign m271_59 =10'b0;

   // m271_60 = W*in
   wire signed [9:0] m271_60;
   assign m271_60 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_61 = W*in
   wire signed [9:0] m271_61;
   assign m271_61 =10'b0;

   // m271_62 = W*in
   wire signed [9:0] m271_62;
   assign m271_62 =10'b0;

   // m271_63 = W*in
   wire signed [9:0] m271_63;
   assign m271_63 ={ {4{in271[5]}} , in271[5:0] };

   // m271_64 = W*in
   wire signed [9:0] m271_64;
   assign m271_64 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_65 = W*in
   wire signed [9:0] m271_65;
   assign m271_65 =10'b0;

   // m271_66 = W*in
   wire signed [9:0] m271_66;
   assign m271_66 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_67 = W*in
   wire signed [9:0] m271_67;
   assign m271_67 =10'b0;

   // m271_68 = W*in
   wire signed [9:0] m271_68;
   assign m271_68 =10'b0;

   // m271_69 = W*in
   wire signed [9:0] m271_69;
   assign m271_69 ={ {4{in271[5]}} , in271[5:0] };

   // m271_70 = W*in
   wire signed [9:0] m271_70;
   assign m271_70 =10'b0;

   // m271_71 = W*in
   wire signed [9:0] m271_71;
   assign m271_71 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_72 = W*in
   wire signed [9:0] m271_72;
   assign m271_72 ={ {4{in271[5]}} , in271[5:0] };

   // m271_73 = W*in
   wire signed [9:0] m271_73;
   assign m271_73 =10'b0;

   // m271_74 = W*in
   wire signed [9:0] m271_74;
   assign m271_74 =10'b0;

   // m271_75 = W*in
   wire signed [9:0] m271_75;
   assign m271_75 =10'b0;

   // m271_76 = W*in
   wire signed [9:0] m271_76;
   assign m271_76 =10'b0;

   // m271_77 = W*in
   wire signed [9:0] m271_77;
   assign m271_77 =10'b0;

   // m271_78 = W*in
   wire signed [9:0] m271_78;
   assign m271_78 ={ {4{in271[5]}} , in271[5:0] };

   // m271_79 = W*in
   wire signed [9:0] m271_79;
   assign m271_79 =10'b0;

   // m271_80 = W*in
   wire signed [9:0] m271_80;
   assign m271_80 =10'b0;

   // m271_81 = W*in
   wire signed [9:0] m271_81;
   assign m271_81 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_82 = W*in
   wire signed [9:0] m271_82;
   assign m271_82 =10'b0;

   // m271_83 = W*in
   wire signed [9:0] m271_83;
   assign m271_83 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_84 = W*in
   wire signed [9:0] m271_84;
   assign m271_84 ={ {4{in271[5]}} , in271[5:0] };

   // m271_85 = W*in
   wire signed [9:0] m271_85;
   assign m271_85 =10'b0;

   // m271_86 = W*in
   wire signed [9:0] m271_86;
   assign m271_86 =10'b0;

   // m271_87 = W*in
   wire signed [9:0] m271_87;
   assign m271_87 =10'b0;

   // m271_88 = W*in
   wire signed [9:0] m271_88;
   assign m271_88 =10'b0;

   // m271_89 = W*in
   wire signed [9:0] m271_89;
   assign m271_89 =10'b0;

   // m271_90 = W*in
   wire signed [9:0] m271_90;
   assign m271_90 =10'b0;

   // m271_91 = W*in
   wire signed [9:0] m271_91;
   assign m271_91 =10'b0;

   // m271_92 = W*in
   wire signed [9:0] m271_92;
   assign m271_92 =10'b0;

   // m271_93 = W*in
   wire signed [9:0] m271_93;
   assign m271_93 ={ {4{in271[5]}} , in271[5:0] };

   // m271_94 = W*in
   wire signed [9:0] m271_94;
   assign m271_94 =10'b0;

   // m271_95 = W*in
   wire signed [9:0] m271_95;
   assign m271_95 =10'b0;

   // m271_96 = W*in
   wire signed [9:0] m271_96;
   assign m271_96 =10'b0;

   // m271_97 = W*in
   wire signed [9:0] m271_97;
   assign m271_97 ={ {4{in271[5]}} , in271[5:0] };

   // m271_98 = W*in
   wire signed [9:0] m271_98;
   assign m271_98 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_99 = W*in
   wire signed [9:0] m271_99;
   assign m271_99 =10'b0;

   // m271_100 = W*in
   wire signed [9:0] m271_100;
   assign m271_100 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_101 = W*in
   wire signed [9:0] m271_101;
   assign m271_101 =10'b0;

   // m271_102 = W*in
   wire signed [9:0] m271_102;
   assign m271_102 ={ {4{in271[5]}} , in271[5:0] };

   // m271_103 = W*in
   wire signed [9:0] m271_103;
   assign m271_103 =10'b0;

   // m271_104 = W*in
   wire signed [9:0] m271_104;
   assign m271_104 =10'b0;

   // m271_105 = W*in
   wire signed [9:0] m271_105;
   assign m271_105 =10'b0;

   // m271_106 = W*in
   wire signed [9:0] m271_106;
   assign m271_106 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_107 = W*in
   wire signed [9:0] m271_107;
   assign m271_107 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_108 = W*in
   wire signed [9:0] m271_108;
   assign m271_108 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_109 = W*in
   wire signed [9:0] m271_109;
   assign m271_109 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_110 = W*in
   wire signed [9:0] m271_110;
   assign m271_110 =10'b0;

   // m271_111 = W*in
   wire signed [9:0] m271_111;
   assign m271_111 ={ {4{in271[5]}} , in271[5:0] };

   // m271_112 = W*in
   wire signed [9:0] m271_112;
   assign m271_112 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_113 = W*in
   wire signed [9:0] m271_113;
   assign m271_113 =10'b0;

   // m271_114 = W*in
   wire signed [9:0] m271_114;
   assign m271_114 ={ {5{neg271[5]}} , neg271[5:1] };

   // m271_115 = W*in
   wire signed [9:0] m271_115;
   assign m271_115 ={ {4{neg271[5]}} , neg271[5:0] };

   // m271_116 = W*in
   wire signed [9:0] m271_116;
   assign m271_116 =10'b0;

   // m271_117 = W*in
   wire signed [9:0] m271_117;
   assign m271_117 ={ {4{neg271[5]}} , neg271[5:0] };

   // m272_1 = W*in
   wire signed [9:0] m272_1;
   assign m272_1 =10'b0;

   // m272_2 = W*in
   wire signed [9:0] m272_2;
   assign m272_2 =10'b0;

   // m272_3 = W*in
   wire signed [9:0] m272_3;
   assign m272_3 =10'b0;

   // m272_4 = W*in
   wire signed [9:0] m272_4;
   assign m272_4 =10'b0;

   // m272_5 = W*in
   wire signed [9:0] m272_5;
   assign m272_5 =10'b0;

   // m272_6 = W*in
   wire signed [9:0] m272_6;
   assign m272_6 =10'b0;

   // m272_7 = W*in
   wire signed [9:0] m272_7;
   assign m272_7 =10'b0;

   // m272_8 = W*in
   wire signed [9:0] m272_8;
   assign m272_8 ={ {4{in272[5]}} , in272[5:0] };

   // m272_9 = W*in
   wire signed [9:0] m272_9;
   assign m272_9 =10'b0;

   // m272_10 = W*in
   wire signed [9:0] m272_10;
   assign m272_10 =10'b0;

   // m272_11 = W*in
   wire signed [9:0] m272_11;
   assign m272_11 =10'b0;

   // m272_12 = W*in
   wire signed [9:0] m272_12;
   assign m272_12 =10'b0;

   // m272_13 = W*in
   wire signed [9:0] m272_13;
   assign m272_13 =10'b0;

   // m272_14 = W*in
   wire signed [9:0] m272_14;
   assign m272_14 =10'b0;

   // m272_15 = W*in
   wire signed [9:0] m272_15;
   assign m272_15 =10'b0;

   // m272_16 = W*in
   wire signed [9:0] m272_16;
   assign m272_16 =10'b0;

   // m272_17 = W*in
   wire signed [9:0] m272_17;
   assign m272_17 =10'b0;

   // m272_18 = W*in
   wire signed [9:0] m272_18;
   assign m272_18 ={ {5{in272[5]}} , in272[5:1] };

   // m272_19 = W*in
   wire signed [9:0] m272_19;
   assign m272_19 ={ {5{in272[5]}} , in272[5:1] };

   // m272_20 = W*in
   wire signed [9:0] m272_20;
   assign m272_20 =10'b0;

   // m272_21 = W*in
   wire signed [9:0] m272_21;
   assign m272_21 ={ {5{neg272[5]}} , neg272[5:1] };

   // m272_22 = W*in
   wire signed [9:0] m272_22;
   assign m272_22 =10'b0;

   // m272_23 = W*in
   wire signed [9:0] m272_23;
   assign m272_23 =10'b0;

   // m272_24 = W*in
   wire signed [9:0] m272_24;
   assign m272_24 =10'b0;

   // m272_25 = W*in
   wire signed [9:0] m272_25;
   assign m272_25 =10'b0;

   // m272_26 = W*in
   wire signed [9:0] m272_26;
   assign m272_26 =10'b0;

   // m272_27 = W*in
   wire signed [9:0] m272_27;
   assign m272_27 ={ {5{neg272[5]}} , neg272[5:1] };

   // m272_28 = W*in
   wire signed [9:0] m272_28;
   assign m272_28 =10'b0;

   // m272_29 = W*in
   wire signed [9:0] m272_29;
   assign m272_29 =10'b0;

   // m272_30 = W*in
   wire signed [9:0] m272_30;
   assign m272_30 =10'b0;

   // m272_31 = W*in
   wire signed [9:0] m272_31;
   assign m272_31 ={ {5{in272[5]}} , in272[5:1] };

   // m272_32 = W*in
   wire signed [9:0] m272_32;
   assign m272_32 =10'b0;

   // m272_33 = W*in
   wire signed [9:0] m272_33;
   assign m272_33 =10'b0;

   // m272_34 = W*in
   wire signed [9:0] m272_34;
   assign m272_34 =10'b0;

   // m272_35 = W*in
   wire signed [9:0] m272_35;
   assign m272_35 =10'b0;

   // m272_36 = W*in
   wire signed [9:0] m272_36;
   assign m272_36 =10'b0;

   // m272_37 = W*in
   wire signed [9:0] m272_37;
   assign m272_37 =10'b0;

   // m272_38 = W*in
   wire signed [9:0] m272_38;
   assign m272_38 =10'b0;

   // m272_39 = W*in
   wire signed [9:0] m272_39;
   assign m272_39 =10'b0;

   // m272_40 = W*in
   wire signed [9:0] m272_40;
   assign m272_40 =10'b0;

   // m272_41 = W*in
   wire signed [9:0] m272_41;
   assign m272_41 =10'b0;

   // m272_42 = W*in
   wire signed [9:0] m272_42;
   assign m272_42 =10'b0;

   // m272_43 = W*in
   wire signed [9:0] m272_43;
   assign m272_43 =10'b0;

   // m272_44 = W*in
   wire signed [9:0] m272_44;
   assign m272_44 =10'b0;

   // m272_45 = W*in
   wire signed [9:0] m272_45;
   assign m272_45 =10'b0;

   // m272_46 = W*in
   wire signed [9:0] m272_46;
   assign m272_46 =10'b0;

   // m272_47 = W*in
   wire signed [9:0] m272_47;
   assign m272_47 =10'b0;

   // m272_48 = W*in
   wire signed [9:0] m272_48;
   assign m272_48 =10'b0;

   // m272_49 = W*in
   wire signed [9:0] m272_49;
   assign m272_49 ={ {4{in272[5]}} , in272[5:0] };

   // m272_50 = W*in
   wire signed [9:0] m272_50;
   assign m272_50 =10'b0;

   // m272_51 = W*in
   wire signed [9:0] m272_51;
   assign m272_51 ={ {4{in272[5]}} , in272[5:0] };

   // m272_52 = W*in
   wire signed [9:0] m272_52;
   assign m272_52 =10'b0;

   // m272_53 = W*in
   wire signed [9:0] m272_53;
   assign m272_53 =10'b0;

   // m272_54 = W*in
   wire signed [9:0] m272_54;
   assign m272_54 =10'b0;

   // m272_55 = W*in
   wire signed [9:0] m272_55;
   assign m272_55 =10'b0;

   // m272_56 = W*in
   wire signed [9:0] m272_56;
   assign m272_56 =10'b0;

   // m272_57 = W*in
   wire signed [9:0] m272_57;
   assign m272_57 =10'b0;

   // m272_58 = W*in
   wire signed [9:0] m272_58;
   assign m272_58 =10'b0;

   // m272_59 = W*in
   wire signed [9:0] m272_59;
   assign m272_59 =10'b0;

   // m272_60 = W*in
   wire signed [9:0] m272_60;
   assign m272_60 =10'b0;

   // m272_61 = W*in
   wire signed [9:0] m272_61;
   assign m272_61 =10'b0;

   // m272_62 = W*in
   wire signed [9:0] m272_62;
   assign m272_62 =10'b0;

   // m272_63 = W*in
   wire signed [9:0] m272_63;
   assign m272_63 =10'b0;

   // m272_64 = W*in
   wire signed [9:0] m272_64;
   assign m272_64 =10'b0;

   // m272_65 = W*in
   wire signed [9:0] m272_65;
   assign m272_65 =10'b0;

   // m272_66 = W*in
   wire signed [9:0] m272_66;
   assign m272_66 =10'b0;

   // m272_67 = W*in
   wire signed [9:0] m272_67;
   assign m272_67 ={ {5{in272[5]}} , in272[5:1] };

   // m272_68 = W*in
   wire signed [9:0] m272_68;
   assign m272_68 ={ {4{in272[5]}} , in272[5:0] };

   // m272_69 = W*in
   wire signed [9:0] m272_69;
   assign m272_69 ={ {4{neg272[5]}} , neg272[5:0] };

   // m272_70 = W*in
   wire signed [9:0] m272_70;
   assign m272_70 ={ {4{neg272[5]}} , neg272[5:0] };

   // m272_71 = W*in
   wire signed [9:0] m272_71;
   assign m272_71 ={ {5{neg272[5]}} , neg272[5:1] };

   // m272_72 = W*in
   wire signed [9:0] m272_72;
   assign m272_72 ={ {5{neg272[5]}} , neg272[5:1] };

   // m272_73 = W*in
   wire signed [9:0] m272_73;
   assign m272_73 ={ {4{in272[5]}} , in272[5:0] };

   // m272_74 = W*in
   wire signed [9:0] m272_74;
   assign m272_74 =10'b0;

   // m272_75 = W*in
   wire signed [9:0] m272_75;
   assign m272_75 =10'b0;

   // m272_76 = W*in
   wire signed [9:0] m272_76;
   assign m272_76 =10'b0;

   // m272_77 = W*in
   wire signed [9:0] m272_77;
   assign m272_77 =10'b0;

   // m272_78 = W*in
   wire signed [9:0] m272_78;
   assign m272_78 =10'b0;

   // m272_79 = W*in
   wire signed [9:0] m272_79;
   assign m272_79 =10'b0;

   // m272_80 = W*in
   wire signed [9:0] m272_80;
   assign m272_80 ={ {4{in272[5]}} , in272[5:0] };

   // m272_81 = W*in
   wire signed [9:0] m272_81;
   assign m272_81 =10'b0;

   // m272_82 = W*in
   wire signed [9:0] m272_82;
   assign m272_82 =10'b0;

   // m272_83 = W*in
   wire signed [9:0] m272_83;
   assign m272_83 =10'b0;

   // m272_84 = W*in
   wire signed [9:0] m272_84;
   assign m272_84 =10'b0;

   // m272_85 = W*in
   wire signed [9:0] m272_85;
   assign m272_85 =10'b0;

   // m272_86 = W*in
   wire signed [9:0] m272_86;
   assign m272_86 =10'b0;

   // m272_87 = W*in
   wire signed [9:0] m272_87;
   assign m272_87 =10'b0;

   // m272_88 = W*in
   wire signed [9:0] m272_88;
   assign m272_88 =10'b0;

   // m272_89 = W*in
   wire signed [9:0] m272_89;
   assign m272_89 =10'b0;

   // m272_90 = W*in
   wire signed [9:0] m272_90;
   assign m272_90 =10'b0;

   // m272_91 = W*in
   wire signed [9:0] m272_91;
   assign m272_91 =10'b0;

   // m272_92 = W*in
   wire signed [9:0] m272_92;
   assign m272_92 =10'b0;

   // m272_93 = W*in
   wire signed [9:0] m272_93;
   assign m272_93 =10'b0;

   // m272_94 = W*in
   wire signed [9:0] m272_94;
   assign m272_94 =10'b0;

   // m272_95 = W*in
   wire signed [9:0] m272_95;
   assign m272_95 =10'b0;

   // m272_96 = W*in
   wire signed [9:0] m272_96;
   assign m272_96 =10'b0;

   // m272_97 = W*in
   wire signed [9:0] m272_97;
   assign m272_97 =10'b0;

   // m272_98 = W*in
   wire signed [9:0] m272_98;
   assign m272_98 =10'b0;

   // m272_99 = W*in
   wire signed [9:0] m272_99;
   assign m272_99 =10'b0;

   // m272_100 = W*in
   wire signed [9:0] m272_100;
   assign m272_100 =10'b0;

   // m272_101 = W*in
   wire signed [9:0] m272_101;
   assign m272_101 =10'b0;

   // m272_102 = W*in
   wire signed [9:0] m272_102;
   assign m272_102 =10'b0;

   // m272_103 = W*in
   wire signed [9:0] m272_103;
   assign m272_103 =10'b0;

   // m272_104 = W*in
   wire signed [9:0] m272_104;
   assign m272_104 =10'b0;

   // m272_105 = W*in
   wire signed [9:0] m272_105;
   assign m272_105 =10'b0;

   // m272_106 = W*in
   wire signed [9:0] m272_106;
   assign m272_106 =10'b0;

   // m272_107 = W*in
   wire signed [9:0] m272_107;
   assign m272_107 =10'b0;

   // m272_108 = W*in
   wire signed [9:0] m272_108;
   assign m272_108 ={ {5{neg272[5]}} , neg272[5:1] };

   // m272_109 = W*in
   wire signed [9:0] m272_109;
   assign m272_109 =10'b0;

   // m272_110 = W*in
   wire signed [9:0] m272_110;
   assign m272_110 =10'b0;

   // m272_111 = W*in
   wire signed [9:0] m272_111;
   assign m272_111 =10'b0;

   // m272_112 = W*in
   wire signed [9:0] m272_112;
   assign m272_112 =10'b0;

   // m272_113 = W*in
   wire signed [9:0] m272_113;
   assign m272_113 =10'b0;

   // m272_114 = W*in
   wire signed [9:0] m272_114;
   assign m272_114 =10'b0;

   // m272_115 = W*in
   wire signed [9:0] m272_115;
   assign m272_115 =10'b0;

   // m272_116 = W*in
   wire signed [9:0] m272_116;
   assign m272_116 =10'b0;

   // m272_117 = W*in
   wire signed [9:0] m272_117;
   assign m272_117 =10'b0;

   // m273_1 = W*in
   wire signed [9:0] m273_1;
   assign m273_1 =10'b0;

   // m273_2 = W*in
   wire signed [9:0] m273_2;
   assign m273_2 =10'b0;

   // m273_3 = W*in
   wire signed [9:0] m273_3;
   assign m273_3 =10'b0;

   // m273_4 = W*in
   wire signed [9:0] m273_4;
   assign m273_4 =10'b0;

   // m273_5 = W*in
   wire signed [9:0] m273_5;
   assign m273_5 =10'b0;

   // m273_6 = W*in
   wire signed [9:0] m273_6;
   assign m273_6 =10'b0;

   // m273_7 = W*in
   wire signed [9:0] m273_7;
   assign m273_7 =10'b0;

   // m273_8 = W*in
   wire signed [9:0] m273_8;
   assign m273_8 =10'b0;

   // m273_9 = W*in
   wire signed [9:0] m273_9;
   assign m273_9 =10'b0;

   // m273_10 = W*in
   wire signed [9:0] m273_10;
   assign m273_10 =10'b0;

   // m273_11 = W*in
   wire signed [9:0] m273_11;
   assign m273_11 =10'b0;

   // m273_12 = W*in
   wire signed [9:0] m273_12;
   assign m273_12 ={ {4{in273[5]}} , in273[5:0] };

   // m273_13 = W*in
   wire signed [9:0] m273_13;
   assign m273_13 =10'b0;

   // m273_14 = W*in
   wire signed [9:0] m273_14;
   assign m273_14 =10'b0;

   // m273_15 = W*in
   wire signed [9:0] m273_15;
   assign m273_15 =10'b0;

   // m273_16 = W*in
   wire signed [9:0] m273_16;
   assign m273_16 =10'b0;

   // m273_17 = W*in
   wire signed [9:0] m273_17;
   assign m273_17 ={ {5{in273[5]}} , in273[5:1] };

   // m273_18 = W*in
   wire signed [9:0] m273_18;
   assign m273_18 =10'b0;

   // m273_19 = W*in
   wire signed [9:0] m273_19;
   assign m273_19 =10'b0;

   // m273_20 = W*in
   wire signed [9:0] m273_20;
   assign m273_20 =10'b0;

   // m273_21 = W*in
   wire signed [9:0] m273_21;
   assign m273_21 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_22 = W*in
   wire signed [9:0] m273_22;
   assign m273_22 =10'b0;

   // m273_23 = W*in
   wire signed [9:0] m273_23;
   assign m273_23 =10'b0;

   // m273_24 = W*in
   wire signed [9:0] m273_24;
   assign m273_24 =10'b0;

   // m273_25 = W*in
   wire signed [9:0] m273_25;
   assign m273_25 ={ {5{in273[5]}} , in273[5:1] };

   // m273_26 = W*in
   wire signed [9:0] m273_26;
   assign m273_26 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_27 = W*in
   wire signed [9:0] m273_27;
   assign m273_27 =10'b0;

   // m273_28 = W*in
   wire signed [9:0] m273_28;
   assign m273_28 ={ {5{in273[5]}} , in273[5:1] };

   // m273_29 = W*in
   wire signed [9:0] m273_29;
   assign m273_29 =10'b0;

   // m273_30 = W*in
   wire signed [9:0] m273_30;
   assign m273_30 =10'b0;

   // m273_31 = W*in
   wire signed [9:0] m273_31;
   assign m273_31 ={ {5{in273[5]}} , in273[5:1] };

   // m273_32 = W*in
   wire signed [9:0] m273_32;
   assign m273_32 =10'b0;

   // m273_33 = W*in
   wire signed [9:0] m273_33;
   assign m273_33 =10'b0;

   // m273_34 = W*in
   wire signed [9:0] m273_34;
   assign m273_34 =10'b0;

   // m273_35 = W*in
   wire signed [9:0] m273_35;
   assign m273_35 =10'b0;

   // m273_36 = W*in
   wire signed [9:0] m273_36;
   assign m273_36 ={ {4{in273[5]}} , in273[5:0] };

   // m273_37 = W*in
   wire signed [9:0] m273_37;
   assign m273_37 =10'b0;

   // m273_38 = W*in
   wire signed [9:0] m273_38;
   assign m273_38 =10'b0;

   // m273_39 = W*in
   wire signed [9:0] m273_39;
   assign m273_39 =10'b0;

   // m273_40 = W*in
   wire signed [9:0] m273_40;
   assign m273_40 =10'b0;

   // m273_41 = W*in
   wire signed [9:0] m273_41;
   assign m273_41 =10'b0;

   // m273_42 = W*in
   wire signed [9:0] m273_42;
   assign m273_42 =10'b0;

   // m273_43 = W*in
   wire signed [9:0] m273_43;
   assign m273_43 =10'b0;

   // m273_44 = W*in
   wire signed [9:0] m273_44;
   assign m273_44 =10'b0;

   // m273_45 = W*in
   wire signed [9:0] m273_45;
   assign m273_45 =10'b0;

   // m273_46 = W*in
   wire signed [9:0] m273_46;
   assign m273_46 =10'b0;

   // m273_47 = W*in
   wire signed [9:0] m273_47;
   assign m273_47 =10'b0;

   // m273_48 = W*in
   wire signed [9:0] m273_48;
   assign m273_48 =10'b0;

   // m273_49 = W*in
   wire signed [9:0] m273_49;
   assign m273_49 =10'b0;

   // m273_50 = W*in
   wire signed [9:0] m273_50;
   assign m273_50 =10'b0;

   // m273_51 = W*in
   wire signed [9:0] m273_51;
   assign m273_51 ={ {4{in273[5]}} , in273[5:0] };

   // m273_52 = W*in
   wire signed [9:0] m273_52;
   assign m273_52 =10'b0;

   // m273_53 = W*in
   wire signed [9:0] m273_53;
   assign m273_53 =10'b0;

   // m273_54 = W*in
   wire signed [9:0] m273_54;
   assign m273_54 =10'b0;

   // m273_55 = W*in
   wire signed [9:0] m273_55;
   assign m273_55 =10'b0;

   // m273_56 = W*in
   wire signed [9:0] m273_56;
   assign m273_56 =10'b0;

   // m273_57 = W*in
   wire signed [9:0] m273_57;
   assign m273_57 =10'b0;

   // m273_58 = W*in
   wire signed [9:0] m273_58;
   assign m273_58 =10'b0;

   // m273_59 = W*in
   wire signed [9:0] m273_59;
   assign m273_59 =10'b0;

   // m273_60 = W*in
   wire signed [9:0] m273_60;
   assign m273_60 =10'b0;

   // m273_61 = W*in
   wire signed [9:0] m273_61;
   assign m273_61 =10'b0;

   // m273_62 = W*in
   wire signed [9:0] m273_62;
   assign m273_62 =10'b0;

   // m273_63 = W*in
   wire signed [9:0] m273_63;
   assign m273_63 =10'b0;

   // m273_64 = W*in
   wire signed [9:0] m273_64;
   assign m273_64 =10'b0;

   // m273_65 = W*in
   wire signed [9:0] m273_65;
   assign m273_65 =10'b0;

   // m273_66 = W*in
   wire signed [9:0] m273_66;
   assign m273_66 ={ {5{in273[5]}} , in273[5:1] };

   // m273_67 = W*in
   wire signed [9:0] m273_67;
   assign m273_67 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_68 = W*in
   wire signed [9:0] m273_68;
   assign m273_68 =10'b0;

   // m273_69 = W*in
   wire signed [9:0] m273_69;
   assign m273_69 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_70 = W*in
   wire signed [9:0] m273_70;
   assign m273_70 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_71 = W*in
   wire signed [9:0] m273_71;
   assign m273_71 =10'b0;

   // m273_72 = W*in
   wire signed [9:0] m273_72;
   assign m273_72 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_73 = W*in
   wire signed [9:0] m273_73;
   assign m273_73 ={ {4{in273[5]}} , in273[5:0] };

   // m273_74 = W*in
   wire signed [9:0] m273_74;
   assign m273_74 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_75 = W*in
   wire signed [9:0] m273_75;
   assign m273_75 =10'b0;

   // m273_76 = W*in
   wire signed [9:0] m273_76;
   assign m273_76 ={ {4{neg273[5]}} , neg273[5:0] };

   // m273_77 = W*in
   wire signed [9:0] m273_77;
   assign m273_77 =10'b0;

   // m273_78 = W*in
   wire signed [9:0] m273_78;
   assign m273_78 =10'b0;

   // m273_79 = W*in
   wire signed [9:0] m273_79;
   assign m273_79 =10'b0;

   // m273_80 = W*in
   wire signed [9:0] m273_80;
   assign m273_80 =10'b0;

   // m273_81 = W*in
   wire signed [9:0] m273_81;
   assign m273_81 ={ {5{neg273[5]}} , neg273[5:1] };

   // m273_82 = W*in
   wire signed [9:0] m273_82;
   assign m273_82 =10'b0;

   // m273_83 = W*in
   wire signed [9:0] m273_83;
   assign m273_83 =10'b0;

   // m273_84 = W*in
   wire signed [9:0] m273_84;
   assign m273_84 =10'b0;

   // m273_85 = W*in
   wire signed [9:0] m273_85;
   assign m273_85 =10'b0;

   // m273_86 = W*in
   wire signed [9:0] m273_86;
   assign m273_86 =10'b0;

   // m273_87 = W*in
   wire signed [9:0] m273_87;
   assign m273_87 =10'b0;

   // m273_88 = W*in
   wire signed [9:0] m273_88;
   assign m273_88 =10'b0;

   // m273_89 = W*in
   wire signed [9:0] m273_89;
   assign m273_89 =10'b0;

   // m273_90 = W*in
   wire signed [9:0] m273_90;
   assign m273_90 =10'b0;

   // m273_91 = W*in
   wire signed [9:0] m273_91;
   assign m273_91 =10'b0;

   // m273_92 = W*in
   wire signed [9:0] m273_92;
   assign m273_92 =10'b0;

   // m273_93 = W*in
   wire signed [9:0] m273_93;
   assign m273_93 =10'b0;

   // m273_94 = W*in
   wire signed [9:0] m273_94;
   assign m273_94 =10'b0;

   // m273_95 = W*in
   wire signed [9:0] m273_95;
   assign m273_95 =10'b0;

   // m273_96 = W*in
   wire signed [9:0] m273_96;
   assign m273_96 =10'b0;

   // m273_97 = W*in
   wire signed [9:0] m273_97;
   assign m273_97 =10'b0;

   // m273_98 = W*in
   wire signed [9:0] m273_98;
   assign m273_98 =10'b0;

   // m273_99 = W*in
   wire signed [9:0] m273_99;
   assign m273_99 =10'b0;

   // m273_100 = W*in
   wire signed [9:0] m273_100;
   assign m273_100 =10'b0;

   // m273_101 = W*in
   wire signed [9:0] m273_101;
   assign m273_101 =10'b0;

   // m273_102 = W*in
   wire signed [9:0] m273_102;
   assign m273_102 =10'b0;

   // m273_103 = W*in
   wire signed [9:0] m273_103;
   assign m273_103 =10'b0;

   // m273_104 = W*in
   wire signed [9:0] m273_104;
   assign m273_104 =10'b0;

   // m273_105 = W*in
   wire signed [9:0] m273_105;
   assign m273_105 =10'b0;

   // m273_106 = W*in
   wire signed [9:0] m273_106;
   assign m273_106 =10'b0;

   // m273_107 = W*in
   wire signed [9:0] m273_107;
   assign m273_107 ={ {4{in273[5]}} , in273[5:0] };

   // m273_108 = W*in
   wire signed [9:0] m273_108;
   assign m273_108 =10'b0;

   // m273_109 = W*in
   wire signed [9:0] m273_109;
   assign m273_109 =10'b0;

   // m273_110 = W*in
   wire signed [9:0] m273_110;
   assign m273_110 =10'b0;

   // m273_111 = W*in
   wire signed [9:0] m273_111;
   assign m273_111 =10'b0;

   // m273_112 = W*in
   wire signed [9:0] m273_112;
   assign m273_112 =10'b0;

   // m273_113 = W*in
   wire signed [9:0] m273_113;
   assign m273_113 =10'b0;

   // m273_114 = W*in
   wire signed [9:0] m273_114;
   assign m273_114 =10'b0;

   // m273_115 = W*in
   wire signed [9:0] m273_115;
   assign m273_115 =10'b0;

   // m273_116 = W*in
   wire signed [9:0] m273_116;
   assign m273_116 =10'b0;

   // m273_117 = W*in
   wire signed [9:0] m273_117;
   assign m273_117 =10'b0;

   // m274_1 = W*in
   wire signed [9:0] m274_1;
   assign m274_1 =10'b0;

   // m274_2 = W*in
   wire signed [9:0] m274_2;
   assign m274_2 =10'b0;

   // m274_3 = W*in
   wire signed [9:0] m274_3;
   assign m274_3 =10'b0;

   // m274_4 = W*in
   wire signed [9:0] m274_4;
   assign m274_4 =10'b0;

   // m274_5 = W*in
   wire signed [9:0] m274_5;
   assign m274_5 =10'b0;

   // m274_6 = W*in
   wire signed [9:0] m274_6;
   assign m274_6 =10'b0;

   // m274_7 = W*in
   wire signed [9:0] m274_7;
   assign m274_7 =10'b0;

   // m274_8 = W*in
   wire signed [9:0] m274_8;
   assign m274_8 =10'b0;

   // m274_9 = W*in
   wire signed [9:0] m274_9;
   assign m274_9 =10'b0;

   // m274_10 = W*in
   wire signed [9:0] m274_10;
   assign m274_10 =10'b0;

   // m274_11 = W*in
   wire signed [9:0] m274_11;
   assign m274_11 =10'b0;

   // m274_12 = W*in
   wire signed [9:0] m274_12;
   assign m274_12 ={ {4{neg274[5]}} , neg274[5:0] };

   // m274_13 = W*in
   wire signed [9:0] m274_13;
   assign m274_13 =10'b0;

   // m274_14 = W*in
   wire signed [9:0] m274_14;
   assign m274_14 =10'b0;

   // m274_15 = W*in
   wire signed [9:0] m274_15;
   assign m274_15 =10'b0;

   // m274_16 = W*in
   wire signed [9:0] m274_16;
   assign m274_16 =10'b0;

   // m274_17 = W*in
   wire signed [9:0] m274_17;
   assign m274_17 =10'b0;

   // m274_18 = W*in
   wire signed [9:0] m274_18;
   assign m274_18 =10'b0;

   // m274_19 = W*in
   wire signed [9:0] m274_19;
   assign m274_19 ={ {5{neg274[5]}} , neg274[5:1] };

   // m274_20 = W*in
   wire signed [9:0] m274_20;
   assign m274_20 =10'b0;

   // m274_21 = W*in
   wire signed [9:0] m274_21;
   assign m274_21 ={ {5{in274[5]}} , in274[5:1] };

   // m274_22 = W*in
   wire signed [9:0] m274_22;
   assign m274_22 =10'b0;

   // m274_23 = W*in
   wire signed [9:0] m274_23;
   assign m274_23 =10'b0;

   // m274_24 = W*in
   wire signed [9:0] m274_24;
   assign m274_24 =10'b0;

   // m274_25 = W*in
   wire signed [9:0] m274_25;
   assign m274_25 =10'b0;

   // m274_26 = W*in
   wire signed [9:0] m274_26;
   assign m274_26 =10'b0;

   // m274_27 = W*in
   wire signed [9:0] m274_27;
   assign m274_27 =10'b0;

   // m274_28 = W*in
   wire signed [9:0] m274_28;
   assign m274_28 ={ {5{neg274[5]}} , neg274[5:1] };

   // m274_29 = W*in
   wire signed [9:0] m274_29;
   assign m274_29 =10'b0;

   // m274_30 = W*in
   wire signed [9:0] m274_30;
   assign m274_30 =10'b0;

   // m274_31 = W*in
   wire signed [9:0] m274_31;
   assign m274_31 =10'b0;

   // m274_32 = W*in
   wire signed [9:0] m274_32;
   assign m274_32 =10'b0;

   // m274_33 = W*in
   wire signed [9:0] m274_33;
   assign m274_33 =10'b0;

   // m274_34 = W*in
   wire signed [9:0] m274_34;
   assign m274_34 =10'b0;

   // m274_35 = W*in
   wire signed [9:0] m274_35;
   assign m274_35 ={ {5{neg274[5]}} , neg274[5:1] };

   // m274_36 = W*in
   wire signed [9:0] m274_36;
   assign m274_36 =10'b0;

   // m274_37 = W*in
   wire signed [9:0] m274_37;
   assign m274_37 =10'b0;

   // m274_38 = W*in
   wire signed [9:0] m274_38;
   assign m274_38 =10'b0;

   // m274_39 = W*in
   wire signed [9:0] m274_39;
   assign m274_39 =10'b0;

   // m274_40 = W*in
   wire signed [9:0] m274_40;
   assign m274_40 =10'b0;

   // m274_41 = W*in
   wire signed [9:0] m274_41;
   assign m274_41 =10'b0;

   // m274_42 = W*in
   wire signed [9:0] m274_42;
   assign m274_42 =10'b0;

   // m274_43 = W*in
   wire signed [9:0] m274_43;
   assign m274_43 =10'b0;

   // m274_44 = W*in
   wire signed [9:0] m274_44;
   assign m274_44 =10'b0;

   // m274_45 = W*in
   wire signed [9:0] m274_45;
   assign m274_45 ={ {4{in274[5]}} , in274[5:0] };

   // m274_46 = W*in
   wire signed [9:0] m274_46;
   assign m274_46 =10'b0;

   // m274_47 = W*in
   wire signed [9:0] m274_47;
   assign m274_47 =10'b0;

   // m274_48 = W*in
   wire signed [9:0] m274_48;
   assign m274_48 =10'b0;

   // m274_49 = W*in
   wire signed [9:0] m274_49;
   assign m274_49 =10'b0;

   // m274_50 = W*in
   wire signed [9:0] m274_50;
   assign m274_50 =10'b0;

   // m274_51 = W*in
   wire signed [9:0] m274_51;
   assign m274_51 ={ {4{in274[5]}} , in274[5:0] };

   // m274_52 = W*in
   wire signed [9:0] m274_52;
   assign m274_52 =10'b0;

   // m274_53 = W*in
   wire signed [9:0] m274_53;
   assign m274_53 =10'b0;

   // m274_54 = W*in
   wire signed [9:0] m274_54;
   assign m274_54 =10'b0;

   // m274_55 = W*in
   wire signed [9:0] m274_55;
   assign m274_55 =10'b0;

   // m274_56 = W*in
   wire signed [9:0] m274_56;
   assign m274_56 =10'b0;

   // m274_57 = W*in
   wire signed [9:0] m274_57;
   assign m274_57 =10'b0;

   // m274_58 = W*in
   wire signed [9:0] m274_58;
   assign m274_58 =10'b0;

   // m274_59 = W*in
   wire signed [9:0] m274_59;
   assign m274_59 =10'b0;

   // m274_60 = W*in
   wire signed [9:0] m274_60;
   assign m274_60 =10'b0;

   // m274_61 = W*in
   wire signed [9:0] m274_61;
   assign m274_61 =10'b0;

   // m274_62 = W*in
   wire signed [9:0] m274_62;
   assign m274_62 =10'b0;

   // m274_63 = W*in
   wire signed [9:0] m274_63;
   assign m274_63 ={ {4{in274[5]}} , in274[5:0] };

   // m274_64 = W*in
   wire signed [9:0] m274_64;
   assign m274_64 ={ {5{neg274[5]}} , neg274[5:1] };

   // m274_65 = W*in
   wire signed [9:0] m274_65;
   assign m274_65 ={ {5{neg274[5]}} , neg274[5:1] };

   // m274_66 = W*in
   wire signed [9:0] m274_66;
   assign m274_66 ={ {5{neg274[5]}} , neg274[5:1] };

   // m274_67 = W*in
   wire signed [9:0] m274_67;
   assign m274_67 =10'b0;

   // m274_68 = W*in
   wire signed [9:0] m274_68;
   assign m274_68 =10'b0;

   // m274_69 = W*in
   wire signed [9:0] m274_69;
   assign m274_69 ={ {5{in274[5]}} , in274[5:1] };

   // m274_70 = W*in
   wire signed [9:0] m274_70;
   assign m274_70 =10'b0;

   // m274_71 = W*in
   wire signed [9:0] m274_71;
   assign m274_71 =10'b0;

   // m274_72 = W*in
   wire signed [9:0] m274_72;
   assign m274_72 =10'b0;

   // m274_73 = W*in
   wire signed [9:0] m274_73;
   assign m274_73 =10'b0;

   // m274_74 = W*in
   wire signed [9:0] m274_74;
   assign m274_74 =10'b0;

   // m274_75 = W*in
   wire signed [9:0] m274_75;
   assign m274_75 =10'b0;

   // m274_76 = W*in
   wire signed [9:0] m274_76;
   assign m274_76 =10'b0;

   // m274_77 = W*in
   wire signed [9:0] m274_77;
   assign m274_77 =10'b0;

   // m274_78 = W*in
   wire signed [9:0] m274_78;
   assign m274_78 ={ {5{in274[5]}} , in274[5:1] };

   // m274_79 = W*in
   wire signed [9:0] m274_79;
   assign m274_79 =10'b0;

   // m274_80 = W*in
   wire signed [9:0] m274_80;
   assign m274_80 =10'b0;

   // m274_81 = W*in
   wire signed [9:0] m274_81;
   assign m274_81 =10'b0;

   // m274_82 = W*in
   wire signed [9:0] m274_82;
   assign m274_82 =10'b0;

   // m274_83 = W*in
   wire signed [9:0] m274_83;
   assign m274_83 =10'b0;

   // m274_84 = W*in
   wire signed [9:0] m274_84;
   assign m274_84 =10'b0;

   // m274_85 = W*in
   wire signed [9:0] m274_85;
   assign m274_85 ={ {4{in274[5]}} , in274[5:0] };

   // m274_86 = W*in
   wire signed [9:0] m274_86;
   assign m274_86 =10'b0;

   // m274_87 = W*in
   wire signed [9:0] m274_87;
   assign m274_87 =10'b0;

   // m274_88 = W*in
   wire signed [9:0] m274_88;
   assign m274_88 =10'b0;

   // m274_89 = W*in
   wire signed [9:0] m274_89;
   assign m274_89 =10'b0;

   // m274_90 = W*in
   wire signed [9:0] m274_90;
   assign m274_90 =10'b0;

   // m274_91 = W*in
   wire signed [9:0] m274_91;
   assign m274_91 =10'b0;

   // m274_92 = W*in
   wire signed [9:0] m274_92;
   assign m274_92 =10'b0;

   // m274_93 = W*in
   wire signed [9:0] m274_93;
   assign m274_93 =10'b0;

   // m274_94 = W*in
   wire signed [9:0] m274_94;
   assign m274_94 =10'b0;

   // m274_95 = W*in
   wire signed [9:0] m274_95;
   assign m274_95 =10'b0;

   // m274_96 = W*in
   wire signed [9:0] m274_96;
   assign m274_96 =10'b0;

   // m274_97 = W*in
   wire signed [9:0] m274_97;
   assign m274_97 =10'b0;

   // m274_98 = W*in
   wire signed [9:0] m274_98;
   assign m274_98 =10'b0;

   // m274_99 = W*in
   wire signed [9:0] m274_99;
   assign m274_99 =10'b0;

   // m274_100 = W*in
   wire signed [9:0] m274_100;
   assign m274_100 =10'b0;

   // m274_101 = W*in
   wire signed [9:0] m274_101;
   assign m274_101 =10'b0;

   // m274_102 = W*in
   wire signed [9:0] m274_102;
   assign m274_102 =10'b0;

   // m274_103 = W*in
   wire signed [9:0] m274_103;
   assign m274_103 =10'b0;

   // m274_104 = W*in
   wire signed [9:0] m274_104;
   assign m274_104 =10'b0;

   // m274_105 = W*in
   wire signed [9:0] m274_105;
   assign m274_105 =10'b0;

   // m274_106 = W*in
   wire signed [9:0] m274_106;
   assign m274_106 =10'b0;

   // m274_107 = W*in
   wire signed [9:0] m274_107;
   assign m274_107 =10'b0;

   // m274_108 = W*in
   wire signed [9:0] m274_108;
   assign m274_108 =10'b0;

   // m274_109 = W*in
   wire signed [9:0] m274_109;
   assign m274_109 =10'b0;

   // m274_110 = W*in
   wire signed [9:0] m274_110;
   assign m274_110 =10'b0;

   // m274_111 = W*in
   wire signed [9:0] m274_111;
   assign m274_111 =10'b0;

   // m274_112 = W*in
   wire signed [9:0] m274_112;
   assign m274_112 =10'b0;

   // m274_113 = W*in
   wire signed [9:0] m274_113;
   assign m274_113 =10'b0;

   // m274_114 = W*in
   wire signed [9:0] m274_114;
   assign m274_114 =10'b0;

   // m274_115 = W*in
   wire signed [9:0] m274_115;
   assign m274_115 =10'b0;

   // m274_116 = W*in
   wire signed [9:0] m274_116;
   assign m274_116 =10'b0;

   // m274_117 = W*in
   wire signed [9:0] m274_117;
   assign m274_117 =10'b0;

   // m275_1 = W*in
   wire signed [9:0] m275_1;
   assign m275_1 =10'b0;

   // m275_2 = W*in
   wire signed [9:0] m275_2;
   assign m275_2 =10'b0;

   // m275_3 = W*in
   wire signed [9:0] m275_3;
   assign m275_3 =10'b0;

   // m275_4 = W*in
   wire signed [9:0] m275_4;
   assign m275_4 =10'b0;

   // m275_5 = W*in
   wire signed [9:0] m275_5;
   assign m275_5 =10'b0;

   // m275_6 = W*in
   wire signed [9:0] m275_6;
   assign m275_6 ={ {4{in275[5]}} , in275[5:0] };

   // m275_7 = W*in
   wire signed [9:0] m275_7;
   assign m275_7 =10'b0;

   // m275_8 = W*in
   wire signed [9:0] m275_8;
   assign m275_8 =10'b0;

   // m275_9 = W*in
   wire signed [9:0] m275_9;
   assign m275_9 =10'b0;

   // m275_10 = W*in
   wire signed [9:0] m275_10;
   assign m275_10 =10'b0;

   // m275_11 = W*in
   wire signed [9:0] m275_11;
   assign m275_11 =10'b0;

   // m275_12 = W*in
   wire signed [9:0] m275_12;
   assign m275_12 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_13 = W*in
   wire signed [9:0] m275_13;
   assign m275_13 =10'b0;

   // m275_14 = W*in
   wire signed [9:0] m275_14;
   assign m275_14 =10'b0;

   // m275_15 = W*in
   wire signed [9:0] m275_15;
   assign m275_15 ={ {4{in275[5]}} , in275[5:0] };

   // m275_16 = W*in
   wire signed [9:0] m275_16;
   assign m275_16 =10'b0;

   // m275_17 = W*in
   wire signed [9:0] m275_17;
   assign m275_17 =10'b0;

   // m275_18 = W*in
   wire signed [9:0] m275_18;
   assign m275_18 =10'b0;

   // m275_19 = W*in
   wire signed [9:0] m275_19;
   assign m275_19 =10'b0;

   // m275_20 = W*in
   wire signed [9:0] m275_20;
   assign m275_20 =10'b0;

   // m275_21 = W*in
   wire signed [9:0] m275_21;
   assign m275_21 ={ {5{in275[5]}} , in275[5:1] };

   // m275_22 = W*in
   wire signed [9:0] m275_22;
   assign m275_22 =10'b0;

   // m275_23 = W*in
   wire signed [9:0] m275_23;
   assign m275_23 =10'b0;

   // m275_24 = W*in
   wire signed [9:0] m275_24;
   assign m275_24 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_25 = W*in
   wire signed [9:0] m275_25;
   assign m275_25 =10'b0;

   // m275_26 = W*in
   wire signed [9:0] m275_26;
   assign m275_26 =10'b0;

   // m275_27 = W*in
   wire signed [9:0] m275_27;
   assign m275_27 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_28 = W*in
   wire signed [9:0] m275_28;
   assign m275_28 =10'b0;

   // m275_29 = W*in
   wire signed [9:0] m275_29;
   assign m275_29 =10'b0;

   // m275_30 = W*in
   wire signed [9:0] m275_30;
   assign m275_30 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_31 = W*in
   wire signed [9:0] m275_31;
   assign m275_31 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_32 = W*in
   wire signed [9:0] m275_32;
   assign m275_32 =10'b0;

   // m275_33 = W*in
   wire signed [9:0] m275_33;
   assign m275_33 =10'b0;

   // m275_34 = W*in
   wire signed [9:0] m275_34;
   assign m275_34 =10'b0;

   // m275_35 = W*in
   wire signed [9:0] m275_35;
   assign m275_35 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_36 = W*in
   wire signed [9:0] m275_36;
   assign m275_36 ={ {5{in275[5]}} , in275[5:1] };

   // m275_37 = W*in
   wire signed [9:0] m275_37;
   assign m275_37 ={ {4{in275[5]}} , in275[5:0] };

   // m275_38 = W*in
   wire signed [9:0] m275_38;
   assign m275_38 ={ {4{in275[5]}} , in275[5:0] };

   // m275_39 = W*in
   wire signed [9:0] m275_39;
   assign m275_39 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_40 = W*in
   wire signed [9:0] m275_40;
   assign m275_40 =10'b0;

   // m275_41 = W*in
   wire signed [9:0] m275_41;
   assign m275_41 =10'b0;

   // m275_42 = W*in
   wire signed [9:0] m275_42;
   assign m275_42 =10'b0;

   // m275_43 = W*in
   wire signed [9:0] m275_43;
   assign m275_43 ={ {4{in275[5]}} , in275[5:0] };

   // m275_44 = W*in
   wire signed [9:0] m275_44;
   assign m275_44 =10'b0;

   // m275_45 = W*in
   wire signed [9:0] m275_45;
   assign m275_45 ={ {4{in275[5]}} , in275[5:0] };

   // m275_46 = W*in
   wire signed [9:0] m275_46;
   assign m275_46 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_47 = W*in
   wire signed [9:0] m275_47;
   assign m275_47 ={ {4{in275[5]}} , in275[5:0] };

   // m275_48 = W*in
   wire signed [9:0] m275_48;
   assign m275_48 ={ {4{in275[5]}} , in275[5:0] };

   // m275_49 = W*in
   wire signed [9:0] m275_49;
   assign m275_49 =10'b0;

   // m275_50 = W*in
   wire signed [9:0] m275_50;
   assign m275_50 ={ {4{in275[5]}} , in275[5:0] };

   // m275_51 = W*in
   wire signed [9:0] m275_51;
   assign m275_51 =10'b0;

   // m275_52 = W*in
   wire signed [9:0] m275_52;
   assign m275_52 =10'b0;

   // m275_53 = W*in
   wire signed [9:0] m275_53;
   assign m275_53 =10'b0;

   // m275_54 = W*in
   wire signed [9:0] m275_54;
   assign m275_54 =10'b0;

   // m275_55 = W*in
   wire signed [9:0] m275_55;
   assign m275_55 =10'b0;

   // m275_56 = W*in
   wire signed [9:0] m275_56;
   assign m275_56 =10'b0;

   // m275_57 = W*in
   wire signed [9:0] m275_57;
   assign m275_57 =10'b0;

   // m275_58 = W*in
   wire signed [9:0] m275_58;
   assign m275_58 =10'b0;

   // m275_59 = W*in
   wire signed [9:0] m275_59;
   assign m275_59 =10'b0;

   // m275_60 = W*in
   wire signed [9:0] m275_60;
   assign m275_60 =10'b0;

   // m275_61 = W*in
   wire signed [9:0] m275_61;
   assign m275_61 =10'b0;

   // m275_62 = W*in
   wire signed [9:0] m275_62;
   assign m275_62 =10'b0;

   // m275_63 = W*in
   wire signed [9:0] m275_63;
   assign m275_63 ={ {4{in275[5]}} , in275[5:0] };

   // m275_64 = W*in
   wire signed [9:0] m275_64;
   assign m275_64 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_65 = W*in
   wire signed [9:0] m275_65;
   assign m275_65 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_66 = W*in
   wire signed [9:0] m275_66;
   assign m275_66 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_67 = W*in
   wire signed [9:0] m275_67;
   assign m275_67 =10'b0;

   // m275_68 = W*in
   wire signed [9:0] m275_68;
   assign m275_68 =10'b0;

   // m275_69 = W*in
   wire signed [9:0] m275_69;
   assign m275_69 ={ {4{in275[5]}} , in275[5:0] };

   // m275_70 = W*in
   wire signed [9:0] m275_70;
   assign m275_70 ={ {5{in275[5]}} , in275[5:1] };

   // m275_71 = W*in
   wire signed [9:0] m275_71;
   assign m275_71 ={ {5{in275[5]}} , in275[5:1] };

   // m275_72 = W*in
   wire signed [9:0] m275_72;
   assign m275_72 ={ {4{in275[5]}} , in275[5:0] };

   // m275_73 = W*in
   wire signed [9:0] m275_73;
   assign m275_73 =10'b0;

   // m275_74 = W*in
   wire signed [9:0] m275_74;
   assign m275_74 =10'b0;

   // m275_75 = W*in
   wire signed [9:0] m275_75;
   assign m275_75 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_76 = W*in
   wire signed [9:0] m275_76;
   assign m275_76 ={ {4{in275[5]}} , in275[5:0] };

   // m275_77 = W*in
   wire signed [9:0] m275_77;
   assign m275_77 =10'b0;

   // m275_78 = W*in
   wire signed [9:0] m275_78;
   assign m275_78 ={ {4{in275[5]}} , in275[5:0] };

   // m275_79 = W*in
   wire signed [9:0] m275_79;
   assign m275_79 =10'b0;

   // m275_80 = W*in
   wire signed [9:0] m275_80;
   assign m275_80 =10'b0;

   // m275_81 = W*in
   wire signed [9:0] m275_81;
   assign m275_81 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_82 = W*in
   wire signed [9:0] m275_82;
   assign m275_82 ={ {4{in275[5]}} , in275[5:0] };

   // m275_83 = W*in
   wire signed [9:0] m275_83;
   assign m275_83 =10'b0;

   // m275_84 = W*in
   wire signed [9:0] m275_84;
   assign m275_84 =10'b0;

   // m275_85 = W*in
   wire signed [9:0] m275_85;
   assign m275_85 ={ {5{in275[5]}} , in275[5:1] };

   // m275_86 = W*in
   wire signed [9:0] m275_86;
   assign m275_86 =10'b0;

   // m275_87 = W*in
   wire signed [9:0] m275_87;
   assign m275_87 ={ {4{in275[5]}} , in275[5:0] };

   // m275_88 = W*in
   wire signed [9:0] m275_88;
   assign m275_88 ={ {4{in275[5]}} , in275[5:0] };

   // m275_89 = W*in
   wire signed [9:0] m275_89;
   assign m275_89 =10'b0;

   // m275_90 = W*in
   wire signed [9:0] m275_90;
   assign m275_90 =10'b0;

   // m275_91 = W*in
   wire signed [9:0] m275_91;
   assign m275_91 =10'b0;

   // m275_92 = W*in
   wire signed [9:0] m275_92;
   assign m275_92 ={ {4{in275[5]}} , in275[5:0] };

   // m275_93 = W*in
   wire signed [9:0] m275_93;
   assign m275_93 =10'b0;

   // m275_94 = W*in
   wire signed [9:0] m275_94;
   assign m275_94 =10'b0;

   // m275_95 = W*in
   wire signed [9:0] m275_95;
   assign m275_95 =10'b0;

   // m275_96 = W*in
   wire signed [9:0] m275_96;
   assign m275_96 =10'b0;

   // m275_97 = W*in
   wire signed [9:0] m275_97;
   assign m275_97 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_98 = W*in
   wire signed [9:0] m275_98;
   assign m275_98 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_99 = W*in
   wire signed [9:0] m275_99;
   assign m275_99 ={ {4{in275[5]}} , in275[5:0] };

   // m275_100 = W*in
   wire signed [9:0] m275_100;
   assign m275_100 =10'b0;

   // m275_101 = W*in
   wire signed [9:0] m275_101;
   assign m275_101 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_102 = W*in
   wire signed [9:0] m275_102;
   assign m275_102 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_103 = W*in
   wire signed [9:0] m275_103;
   assign m275_103 =10'b0;

   // m275_104 = W*in
   wire signed [9:0] m275_104;
   assign m275_104 =10'b0;

   // m275_105 = W*in
   wire signed [9:0] m275_105;
   assign m275_105 =10'b0;

   // m275_106 = W*in
   wire signed [9:0] m275_106;
   assign m275_106 ={ {4{neg275[5]}} , neg275[5:0] };

   // m275_107 = W*in
   wire signed [9:0] m275_107;
   assign m275_107 =10'b0;

   // m275_108 = W*in
   wire signed [9:0] m275_108;
   assign m275_108 =10'b0;

   // m275_109 = W*in
   wire signed [9:0] m275_109;
   assign m275_109 ={ {5{neg275[5]}} , neg275[5:1] };

   // m275_110 = W*in
   wire signed [9:0] m275_110;
   assign m275_110 =10'b0;

   // m275_111 = W*in
   wire signed [9:0] m275_111;
   assign m275_111 =10'b0;

   // m275_112 = W*in
   wire signed [9:0] m275_112;
   assign m275_112 =10'b0;

   // m275_113 = W*in
   wire signed [9:0] m275_113;
   assign m275_113 ={ {4{in275[5]}} , in275[5:0] };

   // m275_114 = W*in
   wire signed [9:0] m275_114;
   assign m275_114 =10'b0;

   // m275_115 = W*in
   wire signed [9:0] m275_115;
   assign m275_115 =10'b0;

   // m275_116 = W*in
   wire signed [9:0] m275_116;
   assign m275_116 =10'b0;

   // m275_117 = W*in
   wire signed [9:0] m275_117;
   assign m275_117 ={ {4{neg275[5]}} , neg275[5:0] };

   // m276_1 = W*in
   wire signed [9:0] m276_1;
   assign m276_1 =10'b0;

   // m276_2 = W*in
   wire signed [9:0] m276_2;
   assign m276_2 =10'b0;

   // m276_3 = W*in
   wire signed [9:0] m276_3;
   assign m276_3 =10'b0;

   // m276_4 = W*in
   wire signed [9:0] m276_4;
   assign m276_4 =10'b0;

   // m276_5 = W*in
   wire signed [9:0] m276_5;
   assign m276_5 =10'b0;

   // m276_6 = W*in
   wire signed [9:0] m276_6;
   assign m276_6 =10'b0;

   // m276_7 = W*in
   wire signed [9:0] m276_7;
   assign m276_7 =10'b0;

   // m276_8 = W*in
   wire signed [9:0] m276_8;
   assign m276_8 =10'b0;

   // m276_9 = W*in
   wire signed [9:0] m276_9;
   assign m276_9 =10'b0;

   // m276_10 = W*in
   wire signed [9:0] m276_10;
   assign m276_10 =10'b0;

   // m276_11 = W*in
   wire signed [9:0] m276_11;
   assign m276_11 =10'b0;

   // m276_12 = W*in
   wire signed [9:0] m276_12;
   assign m276_12 =10'b0;

   // m276_13 = W*in
   wire signed [9:0] m276_13;
   assign m276_13 =10'b0;

   // m276_14 = W*in
   wire signed [9:0] m276_14;
   assign m276_14 =10'b0;

   // m276_15 = W*in
   wire signed [9:0] m276_15;
   assign m276_15 =10'b0;

   // m276_16 = W*in
   wire signed [9:0] m276_16;
   assign m276_16 =10'b0;

   // m276_17 = W*in
   wire signed [9:0] m276_17;
   assign m276_17 =10'b0;

   // m276_18 = W*in
   wire signed [9:0] m276_18;
   assign m276_18 ={ {5{in276[5]}} , in276[5:1] };

   // m276_19 = W*in
   wire signed [9:0] m276_19;
   assign m276_19 =10'b0;

   // m276_20 = W*in
   wire signed [9:0] m276_20;
   assign m276_20 ={ {5{in276[5]}} , in276[5:1] };

   // m276_21 = W*in
   wire signed [9:0] m276_21;
   assign m276_21 =10'b0;

   // m276_22 = W*in
   wire signed [9:0] m276_22;
   assign m276_22 =10'b0;

   // m276_23 = W*in
   wire signed [9:0] m276_23;
   assign m276_23 =10'b0;

   // m276_24 = W*in
   wire signed [9:0] m276_24;
   assign m276_24 ={ {4{neg276[5]}} , neg276[5:0] };

   // m276_25 = W*in
   wire signed [9:0] m276_25;
   assign m276_25 =10'b0;

   // m276_26 = W*in
   wire signed [9:0] m276_26;
   assign m276_26 =10'b0;

   // m276_27 = W*in
   wire signed [9:0] m276_27;
   assign m276_27 =10'b0;

   // m276_28 = W*in
   wire signed [9:0] m276_28;
   assign m276_28 =10'b0;

   // m276_29 = W*in
   wire signed [9:0] m276_29;
   assign m276_29 =10'b0;

   // m276_30 = W*in
   wire signed [9:0] m276_30;
   assign m276_30 =10'b0;

   // m276_31 = W*in
   wire signed [9:0] m276_31;
   assign m276_31 ={ {5{neg276[5]}} , neg276[5:1] };

   // m276_32 = W*in
   wire signed [9:0] m276_32;
   assign m276_32 =10'b0;

   // m276_33 = W*in
   wire signed [9:0] m276_33;
   assign m276_33 =10'b0;

   // m276_34 = W*in
   wire signed [9:0] m276_34;
   assign m276_34 =10'b0;

   // m276_35 = W*in
   wire signed [9:0] m276_35;
   assign m276_35 ={ {5{in276[5]}} , in276[5:1] };

   // m276_36 = W*in
   wire signed [9:0] m276_36;
   assign m276_36 ={ {4{in276[5]}} , in276[5:0] };

   // m276_37 = W*in
   wire signed [9:0] m276_37;
   assign m276_37 =10'b0;

   // m276_38 = W*in
   wire signed [9:0] m276_38;
   assign m276_38 =10'b0;

   // m276_39 = W*in
   wire signed [9:0] m276_39;
   assign m276_39 ={ {4{neg276[5]}} , neg276[5:0] };

   // m276_40 = W*in
   wire signed [9:0] m276_40;
   assign m276_40 =10'b0;

   // m276_41 = W*in
   wire signed [9:0] m276_41;
   assign m276_41 =10'b0;

   // m276_42 = W*in
   wire signed [9:0] m276_42;
   assign m276_42 =10'b0;

   // m276_43 = W*in
   wire signed [9:0] m276_43;
   assign m276_43 =10'b0;

   // m276_44 = W*in
   wire signed [9:0] m276_44;
   assign m276_44 =10'b0;

   // m276_45 = W*in
   wire signed [9:0] m276_45;
   assign m276_45 =10'b0;

   // m276_46 = W*in
   wire signed [9:0] m276_46;
   assign m276_46 =10'b0;

   // m276_47 = W*in
   wire signed [9:0] m276_47;
   assign m276_47 =10'b0;

   // m276_48 = W*in
   wire signed [9:0] m276_48;
   assign m276_48 ={ {4{in276[5]}} , in276[5:0] };

   // m276_49 = W*in
   wire signed [9:0] m276_49;
   assign m276_49 =10'b0;

   // m276_50 = W*in
   wire signed [9:0] m276_50;
   assign m276_50 =10'b0;

   // m276_51 = W*in
   wire signed [9:0] m276_51;
   assign m276_51 ={ {4{neg276[5]}} , neg276[5:0] };

   // m276_52 = W*in
   wire signed [9:0] m276_52;
   assign m276_52 =10'b0;

   // m276_53 = W*in
   wire signed [9:0] m276_53;
   assign m276_53 =10'b0;

   // m276_54 = W*in
   wire signed [9:0] m276_54;
   assign m276_54 =10'b0;

   // m276_55 = W*in
   wire signed [9:0] m276_55;
   assign m276_55 =10'b0;

   // m276_56 = W*in
   wire signed [9:0] m276_56;
   assign m276_56 =10'b0;

   // m276_57 = W*in
   wire signed [9:0] m276_57;
   assign m276_57 ={ {4{in276[5]}} , in276[5:0] };

   // m276_58 = W*in
   wire signed [9:0] m276_58;
   assign m276_58 =10'b0;

   // m276_59 = W*in
   wire signed [9:0] m276_59;
   assign m276_59 =10'b0;

   // m276_60 = W*in
   wire signed [9:0] m276_60;
   assign m276_60 =10'b0;

   // m276_61 = W*in
   wire signed [9:0] m276_61;
   assign m276_61 =10'b0;

   // m276_62 = W*in
   wire signed [9:0] m276_62;
   assign m276_62 =10'b0;

   // m276_63 = W*in
   wire signed [9:0] m276_63;
   assign m276_63 ={ {4{in276[5]}} , in276[5:0] };

   // m276_64 = W*in
   wire signed [9:0] m276_64;
   assign m276_64 =10'b0;

   // m276_65 = W*in
   wire signed [9:0] m276_65;
   assign m276_65 =10'b0;

   // m276_66 = W*in
   wire signed [9:0] m276_66;
   assign m276_66 =10'b0;

   // m276_67 = W*in
   wire signed [9:0] m276_67;
   assign m276_67 =10'b0;

   // m276_68 = W*in
   wire signed [9:0] m276_68;
   assign m276_68 =10'b0;

   // m276_69 = W*in
   wire signed [9:0] m276_69;
   assign m276_69 ={ {4{in276[5]}} , in276[5:0] };

   // m276_70 = W*in
   wire signed [9:0] m276_70;
   assign m276_70 ={ {4{in276[5]}} , in276[5:0] };

   // m276_71 = W*in
   wire signed [9:0] m276_71;
   assign m276_71 =10'b0;

   // m276_72 = W*in
   wire signed [9:0] m276_72;
   assign m276_72 ={ {4{in276[5]}} , in276[5:0] };

   // m276_73 = W*in
   wire signed [9:0] m276_73;
   assign m276_73 =10'b0;

   // m276_74 = W*in
   wire signed [9:0] m276_74;
   assign m276_74 =10'b0;

   // m276_75 = W*in
   wire signed [9:0] m276_75;
   assign m276_75 =10'b0;

   // m276_76 = W*in
   wire signed [9:0] m276_76;
   assign m276_76 =10'b0;

   // m276_77 = W*in
   wire signed [9:0] m276_77;
   assign m276_77 =10'b0;

   // m276_78 = W*in
   wire signed [9:0] m276_78;
   assign m276_78 =10'b0;

   // m276_79 = W*in
   wire signed [9:0] m276_79;
   assign m276_79 =10'b0;

   // m276_80 = W*in
   wire signed [9:0] m276_80;
   assign m276_80 =10'b0;

   // m276_81 = W*in
   wire signed [9:0] m276_81;
   assign m276_81 =10'b0;

   // m276_82 = W*in
   wire signed [9:0] m276_82;
   assign m276_82 =10'b0;

   // m276_83 = W*in
   wire signed [9:0] m276_83;
   assign m276_83 =10'b0;

   // m276_84 = W*in
   wire signed [9:0] m276_84;
   assign m276_84 =10'b0;

   // m276_85 = W*in
   wire signed [9:0] m276_85;
   assign m276_85 =10'b0;

   // m276_86 = W*in
   wire signed [9:0] m276_86;
   assign m276_86 =10'b0;

   // m276_87 = W*in
   wire signed [9:0] m276_87;
   assign m276_87 =10'b0;

   // m276_88 = W*in
   wire signed [9:0] m276_88;
   assign m276_88 =10'b0;

   // m276_89 = W*in
   wire signed [9:0] m276_89;
   assign m276_89 =10'b0;

   // m276_90 = W*in
   wire signed [9:0] m276_90;
   assign m276_90 =10'b0;

   // m276_91 = W*in
   wire signed [9:0] m276_91;
   assign m276_91 =10'b0;

   // m276_92 = W*in
   wire signed [9:0] m276_92;
   assign m276_92 =10'b0;

   // m276_93 = W*in
   wire signed [9:0] m276_93;
   assign m276_93 =10'b0;

   // m276_94 = W*in
   wire signed [9:0] m276_94;
   assign m276_94 =10'b0;

   // m276_95 = W*in
   wire signed [9:0] m276_95;
   assign m276_95 =10'b0;

   // m276_96 = W*in
   wire signed [9:0] m276_96;
   assign m276_96 =10'b0;

   // m276_97 = W*in
   wire signed [9:0] m276_97;
   assign m276_97 =10'b0;

   // m276_98 = W*in
   wire signed [9:0] m276_98;
   assign m276_98 =10'b0;

   // m276_99 = W*in
   wire signed [9:0] m276_99;
   assign m276_99 =10'b0;

   // m276_100 = W*in
   wire signed [9:0] m276_100;
   assign m276_100 =10'b0;

   // m276_101 = W*in
   wire signed [9:0] m276_101;
   assign m276_101 =10'b0;

   // m276_102 = W*in
   wire signed [9:0] m276_102;
   assign m276_102 =10'b0;

   // m276_103 = W*in
   wire signed [9:0] m276_103;
   assign m276_103 =10'b0;

   // m276_104 = W*in
   wire signed [9:0] m276_104;
   assign m276_104 =10'b0;

   // m276_105 = W*in
   wire signed [9:0] m276_105;
   assign m276_105 =10'b0;

   // m276_106 = W*in
   wire signed [9:0] m276_106;
   assign m276_106 =10'b0;

   // m276_107 = W*in
   wire signed [9:0] m276_107;
   assign m276_107 =10'b0;

   // m276_108 = W*in
   wire signed [9:0] m276_108;
   assign m276_108 =10'b0;

   // m276_109 = W*in
   wire signed [9:0] m276_109;
   assign m276_109 =10'b0;

   // m276_110 = W*in
   wire signed [9:0] m276_110;
   assign m276_110 =10'b0;

   // m276_111 = W*in
   wire signed [9:0] m276_111;
   assign m276_111 =10'b0;

   // m276_112 = W*in
   wire signed [9:0] m276_112;
   assign m276_112 =10'b0;

   // m276_113 = W*in
   wire signed [9:0] m276_113;
   assign m276_113 =10'b0;

   // m276_114 = W*in
   wire signed [9:0] m276_114;
   assign m276_114 =10'b0;

   // m276_115 = W*in
   wire signed [9:0] m276_115;
   assign m276_115 =10'b0;

   // m276_116 = W*in
   wire signed [9:0] m276_116;
   assign m276_116 =10'b0;

   // m276_117 = W*in
   wire signed [9:0] m276_117;
   assign m276_117 =10'b0;

   // m277_1 = W*in
   wire signed [9:0] m277_1;
   assign m277_1 =10'b0;

   // m277_2 = W*in
   wire signed [9:0] m277_2;
   assign m277_2 =10'b0;

   // m277_3 = W*in
   wire signed [9:0] m277_3;
   assign m277_3 =10'b0;

   // m277_4 = W*in
   wire signed [9:0] m277_4;
   assign m277_4 =10'b0;

   // m277_5 = W*in
   wire signed [9:0] m277_5;
   assign m277_5 =10'b0;

   // m277_6 = W*in
   wire signed [9:0] m277_6;
   assign m277_6 =10'b0;

   // m277_7 = W*in
   wire signed [9:0] m277_7;
   assign m277_7 =10'b0;

   // m277_8 = W*in
   wire signed [9:0] m277_8;
   assign m277_8 =10'b0;

   // m277_9 = W*in
   wire signed [9:0] m277_9;
   assign m277_9 =10'b0;

   // m277_10 = W*in
   wire signed [9:0] m277_10;
   assign m277_10 =10'b0;

   // m277_11 = W*in
   wire signed [9:0] m277_11;
   assign m277_11 =10'b0;

   // m277_12 = W*in
   wire signed [9:0] m277_12;
   assign m277_12 =10'b0;

   // m277_13 = W*in
   wire signed [9:0] m277_13;
   assign m277_13 =10'b0;

   // m277_14 = W*in
   wire signed [9:0] m277_14;
   assign m277_14 =10'b0;

   // m277_15 = W*in
   wire signed [9:0] m277_15;
   assign m277_15 =10'b0;

   // m277_16 = W*in
   wire signed [9:0] m277_16;
   assign m277_16 =10'b0;

   // m277_17 = W*in
   wire signed [9:0] m277_17;
   assign m277_17 ={ {5{in277[5]}} , in277[5:1] };

   // m277_18 = W*in
   wire signed [9:0] m277_18;
   assign m277_18 =10'b0;

   // m277_19 = W*in
   wire signed [9:0] m277_19;
   assign m277_19 =10'b0;

   // m277_20 = W*in
   wire signed [9:0] m277_20;
   assign m277_20 =10'b0;

   // m277_21 = W*in
   wire signed [9:0] m277_21;
   assign m277_21 =10'b0;

   // m277_22 = W*in
   wire signed [9:0] m277_22;
   assign m277_22 =10'b0;

   // m277_23 = W*in
   wire signed [9:0] m277_23;
   assign m277_23 =10'b0;

   // m277_24 = W*in
   wire signed [9:0] m277_24;
   assign m277_24 =10'b0;

   // m277_25 = W*in
   wire signed [9:0] m277_25;
   assign m277_25 =10'b0;

   // m277_26 = W*in
   wire signed [9:0] m277_26;
   assign m277_26 ={ {5{neg277[5]}} , neg277[5:1] };

   // m277_27 = W*in
   wire signed [9:0] m277_27;
   assign m277_27 =10'b0;

   // m277_28 = W*in
   wire signed [9:0] m277_28;
   assign m277_28 =10'b0;

   // m277_29 = W*in
   wire signed [9:0] m277_29;
   assign m277_29 =10'b0;

   // m277_30 = W*in
   wire signed [9:0] m277_30;
   assign m277_30 =10'b0;

   // m277_31 = W*in
   wire signed [9:0] m277_31;
   assign m277_31 =10'b0;

   // m277_32 = W*in
   wire signed [9:0] m277_32;
   assign m277_32 =10'b0;

   // m277_33 = W*in
   wire signed [9:0] m277_33;
   assign m277_33 =10'b0;

   // m277_34 = W*in
   wire signed [9:0] m277_34;
   assign m277_34 =10'b0;

   // m277_35 = W*in
   wire signed [9:0] m277_35;
   assign m277_35 =10'b0;

   // m277_36 = W*in
   wire signed [9:0] m277_36;
   assign m277_36 =10'b0;

   // m277_37 = W*in
   wire signed [9:0] m277_37;
   assign m277_37 =10'b0;

   // m277_38 = W*in
   wire signed [9:0] m277_38;
   assign m277_38 =10'b0;

   // m277_39 = W*in
   wire signed [9:0] m277_39;
   assign m277_39 =10'b0;

   // m277_40 = W*in
   wire signed [9:0] m277_40;
   assign m277_40 =10'b0;

   // m277_41 = W*in
   wire signed [9:0] m277_41;
   assign m277_41 =10'b0;

   // m277_42 = W*in
   wire signed [9:0] m277_42;
   assign m277_42 =10'b0;

   // m277_43 = W*in
   wire signed [9:0] m277_43;
   assign m277_43 =10'b0;

   // m277_44 = W*in
   wire signed [9:0] m277_44;
   assign m277_44 =10'b0;

   // m277_45 = W*in
   wire signed [9:0] m277_45;
   assign m277_45 =10'b0;

   // m277_46 = W*in
   wire signed [9:0] m277_46;
   assign m277_46 =10'b0;

   // m277_47 = W*in
   wire signed [9:0] m277_47;
   assign m277_47 =10'b0;

   // m277_48 = W*in
   wire signed [9:0] m277_48;
   assign m277_48 =10'b0;

   // m277_49 = W*in
   wire signed [9:0] m277_49;
   assign m277_49 =10'b0;

   // m277_50 = W*in
   wire signed [9:0] m277_50;
   assign m277_50 =10'b0;

   // m277_51 = W*in
   wire signed [9:0] m277_51;
   assign m277_51 ={ {4{in277[5]}} , in277[5:0] };

   // m277_52 = W*in
   wire signed [9:0] m277_52;
   assign m277_52 =10'b0;

   // m277_53 = W*in
   wire signed [9:0] m277_53;
   assign m277_53 =10'b0;

   // m277_54 = W*in
   wire signed [9:0] m277_54;
   assign m277_54 =10'b0;

   // m277_55 = W*in
   wire signed [9:0] m277_55;
   assign m277_55 =10'b0;

   // m277_56 = W*in
   wire signed [9:0] m277_56;
   assign m277_56 =10'b0;

   // m277_57 = W*in
   wire signed [9:0] m277_57;
   assign m277_57 =10'b0;

   // m277_58 = W*in
   wire signed [9:0] m277_58;
   assign m277_58 =10'b0;

   // m277_59 = W*in
   wire signed [9:0] m277_59;
   assign m277_59 =10'b0;

   // m277_60 = W*in
   wire signed [9:0] m277_60;
   assign m277_60 =10'b0;

   // m277_61 = W*in
   wire signed [9:0] m277_61;
   assign m277_61 =10'b0;

   // m277_62 = W*in
   wire signed [9:0] m277_62;
   assign m277_62 =10'b0;

   // m277_63 = W*in
   wire signed [9:0] m277_63;
   assign m277_63 =10'b0;

   // m277_64 = W*in
   wire signed [9:0] m277_64;
   assign m277_64 =10'b0;

   // m277_65 = W*in
   wire signed [9:0] m277_65;
   assign m277_65 =10'b0;

   // m277_66 = W*in
   wire signed [9:0] m277_66;
   assign m277_66 =10'b0;

   // m277_67 = W*in
   wire signed [9:0] m277_67;
   assign m277_67 =10'b0;

   // m277_68 = W*in
   wire signed [9:0] m277_68;
   assign m277_68 =10'b0;

   // m277_69 = W*in
   wire signed [9:0] m277_69;
   assign m277_69 =10'b0;

   // m277_70 = W*in
   wire signed [9:0] m277_70;
   assign m277_70 ={ {5{neg277[5]}} , neg277[5:1] };

   // m277_71 = W*in
   wire signed [9:0] m277_71;
   assign m277_71 =10'b0;

   // m277_72 = W*in
   wire signed [9:0] m277_72;
   assign m277_72 ={ {5{neg277[5]}} , neg277[5:1] };

   // m277_73 = W*in
   wire signed [9:0] m277_73;
   assign m277_73 ={ {5{in277[5]}} , in277[5:1] };

   // m277_74 = W*in
   wire signed [9:0] m277_74;
   assign m277_74 =10'b0;

   // m277_75 = W*in
   wire signed [9:0] m277_75;
   assign m277_75 =10'b0;

   // m277_76 = W*in
   wire signed [9:0] m277_76;
   assign m277_76 =10'b0;

   // m277_77 = W*in
   wire signed [9:0] m277_77;
   assign m277_77 =10'b0;

   // m277_78 = W*in
   wire signed [9:0] m277_78;
   assign m277_78 ={ {5{neg277[5]}} , neg277[5:1] };

   // m277_79 = W*in
   wire signed [9:0] m277_79;
   assign m277_79 =10'b0;

   // m277_80 = W*in
   wire signed [9:0] m277_80;
   assign m277_80 =10'b0;

   // m277_81 = W*in
   wire signed [9:0] m277_81;
   assign m277_81 =10'b0;

   // m277_82 = W*in
   wire signed [9:0] m277_82;
   assign m277_82 =10'b0;

   // m277_83 = W*in
   wire signed [9:0] m277_83;
   assign m277_83 =10'b0;

   // m277_84 = W*in
   wire signed [9:0] m277_84;
   assign m277_84 =10'b0;

   // m277_85 = W*in
   wire signed [9:0] m277_85;
   assign m277_85 =10'b0;

   // m277_86 = W*in
   wire signed [9:0] m277_86;
   assign m277_86 =10'b0;

   // m277_87 = W*in
   wire signed [9:0] m277_87;
   assign m277_87 =10'b0;

   // m277_88 = W*in
   wire signed [9:0] m277_88;
   assign m277_88 =10'b0;

   // m277_89 = W*in
   wire signed [9:0] m277_89;
   assign m277_89 =10'b0;

   // m277_90 = W*in
   wire signed [9:0] m277_90;
   assign m277_90 =10'b0;

   // m277_91 = W*in
   wire signed [9:0] m277_91;
   assign m277_91 =10'b0;

   // m277_92 = W*in
   wire signed [9:0] m277_92;
   assign m277_92 =10'b0;

   // m277_93 = W*in
   wire signed [9:0] m277_93;
   assign m277_93 =10'b0;

   // m277_94 = W*in
   wire signed [9:0] m277_94;
   assign m277_94 =10'b0;

   // m277_95 = W*in
   wire signed [9:0] m277_95;
   assign m277_95 =10'b0;

   // m277_96 = W*in
   wire signed [9:0] m277_96;
   assign m277_96 =10'b0;

   // m277_97 = W*in
   wire signed [9:0] m277_97;
   assign m277_97 =10'b0;

   // m277_98 = W*in
   wire signed [9:0] m277_98;
   assign m277_98 =10'b0;

   // m277_99 = W*in
   wire signed [9:0] m277_99;
   assign m277_99 =10'b0;

   // m277_100 = W*in
   wire signed [9:0] m277_100;
   assign m277_100 =10'b0;

   // m277_101 = W*in
   wire signed [9:0] m277_101;
   assign m277_101 =10'b0;

   // m277_102 = W*in
   wire signed [9:0] m277_102;
   assign m277_102 =10'b0;

   // m277_103 = W*in
   wire signed [9:0] m277_103;
   assign m277_103 =10'b0;

   // m277_104 = W*in
   wire signed [9:0] m277_104;
   assign m277_104 =10'b0;

   // m277_105 = W*in
   wire signed [9:0] m277_105;
   assign m277_105 =10'b0;

   // m277_106 = W*in
   wire signed [9:0] m277_106;
   assign m277_106 =10'b0;

   // m277_107 = W*in
   wire signed [9:0] m277_107;
   assign m277_107 =10'b0;

   // m277_108 = W*in
   wire signed [9:0] m277_108;
   assign m277_108 =10'b0;

   // m277_109 = W*in
   wire signed [9:0] m277_109;
   assign m277_109 =10'b0;

   // m277_110 = W*in
   wire signed [9:0] m277_110;
   assign m277_110 =10'b0;

   // m277_111 = W*in
   wire signed [9:0] m277_111;
   assign m277_111 =10'b0;

   // m277_112 = W*in
   wire signed [9:0] m277_112;
   assign m277_112 =10'b0;

   // m277_113 = W*in
   wire signed [9:0] m277_113;
   assign m277_113 =10'b0;

   // m277_114 = W*in
   wire signed [9:0] m277_114;
   assign m277_114 =10'b0;

   // m277_115 = W*in
   wire signed [9:0] m277_115;
   assign m277_115 =10'b0;

   // m277_116 = W*in
   wire signed [9:0] m277_116;
   assign m277_116 =10'b0;

   // m277_117 = W*in
   wire signed [9:0] m277_117;
   assign m277_117 =10'b0;

   // m278_1 = W*in
   wire signed [9:0] m278_1;
   assign m278_1 =10'b0;

   // m278_2 = W*in
   wire signed [9:0] m278_2;
   assign m278_2 =10'b0;

   // m278_3 = W*in
   wire signed [9:0] m278_3;
   assign m278_3 =10'b0;

   // m278_4 = W*in
   wire signed [9:0] m278_4;
   assign m278_4 =10'b0;

   // m278_5 = W*in
   wire signed [9:0] m278_5;
   assign m278_5 =10'b0;

   // m278_6 = W*in
   wire signed [9:0] m278_6;
   assign m278_6 =10'b0;

   // m278_7 = W*in
   wire signed [9:0] m278_7;
   assign m278_7 ={ {4{in278[5]}} , in278[5:0] };

   // m278_8 = W*in
   wire signed [9:0] m278_8;
   assign m278_8 =10'b0;

   // m278_9 = W*in
   wire signed [9:0] m278_9;
   assign m278_9 =10'b0;

   // m278_10 = W*in
   wire signed [9:0] m278_10;
   assign m278_10 =10'b0;

   // m278_11 = W*in
   wire signed [9:0] m278_11;
   assign m278_11 =10'b0;

   // m278_12 = W*in
   wire signed [9:0] m278_12;
   assign m278_12 =10'b0;

   // m278_13 = W*in
   wire signed [9:0] m278_13;
   assign m278_13 =10'b0;

   // m278_14 = W*in
   wire signed [9:0] m278_14;
   assign m278_14 =10'b0;

   // m278_15 = W*in
   wire signed [9:0] m278_15;
   assign m278_15 =10'b0;

   // m278_16 = W*in
   wire signed [9:0] m278_16;
   assign m278_16 =10'b0;

   // m278_17 = W*in
   wire signed [9:0] m278_17;
   assign m278_17 =10'b0;

   // m278_18 = W*in
   wire signed [9:0] m278_18;
   assign m278_18 =10'b0;

   // m278_19 = W*in
   wire signed [9:0] m278_19;
   assign m278_19 =10'b0;

   // m278_20 = W*in
   wire signed [9:0] m278_20;
   assign m278_20 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_21 = W*in
   wire signed [9:0] m278_21;
   assign m278_21 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_22 = W*in
   wire signed [9:0] m278_22;
   assign m278_22 =10'b0;

   // m278_23 = W*in
   wire signed [9:0] m278_23;
   assign m278_23 =10'b0;

   // m278_24 = W*in
   wire signed [9:0] m278_24;
   assign m278_24 =10'b0;

   // m278_25 = W*in
   wire signed [9:0] m278_25;
   assign m278_25 ={ {4{in278[5]}} , in278[5:0] };

   // m278_26 = W*in
   wire signed [9:0] m278_26;
   assign m278_26 =10'b0;

   // m278_27 = W*in
   wire signed [9:0] m278_27;
   assign m278_27 ={ {4{in278[5]}} , in278[5:0] };

   // m278_28 = W*in
   wire signed [9:0] m278_28;
   assign m278_28 ={ {4{in278[5]}} , in278[5:0] };

   // m278_29 = W*in
   wire signed [9:0] m278_29;
   assign m278_29 =10'b0;

   // m278_30 = W*in
   wire signed [9:0] m278_30;
   assign m278_30 =10'b0;

   // m278_31 = W*in
   wire signed [9:0] m278_31;
   assign m278_31 =10'b0;

   // m278_32 = W*in
   wire signed [9:0] m278_32;
   assign m278_32 =10'b0;

   // m278_33 = W*in
   wire signed [9:0] m278_33;
   assign m278_33 =10'b0;

   // m278_34 = W*in
   wire signed [9:0] m278_34;
   assign m278_34 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_35 = W*in
   wire signed [9:0] m278_35;
   assign m278_35 =10'b0;

   // m278_36 = W*in
   wire signed [9:0] m278_36;
   assign m278_36 ={ {5{in278[5]}} , in278[5:1] };

   // m278_37 = W*in
   wire signed [9:0] m278_37;
   assign m278_37 =10'b0;

   // m278_38 = W*in
   wire signed [9:0] m278_38;
   assign m278_38 =10'b0;

   // m278_39 = W*in
   wire signed [9:0] m278_39;
   assign m278_39 =10'b0;

   // m278_40 = W*in
   wire signed [9:0] m278_40;
   assign m278_40 =10'b0;

   // m278_41 = W*in
   wire signed [9:0] m278_41;
   assign m278_41 =10'b0;

   // m278_42 = W*in
   wire signed [9:0] m278_42;
   assign m278_42 =10'b0;

   // m278_43 = W*in
   wire signed [9:0] m278_43;
   assign m278_43 =10'b0;

   // m278_44 = W*in
   wire signed [9:0] m278_44;
   assign m278_44 =10'b0;

   // m278_45 = W*in
   wire signed [9:0] m278_45;
   assign m278_45 =10'b0;

   // m278_46 = W*in
   wire signed [9:0] m278_46;
   assign m278_46 =10'b0;

   // m278_47 = W*in
   wire signed [9:0] m278_47;
   assign m278_47 =10'b0;

   // m278_48 = W*in
   wire signed [9:0] m278_48;
   assign m278_48 =10'b0;

   // m278_49 = W*in
   wire signed [9:0] m278_49;
   assign m278_49 =10'b0;

   // m278_50 = W*in
   wire signed [9:0] m278_50;
   assign m278_50 =10'b0;

   // m278_51 = W*in
   wire signed [9:0] m278_51;
   assign m278_51 ={ {4{in278[5]}} , in278[5:0] };

   // m278_52 = W*in
   wire signed [9:0] m278_52;
   assign m278_52 =10'b0;

   // m278_53 = W*in
   wire signed [9:0] m278_53;
   assign m278_53 =10'b0;

   // m278_54 = W*in
   wire signed [9:0] m278_54;
   assign m278_54 =10'b0;

   // m278_55 = W*in
   wire signed [9:0] m278_55;
   assign m278_55 =10'b0;

   // m278_56 = W*in
   wire signed [9:0] m278_56;
   assign m278_56 =10'b0;

   // m278_57 = W*in
   wire signed [9:0] m278_57;
   assign m278_57 =10'b0;

   // m278_58 = W*in
   wire signed [9:0] m278_58;
   assign m278_58 =10'b0;

   // m278_59 = W*in
   wire signed [9:0] m278_59;
   assign m278_59 ={ {4{in278[5]}} , in278[5:0] };

   // m278_60 = W*in
   wire signed [9:0] m278_60;
   assign m278_60 =10'b0;

   // m278_61 = W*in
   wire signed [9:0] m278_61;
   assign m278_61 =10'b0;

   // m278_62 = W*in
   wire signed [9:0] m278_62;
   assign m278_62 =10'b0;

   // m278_63 = W*in
   wire signed [9:0] m278_63;
   assign m278_63 =10'b0;

   // m278_64 = W*in
   wire signed [9:0] m278_64;
   assign m278_64 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_65 = W*in
   wire signed [9:0] m278_65;
   assign m278_65 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_66 = W*in
   wire signed [9:0] m278_66;
   assign m278_66 =10'b0;

   // m278_67 = W*in
   wire signed [9:0] m278_67;
   assign m278_67 =10'b0;

   // m278_68 = W*in
   wire signed [9:0] m278_68;
   assign m278_68 =10'b0;

   // m278_69 = W*in
   wire signed [9:0] m278_69;
   assign m278_69 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_70 = W*in
   wire signed [9:0] m278_70;
   assign m278_70 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_71 = W*in
   wire signed [9:0] m278_71;
   assign m278_71 ={ {5{in278[5]}} , in278[5:1] };

   // m278_72 = W*in
   wire signed [9:0] m278_72;
   assign m278_72 =10'b0;

   // m278_73 = W*in
   wire signed [9:0] m278_73;
   assign m278_73 ={ {5{in278[5]}} , in278[5:1] };

   // m278_74 = W*in
   wire signed [9:0] m278_74;
   assign m278_74 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_75 = W*in
   wire signed [9:0] m278_75;
   assign m278_75 =10'b0;

   // m278_76 = W*in
   wire signed [9:0] m278_76;
   assign m278_76 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_77 = W*in
   wire signed [9:0] m278_77;
   assign m278_77 =10'b0;

   // m278_78 = W*in
   wire signed [9:0] m278_78;
   assign m278_78 =10'b0;

   // m278_79 = W*in
   wire signed [9:0] m278_79;
   assign m278_79 =10'b0;

   // m278_80 = W*in
   wire signed [9:0] m278_80;
   assign m278_80 =10'b0;

   // m278_81 = W*in
   wire signed [9:0] m278_81;
   assign m278_81 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_82 = W*in
   wire signed [9:0] m278_82;
   assign m278_82 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_83 = W*in
   wire signed [9:0] m278_83;
   assign m278_83 =10'b0;

   // m278_84 = W*in
   wire signed [9:0] m278_84;
   assign m278_84 =10'b0;

   // m278_85 = W*in
   wire signed [9:0] m278_85;
   assign m278_85 =10'b0;

   // m278_86 = W*in
   wire signed [9:0] m278_86;
   assign m278_86 =10'b0;

   // m278_87 = W*in
   wire signed [9:0] m278_87;
   assign m278_87 =10'b0;

   // m278_88 = W*in
   wire signed [9:0] m278_88;
   assign m278_88 =10'b0;

   // m278_89 = W*in
   wire signed [9:0] m278_89;
   assign m278_89 =10'b0;

   // m278_90 = W*in
   wire signed [9:0] m278_90;
   assign m278_90 =10'b0;

   // m278_91 = W*in
   wire signed [9:0] m278_91;
   assign m278_91 =10'b0;

   // m278_92 = W*in
   wire signed [9:0] m278_92;
   assign m278_92 =10'b0;

   // m278_93 = W*in
   wire signed [9:0] m278_93;
   assign m278_93 =10'b0;

   // m278_94 = W*in
   wire signed [9:0] m278_94;
   assign m278_94 =10'b0;

   // m278_95 = W*in
   wire signed [9:0] m278_95;
   assign m278_95 =10'b0;

   // m278_96 = W*in
   wire signed [9:0] m278_96;
   assign m278_96 =10'b0;

   // m278_97 = W*in
   wire signed [9:0] m278_97;
   assign m278_97 =10'b0;

   // m278_98 = W*in
   wire signed [9:0] m278_98;
   assign m278_98 =10'b0;

   // m278_99 = W*in
   wire signed [9:0] m278_99;
   assign m278_99 ={ {4{neg278[5]}} , neg278[5:0] };

   // m278_100 = W*in
   wire signed [9:0] m278_100;
   assign m278_100 =10'b0;

   // m278_101 = W*in
   wire signed [9:0] m278_101;
   assign m278_101 =10'b0;

   // m278_102 = W*in
   wire signed [9:0] m278_102;
   assign m278_102 =10'b0;

   // m278_103 = W*in
   wire signed [9:0] m278_103;
   assign m278_103 =10'b0;

   // m278_104 = W*in
   wire signed [9:0] m278_104;
   assign m278_104 =10'b0;

   // m278_105 = W*in
   wire signed [9:0] m278_105;
   assign m278_105 =10'b0;

   // m278_106 = W*in
   wire signed [9:0] m278_106;
   assign m278_106 =10'b0;

   // m278_107 = W*in
   wire signed [9:0] m278_107;
   assign m278_107 ={ {4{in278[5]}} , in278[5:0] };

   // m278_108 = W*in
   wire signed [9:0] m278_108;
   assign m278_108 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_109 = W*in
   wire signed [9:0] m278_109;
   assign m278_109 =10'b0;

   // m278_110 = W*in
   wire signed [9:0] m278_110;
   assign m278_110 =10'b0;

   // m278_111 = W*in
   wire signed [9:0] m278_111;
   assign m278_111 =10'b0;

   // m278_112 = W*in
   wire signed [9:0] m278_112;
   assign m278_112 =10'b0;

   // m278_113 = W*in
   wire signed [9:0] m278_113;
   assign m278_113 =10'b0;

   // m278_114 = W*in
   wire signed [9:0] m278_114;
   assign m278_114 =10'b0;

   // m278_115 = W*in
   wire signed [9:0] m278_115;
   assign m278_115 ={ {5{neg278[5]}} , neg278[5:1] };

   // m278_116 = W*in
   wire signed [9:0] m278_116;
   assign m278_116 =10'b0;

   // m278_117 = W*in
   wire signed [9:0] m278_117;
   assign m278_117 =10'b0;

   // m279_1 = W*in
   wire signed [9:0] m279_1;
   assign m279_1 =10'b0;

   // m279_2 = W*in
   wire signed [9:0] m279_2;
   assign m279_2 =10'b0;

   // m279_3 = W*in
   wire signed [9:0] m279_3;
   assign m279_3 =10'b0;

   // m279_4 = W*in
   wire signed [9:0] m279_4;
   assign m279_4 =10'b0;

   // m279_5 = W*in
   wire signed [9:0] m279_5;
   assign m279_5 =10'b0;

   // m279_6 = W*in
   wire signed [9:0] m279_6;
   assign m279_6 =10'b0;

   // m279_7 = W*in
   wire signed [9:0] m279_7;
   assign m279_7 =10'b0;

   // m279_8 = W*in
   wire signed [9:0] m279_8;
   assign m279_8 =10'b0;

   // m279_9 = W*in
   wire signed [9:0] m279_9;
   assign m279_9 =10'b0;

   // m279_10 = W*in
   wire signed [9:0] m279_10;
   assign m279_10 =10'b0;

   // m279_11 = W*in
   wire signed [9:0] m279_11;
   assign m279_11 =10'b0;

   // m279_12 = W*in
   wire signed [9:0] m279_12;
   assign m279_12 =10'b0;

   // m279_13 = W*in
   wire signed [9:0] m279_13;
   assign m279_13 =10'b0;

   // m279_14 = W*in
   wire signed [9:0] m279_14;
   assign m279_14 =10'b0;

   // m279_15 = W*in
   wire signed [9:0] m279_15;
   assign m279_15 =10'b0;

   // m279_16 = W*in
   wire signed [9:0] m279_16;
   assign m279_16 =10'b0;

   // m279_17 = W*in
   wire signed [9:0] m279_17;
   assign m279_17 =10'b0;

   // m279_18 = W*in
   wire signed [9:0] m279_18;
   assign m279_18 ={ {5{in279[5]}} , in279[5:1] };

   // m279_19 = W*in
   wire signed [9:0] m279_19;
   assign m279_19 =10'b0;

   // m279_20 = W*in
   wire signed [9:0] m279_20;
   assign m279_20 =10'b0;

   // m279_21 = W*in
   wire signed [9:0] m279_21;
   assign m279_21 ={ {5{neg279[5]}} , neg279[5:1] };

   // m279_22 = W*in
   wire signed [9:0] m279_22;
   assign m279_22 ={ {4{in279[5]}} , in279[5:0] };

   // m279_23 = W*in
   wire signed [9:0] m279_23;
   assign m279_23 =10'b0;

   // m279_24 = W*in
   wire signed [9:0] m279_24;
   assign m279_24 =10'b0;

   // m279_25 = W*in
   wire signed [9:0] m279_25;
   assign m279_25 =10'b0;

   // m279_26 = W*in
   wire signed [9:0] m279_26;
   assign m279_26 =10'b0;

   // m279_27 = W*in
   wire signed [9:0] m279_27;
   assign m279_27 =10'b0;

   // m279_28 = W*in
   wire signed [9:0] m279_28;
   assign m279_28 =10'b0;

   // m279_29 = W*in
   wire signed [9:0] m279_29;
   assign m279_29 =10'b0;

   // m279_30 = W*in
   wire signed [9:0] m279_30;
   assign m279_30 =10'b0;

   // m279_31 = W*in
   wire signed [9:0] m279_31;
   assign m279_31 =10'b0;

   // m279_32 = W*in
   wire signed [9:0] m279_32;
   assign m279_32 =10'b0;

   // m279_33 = W*in
   wire signed [9:0] m279_33;
   assign m279_33 =10'b0;

   // m279_34 = W*in
   wire signed [9:0] m279_34;
   assign m279_34 ={ {5{in279[5]}} , in279[5:1] };

   // m279_35 = W*in
   wire signed [9:0] m279_35;
   assign m279_35 =10'b0;

   // m279_36 = W*in
   wire signed [9:0] m279_36;
   assign m279_36 =10'b0;

   // m279_37 = W*in
   wire signed [9:0] m279_37;
   assign m279_37 =10'b0;

   // m279_38 = W*in
   wire signed [9:0] m279_38;
   assign m279_38 =10'b0;

   // m279_39 = W*in
   wire signed [9:0] m279_39;
   assign m279_39 =10'b0;

   // m279_40 = W*in
   wire signed [9:0] m279_40;
   assign m279_40 =10'b0;

   // m279_41 = W*in
   wire signed [9:0] m279_41;
   assign m279_41 =10'b0;

   // m279_42 = W*in
   wire signed [9:0] m279_42;
   assign m279_42 =10'b0;

   // m279_43 = W*in
   wire signed [9:0] m279_43;
   assign m279_43 =10'b0;

   // m279_44 = W*in
   wire signed [9:0] m279_44;
   assign m279_44 ={ {4{neg279[5]}} , neg279[5:0] };

   // m279_45 = W*in
   wire signed [9:0] m279_45;
   assign m279_45 =10'b0;

   // m279_46 = W*in
   wire signed [9:0] m279_46;
   assign m279_46 =10'b0;

   // m279_47 = W*in
   wire signed [9:0] m279_47;
   assign m279_47 =10'b0;

   // m279_48 = W*in
   wire signed [9:0] m279_48;
   assign m279_48 =10'b0;

   // m279_49 = W*in
   wire signed [9:0] m279_49;
   assign m279_49 =10'b0;

   // m279_50 = W*in
   wire signed [9:0] m279_50;
   assign m279_50 =10'b0;

   // m279_51 = W*in
   wire signed [9:0] m279_51;
   assign m279_51 =10'b0;

   // m279_52 = W*in
   wire signed [9:0] m279_52;
   assign m279_52 =10'b0;

   // m279_53 = W*in
   wire signed [9:0] m279_53;
   assign m279_53 =10'b0;

   // m279_54 = W*in
   wire signed [9:0] m279_54;
   assign m279_54 =10'b0;

   // m279_55 = W*in
   wire signed [9:0] m279_55;
   assign m279_55 =10'b0;

   // m279_56 = W*in
   wire signed [9:0] m279_56;
   assign m279_56 =10'b0;

   // m279_57 = W*in
   wire signed [9:0] m279_57;
   assign m279_57 =10'b0;

   // m279_58 = W*in
   wire signed [9:0] m279_58;
   assign m279_58 =10'b0;

   // m279_59 = W*in
   wire signed [9:0] m279_59;
   assign m279_59 =10'b0;

   // m279_60 = W*in
   wire signed [9:0] m279_60;
   assign m279_60 =10'b0;

   // m279_61 = W*in
   wire signed [9:0] m279_61;
   assign m279_61 =10'b0;

   // m279_62 = W*in
   wire signed [9:0] m279_62;
   assign m279_62 =10'b0;

   // m279_63 = W*in
   wire signed [9:0] m279_63;
   assign m279_63 =10'b0;

   // m279_64 = W*in
   wire signed [9:0] m279_64;
   assign m279_64 =10'b0;

   // m279_65 = W*in
   wire signed [9:0] m279_65;
   assign m279_65 =10'b0;

   // m279_66 = W*in
   wire signed [9:0] m279_66;
   assign m279_66 =10'b0;

   // m279_67 = W*in
   wire signed [9:0] m279_67;
   assign m279_67 ={ {4{neg279[5]}} , neg279[5:0] };

   // m279_68 = W*in
   wire signed [9:0] m279_68;
   assign m279_68 =10'b0;

   // m279_69 = W*in
   wire signed [9:0] m279_69;
   assign m279_69 =10'b0;

   // m279_70 = W*in
   wire signed [9:0] m279_70;
   assign m279_70 =10'b0;

   // m279_71 = W*in
   wire signed [9:0] m279_71;
   assign m279_71 =10'b0;

   // m279_72 = W*in
   wire signed [9:0] m279_72;
   assign m279_72 =10'b0;

   // m279_73 = W*in
   wire signed [9:0] m279_73;
   assign m279_73 =10'b0;

   // m279_74 = W*in
   wire signed [9:0] m279_74;
   assign m279_74 ={ {5{neg279[5]}} , neg279[5:1] };

   // m279_75 = W*in
   wire signed [9:0] m279_75;
   assign m279_75 =10'b0;

   // m279_76 = W*in
   wire signed [9:0] m279_76;
   assign m279_76 =10'b0;

   // m279_77 = W*in
   wire signed [9:0] m279_77;
   assign m279_77 =10'b0;

   // m279_78 = W*in
   wire signed [9:0] m279_78;
   assign m279_78 =10'b0;

   // m279_79 = W*in
   wire signed [9:0] m279_79;
   assign m279_79 =10'b0;

   // m279_80 = W*in
   wire signed [9:0] m279_80;
   assign m279_80 =10'b0;

   // m279_81 = W*in
   wire signed [9:0] m279_81;
   assign m279_81 ={ {5{in279[5]}} , in279[5:1] };

   // m279_82 = W*in
   wire signed [9:0] m279_82;
   assign m279_82 =10'b0;

   // m279_83 = W*in
   wire signed [9:0] m279_83;
   assign m279_83 ={ {5{in279[5]}} , in279[5:1] };

   // m279_84 = W*in
   wire signed [9:0] m279_84;
   assign m279_84 =10'b0;

   // m279_85 = W*in
   wire signed [9:0] m279_85;
   assign m279_85 =10'b0;

   // m279_86 = W*in
   wire signed [9:0] m279_86;
   assign m279_86 ={ {5{in279[5]}} , in279[5:1] };

   // m279_87 = W*in
   wire signed [9:0] m279_87;
   assign m279_87 =10'b0;

   // m279_88 = W*in
   wire signed [9:0] m279_88;
   assign m279_88 =10'b0;

   // m279_89 = W*in
   wire signed [9:0] m279_89;
   assign m279_89 =10'b0;

   // m279_90 = W*in
   wire signed [9:0] m279_90;
   assign m279_90 =10'b0;

   // m279_91 = W*in
   wire signed [9:0] m279_91;
   assign m279_91 =10'b0;

   // m279_92 = W*in
   wire signed [9:0] m279_92;
   assign m279_92 =10'b0;

   // m279_93 = W*in
   wire signed [9:0] m279_93;
   assign m279_93 =10'b0;

   // m279_94 = W*in
   wire signed [9:0] m279_94;
   assign m279_94 =10'b0;

   // m279_95 = W*in
   wire signed [9:0] m279_95;
   assign m279_95 =10'b0;

   // m279_96 = W*in
   wire signed [9:0] m279_96;
   assign m279_96 =10'b0;

   // m279_97 = W*in
   wire signed [9:0] m279_97;
   assign m279_97 =10'b0;

   // m279_98 = W*in
   wire signed [9:0] m279_98;
   assign m279_98 =10'b0;

   // m279_99 = W*in
   wire signed [9:0] m279_99;
   assign m279_99 =10'b0;

   // m279_100 = W*in
   wire signed [9:0] m279_100;
   assign m279_100 =10'b0;

   // m279_101 = W*in
   wire signed [9:0] m279_101;
   assign m279_101 =10'b0;

   // m279_102 = W*in
   wire signed [9:0] m279_102;
   assign m279_102 =10'b0;

   // m279_103 = W*in
   wire signed [9:0] m279_103;
   assign m279_103 =10'b0;

   // m279_104 = W*in
   wire signed [9:0] m279_104;
   assign m279_104 =10'b0;

   // m279_105 = W*in
   wire signed [9:0] m279_105;
   assign m279_105 =10'b0;

   // m279_106 = W*in
   wire signed [9:0] m279_106;
   assign m279_106 =10'b0;

   // m279_107 = W*in
   wire signed [9:0] m279_107;
   assign m279_107 =10'b0;

   // m279_108 = W*in
   wire signed [9:0] m279_108;
   assign m279_108 =10'b0;

   // m279_109 = W*in
   wire signed [9:0] m279_109;
   assign m279_109 =10'b0;

   // m279_110 = W*in
   wire signed [9:0] m279_110;
   assign m279_110 =10'b0;

   // m279_111 = W*in
   wire signed [9:0] m279_111;
   assign m279_111 =10'b0;

   // m279_112 = W*in
   wire signed [9:0] m279_112;
   assign m279_112 =10'b0;

   // m279_113 = W*in
   wire signed [9:0] m279_113;
   assign m279_113 =10'b0;

   // m279_114 = W*in
   wire signed [9:0] m279_114;
   assign m279_114 =10'b0;

   // m279_115 = W*in
   wire signed [9:0] m279_115;
   assign m279_115 ={ {5{in279[5]}} , in279[5:1] };

   // m279_116 = W*in
   wire signed [9:0] m279_116;
   assign m279_116 =10'b0;

   // m279_117 = W*in
   wire signed [9:0] m279_117;
   assign m279_117 =10'b0;

   // m280_1 = W*in
   wire signed [9:0] m280_1;
   assign m280_1 =10'b0;

   // m280_2 = W*in
   wire signed [9:0] m280_2;
   assign m280_2 =10'b0;

   // m280_3 = W*in
   wire signed [9:0] m280_3;
   assign m280_3 =10'b0;

   // m280_4 = W*in
   wire signed [9:0] m280_4;
   assign m280_4 =10'b0;

   // m280_5 = W*in
   wire signed [9:0] m280_5;
   assign m280_5 =10'b0;

   // m280_6 = W*in
   wire signed [9:0] m280_6;
   assign m280_6 =10'b0;

   // m280_7 = W*in
   wire signed [9:0] m280_7;
   assign m280_7 =10'b0;

   // m280_8 = W*in
   wire signed [9:0] m280_8;
   assign m280_8 =10'b0;

   // m280_9 = W*in
   wire signed [9:0] m280_9;
   assign m280_9 =10'b0;

   // m280_10 = W*in
   wire signed [9:0] m280_10;
   assign m280_10 =10'b0;

   // m280_11 = W*in
   wire signed [9:0] m280_11;
   assign m280_11 =10'b0;

   // m280_12 = W*in
   wire signed [9:0] m280_12;
   assign m280_12 ={ {4{in280[5]}} , in280[5:0] };

   // m280_13 = W*in
   wire signed [9:0] m280_13;
   assign m280_13 =10'b0;

   // m280_14 = W*in
   wire signed [9:0] m280_14;
   assign m280_14 =10'b0;

   // m280_15 = W*in
   wire signed [9:0] m280_15;
   assign m280_15 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_16 = W*in
   wire signed [9:0] m280_16;
   assign m280_16 =10'b0;

   // m280_17 = W*in
   wire signed [9:0] m280_17;
   assign m280_17 =10'b0;

   // m280_18 = W*in
   wire signed [9:0] m280_18;
   assign m280_18 ={ {5{in280[5]}} , in280[5:1] };

   // m280_19 = W*in
   wire signed [9:0] m280_19;
   assign m280_19 =10'b0;

   // m280_20 = W*in
   wire signed [9:0] m280_20;
   assign m280_20 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_21 = W*in
   wire signed [9:0] m280_21;
   assign m280_21 =10'b0;

   // m280_22 = W*in
   wire signed [9:0] m280_22;
   assign m280_22 =10'b0;

   // m280_23 = W*in
   wire signed [9:0] m280_23;
   assign m280_23 =10'b0;

   // m280_24 = W*in
   wire signed [9:0] m280_24;
   assign m280_24 =10'b0;

   // m280_25 = W*in
   wire signed [9:0] m280_25;
   assign m280_25 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_26 = W*in
   wire signed [9:0] m280_26;
   assign m280_26 =10'b0;

   // m280_27 = W*in
   wire signed [9:0] m280_27;
   assign m280_27 ={ {5{neg280[5]}} , neg280[5:1] };

   // m280_28 = W*in
   wire signed [9:0] m280_28;
   assign m280_28 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_29 = W*in
   wire signed [9:0] m280_29;
   assign m280_29 =10'b0;

   // m280_30 = W*in
   wire signed [9:0] m280_30;
   assign m280_30 =10'b0;

   // m280_31 = W*in
   wire signed [9:0] m280_31;
   assign m280_31 ={ {5{neg280[5]}} , neg280[5:1] };

   // m280_32 = W*in
   wire signed [9:0] m280_32;
   assign m280_32 ={ {5{in280[5]}} , in280[5:1] };

   // m280_33 = W*in
   wire signed [9:0] m280_33;
   assign m280_33 =10'b0;

   // m280_34 = W*in
   wire signed [9:0] m280_34;
   assign m280_34 ={ {5{neg280[5]}} , neg280[5:1] };

   // m280_35 = W*in
   wire signed [9:0] m280_35;
   assign m280_35 =10'b0;

   // m280_36 = W*in
   wire signed [9:0] m280_36;
   assign m280_36 ={ {5{neg280[5]}} , neg280[5:1] };

   // m280_37 = W*in
   wire signed [9:0] m280_37;
   assign m280_37 =10'b0;

   // m280_38 = W*in
   wire signed [9:0] m280_38;
   assign m280_38 =10'b0;

   // m280_39 = W*in
   wire signed [9:0] m280_39;
   assign m280_39 =10'b0;

   // m280_40 = W*in
   wire signed [9:0] m280_40;
   assign m280_40 =10'b0;

   // m280_41 = W*in
   wire signed [9:0] m280_41;
   assign m280_41 =10'b0;

   // m280_42 = W*in
   wire signed [9:0] m280_42;
   assign m280_42 =10'b0;

   // m280_43 = W*in
   wire signed [9:0] m280_43;
   assign m280_43 =10'b0;

   // m280_44 = W*in
   wire signed [9:0] m280_44;
   assign m280_44 =10'b0;

   // m280_45 = W*in
   wire signed [9:0] m280_45;
   assign m280_45 =10'b0;

   // m280_46 = W*in
   wire signed [9:0] m280_46;
   assign m280_46 =10'b0;

   // m280_47 = W*in
   wire signed [9:0] m280_47;
   assign m280_47 =10'b0;

   // m280_48 = W*in
   wire signed [9:0] m280_48;
   assign m280_48 =10'b0;

   // m280_49 = W*in
   wire signed [9:0] m280_49;
   assign m280_49 =10'b0;

   // m280_50 = W*in
   wire signed [9:0] m280_50;
   assign m280_50 =10'b0;

   // m280_51 = W*in
   wire signed [9:0] m280_51;
   assign m280_51 =10'b0;

   // m280_52 = W*in
   wire signed [9:0] m280_52;
   assign m280_52 =10'b0;

   // m280_53 = W*in
   wire signed [9:0] m280_53;
   assign m280_53 =10'b0;

   // m280_54 = W*in
   wire signed [9:0] m280_54;
   assign m280_54 =10'b0;

   // m280_55 = W*in
   wire signed [9:0] m280_55;
   assign m280_55 =10'b0;

   // m280_56 = W*in
   wire signed [9:0] m280_56;
   assign m280_56 =10'b0;

   // m280_57 = W*in
   wire signed [9:0] m280_57;
   assign m280_57 =10'b0;

   // m280_58 = W*in
   wire signed [9:0] m280_58;
   assign m280_58 =10'b0;

   // m280_59 = W*in
   wire signed [9:0] m280_59;
   assign m280_59 =10'b0;

   // m280_60 = W*in
   wire signed [9:0] m280_60;
   assign m280_60 =10'b0;

   // m280_61 = W*in
   wire signed [9:0] m280_61;
   assign m280_61 ={ {4{in280[5]}} , in280[5:0] };

   // m280_62 = W*in
   wire signed [9:0] m280_62;
   assign m280_62 =10'b0;

   // m280_63 = W*in
   wire signed [9:0] m280_63;
   assign m280_63 =10'b0;

   // m280_64 = W*in
   wire signed [9:0] m280_64;
   assign m280_64 ={ {4{in280[5]}} , in280[5:0] };

   // m280_65 = W*in
   wire signed [9:0] m280_65;
   assign m280_65 ={ {5{in280[5]}} , in280[5:1] };

   // m280_66 = W*in
   wire signed [9:0] m280_66;
   assign m280_66 ={ {5{in280[5]}} , in280[5:1] };

   // m280_67 = W*in
   wire signed [9:0] m280_67;
   assign m280_67 =10'b0;

   // m280_68 = W*in
   wire signed [9:0] m280_68;
   assign m280_68 =10'b0;

   // m280_69 = W*in
   wire signed [9:0] m280_69;
   assign m280_69 =10'b0;

   // m280_70 = W*in
   wire signed [9:0] m280_70;
   assign m280_70 ={ {4{in280[5]}} , in280[5:0] };

   // m280_71 = W*in
   wire signed [9:0] m280_71;
   assign m280_71 =10'b0;

   // m280_72 = W*in
   wire signed [9:0] m280_72;
   assign m280_72 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_73 = W*in
   wire signed [9:0] m280_73;
   assign m280_73 =10'b0;

   // m280_74 = W*in
   wire signed [9:0] m280_74;
   assign m280_74 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_75 = W*in
   wire signed [9:0] m280_75;
   assign m280_75 =10'b0;

   // m280_76 = W*in
   wire signed [9:0] m280_76;
   assign m280_76 ={ {4{in280[5]}} , in280[5:0] };

   // m280_77 = W*in
   wire signed [9:0] m280_77;
   assign m280_77 =10'b0;

   // m280_78 = W*in
   wire signed [9:0] m280_78;
   assign m280_78 =10'b0;

   // m280_79 = W*in
   wire signed [9:0] m280_79;
   assign m280_79 =10'b0;

   // m280_80 = W*in
   wire signed [9:0] m280_80;
   assign m280_80 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_81 = W*in
   wire signed [9:0] m280_81;
   assign m280_81 ={ {4{in280[5]}} , in280[5:0] };

   // m280_82 = W*in
   wire signed [9:0] m280_82;
   assign m280_82 =10'b0;

   // m280_83 = W*in
   wire signed [9:0] m280_83;
   assign m280_83 =10'b0;

   // m280_84 = W*in
   wire signed [9:0] m280_84;
   assign m280_84 ={ {5{neg280[5]}} , neg280[5:1] };

   // m280_85 = W*in
   wire signed [9:0] m280_85;
   assign m280_85 =10'b0;

   // m280_86 = W*in
   wire signed [9:0] m280_86;
   assign m280_86 ={ {5{in280[5]}} , in280[5:1] };

   // m280_87 = W*in
   wire signed [9:0] m280_87;
   assign m280_87 =10'b0;

   // m280_88 = W*in
   wire signed [9:0] m280_88;
   assign m280_88 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_89 = W*in
   wire signed [9:0] m280_89;
   assign m280_89 =10'b0;

   // m280_90 = W*in
   wire signed [9:0] m280_90;
   assign m280_90 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_91 = W*in
   wire signed [9:0] m280_91;
   assign m280_91 =10'b0;

   // m280_92 = W*in
   wire signed [9:0] m280_92;
   assign m280_92 =10'b0;

   // m280_93 = W*in
   wire signed [9:0] m280_93;
   assign m280_93 =10'b0;

   // m280_94 = W*in
   wire signed [9:0] m280_94;
   assign m280_94 ={ {4{in280[5]}} , in280[5:0] };

   // m280_95 = W*in
   wire signed [9:0] m280_95;
   assign m280_95 ={ {4{in280[5]}} , in280[5:0] };

   // m280_96 = W*in
   wire signed [9:0] m280_96;
   assign m280_96 =10'b0;

   // m280_97 = W*in
   wire signed [9:0] m280_97;
   assign m280_97 =10'b0;

   // m280_98 = W*in
   wire signed [9:0] m280_98;
   assign m280_98 =10'b0;

   // m280_99 = W*in
   wire signed [9:0] m280_99;
   assign m280_99 =10'b0;

   // m280_100 = W*in
   wire signed [9:0] m280_100;
   assign m280_100 ={ {4{in280[5]}} , in280[5:0] };

   // m280_101 = W*in
   wire signed [9:0] m280_101;
   assign m280_101 =10'b0;

   // m280_102 = W*in
   wire signed [9:0] m280_102;
   assign m280_102 =10'b0;

   // m280_103 = W*in
   wire signed [9:0] m280_103;
   assign m280_103 =10'b0;

   // m280_104 = W*in
   wire signed [9:0] m280_104;
   assign m280_104 =10'b0;

   // m280_105 = W*in
   wire signed [9:0] m280_105;
   assign m280_105 =10'b0;

   // m280_106 = W*in
   wire signed [9:0] m280_106;
   assign m280_106 ={ {5{neg280[5]}} , neg280[5:1] };

   // m280_107 = W*in
   wire signed [9:0] m280_107;
   assign m280_107 =10'b0;

   // m280_108 = W*in
   wire signed [9:0] m280_108;
   assign m280_108 =10'b0;

   // m280_109 = W*in
   wire signed [9:0] m280_109;
   assign m280_109 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_110 = W*in
   wire signed [9:0] m280_110;
   assign m280_110 =10'b0;

   // m280_111 = W*in
   wire signed [9:0] m280_111;
   assign m280_111 ={ {4{neg280[5]}} , neg280[5:0] };

   // m280_112 = W*in
   wire signed [9:0] m280_112;
   assign m280_112 ={ {4{in280[5]}} , in280[5:0] };

   // m280_113 = W*in
   wire signed [9:0] m280_113;
   assign m280_113 =10'b0;

   // m280_114 = W*in
   wire signed [9:0] m280_114;
   assign m280_114 =10'b0;

   // m280_115 = W*in
   wire signed [9:0] m280_115;
   assign m280_115 =10'b0;

   // m280_116 = W*in
   wire signed [9:0] m280_116;
   assign m280_116 =10'b0;

   // m280_117 = W*in
   wire signed [9:0] m280_117;
   assign m280_117 =10'b0;

   // m281_1 = W*in
   wire signed [9:0] m281_1;
   assign m281_1 =10'b0;

   // m281_2 = W*in
   wire signed [9:0] m281_2;
   assign m281_2 =10'b0;

   // m281_3 = W*in
   wire signed [9:0] m281_3;
   assign m281_3 =10'b0;

   // m281_4 = W*in
   wire signed [9:0] m281_4;
   assign m281_4 =10'b0;

   // m281_5 = W*in
   wire signed [9:0] m281_5;
   assign m281_5 =10'b0;

   // m281_6 = W*in
   wire signed [9:0] m281_6;
   assign m281_6 =10'b0;

   // m281_7 = W*in
   wire signed [9:0] m281_7;
   assign m281_7 =10'b0;

   // m281_8 = W*in
   wire signed [9:0] m281_8;
   assign m281_8 =10'b0;

   // m281_9 = W*in
   wire signed [9:0] m281_9;
   assign m281_9 =10'b0;

   // m281_10 = W*in
   wire signed [9:0] m281_10;
   assign m281_10 ={ {4{in281[5]}} , in281[5:0] };

   // m281_11 = W*in
   wire signed [9:0] m281_11;
   assign m281_11 =10'b0;

   // m281_12 = W*in
   wire signed [9:0] m281_12;
   assign m281_12 =10'b0;

   // m281_13 = W*in
   wire signed [9:0] m281_13;
   assign m281_13 =10'b0;

   // m281_14 = W*in
   wire signed [9:0] m281_14;
   assign m281_14 ={ {4{in281[5]}} , in281[5:0] };

   // m281_15 = W*in
   wire signed [9:0] m281_15;
   assign m281_15 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_16 = W*in
   wire signed [9:0] m281_16;
   assign m281_16 =10'b0;

   // m281_17 = W*in
   wire signed [9:0] m281_17;
   assign m281_17 =10'b0;

   // m281_18 = W*in
   wire signed [9:0] m281_18;
   assign m281_18 =10'b0;

   // m281_19 = W*in
   wire signed [9:0] m281_19;
   assign m281_19 =10'b0;

   // m281_20 = W*in
   wire signed [9:0] m281_20;
   assign m281_20 =10'b0;

   // m281_21 = W*in
   wire signed [9:0] m281_21;
   assign m281_21 ={ {4{in281[5]}} , in281[5:0] };

   // m281_22 = W*in
   wire signed [9:0] m281_22;
   assign m281_22 =10'b0;

   // m281_23 = W*in
   wire signed [9:0] m281_23;
   assign m281_23 =10'b0;

   // m281_24 = W*in
   wire signed [9:0] m281_24;
   assign m281_24 =10'b0;

   // m281_25 = W*in
   wire signed [9:0] m281_25;
   assign m281_25 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_26 = W*in
   wire signed [9:0] m281_26;
   assign m281_26 =10'b0;

   // m281_27 = W*in
   wire signed [9:0] m281_27;
   assign m281_27 ={ {5{neg281[5]}} , neg281[5:1] };

   // m281_28 = W*in
   wire signed [9:0] m281_28;
   assign m281_28 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_29 = W*in
   wire signed [9:0] m281_29;
   assign m281_29 =10'b0;

   // m281_30 = W*in
   wire signed [9:0] m281_30;
   assign m281_30 =10'b0;

   // m281_31 = W*in
   wire signed [9:0] m281_31;
   assign m281_31 ={ {5{neg281[5]}} , neg281[5:1] };

   // m281_32 = W*in
   wire signed [9:0] m281_32;
   assign m281_32 ={ {5{in281[5]}} , in281[5:1] };

   // m281_33 = W*in
   wire signed [9:0] m281_33;
   assign m281_33 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_34 = W*in
   wire signed [9:0] m281_34;
   assign m281_34 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_35 = W*in
   wire signed [9:0] m281_35;
   assign m281_35 =10'b0;

   // m281_36 = W*in
   wire signed [9:0] m281_36;
   assign m281_36 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_37 = W*in
   wire signed [9:0] m281_37;
   assign m281_37 =10'b0;

   // m281_38 = W*in
   wire signed [9:0] m281_38;
   assign m281_38 =10'b0;

   // m281_39 = W*in
   wire signed [9:0] m281_39;
   assign m281_39 =10'b0;

   // m281_40 = W*in
   wire signed [9:0] m281_40;
   assign m281_40 =10'b0;

   // m281_41 = W*in
   wire signed [9:0] m281_41;
   assign m281_41 =10'b0;

   // m281_42 = W*in
   wire signed [9:0] m281_42;
   assign m281_42 ={ {4{in281[5]}} , in281[5:0] };

   // m281_43 = W*in
   wire signed [9:0] m281_43;
   assign m281_43 =10'b0;

   // m281_44 = W*in
   wire signed [9:0] m281_44;
   assign m281_44 =10'b0;

   // m281_45 = W*in
   wire signed [9:0] m281_45;
   assign m281_45 =10'b0;

   // m281_46 = W*in
   wire signed [9:0] m281_46;
   assign m281_46 =10'b0;

   // m281_47 = W*in
   wire signed [9:0] m281_47;
   assign m281_47 =10'b0;

   // m281_48 = W*in
   wire signed [9:0] m281_48;
   assign m281_48 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_49 = W*in
   wire signed [9:0] m281_49;
   assign m281_49 =10'b0;

   // m281_50 = W*in
   wire signed [9:0] m281_50;
   assign m281_50 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_51 = W*in
   wire signed [9:0] m281_51;
   assign m281_51 =10'b0;

   // m281_52 = W*in
   wire signed [9:0] m281_52;
   assign m281_52 =10'b0;

   // m281_53 = W*in
   wire signed [9:0] m281_53;
   assign m281_53 =10'b0;

   // m281_54 = W*in
   wire signed [9:0] m281_54;
   assign m281_54 =10'b0;

   // m281_55 = W*in
   wire signed [9:0] m281_55;
   assign m281_55 =10'b0;

   // m281_56 = W*in
   wire signed [9:0] m281_56;
   assign m281_56 =10'b0;

   // m281_57 = W*in
   wire signed [9:0] m281_57;
   assign m281_57 =10'b0;

   // m281_58 = W*in
   wire signed [9:0] m281_58;
   assign m281_58 =10'b0;

   // m281_59 = W*in
   wire signed [9:0] m281_59;
   assign m281_59 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_60 = W*in
   wire signed [9:0] m281_60;
   assign m281_60 =10'b0;

   // m281_61 = W*in
   wire signed [9:0] m281_61;
   assign m281_61 =10'b0;

   // m281_62 = W*in
   wire signed [9:0] m281_62;
   assign m281_62 =10'b0;

   // m281_63 = W*in
   wire signed [9:0] m281_63;
   assign m281_63 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_64 = W*in
   wire signed [9:0] m281_64;
   assign m281_64 ={ {4{in281[5]}} , in281[5:0] };

   // m281_65 = W*in
   wire signed [9:0] m281_65;
   assign m281_65 ={ {4{in281[5]}} , in281[5:0] };

   // m281_66 = W*in
   wire signed [9:0] m281_66;
   assign m281_66 ={ {4{in281[5]}} , in281[5:0] };

   // m281_67 = W*in
   wire signed [9:0] m281_67;
   assign m281_67 =10'b0;

   // m281_68 = W*in
   wire signed [9:0] m281_68;
   assign m281_68 =10'b0;

   // m281_69 = W*in
   wire signed [9:0] m281_69;
   assign m281_69 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_70 = W*in
   wire signed [9:0] m281_70;
   assign m281_70 =10'b0;

   // m281_71 = W*in
   wire signed [9:0] m281_71;
   assign m281_71 =10'b0;

   // m281_72 = W*in
   wire signed [9:0] m281_72;
   assign m281_72 =10'b0;

   // m281_73 = W*in
   wire signed [9:0] m281_73;
   assign m281_73 ={ {5{neg281[5]}} , neg281[5:1] };

   // m281_74 = W*in
   wire signed [9:0] m281_74;
   assign m281_74 ={ {4{in281[5]}} , in281[5:0] };

   // m281_75 = W*in
   wire signed [9:0] m281_75;
   assign m281_75 =10'b0;

   // m281_76 = W*in
   wire signed [9:0] m281_76;
   assign m281_76 =10'b0;

   // m281_77 = W*in
   wire signed [9:0] m281_77;
   assign m281_77 =10'b0;

   // m281_78 = W*in
   wire signed [9:0] m281_78;
   assign m281_78 =10'b0;

   // m281_79 = W*in
   wire signed [9:0] m281_79;
   assign m281_79 ={ {4{in281[5]}} , in281[5:0] };

   // m281_80 = W*in
   wire signed [9:0] m281_80;
   assign m281_80 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_81 = W*in
   wire signed [9:0] m281_81;
   assign m281_81 ={ {4{in281[5]}} , in281[5:0] };

   // m281_82 = W*in
   wire signed [9:0] m281_82;
   assign m281_82 =10'b0;

   // m281_83 = W*in
   wire signed [9:0] m281_83;
   assign m281_83 ={ {5{neg281[5]}} , neg281[5:1] };

   // m281_84 = W*in
   wire signed [9:0] m281_84;
   assign m281_84 ={ {5{neg281[5]}} , neg281[5:1] };

   // m281_85 = W*in
   wire signed [9:0] m281_85;
   assign m281_85 =10'b0;

   // m281_86 = W*in
   wire signed [9:0] m281_86;
   assign m281_86 =10'b0;

   // m281_87 = W*in
   wire signed [9:0] m281_87;
   assign m281_87 =10'b0;

   // m281_88 = W*in
   wire signed [9:0] m281_88;
   assign m281_88 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_89 = W*in
   wire signed [9:0] m281_89;
   assign m281_89 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_90 = W*in
   wire signed [9:0] m281_90;
   assign m281_90 =10'b0;

   // m281_91 = W*in
   wire signed [9:0] m281_91;
   assign m281_91 =10'b0;

   // m281_92 = W*in
   wire signed [9:0] m281_92;
   assign m281_92 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_93 = W*in
   wire signed [9:0] m281_93;
   assign m281_93 =10'b0;

   // m281_94 = W*in
   wire signed [9:0] m281_94;
   assign m281_94 =10'b0;

   // m281_95 = W*in
   wire signed [9:0] m281_95;
   assign m281_95 =10'b0;

   // m281_96 = W*in
   wire signed [9:0] m281_96;
   assign m281_96 =10'b0;

   // m281_97 = W*in
   wire signed [9:0] m281_97;
   assign m281_97 =10'b0;

   // m281_98 = W*in
   wire signed [9:0] m281_98;
   assign m281_98 =10'b0;

   // m281_99 = W*in
   wire signed [9:0] m281_99;
   assign m281_99 =10'b0;

   // m281_100 = W*in
   wire signed [9:0] m281_100;
   assign m281_100 =10'b0;

   // m281_101 = W*in
   wire signed [9:0] m281_101;
   assign m281_101 =10'b0;

   // m281_102 = W*in
   wire signed [9:0] m281_102;
   assign m281_102 =10'b0;

   // m281_103 = W*in
   wire signed [9:0] m281_103;
   assign m281_103 =10'b0;

   // m281_104 = W*in
   wire signed [9:0] m281_104;
   assign m281_104 =10'b0;

   // m281_105 = W*in
   wire signed [9:0] m281_105;
   assign m281_105 =10'b0;

   // m281_106 = W*in
   wire signed [9:0] m281_106;
   assign m281_106 =10'b0;

   // m281_107 = W*in
   wire signed [9:0] m281_107;
   assign m281_107 ={ {4{in281[5]}} , in281[5:0] };

   // m281_108 = W*in
   wire signed [9:0] m281_108;
   assign m281_108 =10'b0;

   // m281_109 = W*in
   wire signed [9:0] m281_109;
   assign m281_109 =10'b0;

   // m281_110 = W*in
   wire signed [9:0] m281_110;
   assign m281_110 ={ {4{in281[5]}} , in281[5:0] };

   // m281_111 = W*in
   wire signed [9:0] m281_111;
   assign m281_111 ={ {4{neg281[5]}} , neg281[5:0] };

   // m281_112 = W*in
   wire signed [9:0] m281_112;
   assign m281_112 =10'b0;

   // m281_113 = W*in
   wire signed [9:0] m281_113;
   assign m281_113 =10'b0;

   // m281_114 = W*in
   wire signed [9:0] m281_114;
   assign m281_114 =10'b0;

   // m281_115 = W*in
   wire signed [9:0] m281_115;
   assign m281_115 =10'b0;

   // m281_116 = W*in
   wire signed [9:0] m281_116;
   assign m281_116 =10'b0;

   // m281_117 = W*in
   wire signed [9:0] m281_117;
   assign m281_117 =10'b0;

   // m282_1 = W*in
   wire signed [9:0] m282_1;
   assign m282_1 ={ {4{in282[5]}} , in282[5:0] };

   // m282_2 = W*in
   wire signed [9:0] m282_2;
   assign m282_2 =10'b0;

   // m282_3 = W*in
   wire signed [9:0] m282_3;
   assign m282_3 =10'b0;

   // m282_4 = W*in
   wire signed [9:0] m282_4;
   assign m282_4 =10'b0;

   // m282_5 = W*in
   wire signed [9:0] m282_5;
   assign m282_5 =10'b0;

   // m282_6 = W*in
   wire signed [9:0] m282_6;
   assign m282_6 =10'b0;

   // m282_7 = W*in
   wire signed [9:0] m282_7;
   assign m282_7 =10'b0;

   // m282_8 = W*in
   wire signed [9:0] m282_8;
   assign m282_8 =10'b0;

   // m282_9 = W*in
   wire signed [9:0] m282_9;
   assign m282_9 =10'b0;

   // m282_10 = W*in
   wire signed [9:0] m282_10;
   assign m282_10 =10'b0;

   // m282_11 = W*in
   wire signed [9:0] m282_11;
   assign m282_11 ={ {4{in282[5]}} , in282[5:0] };

   // m282_12 = W*in
   wire signed [9:0] m282_12;
   assign m282_12 =10'b0;

   // m282_13 = W*in
   wire signed [9:0] m282_13;
   assign m282_13 =10'b0;

   // m282_14 = W*in
   wire signed [9:0] m282_14;
   assign m282_14 =10'b0;

   // m282_15 = W*in
   wire signed [9:0] m282_15;
   assign m282_15 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_16 = W*in
   wire signed [9:0] m282_16;
   assign m282_16 =10'b0;

   // m282_17 = W*in
   wire signed [9:0] m282_17;
   assign m282_17 =10'b0;

   // m282_18 = W*in
   wire signed [9:0] m282_18;
   assign m282_18 =10'b0;

   // m282_19 = W*in
   wire signed [9:0] m282_19;
   assign m282_19 =10'b0;

   // m282_20 = W*in
   wire signed [9:0] m282_20;
   assign m282_20 =10'b0;

   // m282_21 = W*in
   wire signed [9:0] m282_21;
   assign m282_21 ={ {5{neg282[5]}} , neg282[5:1] };

   // m282_22 = W*in
   wire signed [9:0] m282_22;
   assign m282_22 =10'b0;

   // m282_23 = W*in
   wire signed [9:0] m282_23;
   assign m282_23 =10'b0;

   // m282_24 = W*in
   wire signed [9:0] m282_24;
   assign m282_24 =10'b0;

   // m282_25 = W*in
   wire signed [9:0] m282_25;
   assign m282_25 =10'b0;

   // m282_26 = W*in
   wire signed [9:0] m282_26;
   assign m282_26 ={ {4{in282[5]}} , in282[5:0] };

   // m282_27 = W*in
   wire signed [9:0] m282_27;
   assign m282_27 ={ {5{neg282[5]}} , neg282[5:1] };

   // m282_28 = W*in
   wire signed [9:0] m282_28;
   assign m282_28 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_29 = W*in
   wire signed [9:0] m282_29;
   assign m282_29 =10'b0;

   // m282_30 = W*in
   wire signed [9:0] m282_30;
   assign m282_30 =10'b0;

   // m282_31 = W*in
   wire signed [9:0] m282_31;
   assign m282_31 ={ {5{neg282[5]}} , neg282[5:1] };

   // m282_32 = W*in
   wire signed [9:0] m282_32;
   assign m282_32 ={ {4{in282[5]}} , in282[5:0] };

   // m282_33 = W*in
   wire signed [9:0] m282_33;
   assign m282_33 =10'b0;

   // m282_34 = W*in
   wire signed [9:0] m282_34;
   assign m282_34 =10'b0;

   // m282_35 = W*in
   wire signed [9:0] m282_35;
   assign m282_35 =10'b0;

   // m282_36 = W*in
   wire signed [9:0] m282_36;
   assign m282_36 =10'b0;

   // m282_37 = W*in
   wire signed [9:0] m282_37;
   assign m282_37 =10'b0;

   // m282_38 = W*in
   wire signed [9:0] m282_38;
   assign m282_38 =10'b0;

   // m282_39 = W*in
   wire signed [9:0] m282_39;
   assign m282_39 =10'b0;

   // m282_40 = W*in
   wire signed [9:0] m282_40;
   assign m282_40 =10'b0;

   // m282_41 = W*in
   wire signed [9:0] m282_41;
   assign m282_41 =10'b0;

   // m282_42 = W*in
   wire signed [9:0] m282_42;
   assign m282_42 =10'b0;

   // m282_43 = W*in
   wire signed [9:0] m282_43;
   assign m282_43 =10'b0;

   // m282_44 = W*in
   wire signed [9:0] m282_44;
   assign m282_44 =10'b0;

   // m282_45 = W*in
   wire signed [9:0] m282_45;
   assign m282_45 ={ {4{in282[5]}} , in282[5:0] };

   // m282_46 = W*in
   wire signed [9:0] m282_46;
   assign m282_46 =10'b0;

   // m282_47 = W*in
   wire signed [9:0] m282_47;
   assign m282_47 =10'b0;

   // m282_48 = W*in
   wire signed [9:0] m282_48;
   assign m282_48 =10'b0;

   // m282_49 = W*in
   wire signed [9:0] m282_49;
   assign m282_49 =10'b0;

   // m282_50 = W*in
   wire signed [9:0] m282_50;
   assign m282_50 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_51 = W*in
   wire signed [9:0] m282_51;
   assign m282_51 =10'b0;

   // m282_52 = W*in
   wire signed [9:0] m282_52;
   assign m282_52 =10'b0;

   // m282_53 = W*in
   wire signed [9:0] m282_53;
   assign m282_53 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_54 = W*in
   wire signed [9:0] m282_54;
   assign m282_54 =10'b0;

   // m282_55 = W*in
   wire signed [9:0] m282_55;
   assign m282_55 =10'b0;

   // m282_56 = W*in
   wire signed [9:0] m282_56;
   assign m282_56 =10'b0;

   // m282_57 = W*in
   wire signed [9:0] m282_57;
   assign m282_57 =10'b0;

   // m282_58 = W*in
   wire signed [9:0] m282_58;
   assign m282_58 =10'b0;

   // m282_59 = W*in
   wire signed [9:0] m282_59;
   assign m282_59 =10'b0;

   // m282_60 = W*in
   wire signed [9:0] m282_60;
   assign m282_60 =10'b0;

   // m282_61 = W*in
   wire signed [9:0] m282_61;
   assign m282_61 =10'b0;

   // m282_62 = W*in
   wire signed [9:0] m282_62;
   assign m282_62 =10'b0;

   // m282_63 = W*in
   wire signed [9:0] m282_63;
   assign m282_63 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_64 = W*in
   wire signed [9:0] m282_64;
   assign m282_64 =10'b0;

   // m282_65 = W*in
   wire signed [9:0] m282_65;
   assign m282_65 =10'b0;

   // m282_66 = W*in
   wire signed [9:0] m282_66;
   assign m282_66 =10'b0;

   // m282_67 = W*in
   wire signed [9:0] m282_67;
   assign m282_67 =10'b0;

   // m282_68 = W*in
   wire signed [9:0] m282_68;
   assign m282_68 =10'b0;

   // m282_69 = W*in
   wire signed [9:0] m282_69;
   assign m282_69 ={ {3{neg282[5]}} , neg282 , {1{1'b0}} };

   // m282_70 = W*in
   wire signed [9:0] m282_70;
   assign m282_70 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_71 = W*in
   wire signed [9:0] m282_71;
   assign m282_71 =10'b0;

   // m282_72 = W*in
   wire signed [9:0] m282_72;
   assign m282_72 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_73 = W*in
   wire signed [9:0] m282_73;
   assign m282_73 =10'b0;

   // m282_74 = W*in
   wire signed [9:0] m282_74;
   assign m282_74 ={ {5{in282[5]}} , in282[5:1] };

   // m282_75 = W*in
   wire signed [9:0] m282_75;
   assign m282_75 =10'b0;

   // m282_76 = W*in
   wire signed [9:0] m282_76;
   assign m282_76 =10'b0;

   // m282_77 = W*in
   wire signed [9:0] m282_77;
   assign m282_77 =10'b0;

   // m282_78 = W*in
   wire signed [9:0] m282_78;
   assign m282_78 =10'b0;

   // m282_79 = W*in
   wire signed [9:0] m282_79;
   assign m282_79 =10'b0;

   // m282_80 = W*in
   wire signed [9:0] m282_80;
   assign m282_80 =10'b0;

   // m282_81 = W*in
   wire signed [9:0] m282_81;
   assign m282_81 =10'b0;

   // m282_82 = W*in
   wire signed [9:0] m282_82;
   assign m282_82 ={ {3{neg282[5]}} , neg282 , {1{1'b0}} };

   // m282_83 = W*in
   wire signed [9:0] m282_83;
   assign m282_83 ={ {5{in282[5]}} , in282[5:1] };

   // m282_84 = W*in
   wire signed [9:0] m282_84;
   assign m282_84 =10'b0;

   // m282_85 = W*in
   wire signed [9:0] m282_85;
   assign m282_85 =10'b0;

   // m282_86 = W*in
   wire signed [9:0] m282_86;
   assign m282_86 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_87 = W*in
   wire signed [9:0] m282_87;
   assign m282_87 =10'b0;

   // m282_88 = W*in
   wire signed [9:0] m282_88;
   assign m282_88 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_89 = W*in
   wire signed [9:0] m282_89;
   assign m282_89 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_90 = W*in
   wire signed [9:0] m282_90;
   assign m282_90 =10'b0;

   // m282_91 = W*in
   wire signed [9:0] m282_91;
   assign m282_91 =10'b0;

   // m282_92 = W*in
   wire signed [9:0] m282_92;
   assign m282_92 ={ {4{neg282[5]}} , neg282[5:0] };

   // m282_93 = W*in
   wire signed [9:0] m282_93;
   assign m282_93 =10'b0;

   // m282_94 = W*in
   wire signed [9:0] m282_94;
   assign m282_94 =10'b0;

   // m282_95 = W*in
   wire signed [9:0] m282_95;
   assign m282_95 =10'b0;

   // m282_96 = W*in
   wire signed [9:0] m282_96;
   assign m282_96 =10'b0;

   // m282_97 = W*in
   wire signed [9:0] m282_97;
   assign m282_97 =10'b0;

   // m282_98 = W*in
   wire signed [9:0] m282_98;
   assign m282_98 =10'b0;

   // m282_99 = W*in
   wire signed [9:0] m282_99;
   assign m282_99 =10'b0;

   // m282_100 = W*in
   wire signed [9:0] m282_100;
   assign m282_100 =10'b0;

   // m282_101 = W*in
   wire signed [9:0] m282_101;
   assign m282_101 =10'b0;

   // m282_102 = W*in
   wire signed [9:0] m282_102;
   assign m282_102 =10'b0;

   // m282_103 = W*in
   wire signed [9:0] m282_103;
   assign m282_103 =10'b0;

   // m282_104 = W*in
   wire signed [9:0] m282_104;
   assign m282_104 ={ {4{in282[5]}} , in282[5:0] };

   // m282_105 = W*in
   wire signed [9:0] m282_105;
   assign m282_105 =10'b0;

   // m282_106 = W*in
   wire signed [9:0] m282_106;
   assign m282_106 =10'b0;

   // m282_107 = W*in
   wire signed [9:0] m282_107;
   assign m282_107 ={ {4{in282[5]}} , in282[5:0] };

   // m282_108 = W*in
   wire signed [9:0] m282_108;
   assign m282_108 =10'b0;

   // m282_109 = W*in
   wire signed [9:0] m282_109;
   assign m282_109 ={ {5{neg282[5]}} , neg282[5:1] };

   // m282_110 = W*in
   wire signed [9:0] m282_110;
   assign m282_110 =10'b0;

   // m282_111 = W*in
   wire signed [9:0] m282_111;
   assign m282_111 =10'b0;

   // m282_112 = W*in
   wire signed [9:0] m282_112;
   assign m282_112 =10'b0;

   // m282_113 = W*in
   wire signed [9:0] m282_113;
   assign m282_113 =10'b0;

   // m282_114 = W*in
   wire signed [9:0] m282_114;
   assign m282_114 ={ {5{neg282[5]}} , neg282[5:1] };

   // m282_115 = W*in
   wire signed [9:0] m282_115;
   assign m282_115 ={ {4{in282[5]}} , in282[5:0] };

   // m282_116 = W*in
   wire signed [9:0] m282_116;
   assign m282_116 =10'b0;

   // m282_117 = W*in
   wire signed [9:0] m282_117;
   assign m282_117 =10'b0;

   // m283_1 = W*in
   wire signed [9:0] m283_1;
   assign m283_1 =10'b0;

   // m283_2 = W*in
   wire signed [9:0] m283_2;
   assign m283_2 =10'b0;

   // m283_3 = W*in
   wire signed [9:0] m283_3;
   assign m283_3 =10'b0;

   // m283_4 = W*in
   wire signed [9:0] m283_4;
   assign m283_4 =10'b0;

   // m283_5 = W*in
   wire signed [9:0] m283_5;
   assign m283_5 =10'b0;

   // m283_6 = W*in
   wire signed [9:0] m283_6;
   assign m283_6 =10'b0;

   // m283_7 = W*in
   wire signed [9:0] m283_7;
   assign m283_7 =10'b0;

   // m283_8 = W*in
   wire signed [9:0] m283_8;
   assign m283_8 =10'b0;

   // m283_9 = W*in
   wire signed [9:0] m283_9;
   assign m283_9 =10'b0;

   // m283_10 = W*in
   wire signed [9:0] m283_10;
   assign m283_10 =10'b0;

   // m283_11 = W*in
   wire signed [9:0] m283_11;
   assign m283_11 =10'b0;

   // m283_12 = W*in
   wire signed [9:0] m283_12;
   assign m283_12 =10'b0;

   // m283_13 = W*in
   wire signed [9:0] m283_13;
   assign m283_13 =10'b0;

   // m283_14 = W*in
   wire signed [9:0] m283_14;
   assign m283_14 =10'b0;

   // m283_15 = W*in
   wire signed [9:0] m283_15;
   assign m283_15 =10'b0;

   // m283_16 = W*in
   wire signed [9:0] m283_16;
   assign m283_16 =10'b0;

   // m283_17 = W*in
   wire signed [9:0] m283_17;
   assign m283_17 =10'b0;

   // m283_18 = W*in
   wire signed [9:0] m283_18;
   assign m283_18 =10'b0;

   // m283_19 = W*in
   wire signed [9:0] m283_19;
   assign m283_19 =10'b0;

   // m283_20 = W*in
   wire signed [9:0] m283_20;
   assign m283_20 =10'b0;

   // m283_21 = W*in
   wire signed [9:0] m283_21;
   assign m283_21 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_22 = W*in
   wire signed [9:0] m283_22;
   assign m283_22 =10'b0;

   // m283_23 = W*in
   wire signed [9:0] m283_23;
   assign m283_23 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_24 = W*in
   wire signed [9:0] m283_24;
   assign m283_24 =10'b0;

   // m283_25 = W*in
   wire signed [9:0] m283_25;
   assign m283_25 ={ {5{in283[5]}} , in283[5:1] };

   // m283_26 = W*in
   wire signed [9:0] m283_26;
   assign m283_26 =10'b0;

   // m283_27 = W*in
   wire signed [9:0] m283_27;
   assign m283_27 =10'b0;

   // m283_28 = W*in
   wire signed [9:0] m283_28;
   assign m283_28 ={ {5{in283[5]}} , in283[5:1] };

   // m283_29 = W*in
   wire signed [9:0] m283_29;
   assign m283_29 =10'b0;

   // m283_30 = W*in
   wire signed [9:0] m283_30;
   assign m283_30 =10'b0;

   // m283_31 = W*in
   wire signed [9:0] m283_31;
   assign m283_31 =10'b0;

   // m283_32 = W*in
   wire signed [9:0] m283_32;
   assign m283_32 =10'b0;

   // m283_33 = W*in
   wire signed [9:0] m283_33;
   assign m283_33 =10'b0;

   // m283_34 = W*in
   wire signed [9:0] m283_34;
   assign m283_34 ={ {5{neg283[5]}} , neg283[5:1] };

   // m283_35 = W*in
   wire signed [9:0] m283_35;
   assign m283_35 ={ {5{neg283[5]}} , neg283[5:1] };

   // m283_36 = W*in
   wire signed [9:0] m283_36;
   assign m283_36 ={ {5{in283[5]}} , in283[5:1] };

   // m283_37 = W*in
   wire signed [9:0] m283_37;
   assign m283_37 =10'b0;

   // m283_38 = W*in
   wire signed [9:0] m283_38;
   assign m283_38 =10'b0;

   // m283_39 = W*in
   wire signed [9:0] m283_39;
   assign m283_39 =10'b0;

   // m283_40 = W*in
   wire signed [9:0] m283_40;
   assign m283_40 =10'b0;

   // m283_41 = W*in
   wire signed [9:0] m283_41;
   assign m283_41 =10'b0;

   // m283_42 = W*in
   wire signed [9:0] m283_42;
   assign m283_42 =10'b0;

   // m283_43 = W*in
   wire signed [9:0] m283_43;
   assign m283_43 ={ {4{in283[5]}} , in283[5:0] };

   // m283_44 = W*in
   wire signed [9:0] m283_44;
   assign m283_44 =10'b0;

   // m283_45 = W*in
   wire signed [9:0] m283_45;
   assign m283_45 ={ {4{in283[5]}} , in283[5:0] };

   // m283_46 = W*in
   wire signed [9:0] m283_46;
   assign m283_46 =10'b0;

   // m283_47 = W*in
   wire signed [9:0] m283_47;
   assign m283_47 =10'b0;

   // m283_48 = W*in
   wire signed [9:0] m283_48;
   assign m283_48 ={ {4{in283[5]}} , in283[5:0] };

   // m283_49 = W*in
   wire signed [9:0] m283_49;
   assign m283_49 =10'b0;

   // m283_50 = W*in
   wire signed [9:0] m283_50;
   assign m283_50 =10'b0;

   // m283_51 = W*in
   wire signed [9:0] m283_51;
   assign m283_51 =10'b0;

   // m283_52 = W*in
   wire signed [9:0] m283_52;
   assign m283_52 =10'b0;

   // m283_53 = W*in
   wire signed [9:0] m283_53;
   assign m283_53 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_54 = W*in
   wire signed [9:0] m283_54;
   assign m283_54 =10'b0;

   // m283_55 = W*in
   wire signed [9:0] m283_55;
   assign m283_55 =10'b0;

   // m283_56 = W*in
   wire signed [9:0] m283_56;
   assign m283_56 =10'b0;

   // m283_57 = W*in
   wire signed [9:0] m283_57;
   assign m283_57 =10'b0;

   // m283_58 = W*in
   wire signed [9:0] m283_58;
   assign m283_58 =10'b0;

   // m283_59 = W*in
   wire signed [9:0] m283_59;
   assign m283_59 =10'b0;

   // m283_60 = W*in
   wire signed [9:0] m283_60;
   assign m283_60 =10'b0;

   // m283_61 = W*in
   wire signed [9:0] m283_61;
   assign m283_61 =10'b0;

   // m283_62 = W*in
   wire signed [9:0] m283_62;
   assign m283_62 =10'b0;

   // m283_63 = W*in
   wire signed [9:0] m283_63;
   assign m283_63 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_64 = W*in
   wire signed [9:0] m283_64;
   assign m283_64 =10'b0;

   // m283_65 = W*in
   wire signed [9:0] m283_65;
   assign m283_65 ={ {5{neg283[5]}} , neg283[5:1] };

   // m283_66 = W*in
   wire signed [9:0] m283_66;
   assign m283_66 =10'b0;

   // m283_67 = W*in
   wire signed [9:0] m283_67;
   assign m283_67 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_68 = W*in
   wire signed [9:0] m283_68;
   assign m283_68 =10'b0;

   // m283_69 = W*in
   wire signed [9:0] m283_69;
   assign m283_69 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_70 = W*in
   wire signed [9:0] m283_70;
   assign m283_70 ={ {5{neg283[5]}} , neg283[5:1] };

   // m283_71 = W*in
   wire signed [9:0] m283_71;
   assign m283_71 ={ {5{in283[5]}} , in283[5:1] };

   // m283_72 = W*in
   wire signed [9:0] m283_72;
   assign m283_72 =10'b0;

   // m283_73 = W*in
   wire signed [9:0] m283_73;
   assign m283_73 =10'b0;

   // m283_74 = W*in
   wire signed [9:0] m283_74;
   assign m283_74 =10'b0;

   // m283_75 = W*in
   wire signed [9:0] m283_75;
   assign m283_75 =10'b0;

   // m283_76 = W*in
   wire signed [9:0] m283_76;
   assign m283_76 =10'b0;

   // m283_77 = W*in
   wire signed [9:0] m283_77;
   assign m283_77 =10'b0;

   // m283_78 = W*in
   wire signed [9:0] m283_78;
   assign m283_78 =10'b0;

   // m283_79 = W*in
   wire signed [9:0] m283_79;
   assign m283_79 =10'b0;

   // m283_80 = W*in
   wire signed [9:0] m283_80;
   assign m283_80 =10'b0;

   // m283_81 = W*in
   wire signed [9:0] m283_81;
   assign m283_81 =10'b0;

   // m283_82 = W*in
   wire signed [9:0] m283_82;
   assign m283_82 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_83 = W*in
   wire signed [9:0] m283_83;
   assign m283_83 ={ {5{in283[5]}} , in283[5:1] };

   // m283_84 = W*in
   wire signed [9:0] m283_84;
   assign m283_84 ={ {5{in283[5]}} , in283[5:1] };

   // m283_85 = W*in
   wire signed [9:0] m283_85;
   assign m283_85 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_86 = W*in
   wire signed [9:0] m283_86;
   assign m283_86 =10'b0;

   // m283_87 = W*in
   wire signed [9:0] m283_87;
   assign m283_87 =10'b0;

   // m283_88 = W*in
   wire signed [9:0] m283_88;
   assign m283_88 =10'b0;

   // m283_89 = W*in
   wire signed [9:0] m283_89;
   assign m283_89 =10'b0;

   // m283_90 = W*in
   wire signed [9:0] m283_90;
   assign m283_90 =10'b0;

   // m283_91 = W*in
   wire signed [9:0] m283_91;
   assign m283_91 =10'b0;

   // m283_92 = W*in
   wire signed [9:0] m283_92;
   assign m283_92 =10'b0;

   // m283_93 = W*in
   wire signed [9:0] m283_93;
   assign m283_93 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_94 = W*in
   wire signed [9:0] m283_94;
   assign m283_94 =10'b0;

   // m283_95 = W*in
   wire signed [9:0] m283_95;
   assign m283_95 =10'b0;

   // m283_96 = W*in
   wire signed [9:0] m283_96;
   assign m283_96 =10'b0;

   // m283_97 = W*in
   wire signed [9:0] m283_97;
   assign m283_97 =10'b0;

   // m283_98 = W*in
   wire signed [9:0] m283_98;
   assign m283_98 =10'b0;

   // m283_99 = W*in
   wire signed [9:0] m283_99;
   assign m283_99 =10'b0;

   // m283_100 = W*in
   wire signed [9:0] m283_100;
   assign m283_100 =10'b0;

   // m283_101 = W*in
   wire signed [9:0] m283_101;
   assign m283_101 =10'b0;

   // m283_102 = W*in
   wire signed [9:0] m283_102;
   assign m283_102 =10'b0;

   // m283_103 = W*in
   wire signed [9:0] m283_103;
   assign m283_103 =10'b0;

   // m283_104 = W*in
   wire signed [9:0] m283_104;
   assign m283_104 ={ {4{in283[5]}} , in283[5:0] };

   // m283_105 = W*in
   wire signed [9:0] m283_105;
   assign m283_105 =10'b0;

   // m283_106 = W*in
   wire signed [9:0] m283_106;
   assign m283_106 =10'b0;

   // m283_107 = W*in
   wire signed [9:0] m283_107;
   assign m283_107 =10'b0;

   // m283_108 = W*in
   wire signed [9:0] m283_108;
   assign m283_108 ={ {5{neg283[5]}} , neg283[5:1] };

   // m283_109 = W*in
   wire signed [9:0] m283_109;
   assign m283_109 ={ {4{neg283[5]}} , neg283[5:0] };

   // m283_110 = W*in
   wire signed [9:0] m283_110;
   assign m283_110 =10'b0;

   // m283_111 = W*in
   wire signed [9:0] m283_111;
   assign m283_111 =10'b0;

   // m283_112 = W*in
   wire signed [9:0] m283_112;
   assign m283_112 =10'b0;

   // m283_113 = W*in
   wire signed [9:0] m283_113;
   assign m283_113 =10'b0;

   // m283_114 = W*in
   wire signed [9:0] m283_114;
   assign m283_114 =10'b0;

   // m283_115 = W*in
   wire signed [9:0] m283_115;
   assign m283_115 =10'b0;

   // m283_116 = W*in
   wire signed [9:0] m283_116;
   assign m283_116 =10'b0;

   // m283_117 = W*in
   wire signed [9:0] m283_117;
   assign m283_117 =10'b0;

   // m284_1 = W*in
   wire signed [9:0] m284_1;
   assign m284_1 =10'b0;

   // m284_2 = W*in
   wire signed [9:0] m284_2;
   assign m284_2 =10'b0;

   // m284_3 = W*in
   wire signed [9:0] m284_3;
   assign m284_3 =10'b0;

   // m284_4 = W*in
   wire signed [9:0] m284_4;
   assign m284_4 =10'b0;

   // m284_5 = W*in
   wire signed [9:0] m284_5;
   assign m284_5 =10'b0;

   // m284_6 = W*in
   wire signed [9:0] m284_6;
   assign m284_6 =10'b0;

   // m284_7 = W*in
   wire signed [9:0] m284_7;
   assign m284_7 =10'b0;

   // m284_8 = W*in
   wire signed [9:0] m284_8;
   assign m284_8 =10'b0;

   // m284_9 = W*in
   wire signed [9:0] m284_9;
   assign m284_9 =10'b0;

   // m284_10 = W*in
   wire signed [9:0] m284_10;
   assign m284_10 =10'b0;

   // m284_11 = W*in
   wire signed [9:0] m284_11;
   assign m284_11 =10'b0;

   // m284_12 = W*in
   wire signed [9:0] m284_12;
   assign m284_12 =10'b0;

   // m284_13 = W*in
   wire signed [9:0] m284_13;
   assign m284_13 =10'b0;

   // m284_14 = W*in
   wire signed [9:0] m284_14;
   assign m284_14 =10'b0;

   // m284_15 = W*in
   wire signed [9:0] m284_15;
   assign m284_15 =10'b0;

   // m284_16 = W*in
   wire signed [9:0] m284_16;
   assign m284_16 =10'b0;

   // m284_17 = W*in
   wire signed [9:0] m284_17;
   assign m284_17 =10'b0;

   // m284_18 = W*in
   wire signed [9:0] m284_18;
   assign m284_18 =10'b0;

   // m284_19 = W*in
   wire signed [9:0] m284_19;
   assign m284_19 ={ {5{in284[5]}} , in284[5:1] };

   // m284_20 = W*in
   wire signed [9:0] m284_20;
   assign m284_20 =10'b0;

   // m284_21 = W*in
   wire signed [9:0] m284_21;
   assign m284_21 =10'b0;

   // m284_22 = W*in
   wire signed [9:0] m284_22;
   assign m284_22 =10'b0;

   // m284_23 = W*in
   wire signed [9:0] m284_23;
   assign m284_23 =10'b0;

   // m284_24 = W*in
   wire signed [9:0] m284_24;
   assign m284_24 =10'b0;

   // m284_25 = W*in
   wire signed [9:0] m284_25;
   assign m284_25 =10'b0;

   // m284_26 = W*in
   wire signed [9:0] m284_26;
   assign m284_26 =10'b0;

   // m284_27 = W*in
   wire signed [9:0] m284_27;
   assign m284_27 =10'b0;

   // m284_28 = W*in
   wire signed [9:0] m284_28;
   assign m284_28 =10'b0;

   // m284_29 = W*in
   wire signed [9:0] m284_29;
   assign m284_29 =10'b0;

   // m284_30 = W*in
   wire signed [9:0] m284_30;
   assign m284_30 =10'b0;

   // m284_31 = W*in
   wire signed [9:0] m284_31;
   assign m284_31 =10'b0;

   // m284_32 = W*in
   wire signed [9:0] m284_32;
   assign m284_32 =10'b0;

   // m284_33 = W*in
   wire signed [9:0] m284_33;
   assign m284_33 =10'b0;

   // m284_34 = W*in
   wire signed [9:0] m284_34;
   assign m284_34 =10'b0;

   // m284_35 = W*in
   wire signed [9:0] m284_35;
   assign m284_35 =10'b0;

   // m284_36 = W*in
   wire signed [9:0] m284_36;
   assign m284_36 =10'b0;

   // m284_37 = W*in
   wire signed [9:0] m284_37;
   assign m284_37 =10'b0;

   // m284_38 = W*in
   wire signed [9:0] m284_38;
   assign m284_38 =10'b0;

   // m284_39 = W*in
   wire signed [9:0] m284_39;
   assign m284_39 =10'b0;

   // m284_40 = W*in
   wire signed [9:0] m284_40;
   assign m284_40 =10'b0;

   // m284_41 = W*in
   wire signed [9:0] m284_41;
   assign m284_41 =10'b0;

   // m284_42 = W*in
   wire signed [9:0] m284_42;
   assign m284_42 =10'b0;

   // m284_43 = W*in
   wire signed [9:0] m284_43;
   assign m284_43 =10'b0;

   // m284_44 = W*in
   wire signed [9:0] m284_44;
   assign m284_44 =10'b0;

   // m284_45 = W*in
   wire signed [9:0] m284_45;
   assign m284_45 =10'b0;

   // m284_46 = W*in
   wire signed [9:0] m284_46;
   assign m284_46 =10'b0;

   // m284_47 = W*in
   wire signed [9:0] m284_47;
   assign m284_47 =10'b0;

   // m284_48 = W*in
   wire signed [9:0] m284_48;
   assign m284_48 =10'b0;

   // m284_49 = W*in
   wire signed [9:0] m284_49;
   assign m284_49 =10'b0;

   // m284_50 = W*in
   wire signed [9:0] m284_50;
   assign m284_50 =10'b0;

   // m284_51 = W*in
   wire signed [9:0] m284_51;
   assign m284_51 =10'b0;

   // m284_52 = W*in
   wire signed [9:0] m284_52;
   assign m284_52 =10'b0;

   // m284_53 = W*in
   wire signed [9:0] m284_53;
   assign m284_53 =10'b0;

   // m284_54 = W*in
   wire signed [9:0] m284_54;
   assign m284_54 =10'b0;

   // m284_55 = W*in
   wire signed [9:0] m284_55;
   assign m284_55 =10'b0;

   // m284_56 = W*in
   wire signed [9:0] m284_56;
   assign m284_56 =10'b0;

   // m284_57 = W*in
   wire signed [9:0] m284_57;
   assign m284_57 =10'b0;

   // m284_58 = W*in
   wire signed [9:0] m284_58;
   assign m284_58 =10'b0;

   // m284_59 = W*in
   wire signed [9:0] m284_59;
   assign m284_59 =10'b0;

   // m284_60 = W*in
   wire signed [9:0] m284_60;
   assign m284_60 =10'b0;

   // m284_61 = W*in
   wire signed [9:0] m284_61;
   assign m284_61 =10'b0;

   // m284_62 = W*in
   wire signed [9:0] m284_62;
   assign m284_62 =10'b0;

   // m284_63 = W*in
   wire signed [9:0] m284_63;
   assign m284_63 =10'b0;

   // m284_64 = W*in
   wire signed [9:0] m284_64;
   assign m284_64 =10'b0;

   // m284_65 = W*in
   wire signed [9:0] m284_65;
   assign m284_65 =10'b0;

   // m284_66 = W*in
   wire signed [9:0] m284_66;
   assign m284_66 =10'b0;

   // m284_67 = W*in
   wire signed [9:0] m284_67;
   assign m284_67 =10'b0;

   // m284_68 = W*in
   wire signed [9:0] m284_68;
   assign m284_68 =10'b0;

   // m284_69 = W*in
   wire signed [9:0] m284_69;
   assign m284_69 =10'b0;

   // m284_70 = W*in
   wire signed [9:0] m284_70;
   assign m284_70 =10'b0;

   // m284_71 = W*in
   wire signed [9:0] m284_71;
   assign m284_71 =10'b0;

   // m284_72 = W*in
   wire signed [9:0] m284_72;
   assign m284_72 =10'b0;

   // m284_73 = W*in
   wire signed [9:0] m284_73;
   assign m284_73 =10'b0;

   // m284_74 = W*in
   wire signed [9:0] m284_74;
   assign m284_74 =10'b0;

   // m284_75 = W*in
   wire signed [9:0] m284_75;
   assign m284_75 =10'b0;

   // m284_76 = W*in
   wire signed [9:0] m284_76;
   assign m284_76 =10'b0;

   // m284_77 = W*in
   wire signed [9:0] m284_77;
   assign m284_77 =10'b0;

   // m284_78 = W*in
   wire signed [9:0] m284_78;
   assign m284_78 =10'b0;

   // m284_79 = W*in
   wire signed [9:0] m284_79;
   assign m284_79 =10'b0;

   // m284_80 = W*in
   wire signed [9:0] m284_80;
   assign m284_80 =10'b0;

   // m284_81 = W*in
   wire signed [9:0] m284_81;
   assign m284_81 =10'b0;

   // m284_82 = W*in
   wire signed [9:0] m284_82;
   assign m284_82 =10'b0;

   // m284_83 = W*in
   wire signed [9:0] m284_83;
   assign m284_83 =10'b0;

   // m284_84 = W*in
   wire signed [9:0] m284_84;
   assign m284_84 =10'b0;

   // m284_85 = W*in
   wire signed [9:0] m284_85;
   assign m284_85 =10'b0;

   // m284_86 = W*in
   wire signed [9:0] m284_86;
   assign m284_86 =10'b0;

   // m284_87 = W*in
   wire signed [9:0] m284_87;
   assign m284_87 =10'b0;

   // m284_88 = W*in
   wire signed [9:0] m284_88;
   assign m284_88 =10'b0;

   // m284_89 = W*in
   wire signed [9:0] m284_89;
   assign m284_89 =10'b0;

   // m284_90 = W*in
   wire signed [9:0] m284_90;
   assign m284_90 =10'b0;

   // m284_91 = W*in
   wire signed [9:0] m284_91;
   assign m284_91 =10'b0;

   // m284_92 = W*in
   wire signed [9:0] m284_92;
   assign m284_92 =10'b0;

   // m284_93 = W*in
   wire signed [9:0] m284_93;
   assign m284_93 =10'b0;

   // m284_94 = W*in
   wire signed [9:0] m284_94;
   assign m284_94 =10'b0;

   // m284_95 = W*in
   wire signed [9:0] m284_95;
   assign m284_95 =10'b0;

   // m284_96 = W*in
   wire signed [9:0] m284_96;
   assign m284_96 =10'b0;

   // m284_97 = W*in
   wire signed [9:0] m284_97;
   assign m284_97 =10'b0;

   // m284_98 = W*in
   wire signed [9:0] m284_98;
   assign m284_98 =10'b0;

   // m284_99 = W*in
   wire signed [9:0] m284_99;
   assign m284_99 =10'b0;

   // m284_100 = W*in
   wire signed [9:0] m284_100;
   assign m284_100 =10'b0;

   // m284_101 = W*in
   wire signed [9:0] m284_101;
   assign m284_101 =10'b0;

   // m284_102 = W*in
   wire signed [9:0] m284_102;
   assign m284_102 =10'b0;

   // m284_103 = W*in
   wire signed [9:0] m284_103;
   assign m284_103 =10'b0;

   // m284_104 = W*in
   wire signed [9:0] m284_104;
   assign m284_104 =10'b0;

   // m284_105 = W*in
   wire signed [9:0] m284_105;
   assign m284_105 =10'b0;

   // m284_106 = W*in
   wire signed [9:0] m284_106;
   assign m284_106 =10'b0;

   // m284_107 = W*in
   wire signed [9:0] m284_107;
   assign m284_107 =10'b0;

   // m284_108 = W*in
   wire signed [9:0] m284_108;
   assign m284_108 =10'b0;

   // m284_109 = W*in
   wire signed [9:0] m284_109;
   assign m284_109 =10'b0;

   // m284_110 = W*in
   wire signed [9:0] m284_110;
   assign m284_110 =10'b0;

   // m284_111 = W*in
   wire signed [9:0] m284_111;
   assign m284_111 =10'b0;

   // m284_112 = W*in
   wire signed [9:0] m284_112;
   assign m284_112 =10'b0;

   // m284_113 = W*in
   wire signed [9:0] m284_113;
   assign m284_113 =10'b0;

   // m284_114 = W*in
   wire signed [9:0] m284_114;
   assign m284_114 =10'b0;

   // m284_115 = W*in
   wire signed [9:0] m284_115;
   assign m284_115 =10'b0;

   // m284_116 = W*in
   wire signed [9:0] m284_116;
   assign m284_116 =10'b0;

   // m284_117 = W*in
   wire signed [9:0] m284_117;
   assign m284_117 =10'b0;

   // m285_1 = W*in
   wire signed [9:0] m285_1;
   assign m285_1 =10'b0;

   // m285_2 = W*in
   wire signed [9:0] m285_2;
   assign m285_2 =10'b0;

   // m285_3 = W*in
   wire signed [9:0] m285_3;
   assign m285_3 =10'b0;

   // m285_4 = W*in
   wire signed [9:0] m285_4;
   assign m285_4 =10'b0;

   // m285_5 = W*in
   wire signed [9:0] m285_5;
   assign m285_5 =10'b0;

   // m285_6 = W*in
   wire signed [9:0] m285_6;
   assign m285_6 =10'b0;

   // m285_7 = W*in
   wire signed [9:0] m285_7;
   assign m285_7 =10'b0;

   // m285_8 = W*in
   wire signed [9:0] m285_8;
   assign m285_8 =10'b0;

   // m285_9 = W*in
   wire signed [9:0] m285_9;
   assign m285_9 =10'b0;

   // m285_10 = W*in
   wire signed [9:0] m285_10;
   assign m285_10 =10'b0;

   // m285_11 = W*in
   wire signed [9:0] m285_11;
   assign m285_11 =10'b0;

   // m285_12 = W*in
   wire signed [9:0] m285_12;
   assign m285_12 =10'b0;

   // m285_13 = W*in
   wire signed [9:0] m285_13;
   assign m285_13 =10'b0;

   // m285_14 = W*in
   wire signed [9:0] m285_14;
   assign m285_14 =10'b0;

   // m285_15 = W*in
   wire signed [9:0] m285_15;
   assign m285_15 =10'b0;

   // m285_16 = W*in
   wire signed [9:0] m285_16;
   assign m285_16 =10'b0;

   // m285_17 = W*in
   wire signed [9:0] m285_17;
   assign m285_17 ={ {5{in285[5]}} , in285[5:1] };

   // m285_18 = W*in
   wire signed [9:0] m285_18;
   assign m285_18 =10'b0;

   // m285_19 = W*in
   wire signed [9:0] m285_19;
   assign m285_19 ={ {5{in285[5]}} , in285[5:1] };

   // m285_20 = W*in
   wire signed [9:0] m285_20;
   assign m285_20 =10'b0;

   // m285_21 = W*in
   wire signed [9:0] m285_21;
   assign m285_21 =10'b0;

   // m285_22 = W*in
   wire signed [9:0] m285_22;
   assign m285_22 =10'b0;

   // m285_23 = W*in
   wire signed [9:0] m285_23;
   assign m285_23 =10'b0;

   // m285_24 = W*in
   wire signed [9:0] m285_24;
   assign m285_24 =10'b0;

   // m285_25 = W*in
   wire signed [9:0] m285_25;
   assign m285_25 =10'b0;

   // m285_26 = W*in
   wire signed [9:0] m285_26;
   assign m285_26 =10'b0;

   // m285_27 = W*in
   wire signed [9:0] m285_27;
   assign m285_27 =10'b0;

   // m285_28 = W*in
   wire signed [9:0] m285_28;
   assign m285_28 =10'b0;

   // m285_29 = W*in
   wire signed [9:0] m285_29;
   assign m285_29 =10'b0;

   // m285_30 = W*in
   wire signed [9:0] m285_30;
   assign m285_30 =10'b0;

   // m285_31 = W*in
   wire signed [9:0] m285_31;
   assign m285_31 =10'b0;

   // m285_32 = W*in
   wire signed [9:0] m285_32;
   assign m285_32 =10'b0;

   // m285_33 = W*in
   wire signed [9:0] m285_33;
   assign m285_33 =10'b0;

   // m285_34 = W*in
   wire signed [9:0] m285_34;
   assign m285_34 =10'b0;

   // m285_35 = W*in
   wire signed [9:0] m285_35;
   assign m285_35 =10'b0;

   // m285_36 = W*in
   wire signed [9:0] m285_36;
   assign m285_36 =10'b0;

   // m285_37 = W*in
   wire signed [9:0] m285_37;
   assign m285_37 =10'b0;

   // m285_38 = W*in
   wire signed [9:0] m285_38;
   assign m285_38 =10'b0;

   // m285_39 = W*in
   wire signed [9:0] m285_39;
   assign m285_39 =10'b0;

   // m285_40 = W*in
   wire signed [9:0] m285_40;
   assign m285_40 =10'b0;

   // m285_41 = W*in
   wire signed [9:0] m285_41;
   assign m285_41 =10'b0;

   // m285_42 = W*in
   wire signed [9:0] m285_42;
   assign m285_42 =10'b0;

   // m285_43 = W*in
   wire signed [9:0] m285_43;
   assign m285_43 =10'b0;

   // m285_44 = W*in
   wire signed [9:0] m285_44;
   assign m285_44 =10'b0;

   // m285_45 = W*in
   wire signed [9:0] m285_45;
   assign m285_45 =10'b0;

   // m285_46 = W*in
   wire signed [9:0] m285_46;
   assign m285_46 =10'b0;

   // m285_47 = W*in
   wire signed [9:0] m285_47;
   assign m285_47 =10'b0;

   // m285_48 = W*in
   wire signed [9:0] m285_48;
   assign m285_48 =10'b0;

   // m285_49 = W*in
   wire signed [9:0] m285_49;
   assign m285_49 =10'b0;

   // m285_50 = W*in
   wire signed [9:0] m285_50;
   assign m285_50 =10'b0;

   // m285_51 = W*in
   wire signed [9:0] m285_51;
   assign m285_51 =10'b0;

   // m285_52 = W*in
   wire signed [9:0] m285_52;
   assign m285_52 =10'b0;

   // m285_53 = W*in
   wire signed [9:0] m285_53;
   assign m285_53 =10'b0;

   // m285_54 = W*in
   wire signed [9:0] m285_54;
   assign m285_54 ={ {4{in285[5]}} , in285[5:0] };

   // m285_55 = W*in
   wire signed [9:0] m285_55;
   assign m285_55 =10'b0;

   // m285_56 = W*in
   wire signed [9:0] m285_56;
   assign m285_56 =10'b0;

   // m285_57 = W*in
   wire signed [9:0] m285_57;
   assign m285_57 =10'b0;

   // m285_58 = W*in
   wire signed [9:0] m285_58;
   assign m285_58 =10'b0;

   // m285_59 = W*in
   wire signed [9:0] m285_59;
   assign m285_59 =10'b0;

   // m285_60 = W*in
   wire signed [9:0] m285_60;
   assign m285_60 =10'b0;

   // m285_61 = W*in
   wire signed [9:0] m285_61;
   assign m285_61 =10'b0;

   // m285_62 = W*in
   wire signed [9:0] m285_62;
   assign m285_62 =10'b0;

   // m285_63 = W*in
   wire signed [9:0] m285_63;
   assign m285_63 =10'b0;

   // m285_64 = W*in
   wire signed [9:0] m285_64;
   assign m285_64 ={ {5{neg285[5]}} , neg285[5:1] };

   // m285_65 = W*in
   wire signed [9:0] m285_65;
   assign m285_65 =10'b0;

   // m285_66 = W*in
   wire signed [9:0] m285_66;
   assign m285_66 =10'b0;

   // m285_67 = W*in
   wire signed [9:0] m285_67;
   assign m285_67 ={ {5{in285[5]}} , in285[5:1] };

   // m285_68 = W*in
   wire signed [9:0] m285_68;
   assign m285_68 =10'b0;

   // m285_69 = W*in
   wire signed [9:0] m285_69;
   assign m285_69 =10'b0;

   // m285_70 = W*in
   wire signed [9:0] m285_70;
   assign m285_70 =10'b0;

   // m285_71 = W*in
   wire signed [9:0] m285_71;
   assign m285_71 =10'b0;

   // m285_72 = W*in
   wire signed [9:0] m285_72;
   assign m285_72 =10'b0;

   // m285_73 = W*in
   wire signed [9:0] m285_73;
   assign m285_73 =10'b0;

   // m285_74 = W*in
   wire signed [9:0] m285_74;
   assign m285_74 =10'b0;

   // m285_75 = W*in
   wire signed [9:0] m285_75;
   assign m285_75 =10'b0;

   // m285_76 = W*in
   wire signed [9:0] m285_76;
   assign m285_76 =10'b0;

   // m285_77 = W*in
   wire signed [9:0] m285_77;
   assign m285_77 =10'b0;

   // m285_78 = W*in
   wire signed [9:0] m285_78;
   assign m285_78 =10'b0;

   // m285_79 = W*in
   wire signed [9:0] m285_79;
   assign m285_79 =10'b0;

   // m285_80 = W*in
   wire signed [9:0] m285_80;
   assign m285_80 =10'b0;

   // m285_81 = W*in
   wire signed [9:0] m285_81;
   assign m285_81 ={ {5{neg285[5]}} , neg285[5:1] };

   // m285_82 = W*in
   wire signed [9:0] m285_82;
   assign m285_82 =10'b0;

   // m285_83 = W*in
   wire signed [9:0] m285_83;
   assign m285_83 =10'b0;

   // m285_84 = W*in
   wire signed [9:0] m285_84;
   assign m285_84 =10'b0;

   // m285_85 = W*in
   wire signed [9:0] m285_85;
   assign m285_85 =10'b0;

   // m285_86 = W*in
   wire signed [9:0] m285_86;
   assign m285_86 =10'b0;

   // m285_87 = W*in
   wire signed [9:0] m285_87;
   assign m285_87 =10'b0;

   // m285_88 = W*in
   wire signed [9:0] m285_88;
   assign m285_88 =10'b0;

   // m285_89 = W*in
   wire signed [9:0] m285_89;
   assign m285_89 =10'b0;

   // m285_90 = W*in
   wire signed [9:0] m285_90;
   assign m285_90 =10'b0;

   // m285_91 = W*in
   wire signed [9:0] m285_91;
   assign m285_91 =10'b0;

   // m285_92 = W*in
   wire signed [9:0] m285_92;
   assign m285_92 =10'b0;

   // m285_93 = W*in
   wire signed [9:0] m285_93;
   assign m285_93 =10'b0;

   // m285_94 = W*in
   wire signed [9:0] m285_94;
   assign m285_94 =10'b0;

   // m285_95 = W*in
   wire signed [9:0] m285_95;
   assign m285_95 =10'b0;

   // m285_96 = W*in
   wire signed [9:0] m285_96;
   assign m285_96 =10'b0;

   // m285_97 = W*in
   wire signed [9:0] m285_97;
   assign m285_97 =10'b0;

   // m285_98 = W*in
   wire signed [9:0] m285_98;
   assign m285_98 =10'b0;

   // m285_99 = W*in
   wire signed [9:0] m285_99;
   assign m285_99 =10'b0;

   // m285_100 = W*in
   wire signed [9:0] m285_100;
   assign m285_100 =10'b0;

   // m285_101 = W*in
   wire signed [9:0] m285_101;
   assign m285_101 =10'b0;

   // m285_102 = W*in
   wire signed [9:0] m285_102;
   assign m285_102 =10'b0;

   // m285_103 = W*in
   wire signed [9:0] m285_103;
   assign m285_103 =10'b0;

   // m285_104 = W*in
   wire signed [9:0] m285_104;
   assign m285_104 =10'b0;

   // m285_105 = W*in
   wire signed [9:0] m285_105;
   assign m285_105 =10'b0;

   // m285_106 = W*in
   wire signed [9:0] m285_106;
   assign m285_106 =10'b0;

   // m285_107 = W*in
   wire signed [9:0] m285_107;
   assign m285_107 =10'b0;

   // m285_108 = W*in
   wire signed [9:0] m285_108;
   assign m285_108 ={ {5{neg285[5]}} , neg285[5:1] };

   // m285_109 = W*in
   wire signed [9:0] m285_109;
   assign m285_109 ={ {5{neg285[5]}} , neg285[5:1] };

   // m285_110 = W*in
   wire signed [9:0] m285_110;
   assign m285_110 =10'b0;

   // m285_111 = W*in
   wire signed [9:0] m285_111;
   assign m285_111 =10'b0;

   // m285_112 = W*in
   wire signed [9:0] m285_112;
   assign m285_112 =10'b0;

   // m285_113 = W*in
   wire signed [9:0] m285_113;
   assign m285_113 =10'b0;

   // m285_114 = W*in
   wire signed [9:0] m285_114;
   assign m285_114 =10'b0;

   // m285_115 = W*in
   wire signed [9:0] m285_115;
   assign m285_115 =10'b0;

   // m285_116 = W*in
   wire signed [9:0] m285_116;
   assign m285_116 =10'b0;

   // m285_117 = W*in
   wire signed [9:0] m285_117;
   assign m285_117 =10'b0;

   // m286_1 = W*in
   wire signed [9:0] m286_1;
   assign m286_1 =10'b0;

   // m286_2 = W*in
   wire signed [9:0] m286_2;
   assign m286_2 =10'b0;

   // m286_3 = W*in
   wire signed [9:0] m286_3;
   assign m286_3 =10'b0;

   // m286_4 = W*in
   wire signed [9:0] m286_4;
   assign m286_4 =10'b0;

   // m286_5 = W*in
   wire signed [9:0] m286_5;
   assign m286_5 =10'b0;

   // m286_6 = W*in
   wire signed [9:0] m286_6;
   assign m286_6 =10'b0;

   // m286_7 = W*in
   wire signed [9:0] m286_7;
   assign m286_7 =10'b0;

   // m286_8 = W*in
   wire signed [9:0] m286_8;
   assign m286_8 =10'b0;

   // m286_9 = W*in
   wire signed [9:0] m286_9;
   assign m286_9 =10'b0;

   // m286_10 = W*in
   wire signed [9:0] m286_10;
   assign m286_10 =10'b0;

   // m286_11 = W*in
   wire signed [9:0] m286_11;
   assign m286_11 =10'b0;

   // m286_12 = W*in
   wire signed [9:0] m286_12;
   assign m286_12 =10'b0;

   // m286_13 = W*in
   wire signed [9:0] m286_13;
   assign m286_13 =10'b0;

   // m286_14 = W*in
   wire signed [9:0] m286_14;
   assign m286_14 =10'b0;

   // m286_15 = W*in
   wire signed [9:0] m286_15;
   assign m286_15 =10'b0;

   // m286_16 = W*in
   wire signed [9:0] m286_16;
   assign m286_16 =10'b0;

   // m286_17 = W*in
   wire signed [9:0] m286_17;
   assign m286_17 =10'b0;

   // m286_18 = W*in
   wire signed [9:0] m286_18;
   assign m286_18 =10'b0;

   // m286_19 = W*in
   wire signed [9:0] m286_19;
   assign m286_19 =10'b0;

   // m286_20 = W*in
   wire signed [9:0] m286_20;
   assign m286_20 ={ {5{neg286[5]}} , neg286[5:1] };

   // m286_21 = W*in
   wire signed [9:0] m286_21;
   assign m286_21 =10'b0;

   // m286_22 = W*in
   wire signed [9:0] m286_22;
   assign m286_22 =10'b0;

   // m286_23 = W*in
   wire signed [9:0] m286_23;
   assign m286_23 =10'b0;

   // m286_24 = W*in
   wire signed [9:0] m286_24;
   assign m286_24 =10'b0;

   // m286_25 = W*in
   wire signed [9:0] m286_25;
   assign m286_25 =10'b0;

   // m286_26 = W*in
   wire signed [9:0] m286_26;
   assign m286_26 =10'b0;

   // m286_27 = W*in
   wire signed [9:0] m286_27;
   assign m286_27 ={ {5{in286[5]}} , in286[5:1] };

   // m286_28 = W*in
   wire signed [9:0] m286_28;
   assign m286_28 =10'b0;

   // m286_29 = W*in
   wire signed [9:0] m286_29;
   assign m286_29 =10'b0;

   // m286_30 = W*in
   wire signed [9:0] m286_30;
   assign m286_30 =10'b0;

   // m286_31 = W*in
   wire signed [9:0] m286_31;
   assign m286_31 =10'b0;

   // m286_32 = W*in
   wire signed [9:0] m286_32;
   assign m286_32 =10'b0;

   // m286_33 = W*in
   wire signed [9:0] m286_33;
   assign m286_33 =10'b0;

   // m286_34 = W*in
   wire signed [9:0] m286_34;
   assign m286_34 =10'b0;

   // m286_35 = W*in
   wire signed [9:0] m286_35;
   assign m286_35 =10'b0;

   // m286_36 = W*in
   wire signed [9:0] m286_36;
   assign m286_36 =10'b0;

   // m286_37 = W*in
   wire signed [9:0] m286_37;
   assign m286_37 =10'b0;

   // m286_38 = W*in
   wire signed [9:0] m286_38;
   assign m286_38 =10'b0;

   // m286_39 = W*in
   wire signed [9:0] m286_39;
   assign m286_39 =10'b0;

   // m286_40 = W*in
   wire signed [9:0] m286_40;
   assign m286_40 =10'b0;

   // m286_41 = W*in
   wire signed [9:0] m286_41;
   assign m286_41 =10'b0;

   // m286_42 = W*in
   wire signed [9:0] m286_42;
   assign m286_42 =10'b0;

   // m286_43 = W*in
   wire signed [9:0] m286_43;
   assign m286_43 =10'b0;

   // m286_44 = W*in
   wire signed [9:0] m286_44;
   assign m286_44 =10'b0;

   // m286_45 = W*in
   wire signed [9:0] m286_45;
   assign m286_45 =10'b0;

   // m286_46 = W*in
   wire signed [9:0] m286_46;
   assign m286_46 =10'b0;

   // m286_47 = W*in
   wire signed [9:0] m286_47;
   assign m286_47 =10'b0;

   // m286_48 = W*in
   wire signed [9:0] m286_48;
   assign m286_48 =10'b0;

   // m286_49 = W*in
   wire signed [9:0] m286_49;
   assign m286_49 =10'b0;

   // m286_50 = W*in
   wire signed [9:0] m286_50;
   assign m286_50 =10'b0;

   // m286_51 = W*in
   wire signed [9:0] m286_51;
   assign m286_51 =10'b0;

   // m286_52 = W*in
   wire signed [9:0] m286_52;
   assign m286_52 =10'b0;

   // m286_53 = W*in
   wire signed [9:0] m286_53;
   assign m286_53 =10'b0;

   // m286_54 = W*in
   wire signed [9:0] m286_54;
   assign m286_54 =10'b0;

   // m286_55 = W*in
   wire signed [9:0] m286_55;
   assign m286_55 =10'b0;

   // m286_56 = W*in
   wire signed [9:0] m286_56;
   assign m286_56 =10'b0;

   // m286_57 = W*in
   wire signed [9:0] m286_57;
   assign m286_57 =10'b0;

   // m286_58 = W*in
   wire signed [9:0] m286_58;
   assign m286_58 =10'b0;

   // m286_59 = W*in
   wire signed [9:0] m286_59;
   assign m286_59 =10'b0;

   // m286_60 = W*in
   wire signed [9:0] m286_60;
   assign m286_60 =10'b0;

   // m286_61 = W*in
   wire signed [9:0] m286_61;
   assign m286_61 =10'b0;

   // m286_62 = W*in
   wire signed [9:0] m286_62;
   assign m286_62 =10'b0;

   // m286_63 = W*in
   wire signed [9:0] m286_63;
   assign m286_63 =10'b0;

   // m286_64 = W*in
   wire signed [9:0] m286_64;
   assign m286_64 ={ {5{neg286[5]}} , neg286[5:1] };

   // m286_65 = W*in
   wire signed [9:0] m286_65;
   assign m286_65 =10'b0;

   // m286_66 = W*in
   wire signed [9:0] m286_66;
   assign m286_66 =10'b0;

   // m286_67 = W*in
   wire signed [9:0] m286_67;
   assign m286_67 =10'b0;

   // m286_68 = W*in
   wire signed [9:0] m286_68;
   assign m286_68 =10'b0;

   // m286_69 = W*in
   wire signed [9:0] m286_69;
   assign m286_69 =10'b0;

   // m286_70 = W*in
   wire signed [9:0] m286_70;
   assign m286_70 =10'b0;

   // m286_71 = W*in
   wire signed [9:0] m286_71;
   assign m286_71 =10'b0;

   // m286_72 = W*in
   wire signed [9:0] m286_72;
   assign m286_72 =10'b0;

   // m286_73 = W*in
   wire signed [9:0] m286_73;
   assign m286_73 =10'b0;

   // m286_74 = W*in
   wire signed [9:0] m286_74;
   assign m286_74 =10'b0;

   // m286_75 = W*in
   wire signed [9:0] m286_75;
   assign m286_75 =10'b0;

   // m286_76 = W*in
   wire signed [9:0] m286_76;
   assign m286_76 =10'b0;

   // m286_77 = W*in
   wire signed [9:0] m286_77;
   assign m286_77 =10'b0;

   // m286_78 = W*in
   wire signed [9:0] m286_78;
   assign m286_78 =10'b0;

   // m286_79 = W*in
   wire signed [9:0] m286_79;
   assign m286_79 =10'b0;

   // m286_80 = W*in
   wire signed [9:0] m286_80;
   assign m286_80 =10'b0;

   // m286_81 = W*in
   wire signed [9:0] m286_81;
   assign m286_81 ={ {5{neg286[5]}} , neg286[5:1] };

   // m286_82 = W*in
   wire signed [9:0] m286_82;
   assign m286_82 =10'b0;

   // m286_83 = W*in
   wire signed [9:0] m286_83;
   assign m286_83 =10'b0;

   // m286_84 = W*in
   wire signed [9:0] m286_84;
   assign m286_84 =10'b0;

   // m286_85 = W*in
   wire signed [9:0] m286_85;
   assign m286_85 =10'b0;

   // m286_86 = W*in
   wire signed [9:0] m286_86;
   assign m286_86 =10'b0;

   // m286_87 = W*in
   wire signed [9:0] m286_87;
   assign m286_87 =10'b0;

   // m286_88 = W*in
   wire signed [9:0] m286_88;
   assign m286_88 =10'b0;

   // m286_89 = W*in
   wire signed [9:0] m286_89;
   assign m286_89 =10'b0;

   // m286_90 = W*in
   wire signed [9:0] m286_90;
   assign m286_90 =10'b0;

   // m286_91 = W*in
   wire signed [9:0] m286_91;
   assign m286_91 =10'b0;

   // m286_92 = W*in
   wire signed [9:0] m286_92;
   assign m286_92 =10'b0;

   // m286_93 = W*in
   wire signed [9:0] m286_93;
   assign m286_93 =10'b0;

   // m286_94 = W*in
   wire signed [9:0] m286_94;
   assign m286_94 =10'b0;

   // m286_95 = W*in
   wire signed [9:0] m286_95;
   assign m286_95 =10'b0;

   // m286_96 = W*in
   wire signed [9:0] m286_96;
   assign m286_96 =10'b0;

   // m286_97 = W*in
   wire signed [9:0] m286_97;
   assign m286_97 =10'b0;

   // m286_98 = W*in
   wire signed [9:0] m286_98;
   assign m286_98 =10'b0;

   // m286_99 = W*in
   wire signed [9:0] m286_99;
   assign m286_99 =10'b0;

   // m286_100 = W*in
   wire signed [9:0] m286_100;
   assign m286_100 =10'b0;

   // m286_101 = W*in
   wire signed [9:0] m286_101;
   assign m286_101 =10'b0;

   // m286_102 = W*in
   wire signed [9:0] m286_102;
   assign m286_102 =10'b0;

   // m286_103 = W*in
   wire signed [9:0] m286_103;
   assign m286_103 =10'b0;

   // m286_104 = W*in
   wire signed [9:0] m286_104;
   assign m286_104 =10'b0;

   // m286_105 = W*in
   wire signed [9:0] m286_105;
   assign m286_105 =10'b0;

   // m286_106 = W*in
   wire signed [9:0] m286_106;
   assign m286_106 =10'b0;

   // m286_107 = W*in
   wire signed [9:0] m286_107;
   assign m286_107 =10'b0;

   // m286_108 = W*in
   wire signed [9:0] m286_108;
   assign m286_108 ={ {5{neg286[5]}} , neg286[5:1] };

   // m286_109 = W*in
   wire signed [9:0] m286_109;
   assign m286_109 ={ {5{neg286[5]}} , neg286[5:1] };

   // m286_110 = W*in
   wire signed [9:0] m286_110;
   assign m286_110 =10'b0;

   // m286_111 = W*in
   wire signed [9:0] m286_111;
   assign m286_111 =10'b0;

   // m286_112 = W*in
   wire signed [9:0] m286_112;
   assign m286_112 =10'b0;

   // m286_113 = W*in
   wire signed [9:0] m286_113;
   assign m286_113 =10'b0;

   // m286_114 = W*in
   wire signed [9:0] m286_114;
   assign m286_114 =10'b0;

   // m286_115 = W*in
   wire signed [9:0] m286_115;
   assign m286_115 =10'b0;

   // m286_116 = W*in
   wire signed [9:0] m286_116;
   assign m286_116 =10'b0;

   // m286_117 = W*in
   wire signed [9:0] m286_117;
   assign m286_117 =10'b0;

   // m287_1 = W*in
   wire signed [9:0] m287_1;
   assign m287_1 =10'b0;

   // m287_2 = W*in
   wire signed [9:0] m287_2;
   assign m287_2 =10'b0;

   // m287_3 = W*in
   wire signed [9:0] m287_3;
   assign m287_3 =10'b0;

   // m287_4 = W*in
   wire signed [9:0] m287_4;
   assign m287_4 =10'b0;

   // m287_5 = W*in
   wire signed [9:0] m287_5;
   assign m287_5 =10'b0;

   // m287_6 = W*in
   wire signed [9:0] m287_6;
   assign m287_6 =10'b0;

   // m287_7 = W*in
   wire signed [9:0] m287_7;
   assign m287_7 =10'b0;

   // m287_8 = W*in
   wire signed [9:0] m287_8;
   assign m287_8 =10'b0;

   // m287_9 = W*in
   wire signed [9:0] m287_9;
   assign m287_9 =10'b0;

   // m287_10 = W*in
   wire signed [9:0] m287_10;
   assign m287_10 =10'b0;

   // m287_11 = W*in
   wire signed [9:0] m287_11;
   assign m287_11 =10'b0;

   // m287_12 = W*in
   wire signed [9:0] m287_12;
   assign m287_12 =10'b0;

   // m287_13 = W*in
   wire signed [9:0] m287_13;
   assign m287_13 =10'b0;

   // m287_14 = W*in
   wire signed [9:0] m287_14;
   assign m287_14 =10'b0;

   // m287_15 = W*in
   wire signed [9:0] m287_15;
   assign m287_15 =10'b0;

   // m287_16 = W*in
   wire signed [9:0] m287_16;
   assign m287_16 =10'b0;

   // m287_17 = W*in
   wire signed [9:0] m287_17;
   assign m287_17 =10'b0;

   // m287_18 = W*in
   wire signed [9:0] m287_18;
   assign m287_18 =10'b0;

   // m287_19 = W*in
   wire signed [9:0] m287_19;
   assign m287_19 =10'b0;

   // m287_20 = W*in
   wire signed [9:0] m287_20;
   assign m287_20 ={ {5{neg287[5]}} , neg287[5:1] };

   // m287_21 = W*in
   wire signed [9:0] m287_21;
   assign m287_21 =10'b0;

   // m287_22 = W*in
   wire signed [9:0] m287_22;
   assign m287_22 =10'b0;

   // m287_23 = W*in
   wire signed [9:0] m287_23;
   assign m287_23 =10'b0;

   // m287_24 = W*in
   wire signed [9:0] m287_24;
   assign m287_24 =10'b0;

   // m287_25 = W*in
   wire signed [9:0] m287_25;
   assign m287_25 =10'b0;

   // m287_26 = W*in
   wire signed [9:0] m287_26;
   assign m287_26 =10'b0;

   // m287_27 = W*in
   wire signed [9:0] m287_27;
   assign m287_27 =10'b0;

   // m287_28 = W*in
   wire signed [9:0] m287_28;
   assign m287_28 =10'b0;

   // m287_29 = W*in
   wire signed [9:0] m287_29;
   assign m287_29 =10'b0;

   // m287_30 = W*in
   wire signed [9:0] m287_30;
   assign m287_30 =10'b0;

   // m287_31 = W*in
   wire signed [9:0] m287_31;
   assign m287_31 =10'b0;

   // m287_32 = W*in
   wire signed [9:0] m287_32;
   assign m287_32 =10'b0;

   // m287_33 = W*in
   wire signed [9:0] m287_33;
   assign m287_33 =10'b0;

   // m287_34 = W*in
   wire signed [9:0] m287_34;
   assign m287_34 =10'b0;

   // m287_35 = W*in
   wire signed [9:0] m287_35;
   assign m287_35 ={ {5{neg287[5]}} , neg287[5:1] };

   // m287_36 = W*in
   wire signed [9:0] m287_36;
   assign m287_36 =10'b0;

   // m287_37 = W*in
   wire signed [9:0] m287_37;
   assign m287_37 =10'b0;

   // m287_38 = W*in
   wire signed [9:0] m287_38;
   assign m287_38 =10'b0;

   // m287_39 = W*in
   wire signed [9:0] m287_39;
   assign m287_39 =10'b0;

   // m287_40 = W*in
   wire signed [9:0] m287_40;
   assign m287_40 =10'b0;

   // m287_41 = W*in
   wire signed [9:0] m287_41;
   assign m287_41 =10'b0;

   // m287_42 = W*in
   wire signed [9:0] m287_42;
   assign m287_42 =10'b0;

   // m287_43 = W*in
   wire signed [9:0] m287_43;
   assign m287_43 =10'b0;

   // m287_44 = W*in
   wire signed [9:0] m287_44;
   assign m287_44 =10'b0;

   // m287_45 = W*in
   wire signed [9:0] m287_45;
   assign m287_45 =10'b0;

   // m287_46 = W*in
   wire signed [9:0] m287_46;
   assign m287_46 =10'b0;

   // m287_47 = W*in
   wire signed [9:0] m287_47;
   assign m287_47 =10'b0;

   // m287_48 = W*in
   wire signed [9:0] m287_48;
   assign m287_48 =10'b0;

   // m287_49 = W*in
   wire signed [9:0] m287_49;
   assign m287_49 =10'b0;

   // m287_50 = W*in
   wire signed [9:0] m287_50;
   assign m287_50 =10'b0;

   // m287_51 = W*in
   wire signed [9:0] m287_51;
   assign m287_51 =10'b0;

   // m287_52 = W*in
   wire signed [9:0] m287_52;
   assign m287_52 =10'b0;

   // m287_53 = W*in
   wire signed [9:0] m287_53;
   assign m287_53 =10'b0;

   // m287_54 = W*in
   wire signed [9:0] m287_54;
   assign m287_54 =10'b0;

   // m287_55 = W*in
   wire signed [9:0] m287_55;
   assign m287_55 =10'b0;

   // m287_56 = W*in
   wire signed [9:0] m287_56;
   assign m287_56 =10'b0;

   // m287_57 = W*in
   wire signed [9:0] m287_57;
   assign m287_57 =10'b0;

   // m287_58 = W*in
   wire signed [9:0] m287_58;
   assign m287_58 =10'b0;

   // m287_59 = W*in
   wire signed [9:0] m287_59;
   assign m287_59 =10'b0;

   // m287_60 = W*in
   wire signed [9:0] m287_60;
   assign m287_60 =10'b0;

   // m287_61 = W*in
   wire signed [9:0] m287_61;
   assign m287_61 =10'b0;

   // m287_62 = W*in
   wire signed [9:0] m287_62;
   assign m287_62 =10'b0;

   // m287_63 = W*in
   wire signed [9:0] m287_63;
   assign m287_63 =10'b0;

   // m287_64 = W*in
   wire signed [9:0] m287_64;
   assign m287_64 =10'b0;

   // m287_65 = W*in
   wire signed [9:0] m287_65;
   assign m287_65 =10'b0;

   // m287_66 = W*in
   wire signed [9:0] m287_66;
   assign m287_66 =10'b0;

   // m287_67 = W*in
   wire signed [9:0] m287_67;
   assign m287_67 =10'b0;

   // m287_68 = W*in
   wire signed [9:0] m287_68;
   assign m287_68 =10'b0;

   // m287_69 = W*in
   wire signed [9:0] m287_69;
   assign m287_69 =10'b0;

   // m287_70 = W*in
   wire signed [9:0] m287_70;
   assign m287_70 =10'b0;

   // m287_71 = W*in
   wire signed [9:0] m287_71;
   assign m287_71 =10'b0;

   // m287_72 = W*in
   wire signed [9:0] m287_72;
   assign m287_72 =10'b0;

   // m287_73 = W*in
   wire signed [9:0] m287_73;
   assign m287_73 =10'b0;

   // m287_74 = W*in
   wire signed [9:0] m287_74;
   assign m287_74 =10'b0;

   // m287_75 = W*in
   wire signed [9:0] m287_75;
   assign m287_75 =10'b0;

   // m287_76 = W*in
   wire signed [9:0] m287_76;
   assign m287_76 =10'b0;

   // m287_77 = W*in
   wire signed [9:0] m287_77;
   assign m287_77 =10'b0;

   // m287_78 = W*in
   wire signed [9:0] m287_78;
   assign m287_78 =10'b0;

   // m287_79 = W*in
   wire signed [9:0] m287_79;
   assign m287_79 =10'b0;

   // m287_80 = W*in
   wire signed [9:0] m287_80;
   assign m287_80 =10'b0;

   // m287_81 = W*in
   wire signed [9:0] m287_81;
   assign m287_81 =10'b0;

   // m287_82 = W*in
   wire signed [9:0] m287_82;
   assign m287_82 =10'b0;

   // m287_83 = W*in
   wire signed [9:0] m287_83;
   assign m287_83 =10'b0;

   // m287_84 = W*in
   wire signed [9:0] m287_84;
   assign m287_84 =10'b0;

   // m287_85 = W*in
   wire signed [9:0] m287_85;
   assign m287_85 =10'b0;

   // m287_86 = W*in
   wire signed [9:0] m287_86;
   assign m287_86 =10'b0;

   // m287_87 = W*in
   wire signed [9:0] m287_87;
   assign m287_87 =10'b0;

   // m287_88 = W*in
   wire signed [9:0] m287_88;
   assign m287_88 =10'b0;

   // m287_89 = W*in
   wire signed [9:0] m287_89;
   assign m287_89 =10'b0;

   // m287_90 = W*in
   wire signed [9:0] m287_90;
   assign m287_90 =10'b0;

   // m287_91 = W*in
   wire signed [9:0] m287_91;
   assign m287_91 =10'b0;

   // m287_92 = W*in
   wire signed [9:0] m287_92;
   assign m287_92 =10'b0;

   // m287_93 = W*in
   wire signed [9:0] m287_93;
   assign m287_93 =10'b0;

   // m287_94 = W*in
   wire signed [9:0] m287_94;
   assign m287_94 =10'b0;

   // m287_95 = W*in
   wire signed [9:0] m287_95;
   assign m287_95 =10'b0;

   // m287_96 = W*in
   wire signed [9:0] m287_96;
   assign m287_96 =10'b0;

   // m287_97 = W*in
   wire signed [9:0] m287_97;
   assign m287_97 =10'b0;

   // m287_98 = W*in
   wire signed [9:0] m287_98;
   assign m287_98 =10'b0;

   // m287_99 = W*in
   wire signed [9:0] m287_99;
   assign m287_99 =10'b0;

   // m287_100 = W*in
   wire signed [9:0] m287_100;
   assign m287_100 =10'b0;

   // m287_101 = W*in
   wire signed [9:0] m287_101;
   assign m287_101 =10'b0;

   // m287_102 = W*in
   wire signed [9:0] m287_102;
   assign m287_102 =10'b0;

   // m287_103 = W*in
   wire signed [9:0] m287_103;
   assign m287_103 =10'b0;

   // m287_104 = W*in
   wire signed [9:0] m287_104;
   assign m287_104 =10'b0;

   // m287_105 = W*in
   wire signed [9:0] m287_105;
   assign m287_105 =10'b0;

   // m287_106 = W*in
   wire signed [9:0] m287_106;
   assign m287_106 =10'b0;

   // m287_107 = W*in
   wire signed [9:0] m287_107;
   assign m287_107 =10'b0;

   // m287_108 = W*in
   wire signed [9:0] m287_108;
   assign m287_108 =10'b0;

   // m287_109 = W*in
   wire signed [9:0] m287_109;
   assign m287_109 =10'b0;

   // m287_110 = W*in
   wire signed [9:0] m287_110;
   assign m287_110 =10'b0;

   // m287_111 = W*in
   wire signed [9:0] m287_111;
   assign m287_111 =10'b0;

   // m287_112 = W*in
   wire signed [9:0] m287_112;
   assign m287_112 =10'b0;

   // m287_113 = W*in
   wire signed [9:0] m287_113;
   assign m287_113 =10'b0;

   // m287_114 = W*in
   wire signed [9:0] m287_114;
   assign m287_114 =10'b0;

   // m287_115 = W*in
   wire signed [9:0] m287_115;
   assign m287_115 =10'b0;

   // m287_116 = W*in
   wire signed [9:0] m287_116;
   assign m287_116 =10'b0;

   // m287_117 = W*in
   wire signed [9:0] m287_117;
   assign m287_117 =10'b0;

   // m288_1 = W*in
   wire signed [9:0] m288_1;
   assign m288_1 =10'b0;

   // m288_2 = W*in
   wire signed [9:0] m288_2;
   assign m288_2 =10'b0;

   // m288_3 = W*in
   wire signed [9:0] m288_3;
   assign m288_3 =10'b0;

   // m288_4 = W*in
   wire signed [9:0] m288_4;
   assign m288_4 =10'b0;

   // m288_5 = W*in
   wire signed [9:0] m288_5;
   assign m288_5 =10'b0;

   // m288_6 = W*in
   wire signed [9:0] m288_6;
   assign m288_6 =10'b0;

   // m288_7 = W*in
   wire signed [9:0] m288_7;
   assign m288_7 =10'b0;

   // m288_8 = W*in
   wire signed [9:0] m288_8;
   assign m288_8 =10'b0;

   // m288_9 = W*in
   wire signed [9:0] m288_9;
   assign m288_9 =10'b0;

   // m288_10 = W*in
   wire signed [9:0] m288_10;
   assign m288_10 =10'b0;

   // m288_11 = W*in
   wire signed [9:0] m288_11;
   assign m288_11 =10'b0;

   // m288_12 = W*in
   wire signed [9:0] m288_12;
   assign m288_12 =10'b0;

   // m288_13 = W*in
   wire signed [9:0] m288_13;
   assign m288_13 =10'b0;

   // m288_14 = W*in
   wire signed [9:0] m288_14;
   assign m288_14 =10'b0;

   // m288_15 = W*in
   wire signed [9:0] m288_15;
   assign m288_15 =10'b0;

   // m288_16 = W*in
   wire signed [9:0] m288_16;
   assign m288_16 =10'b0;

   // m288_17 = W*in
   wire signed [9:0] m288_17;
   assign m288_17 =10'b0;

   // m288_18 = W*in
   wire signed [9:0] m288_18;
   assign m288_18 =10'b0;

   // m288_19 = W*in
   wire signed [9:0] m288_19;
   assign m288_19 =10'b0;

   // m288_20 = W*in
   wire signed [9:0] m288_20;
   assign m288_20 ={ {5{neg288[5]}} , neg288[5:1] };

   // m288_21 = W*in
   wire signed [9:0] m288_21;
   assign m288_21 =10'b0;

   // m288_22 = W*in
   wire signed [9:0] m288_22;
   assign m288_22 =10'b0;

   // m288_23 = W*in
   wire signed [9:0] m288_23;
   assign m288_23 =10'b0;

   // m288_24 = W*in
   wire signed [9:0] m288_24;
   assign m288_24 =10'b0;

   // m288_25 = W*in
   wire signed [9:0] m288_25;
   assign m288_25 =10'b0;

   // m288_26 = W*in
   wire signed [9:0] m288_26;
   assign m288_26 =10'b0;

   // m288_27 = W*in
   wire signed [9:0] m288_27;
   assign m288_27 =10'b0;

   // m288_28 = W*in
   wire signed [9:0] m288_28;
   assign m288_28 =10'b0;

   // m288_29 = W*in
   wire signed [9:0] m288_29;
   assign m288_29 =10'b0;

   // m288_30 = W*in
   wire signed [9:0] m288_30;
   assign m288_30 =10'b0;

   // m288_31 = W*in
   wire signed [9:0] m288_31;
   assign m288_31 =10'b0;

   // m288_32 = W*in
   wire signed [9:0] m288_32;
   assign m288_32 =10'b0;

   // m288_33 = W*in
   wire signed [9:0] m288_33;
   assign m288_33 =10'b0;

   // m288_34 = W*in
   wire signed [9:0] m288_34;
   assign m288_34 =10'b0;

   // m288_35 = W*in
   wire signed [9:0] m288_35;
   assign m288_35 =10'b0;

   // m288_36 = W*in
   wire signed [9:0] m288_36;
   assign m288_36 =10'b0;

   // m288_37 = W*in
   wire signed [9:0] m288_37;
   assign m288_37 =10'b0;

   // m288_38 = W*in
   wire signed [9:0] m288_38;
   assign m288_38 =10'b0;

   // m288_39 = W*in
   wire signed [9:0] m288_39;
   assign m288_39 =10'b0;

   // m288_40 = W*in
   wire signed [9:0] m288_40;
   assign m288_40 =10'b0;

   // m288_41 = W*in
   wire signed [9:0] m288_41;
   assign m288_41 =10'b0;

   // m288_42 = W*in
   wire signed [9:0] m288_42;
   assign m288_42 =10'b0;

   // m288_43 = W*in
   wire signed [9:0] m288_43;
   assign m288_43 =10'b0;

   // m288_44 = W*in
   wire signed [9:0] m288_44;
   assign m288_44 =10'b0;

   // m288_45 = W*in
   wire signed [9:0] m288_45;
   assign m288_45 =10'b0;

   // m288_46 = W*in
   wire signed [9:0] m288_46;
   assign m288_46 =10'b0;

   // m288_47 = W*in
   wire signed [9:0] m288_47;
   assign m288_47 =10'b0;

   // m288_48 = W*in
   wire signed [9:0] m288_48;
   assign m288_48 =10'b0;

   // m288_49 = W*in
   wire signed [9:0] m288_49;
   assign m288_49 =10'b0;

   // m288_50 = W*in
   wire signed [9:0] m288_50;
   assign m288_50 =10'b0;

   // m288_51 = W*in
   wire signed [9:0] m288_51;
   assign m288_51 =10'b0;

   // m288_52 = W*in
   wire signed [9:0] m288_52;
   assign m288_52 =10'b0;

   // m288_53 = W*in
   wire signed [9:0] m288_53;
   assign m288_53 =10'b0;

   // m288_54 = W*in
   wire signed [9:0] m288_54;
   assign m288_54 =10'b0;

   // m288_55 = W*in
   wire signed [9:0] m288_55;
   assign m288_55 =10'b0;

   // m288_56 = W*in
   wire signed [9:0] m288_56;
   assign m288_56 =10'b0;

   // m288_57 = W*in
   wire signed [9:0] m288_57;
   assign m288_57 =10'b0;

   // m288_58 = W*in
   wire signed [9:0] m288_58;
   assign m288_58 =10'b0;

   // m288_59 = W*in
   wire signed [9:0] m288_59;
   assign m288_59 =10'b0;

   // m288_60 = W*in
   wire signed [9:0] m288_60;
   assign m288_60 =10'b0;

   // m288_61 = W*in
   wire signed [9:0] m288_61;
   assign m288_61 =10'b0;

   // m288_62 = W*in
   wire signed [9:0] m288_62;
   assign m288_62 =10'b0;

   // m288_63 = W*in
   wire signed [9:0] m288_63;
   assign m288_63 =10'b0;

   // m288_64 = W*in
   wire signed [9:0] m288_64;
   assign m288_64 =10'b0;

   // m288_65 = W*in
   wire signed [9:0] m288_65;
   assign m288_65 =10'b0;

   // m288_66 = W*in
   wire signed [9:0] m288_66;
   assign m288_66 =10'b0;

   // m288_67 = W*in
   wire signed [9:0] m288_67;
   assign m288_67 =10'b0;

   // m288_68 = W*in
   wire signed [9:0] m288_68;
   assign m288_68 =10'b0;

   // m288_69 = W*in
   wire signed [9:0] m288_69;
   assign m288_69 =10'b0;

   // m288_70 = W*in
   wire signed [9:0] m288_70;
   assign m288_70 =10'b0;

   // m288_71 = W*in
   wire signed [9:0] m288_71;
   assign m288_71 =10'b0;

   // m288_72 = W*in
   wire signed [9:0] m288_72;
   assign m288_72 =10'b0;

   // m288_73 = W*in
   wire signed [9:0] m288_73;
   assign m288_73 =10'b0;

   // m288_74 = W*in
   wire signed [9:0] m288_74;
   assign m288_74 =10'b0;

   // m288_75 = W*in
   wire signed [9:0] m288_75;
   assign m288_75 =10'b0;

   // m288_76 = W*in
   wire signed [9:0] m288_76;
   assign m288_76 =10'b0;

   // m288_77 = W*in
   wire signed [9:0] m288_77;
   assign m288_77 =10'b0;

   // m288_78 = W*in
   wire signed [9:0] m288_78;
   assign m288_78 =10'b0;

   // m288_79 = W*in
   wire signed [9:0] m288_79;
   assign m288_79 =10'b0;

   // m288_80 = W*in
   wire signed [9:0] m288_80;
   assign m288_80 =10'b0;

   // m288_81 = W*in
   wire signed [9:0] m288_81;
   assign m288_81 =10'b0;

   // m288_82 = W*in
   wire signed [9:0] m288_82;
   assign m288_82 =10'b0;

   // m288_83 = W*in
   wire signed [9:0] m288_83;
   assign m288_83 =10'b0;

   // m288_84 = W*in
   wire signed [9:0] m288_84;
   assign m288_84 =10'b0;

   // m288_85 = W*in
   wire signed [9:0] m288_85;
   assign m288_85 =10'b0;

   // m288_86 = W*in
   wire signed [9:0] m288_86;
   assign m288_86 =10'b0;

   // m288_87 = W*in
   wire signed [9:0] m288_87;
   assign m288_87 =10'b0;

   // m288_88 = W*in
   wire signed [9:0] m288_88;
   assign m288_88 =10'b0;

   // m288_89 = W*in
   wire signed [9:0] m288_89;
   assign m288_89 =10'b0;

   // m288_90 = W*in
   wire signed [9:0] m288_90;
   assign m288_90 =10'b0;

   // m288_91 = W*in
   wire signed [9:0] m288_91;
   assign m288_91 =10'b0;

   // m288_92 = W*in
   wire signed [9:0] m288_92;
   assign m288_92 =10'b0;

   // m288_93 = W*in
   wire signed [9:0] m288_93;
   assign m288_93 =10'b0;

   // m288_94 = W*in
   wire signed [9:0] m288_94;
   assign m288_94 =10'b0;

   // m288_95 = W*in
   wire signed [9:0] m288_95;
   assign m288_95 =10'b0;

   // m288_96 = W*in
   wire signed [9:0] m288_96;
   assign m288_96 =10'b0;

   // m288_97 = W*in
   wire signed [9:0] m288_97;
   assign m288_97 =10'b0;

   // m288_98 = W*in
   wire signed [9:0] m288_98;
   assign m288_98 =10'b0;

   // m288_99 = W*in
   wire signed [9:0] m288_99;
   assign m288_99 =10'b0;

   // m288_100 = W*in
   wire signed [9:0] m288_100;
   assign m288_100 =10'b0;

   // m288_101 = W*in
   wire signed [9:0] m288_101;
   assign m288_101 =10'b0;

   // m288_102 = W*in
   wire signed [9:0] m288_102;
   assign m288_102 =10'b0;

   // m288_103 = W*in
   wire signed [9:0] m288_103;
   assign m288_103 =10'b0;

   // m288_104 = W*in
   wire signed [9:0] m288_104;
   assign m288_104 =10'b0;

   // m288_105 = W*in
   wire signed [9:0] m288_105;
   assign m288_105 =10'b0;

   // m288_106 = W*in
   wire signed [9:0] m288_106;
   assign m288_106 =10'b0;

   // m288_107 = W*in
   wire signed [9:0] m288_107;
   assign m288_107 =10'b0;

   // m288_108 = W*in
   wire signed [9:0] m288_108;
   assign m288_108 =10'b0;

   // m288_109 = W*in
   wire signed [9:0] m288_109;
   assign m288_109 =10'b0;

   // m288_110 = W*in
   wire signed [9:0] m288_110;
   assign m288_110 =10'b0;

   // m288_111 = W*in
   wire signed [9:0] m288_111;
   assign m288_111 =10'b0;

   // m288_112 = W*in
   wire signed [9:0] m288_112;
   assign m288_112 =10'b0;

   // m288_113 = W*in
   wire signed [9:0] m288_113;
   assign m288_113 =10'b0;

   // m288_114 = W*in
   wire signed [9:0] m288_114;
   assign m288_114 =10'b0;

   // m288_115 = W*in
   wire signed [9:0] m288_115;
   assign m288_115 =10'b0;

   // m288_116 = W*in
   wire signed [9:0] m288_116;
   assign m288_116 =10'b0;

   // m288_117 = W*in
   wire signed [9:0] m288_117;
   assign m288_117 =10'b0;

   // m289_1 = W*in
   wire signed [9:0] m289_1;
   assign m289_1 =10'b0;

   // m289_2 = W*in
   wire signed [9:0] m289_2;
   assign m289_2 =10'b0;

   // m289_3 = W*in
   wire signed [9:0] m289_3;
   assign m289_3 =10'b0;

   // m289_4 = W*in
   wire signed [9:0] m289_4;
   assign m289_4 =10'b0;

   // m289_5 = W*in
   wire signed [9:0] m289_5;
   assign m289_5 =10'b0;

   // m289_6 = W*in
   wire signed [9:0] m289_6;
   assign m289_6 =10'b0;

   // m289_7 = W*in
   wire signed [9:0] m289_7;
   assign m289_7 =10'b0;

   // m289_8 = W*in
   wire signed [9:0] m289_8;
   assign m289_8 =10'b0;

   // m289_9 = W*in
   wire signed [9:0] m289_9;
   assign m289_9 =10'b0;

   // m289_10 = W*in
   wire signed [9:0] m289_10;
   assign m289_10 =10'b0;

   // m289_11 = W*in
   wire signed [9:0] m289_11;
   assign m289_11 =10'b0;

   // m289_12 = W*in
   wire signed [9:0] m289_12;
   assign m289_12 =10'b0;

   // m289_13 = W*in
   wire signed [9:0] m289_13;
   assign m289_13 =10'b0;

   // m289_14 = W*in
   wire signed [9:0] m289_14;
   assign m289_14 =10'b0;

   // m289_15 = W*in
   wire signed [9:0] m289_15;
   assign m289_15 =10'b0;

   // m289_16 = W*in
   wire signed [9:0] m289_16;
   assign m289_16 =10'b0;

   // m289_17 = W*in
   wire signed [9:0] m289_17;
   assign m289_17 =10'b0;

   // m289_18 = W*in
   wire signed [9:0] m289_18;
   assign m289_18 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_19 = W*in
   wire signed [9:0] m289_19;
   assign m289_19 ={ {4{in289[5]}} , in289[5:0] };

   // m289_20 = W*in
   wire signed [9:0] m289_20;
   assign m289_20 =10'b0;

   // m289_21 = W*in
   wire signed [9:0] m289_21;
   assign m289_21 =10'b0;

   // m289_22 = W*in
   wire signed [9:0] m289_22;
   assign m289_22 =10'b0;

   // m289_23 = W*in
   wire signed [9:0] m289_23;
   assign m289_23 =10'b0;

   // m289_24 = W*in
   wire signed [9:0] m289_24;
   assign m289_24 =10'b0;

   // m289_25 = W*in
   wire signed [9:0] m289_25;
   assign m289_25 =10'b0;

   // m289_26 = W*in
   wire signed [9:0] m289_26;
   assign m289_26 ={ {4{neg289[5]}} , neg289[5:0] };

   // m289_27 = W*in
   wire signed [9:0] m289_27;
   assign m289_27 =10'b0;

   // m289_28 = W*in
   wire signed [9:0] m289_28;
   assign m289_28 =10'b0;

   // m289_29 = W*in
   wire signed [9:0] m289_29;
   assign m289_29 ={ {4{in289[5]}} , in289[5:0] };

   // m289_30 = W*in
   wire signed [9:0] m289_30;
   assign m289_30 =10'b0;

   // m289_31 = W*in
   wire signed [9:0] m289_31;
   assign m289_31 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_32 = W*in
   wire signed [9:0] m289_32;
   assign m289_32 =10'b0;

   // m289_33 = W*in
   wire signed [9:0] m289_33;
   assign m289_33 =10'b0;

   // m289_34 = W*in
   wire signed [9:0] m289_34;
   assign m289_34 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_35 = W*in
   wire signed [9:0] m289_35;
   assign m289_35 =10'b0;

   // m289_36 = W*in
   wire signed [9:0] m289_36;
   assign m289_36 =10'b0;

   // m289_37 = W*in
   wire signed [9:0] m289_37;
   assign m289_37 =10'b0;

   // m289_38 = W*in
   wire signed [9:0] m289_38;
   assign m289_38 =10'b0;

   // m289_39 = W*in
   wire signed [9:0] m289_39;
   assign m289_39 =10'b0;

   // m289_40 = W*in
   wire signed [9:0] m289_40;
   assign m289_40 =10'b0;

   // m289_41 = W*in
   wire signed [9:0] m289_41;
   assign m289_41 =10'b0;

   // m289_42 = W*in
   wire signed [9:0] m289_42;
   assign m289_42 =10'b0;

   // m289_43 = W*in
   wire signed [9:0] m289_43;
   assign m289_43 =10'b0;

   // m289_44 = W*in
   wire signed [9:0] m289_44;
   assign m289_44 =10'b0;

   // m289_45 = W*in
   wire signed [9:0] m289_45;
   assign m289_45 =10'b0;

   // m289_46 = W*in
   wire signed [9:0] m289_46;
   assign m289_46 =10'b0;

   // m289_47 = W*in
   wire signed [9:0] m289_47;
   assign m289_47 =10'b0;

   // m289_48 = W*in
   wire signed [9:0] m289_48;
   assign m289_48 =10'b0;

   // m289_49 = W*in
   wire signed [9:0] m289_49;
   assign m289_49 ={ {4{in289[5]}} , in289[5:0] };

   // m289_50 = W*in
   wire signed [9:0] m289_50;
   assign m289_50 =10'b0;

   // m289_51 = W*in
   wire signed [9:0] m289_51;
   assign m289_51 =10'b0;

   // m289_52 = W*in
   wire signed [9:0] m289_52;
   assign m289_52 =10'b0;

   // m289_53 = W*in
   wire signed [9:0] m289_53;
   assign m289_53 ={ {4{in289[5]}} , in289[5:0] };

   // m289_54 = W*in
   wire signed [9:0] m289_54;
   assign m289_54 =10'b0;

   // m289_55 = W*in
   wire signed [9:0] m289_55;
   assign m289_55 =10'b0;

   // m289_56 = W*in
   wire signed [9:0] m289_56;
   assign m289_56 =10'b0;

   // m289_57 = W*in
   wire signed [9:0] m289_57;
   assign m289_57 =10'b0;

   // m289_58 = W*in
   wire signed [9:0] m289_58;
   assign m289_58 =10'b0;

   // m289_59 = W*in
   wire signed [9:0] m289_59;
   assign m289_59 =10'b0;

   // m289_60 = W*in
   wire signed [9:0] m289_60;
   assign m289_60 =10'b0;

   // m289_61 = W*in
   wire signed [9:0] m289_61;
   assign m289_61 =10'b0;

   // m289_62 = W*in
   wire signed [9:0] m289_62;
   assign m289_62 =10'b0;

   // m289_63 = W*in
   wire signed [9:0] m289_63;
   assign m289_63 =10'b0;

   // m289_64 = W*in
   wire signed [9:0] m289_64;
   assign m289_64 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_65 = W*in
   wire signed [9:0] m289_65;
   assign m289_65 =10'b0;

   // m289_66 = W*in
   wire signed [9:0] m289_66;
   assign m289_66 =10'b0;

   // m289_67 = W*in
   wire signed [9:0] m289_67;
   assign m289_67 ={ {4{in289[5]}} , in289[5:0] };

   // m289_68 = W*in
   wire signed [9:0] m289_68;
   assign m289_68 =10'b0;

   // m289_69 = W*in
   wire signed [9:0] m289_69;
   assign m289_69 =10'b0;

   // m289_70 = W*in
   wire signed [9:0] m289_70;
   assign m289_70 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_71 = W*in
   wire signed [9:0] m289_71;
   assign m289_71 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_72 = W*in
   wire signed [9:0] m289_72;
   assign m289_72 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_73 = W*in
   wire signed [9:0] m289_73;
   assign m289_73 =10'b0;

   // m289_74 = W*in
   wire signed [9:0] m289_74;
   assign m289_74 =10'b0;

   // m289_75 = W*in
   wire signed [9:0] m289_75;
   assign m289_75 =10'b0;

   // m289_76 = W*in
   wire signed [9:0] m289_76;
   assign m289_76 =10'b0;

   // m289_77 = W*in
   wire signed [9:0] m289_77;
   assign m289_77 =10'b0;

   // m289_78 = W*in
   wire signed [9:0] m289_78;
   assign m289_78 =10'b0;

   // m289_79 = W*in
   wire signed [9:0] m289_79;
   assign m289_79 =10'b0;

   // m289_80 = W*in
   wire signed [9:0] m289_80;
   assign m289_80 =10'b0;

   // m289_81 = W*in
   wire signed [9:0] m289_81;
   assign m289_81 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_82 = W*in
   wire signed [9:0] m289_82;
   assign m289_82 =10'b0;

   // m289_83 = W*in
   wire signed [9:0] m289_83;
   assign m289_83 =10'b0;

   // m289_84 = W*in
   wire signed [9:0] m289_84;
   assign m289_84 =10'b0;

   // m289_85 = W*in
   wire signed [9:0] m289_85;
   assign m289_85 ={ {5{in289[5]}} , in289[5:1] };

   // m289_86 = W*in
   wire signed [9:0] m289_86;
   assign m289_86 =10'b0;

   // m289_87 = W*in
   wire signed [9:0] m289_87;
   assign m289_87 =10'b0;

   // m289_88 = W*in
   wire signed [9:0] m289_88;
   assign m289_88 =10'b0;

   // m289_89 = W*in
   wire signed [9:0] m289_89;
   assign m289_89 ={ {4{neg289[5]}} , neg289[5:0] };

   // m289_90 = W*in
   wire signed [9:0] m289_90;
   assign m289_90 =10'b0;

   // m289_91 = W*in
   wire signed [9:0] m289_91;
   assign m289_91 =10'b0;

   // m289_92 = W*in
   wire signed [9:0] m289_92;
   assign m289_92 =10'b0;

   // m289_93 = W*in
   wire signed [9:0] m289_93;
   assign m289_93 ={ {4{in289[5]}} , in289[5:0] };

   // m289_94 = W*in
   wire signed [9:0] m289_94;
   assign m289_94 =10'b0;

   // m289_95 = W*in
   wire signed [9:0] m289_95;
   assign m289_95 =10'b0;

   // m289_96 = W*in
   wire signed [9:0] m289_96;
   assign m289_96 =10'b0;

   // m289_97 = W*in
   wire signed [9:0] m289_97;
   assign m289_97 =10'b0;

   // m289_98 = W*in
   wire signed [9:0] m289_98;
   assign m289_98 =10'b0;

   // m289_99 = W*in
   wire signed [9:0] m289_99;
   assign m289_99 =10'b0;

   // m289_100 = W*in
   wire signed [9:0] m289_100;
   assign m289_100 =10'b0;

   // m289_101 = W*in
   wire signed [9:0] m289_101;
   assign m289_101 =10'b0;

   // m289_102 = W*in
   wire signed [9:0] m289_102;
   assign m289_102 =10'b0;

   // m289_103 = W*in
   wire signed [9:0] m289_103;
   assign m289_103 =10'b0;

   // m289_104 = W*in
   wire signed [9:0] m289_104;
   assign m289_104 =10'b0;

   // m289_105 = W*in
   wire signed [9:0] m289_105;
   assign m289_105 =10'b0;

   // m289_106 = W*in
   wire signed [9:0] m289_106;
   assign m289_106 =10'b0;

   // m289_107 = W*in
   wire signed [9:0] m289_107;
   assign m289_107 =10'b0;

   // m289_108 = W*in
   wire signed [9:0] m289_108;
   assign m289_108 ={ {5{neg289[5]}} , neg289[5:1] };

   // m289_109 = W*in
   wire signed [9:0] m289_109;
   assign m289_109 ={ {4{neg289[5]}} , neg289[5:0] };

   // m289_110 = W*in
   wire signed [9:0] m289_110;
   assign m289_110 =10'b0;

   // m289_111 = W*in
   wire signed [9:0] m289_111;
   assign m289_111 =10'b0;

   // m289_112 = W*in
   wire signed [9:0] m289_112;
   assign m289_112 =10'b0;

   // m289_113 = W*in
   wire signed [9:0] m289_113;
   assign m289_113 =10'b0;

   // m289_114 = W*in
   wire signed [9:0] m289_114;
   assign m289_114 =10'b0;

   // m289_115 = W*in
   wire signed [9:0] m289_115;
   assign m289_115 =10'b0;

   // m289_116 = W*in
   wire signed [9:0] m289_116;
   assign m289_116 =10'b0;

   // m289_117 = W*in
   wire signed [9:0] m289_117;
   assign m289_117 =10'b0;

   // m290_1 = W*in
   wire signed [9:0] m290_1;
   assign m290_1 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_2 = W*in
   wire signed [9:0] m290_2;
   assign m290_2 =10'b0;

   // m290_3 = W*in
   wire signed [9:0] m290_3;
   assign m290_3 =10'b0;

   // m290_4 = W*in
   wire signed [9:0] m290_4;
   assign m290_4 =10'b0;

   // m290_5 = W*in
   wire signed [9:0] m290_5;
   assign m290_5 ={ {4{in290[5]}} , in290[5:0] };

   // m290_6 = W*in
   wire signed [9:0] m290_6;
   assign m290_6 ={ {5{in290[5]}} , in290[5:1] };

   // m290_7 = W*in
   wire signed [9:0] m290_7;
   assign m290_7 =10'b0;

   // m290_8 = W*in
   wire signed [9:0] m290_8;
   assign m290_8 ={ {4{in290[5]}} , in290[5:0] };

   // m290_9 = W*in
   wire signed [9:0] m290_9;
   assign m290_9 =10'b0;

   // m290_10 = W*in
   wire signed [9:0] m290_10;
   assign m290_10 =10'b0;

   // m290_11 = W*in
   wire signed [9:0] m290_11;
   assign m290_11 =10'b0;

   // m290_12 = W*in
   wire signed [9:0] m290_12;
   assign m290_12 =10'b0;

   // m290_13 = W*in
   wire signed [9:0] m290_13;
   assign m290_13 =10'b0;

   // m290_14 = W*in
   wire signed [9:0] m290_14;
   assign m290_14 =10'b0;

   // m290_15 = W*in
   wire signed [9:0] m290_15;
   assign m290_15 =10'b0;

   // m290_16 = W*in
   wire signed [9:0] m290_16;
   assign m290_16 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_17 = W*in
   wire signed [9:0] m290_17;
   assign m290_17 =10'b0;

   // m290_18 = W*in
   wire signed [9:0] m290_18;
   assign m290_18 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_19 = W*in
   wire signed [9:0] m290_19;
   assign m290_19 ={ {4{in290[5]}} , in290[5:0] };

   // m290_20 = W*in
   wire signed [9:0] m290_20;
   assign m290_20 =10'b0;

   // m290_21 = W*in
   wire signed [9:0] m290_21;
   assign m290_21 =10'b0;

   // m290_22 = W*in
   wire signed [9:0] m290_22;
   assign m290_22 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_23 = W*in
   wire signed [9:0] m290_23;
   assign m290_23 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_24 = W*in
   wire signed [9:0] m290_24;
   assign m290_24 =10'b0;

   // m290_25 = W*in
   wire signed [9:0] m290_25;
   assign m290_25 =10'b0;

   // m290_26 = W*in
   wire signed [9:0] m290_26;
   assign m290_26 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_27 = W*in
   wire signed [9:0] m290_27;
   assign m290_27 =10'b0;

   // m290_28 = W*in
   wire signed [9:0] m290_28;
   assign m290_28 =10'b0;

   // m290_29 = W*in
   wire signed [9:0] m290_29;
   assign m290_29 =10'b0;

   // m290_30 = W*in
   wire signed [9:0] m290_30;
   assign m290_30 =10'b0;

   // m290_31 = W*in
   wire signed [9:0] m290_31;
   assign m290_31 =10'b0;

   // m290_32 = W*in
   wire signed [9:0] m290_32;
   assign m290_32 ={ {4{in290[5]}} , in290[5:0] };

   // m290_33 = W*in
   wire signed [9:0] m290_33;
   assign m290_33 =10'b0;

   // m290_34 = W*in
   wire signed [9:0] m290_34;
   assign m290_34 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_35 = W*in
   wire signed [9:0] m290_35;
   assign m290_35 =10'b0;

   // m290_36 = W*in
   wire signed [9:0] m290_36;
   assign m290_36 =10'b0;

   // m290_37 = W*in
   wire signed [9:0] m290_37;
   assign m290_37 =10'b0;

   // m290_38 = W*in
   wire signed [9:0] m290_38;
   assign m290_38 =10'b0;

   // m290_39 = W*in
   wire signed [9:0] m290_39;
   assign m290_39 =10'b0;

   // m290_40 = W*in
   wire signed [9:0] m290_40;
   assign m290_40 =10'b0;

   // m290_41 = W*in
   wire signed [9:0] m290_41;
   assign m290_41 =10'b0;

   // m290_42 = W*in
   wire signed [9:0] m290_42;
   assign m290_42 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_43 = W*in
   wire signed [9:0] m290_43;
   assign m290_43 =10'b0;

   // m290_44 = W*in
   wire signed [9:0] m290_44;
   assign m290_44 =10'b0;

   // m290_45 = W*in
   wire signed [9:0] m290_45;
   assign m290_45 =10'b0;

   // m290_46 = W*in
   wire signed [9:0] m290_46;
   assign m290_46 =10'b0;

   // m290_47 = W*in
   wire signed [9:0] m290_47;
   assign m290_47 =10'b0;

   // m290_48 = W*in
   wire signed [9:0] m290_48;
   assign m290_48 =10'b0;

   // m290_49 = W*in
   wire signed [9:0] m290_49;
   assign m290_49 =10'b0;

   // m290_50 = W*in
   wire signed [9:0] m290_50;
   assign m290_50 =10'b0;

   // m290_51 = W*in
   wire signed [9:0] m290_51;
   assign m290_51 ={ {4{in290[5]}} , in290[5:0] };

   // m290_52 = W*in
   wire signed [9:0] m290_52;
   assign m290_52 =10'b0;

   // m290_53 = W*in
   wire signed [9:0] m290_53;
   assign m290_53 ={ {4{in290[5]}} , in290[5:0] };

   // m290_54 = W*in
   wire signed [9:0] m290_54;
   assign m290_54 ={ {4{in290[5]}} , in290[5:0] };

   // m290_55 = W*in
   wire signed [9:0] m290_55;
   assign m290_55 =10'b0;

   // m290_56 = W*in
   wire signed [9:0] m290_56;
   assign m290_56 =10'b0;

   // m290_57 = W*in
   wire signed [9:0] m290_57;
   assign m290_57 =10'b0;

   // m290_58 = W*in
   wire signed [9:0] m290_58;
   assign m290_58 =10'b0;

   // m290_59 = W*in
   wire signed [9:0] m290_59;
   assign m290_59 =10'b0;

   // m290_60 = W*in
   wire signed [9:0] m290_60;
   assign m290_60 =10'b0;

   // m290_61 = W*in
   wire signed [9:0] m290_61;
   assign m290_61 =10'b0;

   // m290_62 = W*in
   wire signed [9:0] m290_62;
   assign m290_62 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_63 = W*in
   wire signed [9:0] m290_63;
   assign m290_63 =10'b0;

   // m290_64 = W*in
   wire signed [9:0] m290_64;
   assign m290_64 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_65 = W*in
   wire signed [9:0] m290_65;
   assign m290_65 =10'b0;

   // m290_66 = W*in
   wire signed [9:0] m290_66;
   assign m290_66 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_67 = W*in
   wire signed [9:0] m290_67;
   assign m290_67 =10'b0;

   // m290_68 = W*in
   wire signed [9:0] m290_68;
   assign m290_68 =10'b0;

   // m290_69 = W*in
   wire signed [9:0] m290_69;
   assign m290_69 =10'b0;

   // m290_70 = W*in
   wire signed [9:0] m290_70;
   assign m290_70 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_71 = W*in
   wire signed [9:0] m290_71;
   assign m290_71 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_72 = W*in
   wire signed [9:0] m290_72;
   assign m290_72 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_73 = W*in
   wire signed [9:0] m290_73;
   assign m290_73 =10'b0;

   // m290_74 = W*in
   wire signed [9:0] m290_74;
   assign m290_74 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_75 = W*in
   wire signed [9:0] m290_75;
   assign m290_75 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_76 = W*in
   wire signed [9:0] m290_76;
   assign m290_76 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_77 = W*in
   wire signed [9:0] m290_77;
   assign m290_77 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_78 = W*in
   wire signed [9:0] m290_78;
   assign m290_78 =10'b0;

   // m290_79 = W*in
   wire signed [9:0] m290_79;
   assign m290_79 =10'b0;

   // m290_80 = W*in
   wire signed [9:0] m290_80;
   assign m290_80 =10'b0;

   // m290_81 = W*in
   wire signed [9:0] m290_81;
   assign m290_81 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_82 = W*in
   wire signed [9:0] m290_82;
   assign m290_82 =10'b0;

   // m290_83 = W*in
   wire signed [9:0] m290_83;
   assign m290_83 =10'b0;

   // m290_84 = W*in
   wire signed [9:0] m290_84;
   assign m290_84 =10'b0;

   // m290_85 = W*in
   wire signed [9:0] m290_85;
   assign m290_85 ={ {4{in290[5]}} , in290[5:0] };

   // m290_86 = W*in
   wire signed [9:0] m290_86;
   assign m290_86 =10'b0;

   // m290_87 = W*in
   wire signed [9:0] m290_87;
   assign m290_87 =10'b0;

   // m290_88 = W*in
   wire signed [9:0] m290_88;
   assign m290_88 =10'b0;

   // m290_89 = W*in
   wire signed [9:0] m290_89;
   assign m290_89 =10'b0;

   // m290_90 = W*in
   wire signed [9:0] m290_90;
   assign m290_90 =10'b0;

   // m290_91 = W*in
   wire signed [9:0] m290_91;
   assign m290_91 =10'b0;

   // m290_92 = W*in
   wire signed [9:0] m290_92;
   assign m290_92 =10'b0;

   // m290_93 = W*in
   wire signed [9:0] m290_93;
   assign m290_93 ={ {4{in290[5]}} , in290[5:0] };

   // m290_94 = W*in
   wire signed [9:0] m290_94;
   assign m290_94 =10'b0;

   // m290_95 = W*in
   wire signed [9:0] m290_95;
   assign m290_95 ={ {5{in290[5]}} , in290[5:1] };

   // m290_96 = W*in
   wire signed [9:0] m290_96;
   assign m290_96 =10'b0;

   // m290_97 = W*in
   wire signed [9:0] m290_97;
   assign m290_97 =10'b0;

   // m290_98 = W*in
   wire signed [9:0] m290_98;
   assign m290_98 =10'b0;

   // m290_99 = W*in
   wire signed [9:0] m290_99;
   assign m290_99 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_100 = W*in
   wire signed [9:0] m290_100;
   assign m290_100 =10'b0;

   // m290_101 = W*in
   wire signed [9:0] m290_101;
   assign m290_101 =10'b0;

   // m290_102 = W*in
   wire signed [9:0] m290_102;
   assign m290_102 =10'b0;

   // m290_103 = W*in
   wire signed [9:0] m290_103;
   assign m290_103 =10'b0;

   // m290_104 = W*in
   wire signed [9:0] m290_104;
   assign m290_104 =10'b0;

   // m290_105 = W*in
   wire signed [9:0] m290_105;
   assign m290_105 =10'b0;

   // m290_106 = W*in
   wire signed [9:0] m290_106;
   assign m290_106 =10'b0;

   // m290_107 = W*in
   wire signed [9:0] m290_107;
   assign m290_107 =10'b0;

   // m290_108 = W*in
   wire signed [9:0] m290_108;
   assign m290_108 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_109 = W*in
   wire signed [9:0] m290_109;
   assign m290_109 ={ {5{neg290[5]}} , neg290[5:1] };

   // m290_110 = W*in
   wire signed [9:0] m290_110;
   assign m290_110 =10'b0;

   // m290_111 = W*in
   wire signed [9:0] m290_111;
   assign m290_111 =10'b0;

   // m290_112 = W*in
   wire signed [9:0] m290_112;
   assign m290_112 ={ {4{neg290[5]}} , neg290[5:0] };

   // m290_113 = W*in
   wire signed [9:0] m290_113;
   assign m290_113 =10'b0;

   // m290_114 = W*in
   wire signed [9:0] m290_114;
   assign m290_114 =10'b0;

   // m290_115 = W*in
   wire signed [9:0] m290_115;
   assign m290_115 =10'b0;

   // m290_116 = W*in
   wire signed [9:0] m290_116;
   assign m290_116 =10'b0;

   // m290_117 = W*in
   wire signed [9:0] m290_117;
   assign m290_117 =10'b0;

   // m291_1 = W*in
   wire signed [9:0] m291_1;
   assign m291_1 =10'b0;

   // m291_2 = W*in
   wire signed [9:0] m291_2;
   assign m291_2 =10'b0;

   // m291_3 = W*in
   wire signed [9:0] m291_3;
   assign m291_3 =10'b0;

   // m291_4 = W*in
   wire signed [9:0] m291_4;
   assign m291_4 =10'b0;

   // m291_5 = W*in
   wire signed [9:0] m291_5;
   assign m291_5 =10'b0;

   // m291_6 = W*in
   wire signed [9:0] m291_6;
   assign m291_6 =10'b0;

   // m291_7 = W*in
   wire signed [9:0] m291_7;
   assign m291_7 =10'b0;

   // m291_8 = W*in
   wire signed [9:0] m291_8;
   assign m291_8 =10'b0;

   // m291_9 = W*in
   wire signed [9:0] m291_9;
   assign m291_9 =10'b0;

   // m291_10 = W*in
   wire signed [9:0] m291_10;
   assign m291_10 =10'b0;

   // m291_11 = W*in
   wire signed [9:0] m291_11;
   assign m291_11 =10'b0;

   // m291_12 = W*in
   wire signed [9:0] m291_12;
   assign m291_12 =10'b0;

   // m291_13 = W*in
   wire signed [9:0] m291_13;
   assign m291_13 =10'b0;

   // m291_14 = W*in
   wire signed [9:0] m291_14;
   assign m291_14 =10'b0;

   // m291_15 = W*in
   wire signed [9:0] m291_15;
   assign m291_15 =10'b0;

   // m291_16 = W*in
   wire signed [9:0] m291_16;
   assign m291_16 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_17 = W*in
   wire signed [9:0] m291_17;
   assign m291_17 ={ {5{in291[5]}} , in291[5:1] };

   // m291_18 = W*in
   wire signed [9:0] m291_18;
   assign m291_18 =10'b0;

   // m291_19 = W*in
   wire signed [9:0] m291_19;
   assign m291_19 =10'b0;

   // m291_20 = W*in
   wire signed [9:0] m291_20;
   assign m291_20 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_21 = W*in
   wire signed [9:0] m291_21;
   assign m291_21 =10'b0;

   // m291_22 = W*in
   wire signed [9:0] m291_22;
   assign m291_22 =10'b0;

   // m291_23 = W*in
   wire signed [9:0] m291_23;
   assign m291_23 =10'b0;

   // m291_24 = W*in
   wire signed [9:0] m291_24;
   assign m291_24 =10'b0;

   // m291_25 = W*in
   wire signed [9:0] m291_25;
   assign m291_25 =10'b0;

   // m291_26 = W*in
   wire signed [9:0] m291_26;
   assign m291_26 =10'b0;

   // m291_27 = W*in
   wire signed [9:0] m291_27;
   assign m291_27 =10'b0;

   // m291_28 = W*in
   wire signed [9:0] m291_28;
   assign m291_28 ={ {5{in291[5]}} , in291[5:1] };

   // m291_29 = W*in
   wire signed [9:0] m291_29;
   assign m291_29 =10'b0;

   // m291_30 = W*in
   wire signed [9:0] m291_30;
   assign m291_30 =10'b0;

   // m291_31 = W*in
   wire signed [9:0] m291_31;
   assign m291_31 ={ {5{in291[5]}} , in291[5:1] };

   // m291_32 = W*in
   wire signed [9:0] m291_32;
   assign m291_32 =10'b0;

   // m291_33 = W*in
   wire signed [9:0] m291_33;
   assign m291_33 =10'b0;

   // m291_34 = W*in
   wire signed [9:0] m291_34;
   assign m291_34 =10'b0;

   // m291_35 = W*in
   wire signed [9:0] m291_35;
   assign m291_35 =10'b0;

   // m291_36 = W*in
   wire signed [9:0] m291_36;
   assign m291_36 =10'b0;

   // m291_37 = W*in
   wire signed [9:0] m291_37;
   assign m291_37 =10'b0;

   // m291_38 = W*in
   wire signed [9:0] m291_38;
   assign m291_38 =10'b0;

   // m291_39 = W*in
   wire signed [9:0] m291_39;
   assign m291_39 =10'b0;

   // m291_40 = W*in
   wire signed [9:0] m291_40;
   assign m291_40 =10'b0;

   // m291_41 = W*in
   wire signed [9:0] m291_41;
   assign m291_41 =10'b0;

   // m291_42 = W*in
   wire signed [9:0] m291_42;
   assign m291_42 =10'b0;

   // m291_43 = W*in
   wire signed [9:0] m291_43;
   assign m291_43 =10'b0;

   // m291_44 = W*in
   wire signed [9:0] m291_44;
   assign m291_44 =10'b0;

   // m291_45 = W*in
   wire signed [9:0] m291_45;
   assign m291_45 =10'b0;

   // m291_46 = W*in
   wire signed [9:0] m291_46;
   assign m291_46 =10'b0;

   // m291_47 = W*in
   wire signed [9:0] m291_47;
   assign m291_47 =10'b0;

   // m291_48 = W*in
   wire signed [9:0] m291_48;
   assign m291_48 =10'b0;

   // m291_49 = W*in
   wire signed [9:0] m291_49;
   assign m291_49 =10'b0;

   // m291_50 = W*in
   wire signed [9:0] m291_50;
   assign m291_50 =10'b0;

   // m291_51 = W*in
   wire signed [9:0] m291_51;
   assign m291_51 ={ {4{in291[5]}} , in291[5:0] };

   // m291_52 = W*in
   wire signed [9:0] m291_52;
   assign m291_52 =10'b0;

   // m291_53 = W*in
   wire signed [9:0] m291_53;
   assign m291_53 =10'b0;

   // m291_54 = W*in
   wire signed [9:0] m291_54;
   assign m291_54 =10'b0;

   // m291_55 = W*in
   wire signed [9:0] m291_55;
   assign m291_55 =10'b0;

   // m291_56 = W*in
   wire signed [9:0] m291_56;
   assign m291_56 =10'b0;

   // m291_57 = W*in
   wire signed [9:0] m291_57;
   assign m291_57 =10'b0;

   // m291_58 = W*in
   wire signed [9:0] m291_58;
   assign m291_58 =10'b0;

   // m291_59 = W*in
   wire signed [9:0] m291_59;
   assign m291_59 =10'b0;

   // m291_60 = W*in
   wire signed [9:0] m291_60;
   assign m291_60 =10'b0;

   // m291_61 = W*in
   wire signed [9:0] m291_61;
   assign m291_61 =10'b0;

   // m291_62 = W*in
   wire signed [9:0] m291_62;
   assign m291_62 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_63 = W*in
   wire signed [9:0] m291_63;
   assign m291_63 =10'b0;

   // m291_64 = W*in
   wire signed [9:0] m291_64;
   assign m291_64 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_65 = W*in
   wire signed [9:0] m291_65;
   assign m291_65 =10'b0;

   // m291_66 = W*in
   wire signed [9:0] m291_66;
   assign m291_66 =10'b0;

   // m291_67 = W*in
   wire signed [9:0] m291_67;
   assign m291_67 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_68 = W*in
   wire signed [9:0] m291_68;
   assign m291_68 =10'b0;

   // m291_69 = W*in
   wire signed [9:0] m291_69;
   assign m291_69 =10'b0;

   // m291_70 = W*in
   wire signed [9:0] m291_70;
   assign m291_70 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_71 = W*in
   wire signed [9:0] m291_71;
   assign m291_71 =10'b0;

   // m291_72 = W*in
   wire signed [9:0] m291_72;
   assign m291_72 =10'b0;

   // m291_73 = W*in
   wire signed [9:0] m291_73;
   assign m291_73 =10'b0;

   // m291_74 = W*in
   wire signed [9:0] m291_74;
   assign m291_74 =10'b0;

   // m291_75 = W*in
   wire signed [9:0] m291_75;
   assign m291_75 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_76 = W*in
   wire signed [9:0] m291_76;
   assign m291_76 =10'b0;

   // m291_77 = W*in
   wire signed [9:0] m291_77;
   assign m291_77 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_78 = W*in
   wire signed [9:0] m291_78;
   assign m291_78 =10'b0;

   // m291_79 = W*in
   wire signed [9:0] m291_79;
   assign m291_79 =10'b0;

   // m291_80 = W*in
   wire signed [9:0] m291_80;
   assign m291_80 =10'b0;

   // m291_81 = W*in
   wire signed [9:0] m291_81;
   assign m291_81 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_82 = W*in
   wire signed [9:0] m291_82;
   assign m291_82 ={ {4{in291[5]}} , in291[5:0] };

   // m291_83 = W*in
   wire signed [9:0] m291_83;
   assign m291_83 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_84 = W*in
   wire signed [9:0] m291_84;
   assign m291_84 =10'b0;

   // m291_85 = W*in
   wire signed [9:0] m291_85;
   assign m291_85 ={ {5{in291[5]}} , in291[5:1] };

   // m291_86 = W*in
   wire signed [9:0] m291_86;
   assign m291_86 =10'b0;

   // m291_87 = W*in
   wire signed [9:0] m291_87;
   assign m291_87 =10'b0;

   // m291_88 = W*in
   wire signed [9:0] m291_88;
   assign m291_88 =10'b0;

   // m291_89 = W*in
   wire signed [9:0] m291_89;
   assign m291_89 =10'b0;

   // m291_90 = W*in
   wire signed [9:0] m291_90;
   assign m291_90 =10'b0;

   // m291_91 = W*in
   wire signed [9:0] m291_91;
   assign m291_91 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_92 = W*in
   wire signed [9:0] m291_92;
   assign m291_92 =10'b0;

   // m291_93 = W*in
   wire signed [9:0] m291_93;
   assign m291_93 =10'b0;

   // m291_94 = W*in
   wire signed [9:0] m291_94;
   assign m291_94 =10'b0;

   // m291_95 = W*in
   wire signed [9:0] m291_95;
   assign m291_95 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_96 = W*in
   wire signed [9:0] m291_96;
   assign m291_96 =10'b0;

   // m291_97 = W*in
   wire signed [9:0] m291_97;
   assign m291_97 =10'b0;

   // m291_98 = W*in
   wire signed [9:0] m291_98;
   assign m291_98 =10'b0;

   // m291_99 = W*in
   wire signed [9:0] m291_99;
   assign m291_99 ={ {4{neg291[5]}} , neg291[5:0] };

   // m291_100 = W*in
   wire signed [9:0] m291_100;
   assign m291_100 =10'b0;

   // m291_101 = W*in
   wire signed [9:0] m291_101;
   assign m291_101 =10'b0;

   // m291_102 = W*in
   wire signed [9:0] m291_102;
   assign m291_102 =10'b0;

   // m291_103 = W*in
   wire signed [9:0] m291_103;
   assign m291_103 =10'b0;

   // m291_104 = W*in
   wire signed [9:0] m291_104;
   assign m291_104 =10'b0;

   // m291_105 = W*in
   wire signed [9:0] m291_105;
   assign m291_105 =10'b0;

   // m291_106 = W*in
   wire signed [9:0] m291_106;
   assign m291_106 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_107 = W*in
   wire signed [9:0] m291_107;
   assign m291_107 =10'b0;

   // m291_108 = W*in
   wire signed [9:0] m291_108;
   assign m291_108 ={ {5{in291[5]}} , in291[5:1] };

   // m291_109 = W*in
   wire signed [9:0] m291_109;
   assign m291_109 ={ {5{in291[5]}} , in291[5:1] };

   // m291_110 = W*in
   wire signed [9:0] m291_110;
   assign m291_110 =10'b0;

   // m291_111 = W*in
   wire signed [9:0] m291_111;
   assign m291_111 =10'b0;

   // m291_112 = W*in
   wire signed [9:0] m291_112;
   assign m291_112 =10'b0;

   // m291_113 = W*in
   wire signed [9:0] m291_113;
   assign m291_113 =10'b0;

   // m291_114 = W*in
   wire signed [9:0] m291_114;
   assign m291_114 ={ {5{neg291[5]}} , neg291[5:1] };

   // m291_115 = W*in
   wire signed [9:0] m291_115;
   assign m291_115 =10'b0;

   // m291_116 = W*in
   wire signed [9:0] m291_116;
   assign m291_116 =10'b0;

   // m291_117 = W*in
   wire signed [9:0] m291_117;
   assign m291_117 =10'b0;

   // m292_1 = W*in
   wire signed [9:0] m292_1;
   assign m292_1 =10'b0;

   // m292_2 = W*in
   wire signed [9:0] m292_2;
   assign m292_2 =10'b0;

   // m292_3 = W*in
   wire signed [9:0] m292_3;
   assign m292_3 =10'b0;

   // m292_4 = W*in
   wire signed [9:0] m292_4;
   assign m292_4 =10'b0;

   // m292_5 = W*in
   wire signed [9:0] m292_5;
   assign m292_5 =10'b0;

   // m292_6 = W*in
   wire signed [9:0] m292_6;
   assign m292_6 =10'b0;

   // m292_7 = W*in
   wire signed [9:0] m292_7;
   assign m292_7 =10'b0;

   // m292_8 = W*in
   wire signed [9:0] m292_8;
   assign m292_8 =10'b0;

   // m292_9 = W*in
   wire signed [9:0] m292_9;
   assign m292_9 =10'b0;

   // m292_10 = W*in
   wire signed [9:0] m292_10;
   assign m292_10 =10'b0;

   // m292_11 = W*in
   wire signed [9:0] m292_11;
   assign m292_11 =10'b0;

   // m292_12 = W*in
   wire signed [9:0] m292_12;
   assign m292_12 =10'b0;

   // m292_13 = W*in
   wire signed [9:0] m292_13;
   assign m292_13 ={ {4{in292[5]}} , in292[5:0] };

   // m292_14 = W*in
   wire signed [9:0] m292_14;
   assign m292_14 =10'b0;

   // m292_15 = W*in
   wire signed [9:0] m292_15;
   assign m292_15 =10'b0;

   // m292_16 = W*in
   wire signed [9:0] m292_16;
   assign m292_16 =10'b0;

   // m292_17 = W*in
   wire signed [9:0] m292_17;
   assign m292_17 =10'b0;

   // m292_18 = W*in
   wire signed [9:0] m292_18;
   assign m292_18 =10'b0;

   // m292_19 = W*in
   wire signed [9:0] m292_19;
   assign m292_19 =10'b0;

   // m292_20 = W*in
   wire signed [9:0] m292_20;
   assign m292_20 =10'b0;

   // m292_21 = W*in
   wire signed [9:0] m292_21;
   assign m292_21 =10'b0;

   // m292_22 = W*in
   wire signed [9:0] m292_22;
   assign m292_22 =10'b0;

   // m292_23 = W*in
   wire signed [9:0] m292_23;
   assign m292_23 =10'b0;

   // m292_24 = W*in
   wire signed [9:0] m292_24;
   assign m292_24 =10'b0;

   // m292_25 = W*in
   wire signed [9:0] m292_25;
   assign m292_25 =10'b0;

   // m292_26 = W*in
   wire signed [9:0] m292_26;
   assign m292_26 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_27 = W*in
   wire signed [9:0] m292_27;
   assign m292_27 =10'b0;

   // m292_28 = W*in
   wire signed [9:0] m292_28;
   assign m292_28 =10'b0;

   // m292_29 = W*in
   wire signed [9:0] m292_29;
   assign m292_29 =10'b0;

   // m292_30 = W*in
   wire signed [9:0] m292_30;
   assign m292_30 =10'b0;

   // m292_31 = W*in
   wire signed [9:0] m292_31;
   assign m292_31 =10'b0;

   // m292_32 = W*in
   wire signed [9:0] m292_32;
   assign m292_32 =10'b0;

   // m292_33 = W*in
   wire signed [9:0] m292_33;
   assign m292_33 =10'b0;

   // m292_34 = W*in
   wire signed [9:0] m292_34;
   assign m292_34 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_35 = W*in
   wire signed [9:0] m292_35;
   assign m292_35 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_36 = W*in
   wire signed [9:0] m292_36;
   assign m292_36 =10'b0;

   // m292_37 = W*in
   wire signed [9:0] m292_37;
   assign m292_37 ={ {4{in292[5]}} , in292[5:0] };

   // m292_38 = W*in
   wire signed [9:0] m292_38;
   assign m292_38 ={ {4{neg292[5]}} , neg292[5:0] };

   // m292_39 = W*in
   wire signed [9:0] m292_39;
   assign m292_39 =10'b0;

   // m292_40 = W*in
   wire signed [9:0] m292_40;
   assign m292_40 =10'b0;

   // m292_41 = W*in
   wire signed [9:0] m292_41;
   assign m292_41 =10'b0;

   // m292_42 = W*in
   wire signed [9:0] m292_42;
   assign m292_42 =10'b0;

   // m292_43 = W*in
   wire signed [9:0] m292_43;
   assign m292_43 =10'b0;

   // m292_44 = W*in
   wire signed [9:0] m292_44;
   assign m292_44 =10'b0;

   // m292_45 = W*in
   wire signed [9:0] m292_45;
   assign m292_45 =10'b0;

   // m292_46 = W*in
   wire signed [9:0] m292_46;
   assign m292_46 =10'b0;

   // m292_47 = W*in
   wire signed [9:0] m292_47;
   assign m292_47 =10'b0;

   // m292_48 = W*in
   wire signed [9:0] m292_48;
   assign m292_48 =10'b0;

   // m292_49 = W*in
   wire signed [9:0] m292_49;
   assign m292_49 =10'b0;

   // m292_50 = W*in
   wire signed [9:0] m292_50;
   assign m292_50 =10'b0;

   // m292_51 = W*in
   wire signed [9:0] m292_51;
   assign m292_51 =10'b0;

   // m292_52 = W*in
   wire signed [9:0] m292_52;
   assign m292_52 =10'b0;

   // m292_53 = W*in
   wire signed [9:0] m292_53;
   assign m292_53 =10'b0;

   // m292_54 = W*in
   wire signed [9:0] m292_54;
   assign m292_54 =10'b0;

   // m292_55 = W*in
   wire signed [9:0] m292_55;
   assign m292_55 =10'b0;

   // m292_56 = W*in
   wire signed [9:0] m292_56;
   assign m292_56 =10'b0;

   // m292_57 = W*in
   wire signed [9:0] m292_57;
   assign m292_57 =10'b0;

   // m292_58 = W*in
   wire signed [9:0] m292_58;
   assign m292_58 =10'b0;

   // m292_59 = W*in
   wire signed [9:0] m292_59;
   assign m292_59 =10'b0;

   // m292_60 = W*in
   wire signed [9:0] m292_60;
   assign m292_60 =10'b0;

   // m292_61 = W*in
   wire signed [9:0] m292_61;
   assign m292_61 =10'b0;

   // m292_62 = W*in
   wire signed [9:0] m292_62;
   assign m292_62 =10'b0;

   // m292_63 = W*in
   wire signed [9:0] m292_63;
   assign m292_63 =10'b0;

   // m292_64 = W*in
   wire signed [9:0] m292_64;
   assign m292_64 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_65 = W*in
   wire signed [9:0] m292_65;
   assign m292_65 =10'b0;

   // m292_66 = W*in
   wire signed [9:0] m292_66;
   assign m292_66 =10'b0;

   // m292_67 = W*in
   wire signed [9:0] m292_67;
   assign m292_67 =10'b0;

   // m292_68 = W*in
   wire signed [9:0] m292_68;
   assign m292_68 =10'b0;

   // m292_69 = W*in
   wire signed [9:0] m292_69;
   assign m292_69 =10'b0;

   // m292_70 = W*in
   wire signed [9:0] m292_70;
   assign m292_70 =10'b0;

   // m292_71 = W*in
   wire signed [9:0] m292_71;
   assign m292_71 =10'b0;

   // m292_72 = W*in
   wire signed [9:0] m292_72;
   assign m292_72 =10'b0;

   // m292_73 = W*in
   wire signed [9:0] m292_73;
   assign m292_73 =10'b0;

   // m292_74 = W*in
   wire signed [9:0] m292_74;
   assign m292_74 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_75 = W*in
   wire signed [9:0] m292_75;
   assign m292_75 =10'b0;

   // m292_76 = W*in
   wire signed [9:0] m292_76;
   assign m292_76 =10'b0;

   // m292_77 = W*in
   wire signed [9:0] m292_77;
   assign m292_77 ={ {4{neg292[5]}} , neg292[5:0] };

   // m292_78 = W*in
   wire signed [9:0] m292_78;
   assign m292_78 =10'b0;

   // m292_79 = W*in
   wire signed [9:0] m292_79;
   assign m292_79 =10'b0;

   // m292_80 = W*in
   wire signed [9:0] m292_80;
   assign m292_80 =10'b0;

   // m292_81 = W*in
   wire signed [9:0] m292_81;
   assign m292_81 ={ {4{neg292[5]}} , neg292[5:0] };

   // m292_82 = W*in
   wire signed [9:0] m292_82;
   assign m292_82 =10'b0;

   // m292_83 = W*in
   wire signed [9:0] m292_83;
   assign m292_83 =10'b0;

   // m292_84 = W*in
   wire signed [9:0] m292_84;
   assign m292_84 =10'b0;

   // m292_85 = W*in
   wire signed [9:0] m292_85;
   assign m292_85 ={ {5{in292[5]}} , in292[5:1] };

   // m292_86 = W*in
   wire signed [9:0] m292_86;
   assign m292_86 =10'b0;

   // m292_87 = W*in
   wire signed [9:0] m292_87;
   assign m292_87 =10'b0;

   // m292_88 = W*in
   wire signed [9:0] m292_88;
   assign m292_88 =10'b0;

   // m292_89 = W*in
   wire signed [9:0] m292_89;
   assign m292_89 ={ {4{in292[5]}} , in292[5:0] };

   // m292_90 = W*in
   wire signed [9:0] m292_90;
   assign m292_90 =10'b0;

   // m292_91 = W*in
   wire signed [9:0] m292_91;
   assign m292_91 ={ {4{neg292[5]}} , neg292[5:0] };

   // m292_92 = W*in
   wire signed [9:0] m292_92;
   assign m292_92 =10'b0;

   // m292_93 = W*in
   wire signed [9:0] m292_93;
   assign m292_93 =10'b0;

   // m292_94 = W*in
   wire signed [9:0] m292_94;
   assign m292_94 =10'b0;

   // m292_95 = W*in
   wire signed [9:0] m292_95;
   assign m292_95 =10'b0;

   // m292_96 = W*in
   wire signed [9:0] m292_96;
   assign m292_96 =10'b0;

   // m292_97 = W*in
   wire signed [9:0] m292_97;
   assign m292_97 ={ {4{neg292[5]}} , neg292[5:0] };

   // m292_98 = W*in
   wire signed [9:0] m292_98;
   assign m292_98 =10'b0;

   // m292_99 = W*in
   wire signed [9:0] m292_99;
   assign m292_99 =10'b0;

   // m292_100 = W*in
   wire signed [9:0] m292_100;
   assign m292_100 =10'b0;

   // m292_101 = W*in
   wire signed [9:0] m292_101;
   assign m292_101 =10'b0;

   // m292_102 = W*in
   wire signed [9:0] m292_102;
   assign m292_102 =10'b0;

   // m292_103 = W*in
   wire signed [9:0] m292_103;
   assign m292_103 =10'b0;

   // m292_104 = W*in
   wire signed [9:0] m292_104;
   assign m292_104 =10'b0;

   // m292_105 = W*in
   wire signed [9:0] m292_105;
   assign m292_105 =10'b0;

   // m292_106 = W*in
   wire signed [9:0] m292_106;
   assign m292_106 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_107 = W*in
   wire signed [9:0] m292_107;
   assign m292_107 =10'b0;

   // m292_108 = W*in
   wire signed [9:0] m292_108;
   assign m292_108 ={ {5{in292[5]}} , in292[5:1] };

   // m292_109 = W*in
   wire signed [9:0] m292_109;
   assign m292_109 ={ {4{in292[5]}} , in292[5:0] };

   // m292_110 = W*in
   wire signed [9:0] m292_110;
   assign m292_110 =10'b0;

   // m292_111 = W*in
   wire signed [9:0] m292_111;
   assign m292_111 =10'b0;

   // m292_112 = W*in
   wire signed [9:0] m292_112;
   assign m292_112 =10'b0;

   // m292_113 = W*in
   wire signed [9:0] m292_113;
   assign m292_113 =10'b0;

   // m292_114 = W*in
   wire signed [9:0] m292_114;
   assign m292_114 =10'b0;

   // m292_115 = W*in
   wire signed [9:0] m292_115;
   assign m292_115 ={ {5{neg292[5]}} , neg292[5:1] };

   // m292_116 = W*in
   wire signed [9:0] m292_116;
   assign m292_116 =10'b0;

   // m292_117 = W*in
   wire signed [9:0] m292_117;
   assign m292_117 =10'b0;

   // m293_1 = W*in
   wire signed [9:0] m293_1;
   assign m293_1 =10'b0;

   // m293_2 = W*in
   wire signed [9:0] m293_2;
   assign m293_2 =10'b0;

   // m293_3 = W*in
   wire signed [9:0] m293_3;
   assign m293_3 =10'b0;

   // m293_4 = W*in
   wire signed [9:0] m293_4;
   assign m293_4 =10'b0;

   // m293_5 = W*in
   wire signed [9:0] m293_5;
   assign m293_5 =10'b0;

   // m293_6 = W*in
   wire signed [9:0] m293_6;
   assign m293_6 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_7 = W*in
   wire signed [9:0] m293_7;
   assign m293_7 =10'b0;

   // m293_8 = W*in
   wire signed [9:0] m293_8;
   assign m293_8 =10'b0;

   // m293_9 = W*in
   wire signed [9:0] m293_9;
   assign m293_9 =10'b0;

   // m293_10 = W*in
   wire signed [9:0] m293_10;
   assign m293_10 =10'b0;

   // m293_11 = W*in
   wire signed [9:0] m293_11;
   assign m293_11 =10'b0;

   // m293_12 = W*in
   wire signed [9:0] m293_12;
   assign m293_12 =10'b0;

   // m293_13 = W*in
   wire signed [9:0] m293_13;
   assign m293_13 ={ {4{in293[5]}} , in293[5:0] };

   // m293_14 = W*in
   wire signed [9:0] m293_14;
   assign m293_14 =10'b0;

   // m293_15 = W*in
   wire signed [9:0] m293_15;
   assign m293_15 =10'b0;

   // m293_16 = W*in
   wire signed [9:0] m293_16;
   assign m293_16 =10'b0;

   // m293_17 = W*in
   wire signed [9:0] m293_17;
   assign m293_17 =10'b0;

   // m293_18 = W*in
   wire signed [9:0] m293_18;
   assign m293_18 ={ {5{neg293[5]}} , neg293[5:1] };

   // m293_19 = W*in
   wire signed [9:0] m293_19;
   assign m293_19 ={ {5{neg293[5]}} , neg293[5:1] };

   // m293_20 = W*in
   wire signed [9:0] m293_20;
   assign m293_20 =10'b0;

   // m293_21 = W*in
   wire signed [9:0] m293_21;
   assign m293_21 =10'b0;

   // m293_22 = W*in
   wire signed [9:0] m293_22;
   assign m293_22 =10'b0;

   // m293_23 = W*in
   wire signed [9:0] m293_23;
   assign m293_23 =10'b0;

   // m293_24 = W*in
   wire signed [9:0] m293_24;
   assign m293_24 =10'b0;

   // m293_25 = W*in
   wire signed [9:0] m293_25;
   assign m293_25 =10'b0;

   // m293_26 = W*in
   wire signed [9:0] m293_26;
   assign m293_26 ={ {5{neg293[5]}} , neg293[5:1] };

   // m293_27 = W*in
   wire signed [9:0] m293_27;
   assign m293_27 =10'b0;

   // m293_28 = W*in
   wire signed [9:0] m293_28;
   assign m293_28 =10'b0;

   // m293_29 = W*in
   wire signed [9:0] m293_29;
   assign m293_29 =10'b0;

   // m293_30 = W*in
   wire signed [9:0] m293_30;
   assign m293_30 =10'b0;

   // m293_31 = W*in
   wire signed [9:0] m293_31;
   assign m293_31 =10'b0;

   // m293_32 = W*in
   wire signed [9:0] m293_32;
   assign m293_32 =10'b0;

   // m293_33 = W*in
   wire signed [9:0] m293_33;
   assign m293_33 =10'b0;

   // m293_34 = W*in
   wire signed [9:0] m293_34;
   assign m293_34 =10'b0;

   // m293_35 = W*in
   wire signed [9:0] m293_35;
   assign m293_35 =10'b0;

   // m293_36 = W*in
   wire signed [9:0] m293_36;
   assign m293_36 =10'b0;

   // m293_37 = W*in
   wire signed [9:0] m293_37;
   assign m293_37 =10'b0;

   // m293_38 = W*in
   wire signed [9:0] m293_38;
   assign m293_38 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_39 = W*in
   wire signed [9:0] m293_39;
   assign m293_39 =10'b0;

   // m293_40 = W*in
   wire signed [9:0] m293_40;
   assign m293_40 =10'b0;

   // m293_41 = W*in
   wire signed [9:0] m293_41;
   assign m293_41 ={ {4{in293[5]}} , in293[5:0] };

   // m293_42 = W*in
   wire signed [9:0] m293_42;
   assign m293_42 =10'b0;

   // m293_43 = W*in
   wire signed [9:0] m293_43;
   assign m293_43 =10'b0;

   // m293_44 = W*in
   wire signed [9:0] m293_44;
   assign m293_44 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_45 = W*in
   wire signed [9:0] m293_45;
   assign m293_45 =10'b0;

   // m293_46 = W*in
   wire signed [9:0] m293_46;
   assign m293_46 =10'b0;

   // m293_47 = W*in
   wire signed [9:0] m293_47;
   assign m293_47 =10'b0;

   // m293_48 = W*in
   wire signed [9:0] m293_48;
   assign m293_48 =10'b0;

   // m293_49 = W*in
   wire signed [9:0] m293_49;
   assign m293_49 =10'b0;

   // m293_50 = W*in
   wire signed [9:0] m293_50;
   assign m293_50 =10'b0;

   // m293_51 = W*in
   wire signed [9:0] m293_51;
   assign m293_51 =10'b0;

   // m293_52 = W*in
   wire signed [9:0] m293_52;
   assign m293_52 =10'b0;

   // m293_53 = W*in
   wire signed [9:0] m293_53;
   assign m293_53 =10'b0;

   // m293_54 = W*in
   wire signed [9:0] m293_54;
   assign m293_54 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_55 = W*in
   wire signed [9:0] m293_55;
   assign m293_55 =10'b0;

   // m293_56 = W*in
   wire signed [9:0] m293_56;
   assign m293_56 =10'b0;

   // m293_57 = W*in
   wire signed [9:0] m293_57;
   assign m293_57 =10'b0;

   // m293_58 = W*in
   wire signed [9:0] m293_58;
   assign m293_58 =10'b0;

   // m293_59 = W*in
   wire signed [9:0] m293_59;
   assign m293_59 =10'b0;

   // m293_60 = W*in
   wire signed [9:0] m293_60;
   assign m293_60 =10'b0;

   // m293_61 = W*in
   wire signed [9:0] m293_61;
   assign m293_61 =10'b0;

   // m293_62 = W*in
   wire signed [9:0] m293_62;
   assign m293_62 =10'b0;

   // m293_63 = W*in
   wire signed [9:0] m293_63;
   assign m293_63 =10'b0;

   // m293_64 = W*in
   wire signed [9:0] m293_64;
   assign m293_64 =10'b0;

   // m293_65 = W*in
   wire signed [9:0] m293_65;
   assign m293_65 ={ {5{in293[5]}} , in293[5:1] };

   // m293_66 = W*in
   wire signed [9:0] m293_66;
   assign m293_66 ={ {5{in293[5]}} , in293[5:1] };

   // m293_67 = W*in
   wire signed [9:0] m293_67;
   assign m293_67 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_68 = W*in
   wire signed [9:0] m293_68;
   assign m293_68 =10'b0;

   // m293_69 = W*in
   wire signed [9:0] m293_69;
   assign m293_69 =10'b0;

   // m293_70 = W*in
   wire signed [9:0] m293_70;
   assign m293_70 =10'b0;

   // m293_71 = W*in
   wire signed [9:0] m293_71;
   assign m293_71 =10'b0;

   // m293_72 = W*in
   wire signed [9:0] m293_72;
   assign m293_72 =10'b0;

   // m293_73 = W*in
   wire signed [9:0] m293_73;
   assign m293_73 =10'b0;

   // m293_74 = W*in
   wire signed [9:0] m293_74;
   assign m293_74 =10'b0;

   // m293_75 = W*in
   wire signed [9:0] m293_75;
   assign m293_75 =10'b0;

   // m293_76 = W*in
   wire signed [9:0] m293_76;
   assign m293_76 =10'b0;

   // m293_77 = W*in
   wire signed [9:0] m293_77;
   assign m293_77 =10'b0;

   // m293_78 = W*in
   wire signed [9:0] m293_78;
   assign m293_78 =10'b0;

   // m293_79 = W*in
   wire signed [9:0] m293_79;
   assign m293_79 =10'b0;

   // m293_80 = W*in
   wire signed [9:0] m293_80;
   assign m293_80 =10'b0;

   // m293_81 = W*in
   wire signed [9:0] m293_81;
   assign m293_81 =10'b0;

   // m293_82 = W*in
   wire signed [9:0] m293_82;
   assign m293_82 =10'b0;

   // m293_83 = W*in
   wire signed [9:0] m293_83;
   assign m293_83 =10'b0;

   // m293_84 = W*in
   wire signed [9:0] m293_84;
   assign m293_84 =10'b0;

   // m293_85 = W*in
   wire signed [9:0] m293_85;
   assign m293_85 =10'b0;

   // m293_86 = W*in
   wire signed [9:0] m293_86;
   assign m293_86 =10'b0;

   // m293_87 = W*in
   wire signed [9:0] m293_87;
   assign m293_87 =10'b0;

   // m293_88 = W*in
   wire signed [9:0] m293_88;
   assign m293_88 =10'b0;

   // m293_89 = W*in
   wire signed [9:0] m293_89;
   assign m293_89 =10'b0;

   // m293_90 = W*in
   wire signed [9:0] m293_90;
   assign m293_90 =10'b0;

   // m293_91 = W*in
   wire signed [9:0] m293_91;
   assign m293_91 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_92 = W*in
   wire signed [9:0] m293_92;
   assign m293_92 =10'b0;

   // m293_93 = W*in
   wire signed [9:0] m293_93;
   assign m293_93 =10'b0;

   // m293_94 = W*in
   wire signed [9:0] m293_94;
   assign m293_94 =10'b0;

   // m293_95 = W*in
   wire signed [9:0] m293_95;
   assign m293_95 =10'b0;

   // m293_96 = W*in
   wire signed [9:0] m293_96;
   assign m293_96 =10'b0;

   // m293_97 = W*in
   wire signed [9:0] m293_97;
   assign m293_97 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_98 = W*in
   wire signed [9:0] m293_98;
   assign m293_98 =10'b0;

   // m293_99 = W*in
   wire signed [9:0] m293_99;
   assign m293_99 =10'b0;

   // m293_100 = W*in
   wire signed [9:0] m293_100;
   assign m293_100 =10'b0;

   // m293_101 = W*in
   wire signed [9:0] m293_101;
   assign m293_101 =10'b0;

   // m293_102 = W*in
   wire signed [9:0] m293_102;
   assign m293_102 =10'b0;

   // m293_103 = W*in
   wire signed [9:0] m293_103;
   assign m293_103 =10'b0;

   // m293_104 = W*in
   wire signed [9:0] m293_104;
   assign m293_104 =10'b0;

   // m293_105 = W*in
   wire signed [9:0] m293_105;
   assign m293_105 =10'b0;

   // m293_106 = W*in
   wire signed [9:0] m293_106;
   assign m293_106 =10'b0;

   // m293_107 = W*in
   wire signed [9:0] m293_107;
   assign m293_107 =10'b0;

   // m293_108 = W*in
   wire signed [9:0] m293_108;
   assign m293_108 ={ {5{in293[5]}} , in293[5:1] };

   // m293_109 = W*in
   wire signed [9:0] m293_109;
   assign m293_109 ={ {5{in293[5]}} , in293[5:1] };

   // m293_110 = W*in
   wire signed [9:0] m293_110;
   assign m293_110 ={ {4{neg293[5]}} , neg293[5:0] };

   // m293_111 = W*in
   wire signed [9:0] m293_111;
   assign m293_111 =10'b0;

   // m293_112 = W*in
   wire signed [9:0] m293_112;
   assign m293_112 =10'b0;

   // m293_113 = W*in
   wire signed [9:0] m293_113;
   assign m293_113 =10'b0;

   // m293_114 = W*in
   wire signed [9:0] m293_114;
   assign m293_114 =10'b0;

   // m293_115 = W*in
   wire signed [9:0] m293_115;
   assign m293_115 =10'b0;

   // m293_116 = W*in
   wire signed [9:0] m293_116;
   assign m293_116 ={ {4{in293[5]}} , in293[5:0] };

   // m293_117 = W*in
   wire signed [9:0] m293_117;
   assign m293_117 =10'b0;

   // m294_1 = W*in
   wire signed [9:0] m294_1;
   assign m294_1 =10'b0;

   // m294_2 = W*in
   wire signed [9:0] m294_2;
   assign m294_2 =10'b0;

   // m294_3 = W*in
   wire signed [9:0] m294_3;
   assign m294_3 =10'b0;

   // m294_4 = W*in
   wire signed [9:0] m294_4;
   assign m294_4 =10'b0;

   // m294_5 = W*in
   wire signed [9:0] m294_5;
   assign m294_5 =10'b0;

   // m294_6 = W*in
   wire signed [9:0] m294_6;
   assign m294_6 =10'b0;

   // m294_7 = W*in
   wire signed [9:0] m294_7;
   assign m294_7 =10'b0;

   // m294_8 = W*in
   wire signed [9:0] m294_8;
   assign m294_8 =10'b0;

   // m294_9 = W*in
   wire signed [9:0] m294_9;
   assign m294_9 =10'b0;

   // m294_10 = W*in
   wire signed [9:0] m294_10;
   assign m294_10 =10'b0;

   // m294_11 = W*in
   wire signed [9:0] m294_11;
   assign m294_11 =10'b0;

   // m294_12 = W*in
   wire signed [9:0] m294_12;
   assign m294_12 =10'b0;

   // m294_13 = W*in
   wire signed [9:0] m294_13;
   assign m294_13 =10'b0;

   // m294_14 = W*in
   wire signed [9:0] m294_14;
   assign m294_14 =10'b0;

   // m294_15 = W*in
   wire signed [9:0] m294_15;
   assign m294_15 =10'b0;

   // m294_16 = W*in
   wire signed [9:0] m294_16;
   assign m294_16 =10'b0;

   // m294_17 = W*in
   wire signed [9:0] m294_17;
   assign m294_17 ={ {5{in294[5]}} , in294[5:1] };

   // m294_18 = W*in
   wire signed [9:0] m294_18;
   assign m294_18 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_19 = W*in
   wire signed [9:0] m294_19;
   assign m294_19 ={ {4{in294[5]}} , in294[5:0] };

   // m294_20 = W*in
   wire signed [9:0] m294_20;
   assign m294_20 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_21 = W*in
   wire signed [9:0] m294_21;
   assign m294_21 =10'b0;

   // m294_22 = W*in
   wire signed [9:0] m294_22;
   assign m294_22 =10'b0;

   // m294_23 = W*in
   wire signed [9:0] m294_23;
   assign m294_23 =10'b0;

   // m294_24 = W*in
   wire signed [9:0] m294_24;
   assign m294_24 =10'b0;

   // m294_25 = W*in
   wire signed [9:0] m294_25;
   assign m294_25 =10'b0;

   // m294_26 = W*in
   wire signed [9:0] m294_26;
   assign m294_26 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_27 = W*in
   wire signed [9:0] m294_27;
   assign m294_27 =10'b0;

   // m294_28 = W*in
   wire signed [9:0] m294_28;
   assign m294_28 =10'b0;

   // m294_29 = W*in
   wire signed [9:0] m294_29;
   assign m294_29 =10'b0;

   // m294_30 = W*in
   wire signed [9:0] m294_30;
   assign m294_30 =10'b0;

   // m294_31 = W*in
   wire signed [9:0] m294_31;
   assign m294_31 =10'b0;

   // m294_32 = W*in
   wire signed [9:0] m294_32;
   assign m294_32 =10'b0;

   // m294_33 = W*in
   wire signed [9:0] m294_33;
   assign m294_33 =10'b0;

   // m294_34 = W*in
   wire signed [9:0] m294_34;
   assign m294_34 =10'b0;

   // m294_35 = W*in
   wire signed [9:0] m294_35;
   assign m294_35 =10'b0;

   // m294_36 = W*in
   wire signed [9:0] m294_36;
   assign m294_36 =10'b0;

   // m294_37 = W*in
   wire signed [9:0] m294_37;
   assign m294_37 =10'b0;

   // m294_38 = W*in
   wire signed [9:0] m294_38;
   assign m294_38 =10'b0;

   // m294_39 = W*in
   wire signed [9:0] m294_39;
   assign m294_39 =10'b0;

   // m294_40 = W*in
   wire signed [9:0] m294_40;
   assign m294_40 =10'b0;

   // m294_41 = W*in
   wire signed [9:0] m294_41;
   assign m294_41 =10'b0;

   // m294_42 = W*in
   wire signed [9:0] m294_42;
   assign m294_42 =10'b0;

   // m294_43 = W*in
   wire signed [9:0] m294_43;
   assign m294_43 =10'b0;

   // m294_44 = W*in
   wire signed [9:0] m294_44;
   assign m294_44 =10'b0;

   // m294_45 = W*in
   wire signed [9:0] m294_45;
   assign m294_45 =10'b0;

   // m294_46 = W*in
   wire signed [9:0] m294_46;
   assign m294_46 =10'b0;

   // m294_47 = W*in
   wire signed [9:0] m294_47;
   assign m294_47 =10'b0;

   // m294_48 = W*in
   wire signed [9:0] m294_48;
   assign m294_48 =10'b0;

   // m294_49 = W*in
   wire signed [9:0] m294_49;
   assign m294_49 =10'b0;

   // m294_50 = W*in
   wire signed [9:0] m294_50;
   assign m294_50 =10'b0;

   // m294_51 = W*in
   wire signed [9:0] m294_51;
   assign m294_51 =10'b0;

   // m294_52 = W*in
   wire signed [9:0] m294_52;
   assign m294_52 =10'b0;

   // m294_53 = W*in
   wire signed [9:0] m294_53;
   assign m294_53 ={ {4{in294[5]}} , in294[5:0] };

   // m294_54 = W*in
   wire signed [9:0] m294_54;
   assign m294_54 =10'b0;

   // m294_55 = W*in
   wire signed [9:0] m294_55;
   assign m294_55 =10'b0;

   // m294_56 = W*in
   wire signed [9:0] m294_56;
   assign m294_56 =10'b0;

   // m294_57 = W*in
   wire signed [9:0] m294_57;
   assign m294_57 =10'b0;

   // m294_58 = W*in
   wire signed [9:0] m294_58;
   assign m294_58 =10'b0;

   // m294_59 = W*in
   wire signed [9:0] m294_59;
   assign m294_59 =10'b0;

   // m294_60 = W*in
   wire signed [9:0] m294_60;
   assign m294_60 =10'b0;

   // m294_61 = W*in
   wire signed [9:0] m294_61;
   assign m294_61 =10'b0;

   // m294_62 = W*in
   wire signed [9:0] m294_62;
   assign m294_62 =10'b0;

   // m294_63 = W*in
   wire signed [9:0] m294_63;
   assign m294_63 =10'b0;

   // m294_64 = W*in
   wire signed [9:0] m294_64;
   assign m294_64 =10'b0;

   // m294_65 = W*in
   wire signed [9:0] m294_65;
   assign m294_65 ={ {5{in294[5]}} , in294[5:1] };

   // m294_66 = W*in
   wire signed [9:0] m294_66;
   assign m294_66 ={ {5{in294[5]}} , in294[5:1] };

   // m294_67 = W*in
   wire signed [9:0] m294_67;
   assign m294_67 ={ {4{in294[5]}} , in294[5:0] };

   // m294_68 = W*in
   wire signed [9:0] m294_68;
   assign m294_68 =10'b0;

   // m294_69 = W*in
   wire signed [9:0] m294_69;
   assign m294_69 =10'b0;

   // m294_70 = W*in
   wire signed [9:0] m294_70;
   assign m294_70 =10'b0;

   // m294_71 = W*in
   wire signed [9:0] m294_71;
   assign m294_71 =10'b0;

   // m294_72 = W*in
   wire signed [9:0] m294_72;
   assign m294_72 ={ {4{neg294[5]}} , neg294[5:0] };

   // m294_73 = W*in
   wire signed [9:0] m294_73;
   assign m294_73 ={ {5{in294[5]}} , in294[5:1] };

   // m294_74 = W*in
   wire signed [9:0] m294_74;
   assign m294_74 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_75 = W*in
   wire signed [9:0] m294_75;
   assign m294_75 =10'b0;

   // m294_76 = W*in
   wire signed [9:0] m294_76;
   assign m294_76 =10'b0;

   // m294_77 = W*in
   wire signed [9:0] m294_77;
   assign m294_77 =10'b0;

   // m294_78 = W*in
   wire signed [9:0] m294_78;
   assign m294_78 =10'b0;

   // m294_79 = W*in
   wire signed [9:0] m294_79;
   assign m294_79 =10'b0;

   // m294_80 = W*in
   wire signed [9:0] m294_80;
   assign m294_80 =10'b0;

   // m294_81 = W*in
   wire signed [9:0] m294_81;
   assign m294_81 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_82 = W*in
   wire signed [9:0] m294_82;
   assign m294_82 =10'b0;

   // m294_83 = W*in
   wire signed [9:0] m294_83;
   assign m294_83 =10'b0;

   // m294_84 = W*in
   wire signed [9:0] m294_84;
   assign m294_84 ={ {4{neg294[5]}} , neg294[5:0] };

   // m294_85 = W*in
   wire signed [9:0] m294_85;
   assign m294_85 =10'b0;

   // m294_86 = W*in
   wire signed [9:0] m294_86;
   assign m294_86 =10'b0;

   // m294_87 = W*in
   wire signed [9:0] m294_87;
   assign m294_87 =10'b0;

   // m294_88 = W*in
   wire signed [9:0] m294_88;
   assign m294_88 =10'b0;

   // m294_89 = W*in
   wire signed [9:0] m294_89;
   assign m294_89 =10'b0;

   // m294_90 = W*in
   wire signed [9:0] m294_90;
   assign m294_90 =10'b0;

   // m294_91 = W*in
   wire signed [9:0] m294_91;
   assign m294_91 =10'b0;

   // m294_92 = W*in
   wire signed [9:0] m294_92;
   assign m294_92 =10'b0;

   // m294_93 = W*in
   wire signed [9:0] m294_93;
   assign m294_93 ={ {4{in294[5]}} , in294[5:0] };

   // m294_94 = W*in
   wire signed [9:0] m294_94;
   assign m294_94 =10'b0;

   // m294_95 = W*in
   wire signed [9:0] m294_95;
   assign m294_95 =10'b0;

   // m294_96 = W*in
   wire signed [9:0] m294_96;
   assign m294_96 =10'b0;

   // m294_97 = W*in
   wire signed [9:0] m294_97;
   assign m294_97 =10'b0;

   // m294_98 = W*in
   wire signed [9:0] m294_98;
   assign m294_98 =10'b0;

   // m294_99 = W*in
   wire signed [9:0] m294_99;
   assign m294_99 =10'b0;

   // m294_100 = W*in
   wire signed [9:0] m294_100;
   assign m294_100 =10'b0;

   // m294_101 = W*in
   wire signed [9:0] m294_101;
   assign m294_101 =10'b0;

   // m294_102 = W*in
   wire signed [9:0] m294_102;
   assign m294_102 =10'b0;

   // m294_103 = W*in
   wire signed [9:0] m294_103;
   assign m294_103 =10'b0;

   // m294_104 = W*in
   wire signed [9:0] m294_104;
   assign m294_104 =10'b0;

   // m294_105 = W*in
   wire signed [9:0] m294_105;
   assign m294_105 =10'b0;

   // m294_106 = W*in
   wire signed [9:0] m294_106;
   assign m294_106 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_107 = W*in
   wire signed [9:0] m294_107;
   assign m294_107 =10'b0;

   // m294_108 = W*in
   wire signed [9:0] m294_108;
   assign m294_108 =10'b0;

   // m294_109 = W*in
   wire signed [9:0] m294_109;
   assign m294_109 ={ {5{in294[5]}} , in294[5:1] };

   // m294_110 = W*in
   wire signed [9:0] m294_110;
   assign m294_110 =10'b0;

   // m294_111 = W*in
   wire signed [9:0] m294_111;
   assign m294_111 =10'b0;

   // m294_112 = W*in
   wire signed [9:0] m294_112;
   assign m294_112 =10'b0;

   // m294_113 = W*in
   wire signed [9:0] m294_113;
   assign m294_113 ={ {4{neg294[5]}} , neg294[5:0] };

   // m294_114 = W*in
   wire signed [9:0] m294_114;
   assign m294_114 =10'b0;

   // m294_115 = W*in
   wire signed [9:0] m294_115;
   assign m294_115 ={ {5{neg294[5]}} , neg294[5:1] };

   // m294_116 = W*in
   wire signed [9:0] m294_116;
   assign m294_116 =10'b0;

   // m294_117 = W*in
   wire signed [9:0] m294_117;
   assign m294_117 =10'b0;

   // m295_1 = W*in
   wire signed [9:0] m295_1;
   assign m295_1 =10'b0;

   // m295_2 = W*in
   wire signed [9:0] m295_2;
   assign m295_2 =10'b0;

   // m295_3 = W*in
   wire signed [9:0] m295_3;
   assign m295_3 =10'b0;

   // m295_4 = W*in
   wire signed [9:0] m295_4;
   assign m295_4 =10'b0;

   // m295_5 = W*in
   wire signed [9:0] m295_5;
   assign m295_5 =10'b0;

   // m295_6 = W*in
   wire signed [9:0] m295_6;
   assign m295_6 =10'b0;

   // m295_7 = W*in
   wire signed [9:0] m295_7;
   assign m295_7 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_8 = W*in
   wire signed [9:0] m295_8;
   assign m295_8 =10'b0;

   // m295_9 = W*in
   wire signed [9:0] m295_9;
   assign m295_9 =10'b0;

   // m295_10 = W*in
   wire signed [9:0] m295_10;
   assign m295_10 =10'b0;

   // m295_11 = W*in
   wire signed [9:0] m295_11;
   assign m295_11 =10'b0;

   // m295_12 = W*in
   wire signed [9:0] m295_12;
   assign m295_12 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_13 = W*in
   wire signed [9:0] m295_13;
   assign m295_13 =10'b0;

   // m295_14 = W*in
   wire signed [9:0] m295_14;
   assign m295_14 =10'b0;

   // m295_15 = W*in
   wire signed [9:0] m295_15;
   assign m295_15 =10'b0;

   // m295_16 = W*in
   wire signed [9:0] m295_16;
   assign m295_16 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_17 = W*in
   wire signed [9:0] m295_17;
   assign m295_17 ={ {5{in295[5]}} , in295[5:1] };

   // m295_18 = W*in
   wire signed [9:0] m295_18;
   assign m295_18 =10'b0;

   // m295_19 = W*in
   wire signed [9:0] m295_19;
   assign m295_19 =10'b0;

   // m295_20 = W*in
   wire signed [9:0] m295_20;
   assign m295_20 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_21 = W*in
   wire signed [9:0] m295_21;
   assign m295_21 =10'b0;

   // m295_22 = W*in
   wire signed [9:0] m295_22;
   assign m295_22 =10'b0;

   // m295_23 = W*in
   wire signed [9:0] m295_23;
   assign m295_23 =10'b0;

   // m295_24 = W*in
   wire signed [9:0] m295_24;
   assign m295_24 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_25 = W*in
   wire signed [9:0] m295_25;
   assign m295_25 =10'b0;

   // m295_26 = W*in
   wire signed [9:0] m295_26;
   assign m295_26 =10'b0;

   // m295_27 = W*in
   wire signed [9:0] m295_27;
   assign m295_27 =10'b0;

   // m295_28 = W*in
   wire signed [9:0] m295_28;
   assign m295_28 =10'b0;

   // m295_29 = W*in
   wire signed [9:0] m295_29;
   assign m295_29 =10'b0;

   // m295_30 = W*in
   wire signed [9:0] m295_30;
   assign m295_30 =10'b0;

   // m295_31 = W*in
   wire signed [9:0] m295_31;
   assign m295_31 =10'b0;

   // m295_32 = W*in
   wire signed [9:0] m295_32;
   assign m295_32 =10'b0;

   // m295_33 = W*in
   wire signed [9:0] m295_33;
   assign m295_33 =10'b0;

   // m295_34 = W*in
   wire signed [9:0] m295_34;
   assign m295_34 =10'b0;

   // m295_35 = W*in
   wire signed [9:0] m295_35;
   assign m295_35 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_36 = W*in
   wire signed [9:0] m295_36;
   assign m295_36 =10'b0;

   // m295_37 = W*in
   wire signed [9:0] m295_37;
   assign m295_37 =10'b0;

   // m295_38 = W*in
   wire signed [9:0] m295_38;
   assign m295_38 =10'b0;

   // m295_39 = W*in
   wire signed [9:0] m295_39;
   assign m295_39 =10'b0;

   // m295_40 = W*in
   wire signed [9:0] m295_40;
   assign m295_40 =10'b0;

   // m295_41 = W*in
   wire signed [9:0] m295_41;
   assign m295_41 =10'b0;

   // m295_42 = W*in
   wire signed [9:0] m295_42;
   assign m295_42 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_43 = W*in
   wire signed [9:0] m295_43;
   assign m295_43 =10'b0;

   // m295_44 = W*in
   wire signed [9:0] m295_44;
   assign m295_44 =10'b0;

   // m295_45 = W*in
   wire signed [9:0] m295_45;
   assign m295_45 =10'b0;

   // m295_46 = W*in
   wire signed [9:0] m295_46;
   assign m295_46 =10'b0;

   // m295_47 = W*in
   wire signed [9:0] m295_47;
   assign m295_47 =10'b0;

   // m295_48 = W*in
   wire signed [9:0] m295_48;
   assign m295_48 =10'b0;

   // m295_49 = W*in
   wire signed [9:0] m295_49;
   assign m295_49 =10'b0;

   // m295_50 = W*in
   wire signed [9:0] m295_50;
   assign m295_50 ={ {4{in295[5]}} , in295[5:0] };

   // m295_51 = W*in
   wire signed [9:0] m295_51;
   assign m295_51 =10'b0;

   // m295_52 = W*in
   wire signed [9:0] m295_52;
   assign m295_52 =10'b0;

   // m295_53 = W*in
   wire signed [9:0] m295_53;
   assign m295_53 =10'b0;

   // m295_54 = W*in
   wire signed [9:0] m295_54;
   assign m295_54 =10'b0;

   // m295_55 = W*in
   wire signed [9:0] m295_55;
   assign m295_55 =10'b0;

   // m295_56 = W*in
   wire signed [9:0] m295_56;
   assign m295_56 =10'b0;

   // m295_57 = W*in
   wire signed [9:0] m295_57;
   assign m295_57 =10'b0;

   // m295_58 = W*in
   wire signed [9:0] m295_58;
   assign m295_58 =10'b0;

   // m295_59 = W*in
   wire signed [9:0] m295_59;
   assign m295_59 =10'b0;

   // m295_60 = W*in
   wire signed [9:0] m295_60;
   assign m295_60 =10'b0;

   // m295_61 = W*in
   wire signed [9:0] m295_61;
   assign m295_61 =10'b0;

   // m295_62 = W*in
   wire signed [9:0] m295_62;
   assign m295_62 =10'b0;

   // m295_63 = W*in
   wire signed [9:0] m295_63;
   assign m295_63 ={ {4{in295[5]}} , in295[5:0] };

   // m295_64 = W*in
   wire signed [9:0] m295_64;
   assign m295_64 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_65 = W*in
   wire signed [9:0] m295_65;
   assign m295_65 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_66 = W*in
   wire signed [9:0] m295_66;
   assign m295_66 =10'b0;

   // m295_67 = W*in
   wire signed [9:0] m295_67;
   assign m295_67 =10'b0;

   // m295_68 = W*in
   wire signed [9:0] m295_68;
   assign m295_68 =10'b0;

   // m295_69 = W*in
   wire signed [9:0] m295_69;
   assign m295_69 ={ {5{in295[5]}} , in295[5:1] };

   // m295_70 = W*in
   wire signed [9:0] m295_70;
   assign m295_70 =10'b0;

   // m295_71 = W*in
   wire signed [9:0] m295_71;
   assign m295_71 ={ {5{in295[5]}} , in295[5:1] };

   // m295_72 = W*in
   wire signed [9:0] m295_72;
   assign m295_72 ={ {4{in295[5]}} , in295[5:0] };

   // m295_73 = W*in
   wire signed [9:0] m295_73;
   assign m295_73 =10'b0;

   // m295_74 = W*in
   wire signed [9:0] m295_74;
   assign m295_74 =10'b0;

   // m295_75 = W*in
   wire signed [9:0] m295_75;
   assign m295_75 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_76 = W*in
   wire signed [9:0] m295_76;
   assign m295_76 =10'b0;

   // m295_77 = W*in
   wire signed [9:0] m295_77;
   assign m295_77 =10'b0;

   // m295_78 = W*in
   wire signed [9:0] m295_78;
   assign m295_78 =10'b0;

   // m295_79 = W*in
   wire signed [9:0] m295_79;
   assign m295_79 =10'b0;

   // m295_80 = W*in
   wire signed [9:0] m295_80;
   assign m295_80 =10'b0;

   // m295_81 = W*in
   wire signed [9:0] m295_81;
   assign m295_81 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_82 = W*in
   wire signed [9:0] m295_82;
   assign m295_82 =10'b0;

   // m295_83 = W*in
   wire signed [9:0] m295_83;
   assign m295_83 =10'b0;

   // m295_84 = W*in
   wire signed [9:0] m295_84;
   assign m295_84 ={ {4{in295[5]}} , in295[5:0] };

   // m295_85 = W*in
   wire signed [9:0] m295_85;
   assign m295_85 =10'b0;

   // m295_86 = W*in
   wire signed [9:0] m295_86;
   assign m295_86 =10'b0;

   // m295_87 = W*in
   wire signed [9:0] m295_87;
   assign m295_87 ={ {4{in295[5]}} , in295[5:0] };

   // m295_88 = W*in
   wire signed [9:0] m295_88;
   assign m295_88 =10'b0;

   // m295_89 = W*in
   wire signed [9:0] m295_89;
   assign m295_89 =10'b0;

   // m295_90 = W*in
   wire signed [9:0] m295_90;
   assign m295_90 =10'b0;

   // m295_91 = W*in
   wire signed [9:0] m295_91;
   assign m295_91 =10'b0;

   // m295_92 = W*in
   wire signed [9:0] m295_92;
   assign m295_92 =10'b0;

   // m295_93 = W*in
   wire signed [9:0] m295_93;
   assign m295_93 =10'b0;

   // m295_94 = W*in
   wire signed [9:0] m295_94;
   assign m295_94 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_95 = W*in
   wire signed [9:0] m295_95;
   assign m295_95 =10'b0;

   // m295_96 = W*in
   wire signed [9:0] m295_96;
   assign m295_96 =10'b0;

   // m295_97 = W*in
   wire signed [9:0] m295_97;
   assign m295_97 =10'b0;

   // m295_98 = W*in
   wire signed [9:0] m295_98;
   assign m295_98 =10'b0;

   // m295_99 = W*in
   wire signed [9:0] m295_99;
   assign m295_99 =10'b0;

   // m295_100 = W*in
   wire signed [9:0] m295_100;
   assign m295_100 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_101 = W*in
   wire signed [9:0] m295_101;
   assign m295_101 =10'b0;

   // m295_102 = W*in
   wire signed [9:0] m295_102;
   assign m295_102 =10'b0;

   // m295_103 = W*in
   wire signed [9:0] m295_103;
   assign m295_103 =10'b0;

   // m295_104 = W*in
   wire signed [9:0] m295_104;
   assign m295_104 =10'b0;

   // m295_105 = W*in
   wire signed [9:0] m295_105;
   assign m295_105 =10'b0;

   // m295_106 = W*in
   wire signed [9:0] m295_106;
   assign m295_106 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_107 = W*in
   wire signed [9:0] m295_107;
   assign m295_107 =10'b0;

   // m295_108 = W*in
   wire signed [9:0] m295_108;
   assign m295_108 =10'b0;

   // m295_109 = W*in
   wire signed [9:0] m295_109;
   assign m295_109 =10'b0;

   // m295_110 = W*in
   wire signed [9:0] m295_110;
   assign m295_110 =10'b0;

   // m295_111 = W*in
   wire signed [9:0] m295_111;
   assign m295_111 =10'b0;

   // m295_112 = W*in
   wire signed [9:0] m295_112;
   assign m295_112 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_113 = W*in
   wire signed [9:0] m295_113;
   assign m295_113 ={ {4{neg295[5]}} , neg295[5:0] };

   // m295_114 = W*in
   wire signed [9:0] m295_114;
   assign m295_114 =10'b0;

   // m295_115 = W*in
   wire signed [9:0] m295_115;
   assign m295_115 ={ {5{neg295[5]}} , neg295[5:1] };

   // m295_116 = W*in
   wire signed [9:0] m295_116;
   assign m295_116 =10'b0;

   // m295_117 = W*in
   wire signed [9:0] m295_117;
   assign m295_117 =10'b0;

   // m296_1 = W*in
   wire signed [9:0] m296_1;
   assign m296_1 =10'b0;

   // m296_2 = W*in
   wire signed [9:0] m296_2;
   assign m296_2 =10'b0;

   // m296_3 = W*in
   wire signed [9:0] m296_3;
   assign m296_3 ={ {4{neg296[5]}} , neg296[5:0] };

   // m296_4 = W*in
   wire signed [9:0] m296_4;
   assign m296_4 =10'b0;

   // m296_5 = W*in
   wire signed [9:0] m296_5;
   assign m296_5 =10'b0;

   // m296_6 = W*in
   wire signed [9:0] m296_6;
   assign m296_6 =10'b0;

   // m296_7 = W*in
   wire signed [9:0] m296_7;
   assign m296_7 =10'b0;

   // m296_8 = W*in
   wire signed [9:0] m296_8;
   assign m296_8 =10'b0;

   // m296_9 = W*in
   wire signed [9:0] m296_9;
   assign m296_9 =10'b0;

   // m296_10 = W*in
   wire signed [9:0] m296_10;
   assign m296_10 ={ {4{in296[5]}} , in296[5:0] };

   // m296_11 = W*in
   wire signed [9:0] m296_11;
   assign m296_11 =10'b0;

   // m296_12 = W*in
   wire signed [9:0] m296_12;
   assign m296_12 ={ {4{neg296[5]}} , neg296[5:0] };

   // m296_13 = W*in
   wire signed [9:0] m296_13;
   assign m296_13 =10'b0;

   // m296_14 = W*in
   wire signed [9:0] m296_14;
   assign m296_14 =10'b0;

   // m296_15 = W*in
   wire signed [9:0] m296_15;
   assign m296_15 =10'b0;

   // m296_16 = W*in
   wire signed [9:0] m296_16;
   assign m296_16 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_17 = W*in
   wire signed [9:0] m296_17;
   assign m296_17 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_18 = W*in
   wire signed [9:0] m296_18;
   assign m296_18 ={ {5{in296[5]}} , in296[5:1] };

   // m296_19 = W*in
   wire signed [9:0] m296_19;
   assign m296_19 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_20 = W*in
   wire signed [9:0] m296_20;
   assign m296_20 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_21 = W*in
   wire signed [9:0] m296_21;
   assign m296_21 ={ {4{in296[5]}} , in296[5:0] };

   // m296_22 = W*in
   wire signed [9:0] m296_22;
   assign m296_22 =10'b0;

   // m296_23 = W*in
   wire signed [9:0] m296_23;
   assign m296_23 ={ {4{neg296[5]}} , neg296[5:0] };

   // m296_24 = W*in
   wire signed [9:0] m296_24;
   assign m296_24 ={ {4{neg296[5]}} , neg296[5:0] };

   // m296_25 = W*in
   wire signed [9:0] m296_25;
   assign m296_25 =10'b0;

   // m296_26 = W*in
   wire signed [9:0] m296_26;
   assign m296_26 ={ {5{in296[5]}} , in296[5:1] };

   // m296_27 = W*in
   wire signed [9:0] m296_27;
   assign m296_27 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_28 = W*in
   wire signed [9:0] m296_28;
   assign m296_28 =10'b0;

   // m296_29 = W*in
   wire signed [9:0] m296_29;
   assign m296_29 =10'b0;

   // m296_30 = W*in
   wire signed [9:0] m296_30;
   assign m296_30 =10'b0;

   // m296_31 = W*in
   wire signed [9:0] m296_31;
   assign m296_31 =10'b0;

   // m296_32 = W*in
   wire signed [9:0] m296_32;
   assign m296_32 =10'b0;

   // m296_33 = W*in
   wire signed [9:0] m296_33;
   assign m296_33 =10'b0;

   // m296_34 = W*in
   wire signed [9:0] m296_34;
   assign m296_34 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_35 = W*in
   wire signed [9:0] m296_35;
   assign m296_35 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_36 = W*in
   wire signed [9:0] m296_36;
   assign m296_36 =10'b0;

   // m296_37 = W*in
   wire signed [9:0] m296_37;
   assign m296_37 =10'b0;

   // m296_38 = W*in
   wire signed [9:0] m296_38;
   assign m296_38 =10'b0;

   // m296_39 = W*in
   wire signed [9:0] m296_39;
   assign m296_39 ={ {4{neg296[5]}} , neg296[5:0] };

   // m296_40 = W*in
   wire signed [9:0] m296_40;
   assign m296_40 =10'b0;

   // m296_41 = W*in
   wire signed [9:0] m296_41;
   assign m296_41 =10'b0;

   // m296_42 = W*in
   wire signed [9:0] m296_42;
   assign m296_42 =10'b0;

   // m296_43 = W*in
   wire signed [9:0] m296_43;
   assign m296_43 =10'b0;

   // m296_44 = W*in
   wire signed [9:0] m296_44;
   assign m296_44 =10'b0;

   // m296_45 = W*in
   wire signed [9:0] m296_45;
   assign m296_45 =10'b0;

   // m296_46 = W*in
   wire signed [9:0] m296_46;
   assign m296_46 =10'b0;

   // m296_47 = W*in
   wire signed [9:0] m296_47;
   assign m296_47 =10'b0;

   // m296_48 = W*in
   wire signed [9:0] m296_48;
   assign m296_48 =10'b0;

   // m296_49 = W*in
   wire signed [9:0] m296_49;
   assign m296_49 =10'b0;

   // m296_50 = W*in
   wire signed [9:0] m296_50;
   assign m296_50 =10'b0;

   // m296_51 = W*in
   wire signed [9:0] m296_51;
   assign m296_51 =10'b0;

   // m296_52 = W*in
   wire signed [9:0] m296_52;
   assign m296_52 =10'b0;

   // m296_53 = W*in
   wire signed [9:0] m296_53;
   assign m296_53 =10'b0;

   // m296_54 = W*in
   wire signed [9:0] m296_54;
   assign m296_54 =10'b0;

   // m296_55 = W*in
   wire signed [9:0] m296_55;
   assign m296_55 =10'b0;

   // m296_56 = W*in
   wire signed [9:0] m296_56;
   assign m296_56 =10'b0;

   // m296_57 = W*in
   wire signed [9:0] m296_57;
   assign m296_57 =10'b0;

   // m296_58 = W*in
   wire signed [9:0] m296_58;
   assign m296_58 =10'b0;

   // m296_59 = W*in
   wire signed [9:0] m296_59;
   assign m296_59 =10'b0;

   // m296_60 = W*in
   wire signed [9:0] m296_60;
   assign m296_60 =10'b0;

   // m296_61 = W*in
   wire signed [9:0] m296_61;
   assign m296_61 =10'b0;

   // m296_62 = W*in
   wire signed [9:0] m296_62;
   assign m296_62 =10'b0;

   // m296_63 = W*in
   wire signed [9:0] m296_63;
   assign m296_63 ={ {4{in296[5]}} , in296[5:0] };

   // m296_64 = W*in
   wire signed [9:0] m296_64;
   assign m296_64 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_65 = W*in
   wire signed [9:0] m296_65;
   assign m296_65 =10'b0;

   // m296_66 = W*in
   wire signed [9:0] m296_66;
   assign m296_66 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_67 = W*in
   wire signed [9:0] m296_67;
   assign m296_67 =10'b0;

   // m296_68 = W*in
   wire signed [9:0] m296_68;
   assign m296_68 =10'b0;

   // m296_69 = W*in
   wire signed [9:0] m296_69;
   assign m296_69 ={ {5{in296[5]}} , in296[5:1] };

   // m296_70 = W*in
   wire signed [9:0] m296_70;
   assign m296_70 ={ {5{in296[5]}} , in296[5:1] };

   // m296_71 = W*in
   wire signed [9:0] m296_71;
   assign m296_71 ={ {5{in296[5]}} , in296[5:1] };

   // m296_72 = W*in
   wire signed [9:0] m296_72;
   assign m296_72 ={ {4{in296[5]}} , in296[5:0] };

   // m296_73 = W*in
   wire signed [9:0] m296_73;
   assign m296_73 =10'b0;

   // m296_74 = W*in
   wire signed [9:0] m296_74;
   assign m296_74 ={ {5{in296[5]}} , in296[5:1] };

   // m296_75 = W*in
   wire signed [9:0] m296_75;
   assign m296_75 =10'b0;

   // m296_76 = W*in
   wire signed [9:0] m296_76;
   assign m296_76 =10'b0;

   // m296_77 = W*in
   wire signed [9:0] m296_77;
   assign m296_77 =10'b0;

   // m296_78 = W*in
   wire signed [9:0] m296_78;
   assign m296_78 =10'b0;

   // m296_79 = W*in
   wire signed [9:0] m296_79;
   assign m296_79 =10'b0;

   // m296_80 = W*in
   wire signed [9:0] m296_80;
   assign m296_80 =10'b0;

   // m296_81 = W*in
   wire signed [9:0] m296_81;
   assign m296_81 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_82 = W*in
   wire signed [9:0] m296_82;
   assign m296_82 =10'b0;

   // m296_83 = W*in
   wire signed [9:0] m296_83;
   assign m296_83 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_84 = W*in
   wire signed [9:0] m296_84;
   assign m296_84 ={ {4{in296[5]}} , in296[5:0] };

   // m296_85 = W*in
   wire signed [9:0] m296_85;
   assign m296_85 =10'b0;

   // m296_86 = W*in
   wire signed [9:0] m296_86;
   assign m296_86 =10'b0;

   // m296_87 = W*in
   wire signed [9:0] m296_87;
   assign m296_87 ={ {4{in296[5]}} , in296[5:0] };

   // m296_88 = W*in
   wire signed [9:0] m296_88;
   assign m296_88 =10'b0;

   // m296_89 = W*in
   wire signed [9:0] m296_89;
   assign m296_89 =10'b0;

   // m296_90 = W*in
   wire signed [9:0] m296_90;
   assign m296_90 =10'b0;

   // m296_91 = W*in
   wire signed [9:0] m296_91;
   assign m296_91 =10'b0;

   // m296_92 = W*in
   wire signed [9:0] m296_92;
   assign m296_92 =10'b0;

   // m296_93 = W*in
   wire signed [9:0] m296_93;
   assign m296_93 =10'b0;

   // m296_94 = W*in
   wire signed [9:0] m296_94;
   assign m296_94 =10'b0;

   // m296_95 = W*in
   wire signed [9:0] m296_95;
   assign m296_95 =10'b0;

   // m296_96 = W*in
   wire signed [9:0] m296_96;
   assign m296_96 =10'b0;

   // m296_97 = W*in
   wire signed [9:0] m296_97;
   assign m296_97 =10'b0;

   // m296_98 = W*in
   wire signed [9:0] m296_98;
   assign m296_98 =10'b0;

   // m296_99 = W*in
   wire signed [9:0] m296_99;
   assign m296_99 =10'b0;

   // m296_100 = W*in
   wire signed [9:0] m296_100;
   assign m296_100 =10'b0;

   // m296_101 = W*in
   wire signed [9:0] m296_101;
   assign m296_101 =10'b0;

   // m296_102 = W*in
   wire signed [9:0] m296_102;
   assign m296_102 =10'b0;

   // m296_103 = W*in
   wire signed [9:0] m296_103;
   assign m296_103 =10'b0;

   // m296_104 = W*in
   wire signed [9:0] m296_104;
   assign m296_104 =10'b0;

   // m296_105 = W*in
   wire signed [9:0] m296_105;
   assign m296_105 =10'b0;

   // m296_106 = W*in
   wire signed [9:0] m296_106;
   assign m296_106 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_107 = W*in
   wire signed [9:0] m296_107;
   assign m296_107 ={ {4{neg296[5]}} , neg296[5:0] };

   // m296_108 = W*in
   wire signed [9:0] m296_108;
   assign m296_108 =10'b0;

   // m296_109 = W*in
   wire signed [9:0] m296_109;
   assign m296_109 =10'b0;

   // m296_110 = W*in
   wire signed [9:0] m296_110;
   assign m296_110 =10'b0;

   // m296_111 = W*in
   wire signed [9:0] m296_111;
   assign m296_111 =10'b0;

   // m296_112 = W*in
   wire signed [9:0] m296_112;
   assign m296_112 =10'b0;

   // m296_113 = W*in
   wire signed [9:0] m296_113;
   assign m296_113 =10'b0;

   // m296_114 = W*in
   wire signed [9:0] m296_114;
   assign m296_114 =10'b0;

   // m296_115 = W*in
   wire signed [9:0] m296_115;
   assign m296_115 ={ {5{neg296[5]}} , neg296[5:1] };

   // m296_116 = W*in
   wire signed [9:0] m296_116;
   assign m296_116 =10'b0;

   // m296_117 = W*in
   wire signed [9:0] m296_117;
   assign m296_117 =10'b0;

   // m297_1 = W*in
   wire signed [9:0] m297_1;
   assign m297_1 =10'b0;

   // m297_2 = W*in
   wire signed [9:0] m297_2;
   assign m297_2 =10'b0;

   // m297_3 = W*in
   wire signed [9:0] m297_3;
   assign m297_3 =10'b0;

   // m297_4 = W*in
   wire signed [9:0] m297_4;
   assign m297_4 =10'b0;

   // m297_5 = W*in
   wire signed [9:0] m297_5;
   assign m297_5 =10'b0;

   // m297_6 = W*in
   wire signed [9:0] m297_6;
   assign m297_6 =10'b0;

   // m297_7 = W*in
   wire signed [9:0] m297_7;
   assign m297_7 =10'b0;

   // m297_8 = W*in
   wire signed [9:0] m297_8;
   assign m297_8 ={ {4{in297[5]}} , in297[5:0] };

   // m297_9 = W*in
   wire signed [9:0] m297_9;
   assign m297_9 =10'b0;

   // m297_10 = W*in
   wire signed [9:0] m297_10;
   assign m297_10 =10'b0;

   // m297_11 = W*in
   wire signed [9:0] m297_11;
   assign m297_11 =10'b0;

   // m297_12 = W*in
   wire signed [9:0] m297_12;
   assign m297_12 =10'b0;

   // m297_13 = W*in
   wire signed [9:0] m297_13;
   assign m297_13 =10'b0;

   // m297_14 = W*in
   wire signed [9:0] m297_14;
   assign m297_14 =10'b0;

   // m297_15 = W*in
   wire signed [9:0] m297_15;
   assign m297_15 =10'b0;

   // m297_16 = W*in
   wire signed [9:0] m297_16;
   assign m297_16 =10'b0;

   // m297_17 = W*in
   wire signed [9:0] m297_17;
   assign m297_17 =10'b0;

   // m297_18 = W*in
   wire signed [9:0] m297_18;
   assign m297_18 ={ {5{neg297[5]}} , neg297[5:1] };

   // m297_19 = W*in
   wire signed [9:0] m297_19;
   assign m297_19 =10'b0;

   // m297_20 = W*in
   wire signed [9:0] m297_20;
   assign m297_20 =10'b0;

   // m297_21 = W*in
   wire signed [9:0] m297_21;
   assign m297_21 =10'b0;

   // m297_22 = W*in
   wire signed [9:0] m297_22;
   assign m297_22 =10'b0;

   // m297_23 = W*in
   wire signed [9:0] m297_23;
   assign m297_23 =10'b0;

   // m297_24 = W*in
   wire signed [9:0] m297_24;
   assign m297_24 =10'b0;

   // m297_25 = W*in
   wire signed [9:0] m297_25;
   assign m297_25 =10'b0;

   // m297_26 = W*in
   wire signed [9:0] m297_26;
   assign m297_26 ={ {4{neg297[5]}} , neg297[5:0] };

   // m297_27 = W*in
   wire signed [9:0] m297_27;
   assign m297_27 =10'b0;

   // m297_28 = W*in
   wire signed [9:0] m297_28;
   assign m297_28 =10'b0;

   // m297_29 = W*in
   wire signed [9:0] m297_29;
   assign m297_29 =10'b0;

   // m297_30 = W*in
   wire signed [9:0] m297_30;
   assign m297_30 =10'b0;

   // m297_31 = W*in
   wire signed [9:0] m297_31;
   assign m297_31 ={ {5{in297[5]}} , in297[5:1] };

   // m297_32 = W*in
   wire signed [9:0] m297_32;
   assign m297_32 =10'b0;

   // m297_33 = W*in
   wire signed [9:0] m297_33;
   assign m297_33 =10'b0;

   // m297_34 = W*in
   wire signed [9:0] m297_34;
   assign m297_34 =10'b0;

   // m297_35 = W*in
   wire signed [9:0] m297_35;
   assign m297_35 =10'b0;

   // m297_36 = W*in
   wire signed [9:0] m297_36;
   assign m297_36 =10'b0;

   // m297_37 = W*in
   wire signed [9:0] m297_37;
   assign m297_37 =10'b0;

   // m297_38 = W*in
   wire signed [9:0] m297_38;
   assign m297_38 =10'b0;

   // m297_39 = W*in
   wire signed [9:0] m297_39;
   assign m297_39 =10'b0;

   // m297_40 = W*in
   wire signed [9:0] m297_40;
   assign m297_40 =10'b0;

   // m297_41 = W*in
   wire signed [9:0] m297_41;
   assign m297_41 =10'b0;

   // m297_42 = W*in
   wire signed [9:0] m297_42;
   assign m297_42 =10'b0;

   // m297_43 = W*in
   wire signed [9:0] m297_43;
   assign m297_43 =10'b0;

   // m297_44 = W*in
   wire signed [9:0] m297_44;
   assign m297_44 =10'b0;

   // m297_45 = W*in
   wire signed [9:0] m297_45;
   assign m297_45 =10'b0;

   // m297_46 = W*in
   wire signed [9:0] m297_46;
   assign m297_46 =10'b0;

   // m297_47 = W*in
   wire signed [9:0] m297_47;
   assign m297_47 =10'b0;

   // m297_48 = W*in
   wire signed [9:0] m297_48;
   assign m297_48 =10'b0;

   // m297_49 = W*in
   wire signed [9:0] m297_49;
   assign m297_49 =10'b0;

   // m297_50 = W*in
   wire signed [9:0] m297_50;
   assign m297_50 =10'b0;

   // m297_51 = W*in
   wire signed [9:0] m297_51;
   assign m297_51 =10'b0;

   // m297_52 = W*in
   wire signed [9:0] m297_52;
   assign m297_52 =10'b0;

   // m297_53 = W*in
   wire signed [9:0] m297_53;
   assign m297_53 =10'b0;

   // m297_54 = W*in
   wire signed [9:0] m297_54;
   assign m297_54 =10'b0;

   // m297_55 = W*in
   wire signed [9:0] m297_55;
   assign m297_55 =10'b0;

   // m297_56 = W*in
   wire signed [9:0] m297_56;
   assign m297_56 =10'b0;

   // m297_57 = W*in
   wire signed [9:0] m297_57;
   assign m297_57 =10'b0;

   // m297_58 = W*in
   wire signed [9:0] m297_58;
   assign m297_58 =10'b0;

   // m297_59 = W*in
   wire signed [9:0] m297_59;
   assign m297_59 =10'b0;

   // m297_60 = W*in
   wire signed [9:0] m297_60;
   assign m297_60 =10'b0;

   // m297_61 = W*in
   wire signed [9:0] m297_61;
   assign m297_61 =10'b0;

   // m297_62 = W*in
   wire signed [9:0] m297_62;
   assign m297_62 =10'b0;

   // m297_63 = W*in
   wire signed [9:0] m297_63;
   assign m297_63 =10'b0;

   // m297_64 = W*in
   wire signed [9:0] m297_64;
   assign m297_64 ={ {5{neg297[5]}} , neg297[5:1] };

   // m297_65 = W*in
   wire signed [9:0] m297_65;
   assign m297_65 =10'b0;

   // m297_66 = W*in
   wire signed [9:0] m297_66;
   assign m297_66 =10'b0;

   // m297_67 = W*in
   wire signed [9:0] m297_67;
   assign m297_67 =10'b0;

   // m297_68 = W*in
   wire signed [9:0] m297_68;
   assign m297_68 =10'b0;

   // m297_69 = W*in
   wire signed [9:0] m297_69;
   assign m297_69 ={ {5{in297[5]}} , in297[5:1] };

   // m297_70 = W*in
   wire signed [9:0] m297_70;
   assign m297_70 =10'b0;

   // m297_71 = W*in
   wire signed [9:0] m297_71;
   assign m297_71 =10'b0;

   // m297_72 = W*in
   wire signed [9:0] m297_72;
   assign m297_72 =10'b0;

   // m297_73 = W*in
   wire signed [9:0] m297_73;
   assign m297_73 ={ {5{in297[5]}} , in297[5:1] };

   // m297_74 = W*in
   wire signed [9:0] m297_74;
   assign m297_74 =10'b0;

   // m297_75 = W*in
   wire signed [9:0] m297_75;
   assign m297_75 =10'b0;

   // m297_76 = W*in
   wire signed [9:0] m297_76;
   assign m297_76 =10'b0;

   // m297_77 = W*in
   wire signed [9:0] m297_77;
   assign m297_77 ={ {4{neg297[5]}} , neg297[5:0] };

   // m297_78 = W*in
   wire signed [9:0] m297_78;
   assign m297_78 =10'b0;

   // m297_79 = W*in
   wire signed [9:0] m297_79;
   assign m297_79 =10'b0;

   // m297_80 = W*in
   wire signed [9:0] m297_80;
   assign m297_80 =10'b0;

   // m297_81 = W*in
   wire signed [9:0] m297_81;
   assign m297_81 =10'b0;

   // m297_82 = W*in
   wire signed [9:0] m297_82;
   assign m297_82 ={ {4{in297[5]}} , in297[5:0] };

   // m297_83 = W*in
   wire signed [9:0] m297_83;
   assign m297_83 =10'b0;

   // m297_84 = W*in
   wire signed [9:0] m297_84;
   assign m297_84 =10'b0;

   // m297_85 = W*in
   wire signed [9:0] m297_85;
   assign m297_85 ={ {4{in297[5]}} , in297[5:0] };

   // m297_86 = W*in
   wire signed [9:0] m297_86;
   assign m297_86 =10'b0;

   // m297_87 = W*in
   wire signed [9:0] m297_87;
   assign m297_87 =10'b0;

   // m297_88 = W*in
   wire signed [9:0] m297_88;
   assign m297_88 =10'b0;

   // m297_89 = W*in
   wire signed [9:0] m297_89;
   assign m297_89 =10'b0;

   // m297_90 = W*in
   wire signed [9:0] m297_90;
   assign m297_90 =10'b0;

   // m297_91 = W*in
   wire signed [9:0] m297_91;
   assign m297_91 =10'b0;

   // m297_92 = W*in
   wire signed [9:0] m297_92;
   assign m297_92 =10'b0;

   // m297_93 = W*in
   wire signed [9:0] m297_93;
   assign m297_93 =10'b0;

   // m297_94 = W*in
   wire signed [9:0] m297_94;
   assign m297_94 =10'b0;

   // m297_95 = W*in
   wire signed [9:0] m297_95;
   assign m297_95 =10'b0;

   // m297_96 = W*in
   wire signed [9:0] m297_96;
   assign m297_96 =10'b0;

   // m297_97 = W*in
   wire signed [9:0] m297_97;
   assign m297_97 ={ {4{neg297[5]}} , neg297[5:0] };

   // m297_98 = W*in
   wire signed [9:0] m297_98;
   assign m297_98 =10'b0;

   // m297_99 = W*in
   wire signed [9:0] m297_99;
   assign m297_99 =10'b0;

   // m297_100 = W*in
   wire signed [9:0] m297_100;
   assign m297_100 =10'b0;

   // m297_101 = W*in
   wire signed [9:0] m297_101;
   assign m297_101 =10'b0;

   // m297_102 = W*in
   wire signed [9:0] m297_102;
   assign m297_102 =10'b0;

   // m297_103 = W*in
   wire signed [9:0] m297_103;
   assign m297_103 =10'b0;

   // m297_104 = W*in
   wire signed [9:0] m297_104;
   assign m297_104 =10'b0;

   // m297_105 = W*in
   wire signed [9:0] m297_105;
   assign m297_105 =10'b0;

   // m297_106 = W*in
   wire signed [9:0] m297_106;
   assign m297_106 =10'b0;

   // m297_107 = W*in
   wire signed [9:0] m297_107;
   assign m297_107 =10'b0;

   // m297_108 = W*in
   wire signed [9:0] m297_108;
   assign m297_108 ={ {5{in297[5]}} , in297[5:1] };

   // m297_109 = W*in
   wire signed [9:0] m297_109;
   assign m297_109 ={ {4{in297[5]}} , in297[5:0] };

   // m297_110 = W*in
   wire signed [9:0] m297_110;
   assign m297_110 =10'b0;

   // m297_111 = W*in
   wire signed [9:0] m297_111;
   assign m297_111 =10'b0;

   // m297_112 = W*in
   wire signed [9:0] m297_112;
   assign m297_112 =10'b0;

   // m297_113 = W*in
   wire signed [9:0] m297_113;
   assign m297_113 =10'b0;

   // m297_114 = W*in
   wire signed [9:0] m297_114;
   assign m297_114 =10'b0;

   // m297_115 = W*in
   wire signed [9:0] m297_115;
   assign m297_115 =10'b0;

   // m297_116 = W*in
   wire signed [9:0] m297_116;
   assign m297_116 =10'b0;

   // m297_117 = W*in
   wire signed [9:0] m297_117;
   assign m297_117 =10'b0;

   // m298_1 = W*in
   wire signed [9:0] m298_1;
   assign m298_1 =10'b0;

   // m298_2 = W*in
   wire signed [9:0] m298_2;
   assign m298_2 =10'b0;

   // m298_3 = W*in
   wire signed [9:0] m298_3;
   assign m298_3 =10'b0;

   // m298_4 = W*in
   wire signed [9:0] m298_4;
   assign m298_4 =10'b0;

   // m298_5 = W*in
   wire signed [9:0] m298_5;
   assign m298_5 =10'b0;

   // m298_6 = W*in
   wire signed [9:0] m298_6;
   assign m298_6 =10'b0;

   // m298_7 = W*in
   wire signed [9:0] m298_7;
   assign m298_7 =10'b0;

   // m298_8 = W*in
   wire signed [9:0] m298_8;
   assign m298_8 =10'b0;

   // m298_9 = W*in
   wire signed [9:0] m298_9;
   assign m298_9 =10'b0;

   // m298_10 = W*in
   wire signed [9:0] m298_10;
   assign m298_10 =10'b0;

   // m298_11 = W*in
   wire signed [9:0] m298_11;
   assign m298_11 =10'b0;

   // m298_12 = W*in
   wire signed [9:0] m298_12;
   assign m298_12 =10'b0;

   // m298_13 = W*in
   wire signed [9:0] m298_13;
   assign m298_13 ={ {4{in298[5]}} , in298[5:0] };

   // m298_14 = W*in
   wire signed [9:0] m298_14;
   assign m298_14 =10'b0;

   // m298_15 = W*in
   wire signed [9:0] m298_15;
   assign m298_15 =10'b0;

   // m298_16 = W*in
   wire signed [9:0] m298_16;
   assign m298_16 =10'b0;

   // m298_17 = W*in
   wire signed [9:0] m298_17;
   assign m298_17 =10'b0;

   // m298_18 = W*in
   wire signed [9:0] m298_18;
   assign m298_18 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_19 = W*in
   wire signed [9:0] m298_19;
   assign m298_19 =10'b0;

   // m298_20 = W*in
   wire signed [9:0] m298_20;
   assign m298_20 ={ {5{neg298[5]}} , neg298[5:1] };

   // m298_21 = W*in
   wire signed [9:0] m298_21;
   assign m298_21 ={ {5{in298[5]}} , in298[5:1] };

   // m298_22 = W*in
   wire signed [9:0] m298_22;
   assign m298_22 =10'b0;

   // m298_23 = W*in
   wire signed [9:0] m298_23;
   assign m298_23 =10'b0;

   // m298_24 = W*in
   wire signed [9:0] m298_24;
   assign m298_24 =10'b0;

   // m298_25 = W*in
   wire signed [9:0] m298_25;
   assign m298_25 =10'b0;

   // m298_26 = W*in
   wire signed [9:0] m298_26;
   assign m298_26 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_27 = W*in
   wire signed [9:0] m298_27;
   assign m298_27 =10'b0;

   // m298_28 = W*in
   wire signed [9:0] m298_28;
   assign m298_28 =10'b0;

   // m298_29 = W*in
   wire signed [9:0] m298_29;
   assign m298_29 =10'b0;

   // m298_30 = W*in
   wire signed [9:0] m298_30;
   assign m298_30 =10'b0;

   // m298_31 = W*in
   wire signed [9:0] m298_31;
   assign m298_31 =10'b0;

   // m298_32 = W*in
   wire signed [9:0] m298_32;
   assign m298_32 =10'b0;

   // m298_33 = W*in
   wire signed [9:0] m298_33;
   assign m298_33 =10'b0;

   // m298_34 = W*in
   wire signed [9:0] m298_34;
   assign m298_34 =10'b0;

   // m298_35 = W*in
   wire signed [9:0] m298_35;
   assign m298_35 =10'b0;

   // m298_36 = W*in
   wire signed [9:0] m298_36;
   assign m298_36 =10'b0;

   // m298_37 = W*in
   wire signed [9:0] m298_37;
   assign m298_37 =10'b0;

   // m298_38 = W*in
   wire signed [9:0] m298_38;
   assign m298_38 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_39 = W*in
   wire signed [9:0] m298_39;
   assign m298_39 =10'b0;

   // m298_40 = W*in
   wire signed [9:0] m298_40;
   assign m298_40 =10'b0;

   // m298_41 = W*in
   wire signed [9:0] m298_41;
   assign m298_41 ={ {4{in298[5]}} , in298[5:0] };

   // m298_42 = W*in
   wire signed [9:0] m298_42;
   assign m298_42 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_43 = W*in
   wire signed [9:0] m298_43;
   assign m298_43 =10'b0;

   // m298_44 = W*in
   wire signed [9:0] m298_44;
   assign m298_44 =10'b0;

   // m298_45 = W*in
   wire signed [9:0] m298_45;
   assign m298_45 =10'b0;

   // m298_46 = W*in
   wire signed [9:0] m298_46;
   assign m298_46 =10'b0;

   // m298_47 = W*in
   wire signed [9:0] m298_47;
   assign m298_47 =10'b0;

   // m298_48 = W*in
   wire signed [9:0] m298_48;
   assign m298_48 =10'b0;

   // m298_49 = W*in
   wire signed [9:0] m298_49;
   assign m298_49 =10'b0;

   // m298_50 = W*in
   wire signed [9:0] m298_50;
   assign m298_50 =10'b0;

   // m298_51 = W*in
   wire signed [9:0] m298_51;
   assign m298_51 =10'b0;

   // m298_52 = W*in
   wire signed [9:0] m298_52;
   assign m298_52 =10'b0;

   // m298_53 = W*in
   wire signed [9:0] m298_53;
   assign m298_53 =10'b0;

   // m298_54 = W*in
   wire signed [9:0] m298_54;
   assign m298_54 =10'b0;

   // m298_55 = W*in
   wire signed [9:0] m298_55;
   assign m298_55 =10'b0;

   // m298_56 = W*in
   wire signed [9:0] m298_56;
   assign m298_56 =10'b0;

   // m298_57 = W*in
   wire signed [9:0] m298_57;
   assign m298_57 =10'b0;

   // m298_58 = W*in
   wire signed [9:0] m298_58;
   assign m298_58 =10'b0;

   // m298_59 = W*in
   wire signed [9:0] m298_59;
   assign m298_59 =10'b0;

   // m298_60 = W*in
   wire signed [9:0] m298_60;
   assign m298_60 =10'b0;

   // m298_61 = W*in
   wire signed [9:0] m298_61;
   assign m298_61 =10'b0;

   // m298_62 = W*in
   wire signed [9:0] m298_62;
   assign m298_62 =10'b0;

   // m298_63 = W*in
   wire signed [9:0] m298_63;
   assign m298_63 =10'b0;

   // m298_64 = W*in
   wire signed [9:0] m298_64;
   assign m298_64 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_65 = W*in
   wire signed [9:0] m298_65;
   assign m298_65 =10'b0;

   // m298_66 = W*in
   wire signed [9:0] m298_66;
   assign m298_66 =10'b0;

   // m298_67 = W*in
   wire signed [9:0] m298_67;
   assign m298_67 =10'b0;

   // m298_68 = W*in
   wire signed [9:0] m298_68;
   assign m298_68 =10'b0;

   // m298_69 = W*in
   wire signed [9:0] m298_69;
   assign m298_69 ={ {4{in298[5]}} , in298[5:0] };

   // m298_70 = W*in
   wire signed [9:0] m298_70;
   assign m298_70 =10'b0;

   // m298_71 = W*in
   wire signed [9:0] m298_71;
   assign m298_71 =10'b0;

   // m298_72 = W*in
   wire signed [9:0] m298_72;
   assign m298_72 =10'b0;

   // m298_73 = W*in
   wire signed [9:0] m298_73;
   assign m298_73 =10'b0;

   // m298_74 = W*in
   wire signed [9:0] m298_74;
   assign m298_74 =10'b0;

   // m298_75 = W*in
   wire signed [9:0] m298_75;
   assign m298_75 =10'b0;

   // m298_76 = W*in
   wire signed [9:0] m298_76;
   assign m298_76 =10'b0;

   // m298_77 = W*in
   wire signed [9:0] m298_77;
   assign m298_77 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_78 = W*in
   wire signed [9:0] m298_78;
   assign m298_78 =10'b0;

   // m298_79 = W*in
   wire signed [9:0] m298_79;
   assign m298_79 =10'b0;

   // m298_80 = W*in
   wire signed [9:0] m298_80;
   assign m298_80 =10'b0;

   // m298_81 = W*in
   wire signed [9:0] m298_81;
   assign m298_81 ={ {5{neg298[5]}} , neg298[5:1] };

   // m298_82 = W*in
   wire signed [9:0] m298_82;
   assign m298_82 =10'b0;

   // m298_83 = W*in
   wire signed [9:0] m298_83;
   assign m298_83 =10'b0;

   // m298_84 = W*in
   wire signed [9:0] m298_84;
   assign m298_84 =10'b0;

   // m298_85 = W*in
   wire signed [9:0] m298_85;
   assign m298_85 ={ {4{in298[5]}} , in298[5:0] };

   // m298_86 = W*in
   wire signed [9:0] m298_86;
   assign m298_86 =10'b0;

   // m298_87 = W*in
   wire signed [9:0] m298_87;
   assign m298_87 =10'b0;

   // m298_88 = W*in
   wire signed [9:0] m298_88;
   assign m298_88 =10'b0;

   // m298_89 = W*in
   wire signed [9:0] m298_89;
   assign m298_89 =10'b0;

   // m298_90 = W*in
   wire signed [9:0] m298_90;
   assign m298_90 =10'b0;

   // m298_91 = W*in
   wire signed [9:0] m298_91;
   assign m298_91 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_92 = W*in
   wire signed [9:0] m298_92;
   assign m298_92 =10'b0;

   // m298_93 = W*in
   wire signed [9:0] m298_93;
   assign m298_93 =10'b0;

   // m298_94 = W*in
   wire signed [9:0] m298_94;
   assign m298_94 =10'b0;

   // m298_95 = W*in
   wire signed [9:0] m298_95;
   assign m298_95 =10'b0;

   // m298_96 = W*in
   wire signed [9:0] m298_96;
   assign m298_96 =10'b0;

   // m298_97 = W*in
   wire signed [9:0] m298_97;
   assign m298_97 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_98 = W*in
   wire signed [9:0] m298_98;
   assign m298_98 =10'b0;

   // m298_99 = W*in
   wire signed [9:0] m298_99;
   assign m298_99 =10'b0;

   // m298_100 = W*in
   wire signed [9:0] m298_100;
   assign m298_100 =10'b0;

   // m298_101 = W*in
   wire signed [9:0] m298_101;
   assign m298_101 =10'b0;

   // m298_102 = W*in
   wire signed [9:0] m298_102;
   assign m298_102 =10'b0;

   // m298_103 = W*in
   wire signed [9:0] m298_103;
   assign m298_103 =10'b0;

   // m298_104 = W*in
   wire signed [9:0] m298_104;
   assign m298_104 =10'b0;

   // m298_105 = W*in
   wire signed [9:0] m298_105;
   assign m298_105 =10'b0;

   // m298_106 = W*in
   wire signed [9:0] m298_106;
   assign m298_106 =10'b0;

   // m298_107 = W*in
   wire signed [9:0] m298_107;
   assign m298_107 =10'b0;

   // m298_108 = W*in
   wire signed [9:0] m298_108;
   assign m298_108 ={ {4{in298[5]}} , in298[5:0] };

   // m298_109 = W*in
   wire signed [9:0] m298_109;
   assign m298_109 ={ {4{in298[5]}} , in298[5:0] };

   // m298_110 = W*in
   wire signed [9:0] m298_110;
   assign m298_110 ={ {4{neg298[5]}} , neg298[5:0] };

   // m298_111 = W*in
   wire signed [9:0] m298_111;
   assign m298_111 =10'b0;

   // m298_112 = W*in
   wire signed [9:0] m298_112;
   assign m298_112 =10'b0;

   // m298_113 = W*in
   wire signed [9:0] m298_113;
   assign m298_113 =10'b0;

   // m298_114 = W*in
   wire signed [9:0] m298_114;
   assign m298_114 =10'b0;

   // m298_115 = W*in
   wire signed [9:0] m298_115;
   assign m298_115 =10'b0;

   // m298_116 = W*in
   wire signed [9:0] m298_116;
   assign m298_116 ={ {4{in298[5]}} , in298[5:0] };

   // m298_117 = W*in
   wire signed [9:0] m298_117;
   assign m298_117 =10'b0;

   // m299_1 = W*in
   wire signed [9:0] m299_1;
   assign m299_1 ={ {4{in299[5]}} , in299[5:0] };

   // m299_2 = W*in
   wire signed [9:0] m299_2;
   assign m299_2 =10'b0;

   // m299_3 = W*in
   wire signed [9:0] m299_3;
   assign m299_3 =10'b0;

   // m299_4 = W*in
   wire signed [9:0] m299_4;
   assign m299_4 =10'b0;

   // m299_5 = W*in
   wire signed [9:0] m299_5;
   assign m299_5 =10'b0;

   // m299_6 = W*in
   wire signed [9:0] m299_6;
   assign m299_6 =10'b0;

   // m299_7 = W*in
   wire signed [9:0] m299_7;
   assign m299_7 ={ {4{in299[5]}} , in299[5:0] };

   // m299_8 = W*in
   wire signed [9:0] m299_8;
   assign m299_8 =10'b0;

   // m299_9 = W*in
   wire signed [9:0] m299_9;
   assign m299_9 =10'b0;

   // m299_10 = W*in
   wire signed [9:0] m299_10;
   assign m299_10 =10'b0;

   // m299_11 = W*in
   wire signed [9:0] m299_11;
   assign m299_11 =10'b0;

   // m299_12 = W*in
   wire signed [9:0] m299_12;
   assign m299_12 =10'b0;

   // m299_13 = W*in
   wire signed [9:0] m299_13;
   assign m299_13 =10'b0;

   // m299_14 = W*in
   wire signed [9:0] m299_14;
   assign m299_14 =10'b0;

   // m299_15 = W*in
   wire signed [9:0] m299_15;
   assign m299_15 =10'b0;

   // m299_16 = W*in
   wire signed [9:0] m299_16;
   assign m299_16 =10'b0;

   // m299_17 = W*in
   wire signed [9:0] m299_17;
   assign m299_17 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_18 = W*in
   wire signed [9:0] m299_18;
   assign m299_18 =10'b0;

   // m299_19 = W*in
   wire signed [9:0] m299_19;
   assign m299_19 ={ {4{neg299[5]}} , neg299[5:0] };

   // m299_20 = W*in
   wire signed [9:0] m299_20;
   assign m299_20 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_21 = W*in
   wire signed [9:0] m299_21;
   assign m299_21 ={ {5{in299[5]}} , in299[5:1] };

   // m299_22 = W*in
   wire signed [9:0] m299_22;
   assign m299_22 =10'b0;

   // m299_23 = W*in
   wire signed [9:0] m299_23;
   assign m299_23 =10'b0;

   // m299_24 = W*in
   wire signed [9:0] m299_24;
   assign m299_24 =10'b0;

   // m299_25 = W*in
   wire signed [9:0] m299_25;
   assign m299_25 =10'b0;

   // m299_26 = W*in
   wire signed [9:0] m299_26;
   assign m299_26 ={ {5{in299[5]}} , in299[5:1] };

   // m299_27 = W*in
   wire signed [9:0] m299_27;
   assign m299_27 =10'b0;

   // m299_28 = W*in
   wire signed [9:0] m299_28;
   assign m299_28 ={ {5{in299[5]}} , in299[5:1] };

   // m299_29 = W*in
   wire signed [9:0] m299_29;
   assign m299_29 =10'b0;

   // m299_30 = W*in
   wire signed [9:0] m299_30;
   assign m299_30 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_31 = W*in
   wire signed [9:0] m299_31;
   assign m299_31 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_32 = W*in
   wire signed [9:0] m299_32;
   assign m299_32 =10'b0;

   // m299_33 = W*in
   wire signed [9:0] m299_33;
   assign m299_33 ={ {4{in299[5]}} , in299[5:0] };

   // m299_34 = W*in
   wire signed [9:0] m299_34;
   assign m299_34 =10'b0;

   // m299_35 = W*in
   wire signed [9:0] m299_35;
   assign m299_35 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_36 = W*in
   wire signed [9:0] m299_36;
   assign m299_36 =10'b0;

   // m299_37 = W*in
   wire signed [9:0] m299_37;
   assign m299_37 =10'b0;

   // m299_38 = W*in
   wire signed [9:0] m299_38;
   assign m299_38 =10'b0;

   // m299_39 = W*in
   wire signed [9:0] m299_39;
   assign m299_39 =10'b0;

   // m299_40 = W*in
   wire signed [9:0] m299_40;
   assign m299_40 =10'b0;

   // m299_41 = W*in
   wire signed [9:0] m299_41;
   assign m299_41 =10'b0;

   // m299_42 = W*in
   wire signed [9:0] m299_42;
   assign m299_42 =10'b0;

   // m299_43 = W*in
   wire signed [9:0] m299_43;
   assign m299_43 =10'b0;

   // m299_44 = W*in
   wire signed [9:0] m299_44;
   assign m299_44 =10'b0;

   // m299_45 = W*in
   wire signed [9:0] m299_45;
   assign m299_45 =10'b0;

   // m299_46 = W*in
   wire signed [9:0] m299_46;
   assign m299_46 =10'b0;

   // m299_47 = W*in
   wire signed [9:0] m299_47;
   assign m299_47 =10'b0;

   // m299_48 = W*in
   wire signed [9:0] m299_48;
   assign m299_48 =10'b0;

   // m299_49 = W*in
   wire signed [9:0] m299_49;
   assign m299_49 =10'b0;

   // m299_50 = W*in
   wire signed [9:0] m299_50;
   assign m299_50 =10'b0;

   // m299_51 = W*in
   wire signed [9:0] m299_51;
   assign m299_51 =10'b0;

   // m299_52 = W*in
   wire signed [9:0] m299_52;
   assign m299_52 =10'b0;

   // m299_53 = W*in
   wire signed [9:0] m299_53;
   assign m299_53 ={ {4{neg299[5]}} , neg299[5:0] };

   // m299_54 = W*in
   wire signed [9:0] m299_54;
   assign m299_54 =10'b0;

   // m299_55 = W*in
   wire signed [9:0] m299_55;
   assign m299_55 =10'b0;

   // m299_56 = W*in
   wire signed [9:0] m299_56;
   assign m299_56 =10'b0;

   // m299_57 = W*in
   wire signed [9:0] m299_57;
   assign m299_57 =10'b0;

   // m299_58 = W*in
   wire signed [9:0] m299_58;
   assign m299_58 =10'b0;

   // m299_59 = W*in
   wire signed [9:0] m299_59;
   assign m299_59 =10'b0;

   // m299_60 = W*in
   wire signed [9:0] m299_60;
   assign m299_60 =10'b0;

   // m299_61 = W*in
   wire signed [9:0] m299_61;
   assign m299_61 ={ {4{neg299[5]}} , neg299[5:0] };

   // m299_62 = W*in
   wire signed [9:0] m299_62;
   assign m299_62 =10'b0;

   // m299_63 = W*in
   wire signed [9:0] m299_63;
   assign m299_63 =10'b0;

   // m299_64 = W*in
   wire signed [9:0] m299_64;
   assign m299_64 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_65 = W*in
   wire signed [9:0] m299_65;
   assign m299_65 =10'b0;

   // m299_66 = W*in
   wire signed [9:0] m299_66;
   assign m299_66 =10'b0;

   // m299_67 = W*in
   wire signed [9:0] m299_67;
   assign m299_67 =10'b0;

   // m299_68 = W*in
   wire signed [9:0] m299_68;
   assign m299_68 =10'b0;

   // m299_69 = W*in
   wire signed [9:0] m299_69;
   assign m299_69 =10'b0;

   // m299_70 = W*in
   wire signed [9:0] m299_70;
   assign m299_70 =10'b0;

   // m299_71 = W*in
   wire signed [9:0] m299_71;
   assign m299_71 =10'b0;

   // m299_72 = W*in
   wire signed [9:0] m299_72;
   assign m299_72 =10'b0;

   // m299_73 = W*in
   wire signed [9:0] m299_73;
   assign m299_73 =10'b0;

   // m299_74 = W*in
   wire signed [9:0] m299_74;
   assign m299_74 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_75 = W*in
   wire signed [9:0] m299_75;
   assign m299_75 =10'b0;

   // m299_76 = W*in
   wire signed [9:0] m299_76;
   assign m299_76 =10'b0;

   // m299_77 = W*in
   wire signed [9:0] m299_77;
   assign m299_77 =10'b0;

   // m299_78 = W*in
   wire signed [9:0] m299_78;
   assign m299_78 ={ {4{in299[5]}} , in299[5:0] };

   // m299_79 = W*in
   wire signed [9:0] m299_79;
   assign m299_79 =10'b0;

   // m299_80 = W*in
   wire signed [9:0] m299_80;
   assign m299_80 =10'b0;

   // m299_81 = W*in
   wire signed [9:0] m299_81;
   assign m299_81 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_82 = W*in
   wire signed [9:0] m299_82;
   assign m299_82 =10'b0;

   // m299_83 = W*in
   wire signed [9:0] m299_83;
   assign m299_83 =10'b0;

   // m299_84 = W*in
   wire signed [9:0] m299_84;
   assign m299_84 ={ {5{in299[5]}} , in299[5:1] };

   // m299_85 = W*in
   wire signed [9:0] m299_85;
   assign m299_85 ={ {5{in299[5]}} , in299[5:1] };

   // m299_86 = W*in
   wire signed [9:0] m299_86;
   assign m299_86 =10'b0;

   // m299_87 = W*in
   wire signed [9:0] m299_87;
   assign m299_87 =10'b0;

   // m299_88 = W*in
   wire signed [9:0] m299_88;
   assign m299_88 =10'b0;

   // m299_89 = W*in
   wire signed [9:0] m299_89;
   assign m299_89 =10'b0;

   // m299_90 = W*in
   wire signed [9:0] m299_90;
   assign m299_90 =10'b0;

   // m299_91 = W*in
   wire signed [9:0] m299_91;
   assign m299_91 =10'b0;

   // m299_92 = W*in
   wire signed [9:0] m299_92;
   assign m299_92 =10'b0;

   // m299_93 = W*in
   wire signed [9:0] m299_93;
   assign m299_93 =10'b0;

   // m299_94 = W*in
   wire signed [9:0] m299_94;
   assign m299_94 =10'b0;

   // m299_95 = W*in
   wire signed [9:0] m299_95;
   assign m299_95 =10'b0;

   // m299_96 = W*in
   wire signed [9:0] m299_96;
   assign m299_96 =10'b0;

   // m299_97 = W*in
   wire signed [9:0] m299_97;
   assign m299_97 =10'b0;

   // m299_98 = W*in
   wire signed [9:0] m299_98;
   assign m299_98 =10'b0;

   // m299_99 = W*in
   wire signed [9:0] m299_99;
   assign m299_99 =10'b0;

   // m299_100 = W*in
   wire signed [9:0] m299_100;
   assign m299_100 =10'b0;

   // m299_101 = W*in
   wire signed [9:0] m299_101;
   assign m299_101 =10'b0;

   // m299_102 = W*in
   wire signed [9:0] m299_102;
   assign m299_102 =10'b0;

   // m299_103 = W*in
   wire signed [9:0] m299_103;
   assign m299_103 =10'b0;

   // m299_104 = W*in
   wire signed [9:0] m299_104;
   assign m299_104 =10'b0;

   // m299_105 = W*in
   wire signed [9:0] m299_105;
   assign m299_105 =10'b0;

   // m299_106 = W*in
   wire signed [9:0] m299_106;
   assign m299_106 =10'b0;

   // m299_107 = W*in
   wire signed [9:0] m299_107;
   assign m299_107 =10'b0;

   // m299_108 = W*in
   wire signed [9:0] m299_108;
   assign m299_108 =10'b0;

   // m299_109 = W*in
   wire signed [9:0] m299_109;
   assign m299_109 =10'b0;

   // m299_110 = W*in
   wire signed [9:0] m299_110;
   assign m299_110 =10'b0;

   // m299_111 = W*in
   wire signed [9:0] m299_111;
   assign m299_111 ={ {4{in299[5]}} , in299[5:0] };

   // m299_112 = W*in
   wire signed [9:0] m299_112;
   assign m299_112 =10'b0;

   // m299_113 = W*in
   wire signed [9:0] m299_113;
   assign m299_113 =10'b0;

   // m299_114 = W*in
   wire signed [9:0] m299_114;
   assign m299_114 =10'b0;

   // m299_115 = W*in
   wire signed [9:0] m299_115;
   assign m299_115 ={ {5{neg299[5]}} , neg299[5:1] };

   // m299_116 = W*in
   wire signed [9:0] m299_116;
   assign m299_116 =10'b0;

   // m299_117 = W*in
   wire signed [9:0] m299_117;
   assign m299_117 =10'b0;

   // m300_1 = W*in
   wire signed [9:0] m300_1;
   assign m300_1 =10'b0;

   // m300_2 = W*in
   wire signed [9:0] m300_2;
   assign m300_2 =10'b0;

   // m300_3 = W*in
   wire signed [9:0] m300_3;
   assign m300_3 =10'b0;

   // m300_4 = W*in
   wire signed [9:0] m300_4;
   assign m300_4 =10'b0;

   // m300_5 = W*in
   wire signed [9:0] m300_5;
   assign m300_5 =10'b0;

   // m300_6 = W*in
   wire signed [9:0] m300_6;
   assign m300_6 ={ {4{in300[5]}} , in300[5:0] };

   // m300_7 = W*in
   wire signed [9:0] m300_7;
   assign m300_7 =10'b0;

   // m300_8 = W*in
   wire signed [9:0] m300_8;
   assign m300_8 =10'b0;

   // m300_9 = W*in
   wire signed [9:0] m300_9;
   assign m300_9 =10'b0;

   // m300_10 = W*in
   wire signed [9:0] m300_10;
   assign m300_10 =10'b0;

   // m300_11 = W*in
   wire signed [9:0] m300_11;
   assign m300_11 =10'b0;

   // m300_12 = W*in
   wire signed [9:0] m300_12;
   assign m300_12 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_13 = W*in
   wire signed [9:0] m300_13;
   assign m300_13 =10'b0;

   // m300_14 = W*in
   wire signed [9:0] m300_14;
   assign m300_14 =10'b0;

   // m300_15 = W*in
   wire signed [9:0] m300_15;
   assign m300_15 ={ {4{in300[5]}} , in300[5:0] };

   // m300_16 = W*in
   wire signed [9:0] m300_16;
   assign m300_16 =10'b0;

   // m300_17 = W*in
   wire signed [9:0] m300_17;
   assign m300_17 =10'b0;

   // m300_18 = W*in
   wire signed [9:0] m300_18;
   assign m300_18 =10'b0;

   // m300_19 = W*in
   wire signed [9:0] m300_19;
   assign m300_19 =10'b0;

   // m300_20 = W*in
   wire signed [9:0] m300_20;
   assign m300_20 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_21 = W*in
   wire signed [9:0] m300_21;
   assign m300_21 ={ {4{in300[5]}} , in300[5:0] };

   // m300_22 = W*in
   wire signed [9:0] m300_22;
   assign m300_22 =10'b0;

   // m300_23 = W*in
   wire signed [9:0] m300_23;
   assign m300_23 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_24 = W*in
   wire signed [9:0] m300_24;
   assign m300_24 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_25 = W*in
   wire signed [9:0] m300_25;
   assign m300_25 ={ {5{in300[5]}} , in300[5:1] };

   // m300_26 = W*in
   wire signed [9:0] m300_26;
   assign m300_26 ={ {4{in300[5]}} , in300[5:0] };

   // m300_27 = W*in
   wire signed [9:0] m300_27;
   assign m300_27 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_28 = W*in
   wire signed [9:0] m300_28;
   assign m300_28 ={ {5{in300[5]}} , in300[5:1] };

   // m300_29 = W*in
   wire signed [9:0] m300_29;
   assign m300_29 =10'b0;

   // m300_30 = W*in
   wire signed [9:0] m300_30;
   assign m300_30 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_31 = W*in
   wire signed [9:0] m300_31;
   assign m300_31 =10'b0;

   // m300_32 = W*in
   wire signed [9:0] m300_32;
   assign m300_32 ={ {4{in300[5]}} , in300[5:0] };

   // m300_33 = W*in
   wire signed [9:0] m300_33;
   assign m300_33 =10'b0;

   // m300_34 = W*in
   wire signed [9:0] m300_34;
   assign m300_34 =10'b0;

   // m300_35 = W*in
   wire signed [9:0] m300_35;
   assign m300_35 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_36 = W*in
   wire signed [9:0] m300_36;
   assign m300_36 =10'b0;

   // m300_37 = W*in
   wire signed [9:0] m300_37;
   assign m300_37 =10'b0;

   // m300_38 = W*in
   wire signed [9:0] m300_38;
   assign m300_38 ={ {4{in300[5]}} , in300[5:0] };

   // m300_39 = W*in
   wire signed [9:0] m300_39;
   assign m300_39 =10'b0;

   // m300_40 = W*in
   wire signed [9:0] m300_40;
   assign m300_40 =10'b0;

   // m300_41 = W*in
   wire signed [9:0] m300_41;
   assign m300_41 =10'b0;

   // m300_42 = W*in
   wire signed [9:0] m300_42;
   assign m300_42 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_43 = W*in
   wire signed [9:0] m300_43;
   assign m300_43 ={ {4{in300[5]}} , in300[5:0] };

   // m300_44 = W*in
   wire signed [9:0] m300_44;
   assign m300_44 =10'b0;

   // m300_45 = W*in
   wire signed [9:0] m300_45;
   assign m300_45 =10'b0;

   // m300_46 = W*in
   wire signed [9:0] m300_46;
   assign m300_46 =10'b0;

   // m300_47 = W*in
   wire signed [9:0] m300_47;
   assign m300_47 ={ {4{in300[5]}} , in300[5:0] };

   // m300_48 = W*in
   wire signed [9:0] m300_48;
   assign m300_48 =10'b0;

   // m300_49 = W*in
   wire signed [9:0] m300_49;
   assign m300_49 =10'b0;

   // m300_50 = W*in
   wire signed [9:0] m300_50;
   assign m300_50 =10'b0;

   // m300_51 = W*in
   wire signed [9:0] m300_51;
   assign m300_51 =10'b0;

   // m300_52 = W*in
   wire signed [9:0] m300_52;
   assign m300_52 =10'b0;

   // m300_53 = W*in
   wire signed [9:0] m300_53;
   assign m300_53 =10'b0;

   // m300_54 = W*in
   wire signed [9:0] m300_54;
   assign m300_54 =10'b0;

   // m300_55 = W*in
   wire signed [9:0] m300_55;
   assign m300_55 ={ {4{in300[5]}} , in300[5:0] };

   // m300_56 = W*in
   wire signed [9:0] m300_56;
   assign m300_56 =10'b0;

   // m300_57 = W*in
   wire signed [9:0] m300_57;
   assign m300_57 =10'b0;

   // m300_58 = W*in
   wire signed [9:0] m300_58;
   assign m300_58 =10'b0;

   // m300_59 = W*in
   wire signed [9:0] m300_59;
   assign m300_59 =10'b0;

   // m300_60 = W*in
   wire signed [9:0] m300_60;
   assign m300_60 =10'b0;

   // m300_61 = W*in
   wire signed [9:0] m300_61;
   assign m300_61 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_62 = W*in
   wire signed [9:0] m300_62;
   assign m300_62 =10'b0;

   // m300_63 = W*in
   wire signed [9:0] m300_63;
   assign m300_63 ={ {4{in300[5]}} , in300[5:0] };

   // m300_64 = W*in
   wire signed [9:0] m300_64;
   assign m300_64 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_65 = W*in
   wire signed [9:0] m300_65;
   assign m300_65 ={ {5{neg300[5]}} , neg300[5:1] };

   // m300_66 = W*in
   wire signed [9:0] m300_66;
   assign m300_66 =10'b0;

   // m300_67 = W*in
   wire signed [9:0] m300_67;
   assign m300_67 ={ {4{in300[5]}} , in300[5:0] };

   // m300_68 = W*in
   wire signed [9:0] m300_68;
   assign m300_68 =10'b0;

   // m300_69 = W*in
   wire signed [9:0] m300_69;
   assign m300_69 ={ {4{in300[5]}} , in300[5:0] };

   // m300_70 = W*in
   wire signed [9:0] m300_70;
   assign m300_70 ={ {5{in300[5]}} , in300[5:1] };

   // m300_71 = W*in
   wire signed [9:0] m300_71;
   assign m300_71 =10'b0;

   // m300_72 = W*in
   wire signed [9:0] m300_72;
   assign m300_72 ={ {4{in300[5]}} , in300[5:0] };

   // m300_73 = W*in
   wire signed [9:0] m300_73;
   assign m300_73 =10'b0;

   // m300_74 = W*in
   wire signed [9:0] m300_74;
   assign m300_74 =10'b0;

   // m300_75 = W*in
   wire signed [9:0] m300_75;
   assign m300_75 =10'b0;

   // m300_76 = W*in
   wire signed [9:0] m300_76;
   assign m300_76 =10'b0;

   // m300_77 = W*in
   wire signed [9:0] m300_77;
   assign m300_77 =10'b0;

   // m300_78 = W*in
   wire signed [9:0] m300_78;
   assign m300_78 ={ {4{in300[5]}} , in300[5:0] };

   // m300_79 = W*in
   wire signed [9:0] m300_79;
   assign m300_79 =10'b0;

   // m300_80 = W*in
   wire signed [9:0] m300_80;
   assign m300_80 =10'b0;

   // m300_81 = W*in
   wire signed [9:0] m300_81;
   assign m300_81 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_82 = W*in
   wire signed [9:0] m300_82;
   assign m300_82 ={ {4{in300[5]}} , in300[5:0] };

   // m300_83 = W*in
   wire signed [9:0] m300_83;
   assign m300_83 =10'b0;

   // m300_84 = W*in
   wire signed [9:0] m300_84;
   assign m300_84 ={ {4{in300[5]}} , in300[5:0] };

   // m300_85 = W*in
   wire signed [9:0] m300_85;
   assign m300_85 ={ {4{in300[5]}} , in300[5:0] };

   // m300_86 = W*in
   wire signed [9:0] m300_86;
   assign m300_86 ={ {4{in300[5]}} , in300[5:0] };

   // m300_87 = W*in
   wire signed [9:0] m300_87;
   assign m300_87 ={ {4{in300[5]}} , in300[5:0] };

   // m300_88 = W*in
   wire signed [9:0] m300_88;
   assign m300_88 ={ {4{in300[5]}} , in300[5:0] };

   // m300_89 = W*in
   wire signed [9:0] m300_89;
   assign m300_89 ={ {4{in300[5]}} , in300[5:0] };

   // m300_90 = W*in
   wire signed [9:0] m300_90;
   assign m300_90 ={ {4{in300[5]}} , in300[5:0] };

   // m300_91 = W*in
   wire signed [9:0] m300_91;
   assign m300_91 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_92 = W*in
   wire signed [9:0] m300_92;
   assign m300_92 ={ {5{in300[5]}} , in300[5:1] };

   // m300_93 = W*in
   wire signed [9:0] m300_93;
   assign m300_93 =10'b0;

   // m300_94 = W*in
   wire signed [9:0] m300_94;
   assign m300_94 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_95 = W*in
   wire signed [9:0] m300_95;
   assign m300_95 =10'b0;

   // m300_96 = W*in
   wire signed [9:0] m300_96;
   assign m300_96 =10'b0;

   // m300_97 = W*in
   wire signed [9:0] m300_97;
   assign m300_97 =10'b0;

   // m300_98 = W*in
   wire signed [9:0] m300_98;
   assign m300_98 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_99 = W*in
   wire signed [9:0] m300_99;
   assign m300_99 =10'b0;

   // m300_100 = W*in
   wire signed [9:0] m300_100;
   assign m300_100 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_101 = W*in
   wire signed [9:0] m300_101;
   assign m300_101 =10'b0;

   // m300_102 = W*in
   wire signed [9:0] m300_102;
   assign m300_102 =10'b0;

   // m300_103 = W*in
   wire signed [9:0] m300_103;
   assign m300_103 =10'b0;

   // m300_104 = W*in
   wire signed [9:0] m300_104;
   assign m300_104 =10'b0;

   // m300_105 = W*in
   wire signed [9:0] m300_105;
   assign m300_105 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_106 = W*in
   wire signed [9:0] m300_106;
   assign m300_106 =10'b0;

   // m300_107 = W*in
   wire signed [9:0] m300_107;
   assign m300_107 =10'b0;

   // m300_108 = W*in
   wire signed [9:0] m300_108;
   assign m300_108 ={ {5{neg300[5]}} , neg300[5:1] };

   // m300_109 = W*in
   wire signed [9:0] m300_109;
   assign m300_109 ={ {5{neg300[5]}} , neg300[5:1] };

   // m300_110 = W*in
   wire signed [9:0] m300_110;
   assign m300_110 =10'b0;

   // m300_111 = W*in
   wire signed [9:0] m300_111;
   assign m300_111 ={ {4{in300[5]}} , in300[5:0] };

   // m300_112 = W*in
   wire signed [9:0] m300_112;
   assign m300_112 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_113 = W*in
   wire signed [9:0] m300_113;
   assign m300_113 =10'b0;

   // m300_114 = W*in
   wire signed [9:0] m300_114;
   assign m300_114 ={ {5{neg300[5]}} , neg300[5:1] };

   // m300_115 = W*in
   wire signed [9:0] m300_115;
   assign m300_115 ={ {4{neg300[5]}} , neg300[5:0] };

   // m300_116 = W*in
   wire signed [9:0] m300_116;
   assign m300_116 =10'b0;

   // m300_117 = W*in
   wire signed [9:0] m300_117;
   assign m300_117 ={ {4{neg300[5]}} , neg300[5:0] };

   // m301_1 = W*in
   wire signed [9:0] m301_1;
   assign m301_1 =10'b0;

   // m301_2 = W*in
   wire signed [9:0] m301_2;
   assign m301_2 =10'b0;

   // m301_3 = W*in
   wire signed [9:0] m301_3;
   assign m301_3 =10'b0;

   // m301_4 = W*in
   wire signed [9:0] m301_4;
   assign m301_4 =10'b0;

   // m301_5 = W*in
   wire signed [9:0] m301_5;
   assign m301_5 =10'b0;

   // m301_6 = W*in
   wire signed [9:0] m301_6;
   assign m301_6 =10'b0;

   // m301_7 = W*in
   wire signed [9:0] m301_7;
   assign m301_7 ={ {4{in301[5]}} , in301[5:0] };

   // m301_8 = W*in
   wire signed [9:0] m301_8;
   assign m301_8 =10'b0;

   // m301_9 = W*in
   wire signed [9:0] m301_9;
   assign m301_9 =10'b0;

   // m301_10 = W*in
   wire signed [9:0] m301_10;
   assign m301_10 =10'b0;

   // m301_11 = W*in
   wire signed [9:0] m301_11;
   assign m301_11 =10'b0;

   // m301_12 = W*in
   wire signed [9:0] m301_12;
   assign m301_12 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_13 = W*in
   wire signed [9:0] m301_13;
   assign m301_13 =10'b0;

   // m301_14 = W*in
   wire signed [9:0] m301_14;
   assign m301_14 =10'b0;

   // m301_15 = W*in
   wire signed [9:0] m301_15;
   assign m301_15 =10'b0;

   // m301_16 = W*in
   wire signed [9:0] m301_16;
   assign m301_16 =10'b0;

   // m301_17 = W*in
   wire signed [9:0] m301_17;
   assign m301_17 =10'b0;

   // m301_18 = W*in
   wire signed [9:0] m301_18;
   assign m301_18 ={ {4{in301[5]}} , in301[5:0] };

   // m301_19 = W*in
   wire signed [9:0] m301_19;
   assign m301_19 =10'b0;

   // m301_20 = W*in
   wire signed [9:0] m301_20;
   assign m301_20 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_21 = W*in
   wire signed [9:0] m301_21;
   assign m301_21 =10'b0;

   // m301_22 = W*in
   wire signed [9:0] m301_22;
   assign m301_22 =10'b0;

   // m301_23 = W*in
   wire signed [9:0] m301_23;
   assign m301_23 =10'b0;

   // m301_24 = W*in
   wire signed [9:0] m301_24;
   assign m301_24 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_25 = W*in
   wire signed [9:0] m301_25;
   assign m301_25 ={ {4{in301[5]}} , in301[5:0] };

   // m301_26 = W*in
   wire signed [9:0] m301_26;
   assign m301_26 =10'b0;

   // m301_27 = W*in
   wire signed [9:0] m301_27;
   assign m301_27 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_28 = W*in
   wire signed [9:0] m301_28;
   assign m301_28 ={ {4{in301[5]}} , in301[5:0] };

   // m301_29 = W*in
   wire signed [9:0] m301_29;
   assign m301_29 =10'b0;

   // m301_30 = W*in
   wire signed [9:0] m301_30;
   assign m301_30 =10'b0;

   // m301_31 = W*in
   wire signed [9:0] m301_31;
   assign m301_31 =10'b0;

   // m301_32 = W*in
   wire signed [9:0] m301_32;
   assign m301_32 =10'b0;

   // m301_33 = W*in
   wire signed [9:0] m301_33;
   assign m301_33 ={ {4{in301[5]}} , in301[5:0] };

   // m301_34 = W*in
   wire signed [9:0] m301_34;
   assign m301_34 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_35 = W*in
   wire signed [9:0] m301_35;
   assign m301_35 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_36 = W*in
   wire signed [9:0] m301_36;
   assign m301_36 =10'b0;

   // m301_37 = W*in
   wire signed [9:0] m301_37;
   assign m301_37 =10'b0;

   // m301_38 = W*in
   wire signed [9:0] m301_38;
   assign m301_38 =10'b0;

   // m301_39 = W*in
   wire signed [9:0] m301_39;
   assign m301_39 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_40 = W*in
   wire signed [9:0] m301_40;
   assign m301_40 =10'b0;

   // m301_41 = W*in
   wire signed [9:0] m301_41;
   assign m301_41 =10'b0;

   // m301_42 = W*in
   wire signed [9:0] m301_42;
   assign m301_42 =10'b0;

   // m301_43 = W*in
   wire signed [9:0] m301_43;
   assign m301_43 ={ {4{in301[5]}} , in301[5:0] };

   // m301_44 = W*in
   wire signed [9:0] m301_44;
   assign m301_44 =10'b0;

   // m301_45 = W*in
   wire signed [9:0] m301_45;
   assign m301_45 =10'b0;

   // m301_46 = W*in
   wire signed [9:0] m301_46;
   assign m301_46 =10'b0;

   // m301_47 = W*in
   wire signed [9:0] m301_47;
   assign m301_47 =10'b0;

   // m301_48 = W*in
   wire signed [9:0] m301_48;
   assign m301_48 ={ {4{in301[5]}} , in301[5:0] };

   // m301_49 = W*in
   wire signed [9:0] m301_49;
   assign m301_49 =10'b0;

   // m301_50 = W*in
   wire signed [9:0] m301_50;
   assign m301_50 =10'b0;

   // m301_51 = W*in
   wire signed [9:0] m301_51;
   assign m301_51 =10'b0;

   // m301_52 = W*in
   wire signed [9:0] m301_52;
   assign m301_52 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_53 = W*in
   wire signed [9:0] m301_53;
   assign m301_53 =10'b0;

   // m301_54 = W*in
   wire signed [9:0] m301_54;
   assign m301_54 =10'b0;

   // m301_55 = W*in
   wire signed [9:0] m301_55;
   assign m301_55 =10'b0;

   // m301_56 = W*in
   wire signed [9:0] m301_56;
   assign m301_56 =10'b0;

   // m301_57 = W*in
   wire signed [9:0] m301_57;
   assign m301_57 =10'b0;

   // m301_58 = W*in
   wire signed [9:0] m301_58;
   assign m301_58 =10'b0;

   // m301_59 = W*in
   wire signed [9:0] m301_59;
   assign m301_59 ={ {4{in301[5]}} , in301[5:0] };

   // m301_60 = W*in
   wire signed [9:0] m301_60;
   assign m301_60 =10'b0;

   // m301_61 = W*in
   wire signed [9:0] m301_61;
   assign m301_61 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_62 = W*in
   wire signed [9:0] m301_62;
   assign m301_62 =10'b0;

   // m301_63 = W*in
   wire signed [9:0] m301_63;
   assign m301_63 =10'b0;

   // m301_64 = W*in
   wire signed [9:0] m301_64;
   assign m301_64 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_65 = W*in
   wire signed [9:0] m301_65;
   assign m301_65 =10'b0;

   // m301_66 = W*in
   wire signed [9:0] m301_66;
   assign m301_66 =10'b0;

   // m301_67 = W*in
   wire signed [9:0] m301_67;
   assign m301_67 ={ {4{in301[5]}} , in301[5:0] };

   // m301_68 = W*in
   wire signed [9:0] m301_68;
   assign m301_68 =10'b0;

   // m301_69 = W*in
   wire signed [9:0] m301_69;
   assign m301_69 =10'b0;

   // m301_70 = W*in
   wire signed [9:0] m301_70;
   assign m301_70 =10'b0;

   // m301_71 = W*in
   wire signed [9:0] m301_71;
   assign m301_71 ={ {5{in301[5]}} , in301[5:1] };

   // m301_72 = W*in
   wire signed [9:0] m301_72;
   assign m301_72 ={ {4{in301[5]}} , in301[5:0] };

   // m301_73 = W*in
   wire signed [9:0] m301_73;
   assign m301_73 =10'b0;

   // m301_74 = W*in
   wire signed [9:0] m301_74;
   assign m301_74 =10'b0;

   // m301_75 = W*in
   wire signed [9:0] m301_75;
   assign m301_75 =10'b0;

   // m301_76 = W*in
   wire signed [9:0] m301_76;
   assign m301_76 =10'b0;

   // m301_77 = W*in
   wire signed [9:0] m301_77;
   assign m301_77 =10'b0;

   // m301_78 = W*in
   wire signed [9:0] m301_78;
   assign m301_78 =10'b0;

   // m301_79 = W*in
   wire signed [9:0] m301_79;
   assign m301_79 =10'b0;

   // m301_80 = W*in
   wire signed [9:0] m301_80;
   assign m301_80 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_81 = W*in
   wire signed [9:0] m301_81;
   assign m301_81 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_82 = W*in
   wire signed [9:0] m301_82;
   assign m301_82 =10'b0;

   // m301_83 = W*in
   wire signed [9:0] m301_83;
   assign m301_83 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_84 = W*in
   wire signed [9:0] m301_84;
   assign m301_84 ={ {4{in301[5]}} , in301[5:0] };

   // m301_85 = W*in
   wire signed [9:0] m301_85;
   assign m301_85 =10'b0;

   // m301_86 = W*in
   wire signed [9:0] m301_86;
   assign m301_86 =10'b0;

   // m301_87 = W*in
   wire signed [9:0] m301_87;
   assign m301_87 =10'b0;

   // m301_88 = W*in
   wire signed [9:0] m301_88;
   assign m301_88 =10'b0;

   // m301_89 = W*in
   wire signed [9:0] m301_89;
   assign m301_89 =10'b0;

   // m301_90 = W*in
   wire signed [9:0] m301_90;
   assign m301_90 =10'b0;

   // m301_91 = W*in
   wire signed [9:0] m301_91;
   assign m301_91 =10'b0;

   // m301_92 = W*in
   wire signed [9:0] m301_92;
   assign m301_92 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_93 = W*in
   wire signed [9:0] m301_93;
   assign m301_93 =10'b0;

   // m301_94 = W*in
   wire signed [9:0] m301_94;
   assign m301_94 =10'b0;

   // m301_95 = W*in
   wire signed [9:0] m301_95;
   assign m301_95 =10'b0;

   // m301_96 = W*in
   wire signed [9:0] m301_96;
   assign m301_96 =10'b0;

   // m301_97 = W*in
   wire signed [9:0] m301_97;
   assign m301_97 =10'b0;

   // m301_98 = W*in
   wire signed [9:0] m301_98;
   assign m301_98 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_99 = W*in
   wire signed [9:0] m301_99;
   assign m301_99 =10'b0;

   // m301_100 = W*in
   wire signed [9:0] m301_100;
   assign m301_100 =10'b0;

   // m301_101 = W*in
   wire signed [9:0] m301_101;
   assign m301_101 =10'b0;

   // m301_102 = W*in
   wire signed [9:0] m301_102;
   assign m301_102 ={ {4{in301[5]}} , in301[5:0] };

   // m301_103 = W*in
   wire signed [9:0] m301_103;
   assign m301_103 =10'b0;

   // m301_104 = W*in
   wire signed [9:0] m301_104;
   assign m301_104 =10'b0;

   // m301_105 = W*in
   wire signed [9:0] m301_105;
   assign m301_105 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_106 = W*in
   wire signed [9:0] m301_106;
   assign m301_106 =10'b0;

   // m301_107 = W*in
   wire signed [9:0] m301_107;
   assign m301_107 =10'b0;

   // m301_108 = W*in
   wire signed [9:0] m301_108;
   assign m301_108 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_109 = W*in
   wire signed [9:0] m301_109;
   assign m301_109 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_110 = W*in
   wire signed [9:0] m301_110;
   assign m301_110 =10'b0;

   // m301_111 = W*in
   wire signed [9:0] m301_111;
   assign m301_111 =10'b0;

   // m301_112 = W*in
   wire signed [9:0] m301_112;
   assign m301_112 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_113 = W*in
   wire signed [9:0] m301_113;
   assign m301_113 =10'b0;

   // m301_114 = W*in
   wire signed [9:0] m301_114;
   assign m301_114 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_115 = W*in
   wire signed [9:0] m301_115;
   assign m301_115 ={ {5{neg301[5]}} , neg301[5:1] };

   // m301_116 = W*in
   wire signed [9:0] m301_116;
   assign m301_116 ={ {4{neg301[5]}} , neg301[5:0] };

   // m301_117 = W*in
   wire signed [9:0] m301_117;
   assign m301_117 =10'b0;

   // m302_1 = W*in
   wire signed [9:0] m302_1;
   assign m302_1 ={ {4{in302[5]}} , in302[5:0] };

   // m302_2 = W*in
   wire signed [9:0] m302_2;
   assign m302_2 =10'b0;

   // m302_3 = W*in
   wire signed [9:0] m302_3;
   assign m302_3 =10'b0;

   // m302_4 = W*in
   wire signed [9:0] m302_4;
   assign m302_4 =10'b0;

   // m302_5 = W*in
   wire signed [9:0] m302_5;
   assign m302_5 =10'b0;

   // m302_6 = W*in
   wire signed [9:0] m302_6;
   assign m302_6 =10'b0;

   // m302_7 = W*in
   wire signed [9:0] m302_7;
   assign m302_7 ={ {4{in302[5]}} , in302[5:0] };

   // m302_8 = W*in
   wire signed [9:0] m302_8;
   assign m302_8 =10'b0;

   // m302_9 = W*in
   wire signed [9:0] m302_9;
   assign m302_9 =10'b0;

   // m302_10 = W*in
   wire signed [9:0] m302_10;
   assign m302_10 =10'b0;

   // m302_11 = W*in
   wire signed [9:0] m302_11;
   assign m302_11 =10'b0;

   // m302_12 = W*in
   wire signed [9:0] m302_12;
   assign m302_12 =10'b0;

   // m302_13 = W*in
   wire signed [9:0] m302_13;
   assign m302_13 =10'b0;

   // m302_14 = W*in
   wire signed [9:0] m302_14;
   assign m302_14 =10'b0;

   // m302_15 = W*in
   wire signed [9:0] m302_15;
   assign m302_15 =10'b0;

   // m302_16 = W*in
   wire signed [9:0] m302_16;
   assign m302_16 =10'b0;

   // m302_17 = W*in
   wire signed [9:0] m302_17;
   assign m302_17 =10'b0;

   // m302_18 = W*in
   wire signed [9:0] m302_18;
   assign m302_18 ={ {5{in302[5]}} , in302[5:1] };

   // m302_19 = W*in
   wire signed [9:0] m302_19;
   assign m302_19 =10'b0;

   // m302_20 = W*in
   wire signed [9:0] m302_20;
   assign m302_20 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_21 = W*in
   wire signed [9:0] m302_21;
   assign m302_21 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_22 = W*in
   wire signed [9:0] m302_22;
   assign m302_22 =10'b0;

   // m302_23 = W*in
   wire signed [9:0] m302_23;
   assign m302_23 =10'b0;

   // m302_24 = W*in
   wire signed [9:0] m302_24;
   assign m302_24 =10'b0;

   // m302_25 = W*in
   wire signed [9:0] m302_25;
   assign m302_25 ={ {5{in302[5]}} , in302[5:1] };

   // m302_26 = W*in
   wire signed [9:0] m302_26;
   assign m302_26 =10'b0;

   // m302_27 = W*in
   wire signed [9:0] m302_27;
   assign m302_27 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_28 = W*in
   wire signed [9:0] m302_28;
   assign m302_28 ={ {4{in302[5]}} , in302[5:0] };

   // m302_29 = W*in
   wire signed [9:0] m302_29;
   assign m302_29 =10'b0;

   // m302_30 = W*in
   wire signed [9:0] m302_30;
   assign m302_30 =10'b0;

   // m302_31 = W*in
   wire signed [9:0] m302_31;
   assign m302_31 =10'b0;

   // m302_32 = W*in
   wire signed [9:0] m302_32;
   assign m302_32 =10'b0;

   // m302_33 = W*in
   wire signed [9:0] m302_33;
   assign m302_33 ={ {4{in302[5]}} , in302[5:0] };

   // m302_34 = W*in
   wire signed [9:0] m302_34;
   assign m302_34 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_35 = W*in
   wire signed [9:0] m302_35;
   assign m302_35 =10'b0;

   // m302_36 = W*in
   wire signed [9:0] m302_36;
   assign m302_36 =10'b0;

   // m302_37 = W*in
   wire signed [9:0] m302_37;
   assign m302_37 =10'b0;

   // m302_38 = W*in
   wire signed [9:0] m302_38;
   assign m302_38 =10'b0;

   // m302_39 = W*in
   wire signed [9:0] m302_39;
   assign m302_39 =10'b0;

   // m302_40 = W*in
   wire signed [9:0] m302_40;
   assign m302_40 =10'b0;

   // m302_41 = W*in
   wire signed [9:0] m302_41;
   assign m302_41 =10'b0;

   // m302_42 = W*in
   wire signed [9:0] m302_42;
   assign m302_42 =10'b0;

   // m302_43 = W*in
   wire signed [9:0] m302_43;
   assign m302_43 =10'b0;

   // m302_44 = W*in
   wire signed [9:0] m302_44;
   assign m302_44 =10'b0;

   // m302_45 = W*in
   wire signed [9:0] m302_45;
   assign m302_45 =10'b0;

   // m302_46 = W*in
   wire signed [9:0] m302_46;
   assign m302_46 =10'b0;

   // m302_47 = W*in
   wire signed [9:0] m302_47;
   assign m302_47 =10'b0;

   // m302_48 = W*in
   wire signed [9:0] m302_48;
   assign m302_48 =10'b0;

   // m302_49 = W*in
   wire signed [9:0] m302_49;
   assign m302_49 =10'b0;

   // m302_50 = W*in
   wire signed [9:0] m302_50;
   assign m302_50 =10'b0;

   // m302_51 = W*in
   wire signed [9:0] m302_51;
   assign m302_51 =10'b0;

   // m302_52 = W*in
   wire signed [9:0] m302_52;
   assign m302_52 =10'b0;

   // m302_53 = W*in
   wire signed [9:0] m302_53;
   assign m302_53 =10'b0;

   // m302_54 = W*in
   wire signed [9:0] m302_54;
   assign m302_54 =10'b0;

   // m302_55 = W*in
   wire signed [9:0] m302_55;
   assign m302_55 =10'b0;

   // m302_56 = W*in
   wire signed [9:0] m302_56;
   assign m302_56 =10'b0;

   // m302_57 = W*in
   wire signed [9:0] m302_57;
   assign m302_57 =10'b0;

   // m302_58 = W*in
   wire signed [9:0] m302_58;
   assign m302_58 =10'b0;

   // m302_59 = W*in
   wire signed [9:0] m302_59;
   assign m302_59 =10'b0;

   // m302_60 = W*in
   wire signed [9:0] m302_60;
   assign m302_60 =10'b0;

   // m302_61 = W*in
   wire signed [9:0] m302_61;
   assign m302_61 =10'b0;

   // m302_62 = W*in
   wire signed [9:0] m302_62;
   assign m302_62 =10'b0;

   // m302_63 = W*in
   wire signed [9:0] m302_63;
   assign m302_63 ={ {4{neg302[5]}} , neg302[5:0] };

   // m302_64 = W*in
   wire signed [9:0] m302_64;
   assign m302_64 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_65 = W*in
   wire signed [9:0] m302_65;
   assign m302_65 =10'b0;

   // m302_66 = W*in
   wire signed [9:0] m302_66;
   assign m302_66 =10'b0;

   // m302_67 = W*in
   wire signed [9:0] m302_67;
   assign m302_67 =10'b0;

   // m302_68 = W*in
   wire signed [9:0] m302_68;
   assign m302_68 =10'b0;

   // m302_69 = W*in
   wire signed [9:0] m302_69;
   assign m302_69 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_70 = W*in
   wire signed [9:0] m302_70;
   assign m302_70 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_71 = W*in
   wire signed [9:0] m302_71;
   assign m302_71 =10'b0;

   // m302_72 = W*in
   wire signed [9:0] m302_72;
   assign m302_72 =10'b0;

   // m302_73 = W*in
   wire signed [9:0] m302_73;
   assign m302_73 ={ {5{in302[5]}} , in302[5:1] };

   // m302_74 = W*in
   wire signed [9:0] m302_74;
   assign m302_74 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_75 = W*in
   wire signed [9:0] m302_75;
   assign m302_75 =10'b0;

   // m302_76 = W*in
   wire signed [9:0] m302_76;
   assign m302_76 =10'b0;

   // m302_77 = W*in
   wire signed [9:0] m302_77;
   assign m302_77 =10'b0;

   // m302_78 = W*in
   wire signed [9:0] m302_78;
   assign m302_78 =10'b0;

   // m302_79 = W*in
   wire signed [9:0] m302_79;
   assign m302_79 =10'b0;

   // m302_80 = W*in
   wire signed [9:0] m302_80;
   assign m302_80 =10'b0;

   // m302_81 = W*in
   wire signed [9:0] m302_81;
   assign m302_81 =10'b0;

   // m302_82 = W*in
   wire signed [9:0] m302_82;
   assign m302_82 ={ {4{neg302[5]}} , neg302[5:0] };

   // m302_83 = W*in
   wire signed [9:0] m302_83;
   assign m302_83 =10'b0;

   // m302_84 = W*in
   wire signed [9:0] m302_84;
   assign m302_84 ={ {5{in302[5]}} , in302[5:1] };

   // m302_85 = W*in
   wire signed [9:0] m302_85;
   assign m302_85 =10'b0;

   // m302_86 = W*in
   wire signed [9:0] m302_86;
   assign m302_86 =10'b0;

   // m302_87 = W*in
   wire signed [9:0] m302_87;
   assign m302_87 =10'b0;

   // m302_88 = W*in
   wire signed [9:0] m302_88;
   assign m302_88 =10'b0;

   // m302_89 = W*in
   wire signed [9:0] m302_89;
   assign m302_89 =10'b0;

   // m302_90 = W*in
   wire signed [9:0] m302_90;
   assign m302_90 =10'b0;

   // m302_91 = W*in
   wire signed [9:0] m302_91;
   assign m302_91 ={ {4{neg302[5]}} , neg302[5:0] };

   // m302_92 = W*in
   wire signed [9:0] m302_92;
   assign m302_92 =10'b0;

   // m302_93 = W*in
   wire signed [9:0] m302_93;
   assign m302_93 =10'b0;

   // m302_94 = W*in
   wire signed [9:0] m302_94;
   assign m302_94 =10'b0;

   // m302_95 = W*in
   wire signed [9:0] m302_95;
   assign m302_95 =10'b0;

   // m302_96 = W*in
   wire signed [9:0] m302_96;
   assign m302_96 =10'b0;

   // m302_97 = W*in
   wire signed [9:0] m302_97;
   assign m302_97 =10'b0;

   // m302_98 = W*in
   wire signed [9:0] m302_98;
   assign m302_98 =10'b0;

   // m302_99 = W*in
   wire signed [9:0] m302_99;
   assign m302_99 =10'b0;

   // m302_100 = W*in
   wire signed [9:0] m302_100;
   assign m302_100 =10'b0;

   // m302_101 = W*in
   wire signed [9:0] m302_101;
   assign m302_101 =10'b0;

   // m302_102 = W*in
   wire signed [9:0] m302_102;
   assign m302_102 =10'b0;

   // m302_103 = W*in
   wire signed [9:0] m302_103;
   assign m302_103 =10'b0;

   // m302_104 = W*in
   wire signed [9:0] m302_104;
   assign m302_104 =10'b0;

   // m302_105 = W*in
   wire signed [9:0] m302_105;
   assign m302_105 =10'b0;

   // m302_106 = W*in
   wire signed [9:0] m302_106;
   assign m302_106 =10'b0;

   // m302_107 = W*in
   wire signed [9:0] m302_107;
   assign m302_107 =10'b0;

   // m302_108 = W*in
   wire signed [9:0] m302_108;
   assign m302_108 ={ {5{neg302[5]}} , neg302[5:1] };

   // m302_109 = W*in
   wire signed [9:0] m302_109;
   assign m302_109 =10'b0;

   // m302_110 = W*in
   wire signed [9:0] m302_110;
   assign m302_110 =10'b0;

   // m302_111 = W*in
   wire signed [9:0] m302_111;
   assign m302_111 =10'b0;

   // m302_112 = W*in
   wire signed [9:0] m302_112;
   assign m302_112 ={ {4{neg302[5]}} , neg302[5:0] };

   // m302_113 = W*in
   wire signed [9:0] m302_113;
   assign m302_113 =10'b0;

   // m302_114 = W*in
   wire signed [9:0] m302_114;
   assign m302_114 =10'b0;

   // m302_115 = W*in
   wire signed [9:0] m302_115;
   assign m302_115 =10'b0;

   // m302_116 = W*in
   wire signed [9:0] m302_116;
   assign m302_116 =10'b0;

   // m302_117 = W*in
   wire signed [9:0] m302_117;
   assign m302_117 =10'b0;

   // m303_1 = W*in
   wire signed [9:0] m303_1;
   assign m303_1 =10'b0;

   // m303_2 = W*in
   wire signed [9:0] m303_2;
   assign m303_2 =10'b0;

   // m303_3 = W*in
   wire signed [9:0] m303_3;
   assign m303_3 ={ {4{in303[5]}} , in303[5:0] };

   // m303_4 = W*in
   wire signed [9:0] m303_4;
   assign m303_4 =10'b0;

   // m303_5 = W*in
   wire signed [9:0] m303_5;
   assign m303_5 =10'b0;

   // m303_6 = W*in
   wire signed [9:0] m303_6;
   assign m303_6 =10'b0;

   // m303_7 = W*in
   wire signed [9:0] m303_7;
   assign m303_7 =10'b0;

   // m303_8 = W*in
   wire signed [9:0] m303_8;
   assign m303_8 =10'b0;

   // m303_9 = W*in
   wire signed [9:0] m303_9;
   assign m303_9 =10'b0;

   // m303_10 = W*in
   wire signed [9:0] m303_10;
   assign m303_10 =10'b0;

   // m303_11 = W*in
   wire signed [9:0] m303_11;
   assign m303_11 =10'b0;

   // m303_12 = W*in
   wire signed [9:0] m303_12;
   assign m303_12 ={ {4{in303[5]}} , in303[5:0] };

   // m303_13 = W*in
   wire signed [9:0] m303_13;
   assign m303_13 =10'b0;

   // m303_14 = W*in
   wire signed [9:0] m303_14;
   assign m303_14 =10'b0;

   // m303_15 = W*in
   wire signed [9:0] m303_15;
   assign m303_15 =10'b0;

   // m303_16 = W*in
   wire signed [9:0] m303_16;
   assign m303_16 =10'b0;

   // m303_17 = W*in
   wire signed [9:0] m303_17;
   assign m303_17 ={ {5{in303[5]}} , in303[5:1] };

   // m303_18 = W*in
   wire signed [9:0] m303_18;
   assign m303_18 =10'b0;

   // m303_19 = W*in
   wire signed [9:0] m303_19;
   assign m303_19 =10'b0;

   // m303_20 = W*in
   wire signed [9:0] m303_20;
   assign m303_20 =10'b0;

   // m303_21 = W*in
   wire signed [9:0] m303_21;
   assign m303_21 ={ {4{neg303[5]}} , neg303[5:0] };

   // m303_22 = W*in
   wire signed [9:0] m303_22;
   assign m303_22 =10'b0;

   // m303_23 = W*in
   wire signed [9:0] m303_23;
   assign m303_23 =10'b0;

   // m303_24 = W*in
   wire signed [9:0] m303_24;
   assign m303_24 =10'b0;

   // m303_25 = W*in
   wire signed [9:0] m303_25;
   assign m303_25 ={ {5{in303[5]}} , in303[5:1] };

   // m303_26 = W*in
   wire signed [9:0] m303_26;
   assign m303_26 =10'b0;

   // m303_27 = W*in
   wire signed [9:0] m303_27;
   assign m303_27 =10'b0;

   // m303_28 = W*in
   wire signed [9:0] m303_28;
   assign m303_28 ={ {5{in303[5]}} , in303[5:1] };

   // m303_29 = W*in
   wire signed [9:0] m303_29;
   assign m303_29 =10'b0;

   // m303_30 = W*in
   wire signed [9:0] m303_30;
   assign m303_30 =10'b0;

   // m303_31 = W*in
   wire signed [9:0] m303_31;
   assign m303_31 =10'b0;

   // m303_32 = W*in
   wire signed [9:0] m303_32;
   assign m303_32 =10'b0;

   // m303_33 = W*in
   wire signed [9:0] m303_33;
   assign m303_33 =10'b0;

   // m303_34 = W*in
   wire signed [9:0] m303_34;
   assign m303_34 =10'b0;

   // m303_35 = W*in
   wire signed [9:0] m303_35;
   assign m303_35 =10'b0;

   // m303_36 = W*in
   wire signed [9:0] m303_36;
   assign m303_36 ={ {4{in303[5]}} , in303[5:0] };

   // m303_37 = W*in
   wire signed [9:0] m303_37;
   assign m303_37 =10'b0;

   // m303_38 = W*in
   wire signed [9:0] m303_38;
   assign m303_38 =10'b0;

   // m303_39 = W*in
   wire signed [9:0] m303_39;
   assign m303_39 =10'b0;

   // m303_40 = W*in
   wire signed [9:0] m303_40;
   assign m303_40 =10'b0;

   // m303_41 = W*in
   wire signed [9:0] m303_41;
   assign m303_41 =10'b0;

   // m303_42 = W*in
   wire signed [9:0] m303_42;
   assign m303_42 =10'b0;

   // m303_43 = W*in
   wire signed [9:0] m303_43;
   assign m303_43 =10'b0;

   // m303_44 = W*in
   wire signed [9:0] m303_44;
   assign m303_44 =10'b0;

   // m303_45 = W*in
   wire signed [9:0] m303_45;
   assign m303_45 =10'b0;

   // m303_46 = W*in
   wire signed [9:0] m303_46;
   assign m303_46 =10'b0;

   // m303_47 = W*in
   wire signed [9:0] m303_47;
   assign m303_47 =10'b0;

   // m303_48 = W*in
   wire signed [9:0] m303_48;
   assign m303_48 =10'b0;

   // m303_49 = W*in
   wire signed [9:0] m303_49;
   assign m303_49 =10'b0;

   // m303_50 = W*in
   wire signed [9:0] m303_50;
   assign m303_50 =10'b0;

   // m303_51 = W*in
   wire signed [9:0] m303_51;
   assign m303_51 =10'b0;

   // m303_52 = W*in
   wire signed [9:0] m303_52;
   assign m303_52 =10'b0;

   // m303_53 = W*in
   wire signed [9:0] m303_53;
   assign m303_53 =10'b0;

   // m303_54 = W*in
   wire signed [9:0] m303_54;
   assign m303_54 =10'b0;

   // m303_55 = W*in
   wire signed [9:0] m303_55;
   assign m303_55 =10'b0;

   // m303_56 = W*in
   wire signed [9:0] m303_56;
   assign m303_56 =10'b0;

   // m303_57 = W*in
   wire signed [9:0] m303_57;
   assign m303_57 =10'b0;

   // m303_58 = W*in
   wire signed [9:0] m303_58;
   assign m303_58 =10'b0;

   // m303_59 = W*in
   wire signed [9:0] m303_59;
   assign m303_59 =10'b0;

   // m303_60 = W*in
   wire signed [9:0] m303_60;
   assign m303_60 =10'b0;

   // m303_61 = W*in
   wire signed [9:0] m303_61;
   assign m303_61 =10'b0;

   // m303_62 = W*in
   wire signed [9:0] m303_62;
   assign m303_62 =10'b0;

   // m303_63 = W*in
   wire signed [9:0] m303_63;
   assign m303_63 =10'b0;

   // m303_64 = W*in
   wire signed [9:0] m303_64;
   assign m303_64 =10'b0;

   // m303_65 = W*in
   wire signed [9:0] m303_65;
   assign m303_65 ={ {5{neg303[5]}} , neg303[5:1] };

   // m303_66 = W*in
   wire signed [9:0] m303_66;
   assign m303_66 ={ {5{in303[5]}} , in303[5:1] };

   // m303_67 = W*in
   wire signed [9:0] m303_67;
   assign m303_67 ={ {4{neg303[5]}} , neg303[5:0] };

   // m303_68 = W*in
   wire signed [9:0] m303_68;
   assign m303_68 =10'b0;

   // m303_69 = W*in
   wire signed [9:0] m303_69;
   assign m303_69 ={ {5{neg303[5]}} , neg303[5:1] };

   // m303_70 = W*in
   wire signed [9:0] m303_70;
   assign m303_70 ={ {5{neg303[5]}} , neg303[5:1] };

   // m303_71 = W*in
   wire signed [9:0] m303_71;
   assign m303_71 ={ {5{in303[5]}} , in303[5:1] };

   // m303_72 = W*in
   wire signed [9:0] m303_72;
   assign m303_72 ={ {5{neg303[5]}} , neg303[5:1] };

   // m303_73 = W*in
   wire signed [9:0] m303_73;
   assign m303_73 ={ {4{in303[5]}} , in303[5:0] };

   // m303_74 = W*in
   wire signed [9:0] m303_74;
   assign m303_74 =10'b0;

   // m303_75 = W*in
   wire signed [9:0] m303_75;
   assign m303_75 =10'b0;

   // m303_76 = W*in
   wire signed [9:0] m303_76;
   assign m303_76 =10'b0;

   // m303_77 = W*in
   wire signed [9:0] m303_77;
   assign m303_77 =10'b0;

   // m303_78 = W*in
   wire signed [9:0] m303_78;
   assign m303_78 =10'b0;

   // m303_79 = W*in
   wire signed [9:0] m303_79;
   assign m303_79 =10'b0;

   // m303_80 = W*in
   wire signed [9:0] m303_80;
   assign m303_80 =10'b0;

   // m303_81 = W*in
   wire signed [9:0] m303_81;
   assign m303_81 =10'b0;

   // m303_82 = W*in
   wire signed [9:0] m303_82;
   assign m303_82 ={ {4{neg303[5]}} , neg303[5:0] };

   // m303_83 = W*in
   wire signed [9:0] m303_83;
   assign m303_83 =10'b0;

   // m303_84 = W*in
   wire signed [9:0] m303_84;
   assign m303_84 ={ {5{neg303[5]}} , neg303[5:1] };

   // m303_85 = W*in
   wire signed [9:0] m303_85;
   assign m303_85 =10'b0;

   // m303_86 = W*in
   wire signed [9:0] m303_86;
   assign m303_86 =10'b0;

   // m303_87 = W*in
   wire signed [9:0] m303_87;
   assign m303_87 =10'b0;

   // m303_88 = W*in
   wire signed [9:0] m303_88;
   assign m303_88 =10'b0;

   // m303_89 = W*in
   wire signed [9:0] m303_89;
   assign m303_89 =10'b0;

   // m303_90 = W*in
   wire signed [9:0] m303_90;
   assign m303_90 =10'b0;

   // m303_91 = W*in
   wire signed [9:0] m303_91;
   assign m303_91 =10'b0;

   // m303_92 = W*in
   wire signed [9:0] m303_92;
   assign m303_92 =10'b0;

   // m303_93 = W*in
   wire signed [9:0] m303_93;
   assign m303_93 =10'b0;

   // m303_94 = W*in
   wire signed [9:0] m303_94;
   assign m303_94 =10'b0;

   // m303_95 = W*in
   wire signed [9:0] m303_95;
   assign m303_95 =10'b0;

   // m303_96 = W*in
   wire signed [9:0] m303_96;
   assign m303_96 =10'b0;

   // m303_97 = W*in
   wire signed [9:0] m303_97;
   assign m303_97 =10'b0;

   // m303_98 = W*in
   wire signed [9:0] m303_98;
   assign m303_98 =10'b0;

   // m303_99 = W*in
   wire signed [9:0] m303_99;
   assign m303_99 =10'b0;

   // m303_100 = W*in
   wire signed [9:0] m303_100;
   assign m303_100 =10'b0;

   // m303_101 = W*in
   wire signed [9:0] m303_101;
   assign m303_101 =10'b0;

   // m303_102 = W*in
   wire signed [9:0] m303_102;
   assign m303_102 =10'b0;

   // m303_103 = W*in
   wire signed [9:0] m303_103;
   assign m303_103 =10'b0;

   // m303_104 = W*in
   wire signed [9:0] m303_104;
   assign m303_104 =10'b0;

   // m303_105 = W*in
   wire signed [9:0] m303_105;
   assign m303_105 =10'b0;

   // m303_106 = W*in
   wire signed [9:0] m303_106;
   assign m303_106 =10'b0;

   // m303_107 = W*in
   wire signed [9:0] m303_107;
   assign m303_107 ={ {4{in303[5]}} , in303[5:0] };

   // m303_108 = W*in
   wire signed [9:0] m303_108;
   assign m303_108 ={ {5{neg303[5]}} , neg303[5:1] };

   // m303_109 = W*in
   wire signed [9:0] m303_109;
   assign m303_109 =10'b0;

   // m303_110 = W*in
   wire signed [9:0] m303_110;
   assign m303_110 =10'b0;

   // m303_111 = W*in
   wire signed [9:0] m303_111;
   assign m303_111 =10'b0;

   // m303_112 = W*in
   wire signed [9:0] m303_112;
   assign m303_112 =10'b0;

   // m303_113 = W*in
   wire signed [9:0] m303_113;
   assign m303_113 =10'b0;

   // m303_114 = W*in
   wire signed [9:0] m303_114;
   assign m303_114 =10'b0;

   // m303_115 = W*in
   wire signed [9:0] m303_115;
   assign m303_115 =10'b0;

   // m303_116 = W*in
   wire signed [9:0] m303_116;
   assign m303_116 =10'b0;

   // m303_117 = W*in
   wire signed [9:0] m303_117;
   assign m303_117 =10'b0;

   // m304_1 = W*in
   wire signed [9:0] m304_1;
   assign m304_1 =10'b0;

   // m304_2 = W*in
   wire signed [9:0] m304_2;
   assign m304_2 =10'b0;

   // m304_3 = W*in
   wire signed [9:0] m304_3;
   assign m304_3 =10'b0;

   // m304_4 = W*in
   wire signed [9:0] m304_4;
   assign m304_4 =10'b0;

   // m304_5 = W*in
   wire signed [9:0] m304_5;
   assign m304_5 =10'b0;

   // m304_6 = W*in
   wire signed [9:0] m304_6;
   assign m304_6 =10'b0;

   // m304_7 = W*in
   wire signed [9:0] m304_7;
   assign m304_7 =10'b0;

   // m304_8 = W*in
   wire signed [9:0] m304_8;
   assign m304_8 =10'b0;

   // m304_9 = W*in
   wire signed [9:0] m304_9;
   assign m304_9 =10'b0;

   // m304_10 = W*in
   wire signed [9:0] m304_10;
   assign m304_10 =10'b0;

   // m304_11 = W*in
   wire signed [9:0] m304_11;
   assign m304_11 =10'b0;

   // m304_12 = W*in
   wire signed [9:0] m304_12;
   assign m304_12 =10'b0;

   // m304_13 = W*in
   wire signed [9:0] m304_13;
   assign m304_13 =10'b0;

   // m304_14 = W*in
   wire signed [9:0] m304_14;
   assign m304_14 =10'b0;

   // m304_15 = W*in
   wire signed [9:0] m304_15;
   assign m304_15 =10'b0;

   // m304_16 = W*in
   wire signed [9:0] m304_16;
   assign m304_16 =10'b0;

   // m304_17 = W*in
   wire signed [9:0] m304_17;
   assign m304_17 =10'b0;

   // m304_18 = W*in
   wire signed [9:0] m304_18;
   assign m304_18 =10'b0;

   // m304_19 = W*in
   wire signed [9:0] m304_19;
   assign m304_19 =10'b0;

   // m304_20 = W*in
   wire signed [9:0] m304_20;
   assign m304_20 ={ {5{in304[5]}} , in304[5:1] };

   // m304_21 = W*in
   wire signed [9:0] m304_21;
   assign m304_21 =10'b0;

   // m304_22 = W*in
   wire signed [9:0] m304_22;
   assign m304_22 =10'b0;

   // m304_23 = W*in
   wire signed [9:0] m304_23;
   assign m304_23 =10'b0;

   // m304_24 = W*in
   wire signed [9:0] m304_24;
   assign m304_24 =10'b0;

   // m304_25 = W*in
   wire signed [9:0] m304_25;
   assign m304_25 ={ {5{in304[5]}} , in304[5:1] };

   // m304_26 = W*in
   wire signed [9:0] m304_26;
   assign m304_26 =10'b0;

   // m304_27 = W*in
   wire signed [9:0] m304_27;
   assign m304_27 =10'b0;

   // m304_28 = W*in
   wire signed [9:0] m304_28;
   assign m304_28 =10'b0;

   // m304_29 = W*in
   wire signed [9:0] m304_29;
   assign m304_29 =10'b0;

   // m304_30 = W*in
   wire signed [9:0] m304_30;
   assign m304_30 =10'b0;

   // m304_31 = W*in
   wire signed [9:0] m304_31;
   assign m304_31 =10'b0;

   // m304_32 = W*in
   wire signed [9:0] m304_32;
   assign m304_32 =10'b0;

   // m304_33 = W*in
   wire signed [9:0] m304_33;
   assign m304_33 =10'b0;

   // m304_34 = W*in
   wire signed [9:0] m304_34;
   assign m304_34 =10'b0;

   // m304_35 = W*in
   wire signed [9:0] m304_35;
   assign m304_35 ={ {5{neg304[5]}} , neg304[5:1] };

   // m304_36 = W*in
   wire signed [9:0] m304_36;
   assign m304_36 =10'b0;

   // m304_37 = W*in
   wire signed [9:0] m304_37;
   assign m304_37 =10'b0;

   // m304_38 = W*in
   wire signed [9:0] m304_38;
   assign m304_38 =10'b0;

   // m304_39 = W*in
   wire signed [9:0] m304_39;
   assign m304_39 =10'b0;

   // m304_40 = W*in
   wire signed [9:0] m304_40;
   assign m304_40 =10'b0;

   // m304_41 = W*in
   wire signed [9:0] m304_41;
   assign m304_41 =10'b0;

   // m304_42 = W*in
   wire signed [9:0] m304_42;
   assign m304_42 =10'b0;

   // m304_43 = W*in
   wire signed [9:0] m304_43;
   assign m304_43 =10'b0;

   // m304_44 = W*in
   wire signed [9:0] m304_44;
   assign m304_44 =10'b0;

   // m304_45 = W*in
   wire signed [9:0] m304_45;
   assign m304_45 =10'b0;

   // m304_46 = W*in
   wire signed [9:0] m304_46;
   assign m304_46 =10'b0;

   // m304_47 = W*in
   wire signed [9:0] m304_47;
   assign m304_47 =10'b0;

   // m304_48 = W*in
   wire signed [9:0] m304_48;
   assign m304_48 ={ {4{in304[5]}} , in304[5:0] };

   // m304_49 = W*in
   wire signed [9:0] m304_49;
   assign m304_49 ={ {4{neg304[5]}} , neg304[5:0] };

   // m304_50 = W*in
   wire signed [9:0] m304_50;
   assign m304_50 =10'b0;

   // m304_51 = W*in
   wire signed [9:0] m304_51;
   assign m304_51 =10'b0;

   // m304_52 = W*in
   wire signed [9:0] m304_52;
   assign m304_52 =10'b0;

   // m304_53 = W*in
   wire signed [9:0] m304_53;
   assign m304_53 =10'b0;

   // m304_54 = W*in
   wire signed [9:0] m304_54;
   assign m304_54 =10'b0;

   // m304_55 = W*in
   wire signed [9:0] m304_55;
   assign m304_55 =10'b0;

   // m304_56 = W*in
   wire signed [9:0] m304_56;
   assign m304_56 =10'b0;

   // m304_57 = W*in
   wire signed [9:0] m304_57;
   assign m304_57 =10'b0;

   // m304_58 = W*in
   wire signed [9:0] m304_58;
   assign m304_58 =10'b0;

   // m304_59 = W*in
   wire signed [9:0] m304_59;
   assign m304_59 =10'b0;

   // m304_60 = W*in
   wire signed [9:0] m304_60;
   assign m304_60 =10'b0;

   // m304_61 = W*in
   wire signed [9:0] m304_61;
   assign m304_61 =10'b0;

   // m304_62 = W*in
   wire signed [9:0] m304_62;
   assign m304_62 =10'b0;

   // m304_63 = W*in
   wire signed [9:0] m304_63;
   assign m304_63 =10'b0;

   // m304_64 = W*in
   wire signed [9:0] m304_64;
   assign m304_64 =10'b0;

   // m304_65 = W*in
   wire signed [9:0] m304_65;
   assign m304_65 ={ {5{neg304[5]}} , neg304[5:1] };

   // m304_66 = W*in
   wire signed [9:0] m304_66;
   assign m304_66 ={ {5{neg304[5]}} , neg304[5:1] };

   // m304_67 = W*in
   wire signed [9:0] m304_67;
   assign m304_67 =10'b0;

   // m304_68 = W*in
   wire signed [9:0] m304_68;
   assign m304_68 =10'b0;

   // m304_69 = W*in
   wire signed [9:0] m304_69;
   assign m304_69 =10'b0;

   // m304_70 = W*in
   wire signed [9:0] m304_70;
   assign m304_70 ={ {4{in304[5]}} , in304[5:0] };

   // m304_71 = W*in
   wire signed [9:0] m304_71;
   assign m304_71 =10'b0;

   // m304_72 = W*in
   wire signed [9:0] m304_72;
   assign m304_72 =10'b0;

   // m304_73 = W*in
   wire signed [9:0] m304_73;
   assign m304_73 =10'b0;

   // m304_74 = W*in
   wire signed [9:0] m304_74;
   assign m304_74 =10'b0;

   // m304_75 = W*in
   wire signed [9:0] m304_75;
   assign m304_75 =10'b0;

   // m304_76 = W*in
   wire signed [9:0] m304_76;
   assign m304_76 =10'b0;

   // m304_77 = W*in
   wire signed [9:0] m304_77;
   assign m304_77 =10'b0;

   // m304_78 = W*in
   wire signed [9:0] m304_78;
   assign m304_78 =10'b0;

   // m304_79 = W*in
   wire signed [9:0] m304_79;
   assign m304_79 =10'b0;

   // m304_80 = W*in
   wire signed [9:0] m304_80;
   assign m304_80 =10'b0;

   // m304_81 = W*in
   wire signed [9:0] m304_81;
   assign m304_81 =10'b0;

   // m304_82 = W*in
   wire signed [9:0] m304_82;
   assign m304_82 =10'b0;

   // m304_83 = W*in
   wire signed [9:0] m304_83;
   assign m304_83 =10'b0;

   // m304_84 = W*in
   wire signed [9:0] m304_84;
   assign m304_84 =10'b0;

   // m304_85 = W*in
   wire signed [9:0] m304_85;
   assign m304_85 =10'b0;

   // m304_86 = W*in
   wire signed [9:0] m304_86;
   assign m304_86 =10'b0;

   // m304_87 = W*in
   wire signed [9:0] m304_87;
   assign m304_87 =10'b0;

   // m304_88 = W*in
   wire signed [9:0] m304_88;
   assign m304_88 =10'b0;

   // m304_89 = W*in
   wire signed [9:0] m304_89;
   assign m304_89 =10'b0;

   // m304_90 = W*in
   wire signed [9:0] m304_90;
   assign m304_90 =10'b0;

   // m304_91 = W*in
   wire signed [9:0] m304_91;
   assign m304_91 =10'b0;

   // m304_92 = W*in
   wire signed [9:0] m304_92;
   assign m304_92 =10'b0;

   // m304_93 = W*in
   wire signed [9:0] m304_93;
   assign m304_93 =10'b0;

   // m304_94 = W*in
   wire signed [9:0] m304_94;
   assign m304_94 =10'b0;

   // m304_95 = W*in
   wire signed [9:0] m304_95;
   assign m304_95 =10'b0;

   // m304_96 = W*in
   wire signed [9:0] m304_96;
   assign m304_96 =10'b0;

   // m304_97 = W*in
   wire signed [9:0] m304_97;
   assign m304_97 =10'b0;

   // m304_98 = W*in
   wire signed [9:0] m304_98;
   assign m304_98 =10'b0;

   // m304_99 = W*in
   wire signed [9:0] m304_99;
   assign m304_99 =10'b0;

   // m304_100 = W*in
   wire signed [9:0] m304_100;
   assign m304_100 =10'b0;

   // m304_101 = W*in
   wire signed [9:0] m304_101;
   assign m304_101 =10'b0;

   // m304_102 = W*in
   wire signed [9:0] m304_102;
   assign m304_102 =10'b0;

   // m304_103 = W*in
   wire signed [9:0] m304_103;
   assign m304_103 =10'b0;

   // m304_104 = W*in
   wire signed [9:0] m304_104;
   assign m304_104 =10'b0;

   // m304_105 = W*in
   wire signed [9:0] m304_105;
   assign m304_105 =10'b0;

   // m304_106 = W*in
   wire signed [9:0] m304_106;
   assign m304_106 =10'b0;

   // m304_107 = W*in
   wire signed [9:0] m304_107;
   assign m304_107 =10'b0;

   // m304_108 = W*in
   wire signed [9:0] m304_108;
   assign m304_108 =10'b0;

   // m304_109 = W*in
   wire signed [9:0] m304_109;
   assign m304_109 ={ {5{neg304[5]}} , neg304[5:1] };

   // m304_110 = W*in
   wire signed [9:0] m304_110;
   assign m304_110 =10'b0;

   // m304_111 = W*in
   wire signed [9:0] m304_111;
   assign m304_111 =10'b0;

   // m304_112 = W*in
   wire signed [9:0] m304_112;
   assign m304_112 =10'b0;

   // m304_113 = W*in
   wire signed [9:0] m304_113;
   assign m304_113 ={ {4{in304[5]}} , in304[5:0] };

   // m304_114 = W*in
   wire signed [9:0] m304_114;
   assign m304_114 =10'b0;

   // m304_115 = W*in
   wire signed [9:0] m304_115;
   assign m304_115 =10'b0;

   // m304_116 = W*in
   wire signed [9:0] m304_116;
   assign m304_116 =10'b0;

   // m304_117 = W*in
   wire signed [9:0] m304_117;
   assign m304_117 =10'b0;

   // m305_1 = W*in
   wire signed [9:0] m305_1;
   assign m305_1 =10'b0;

   // m305_2 = W*in
   wire signed [9:0] m305_2;
   assign m305_2 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_3 = W*in
   wire signed [9:0] m305_3;
   assign m305_3 =10'b0;

   // m305_4 = W*in
   wire signed [9:0] m305_4;
   assign m305_4 =10'b0;

   // m305_5 = W*in
   wire signed [9:0] m305_5;
   assign m305_5 =10'b0;

   // m305_6 = W*in
   wire signed [9:0] m305_6;
   assign m305_6 =10'b0;

   // m305_7 = W*in
   wire signed [9:0] m305_7;
   assign m305_7 =10'b0;

   // m305_8 = W*in
   wire signed [9:0] m305_8;
   assign m305_8 =10'b0;

   // m305_9 = W*in
   wire signed [9:0] m305_9;
   assign m305_9 =10'b0;

   // m305_10 = W*in
   wire signed [9:0] m305_10;
   assign m305_10 =10'b0;

   // m305_11 = W*in
   wire signed [9:0] m305_11;
   assign m305_11 =10'b0;

   // m305_12 = W*in
   wire signed [9:0] m305_12;
   assign m305_12 =10'b0;

   // m305_13 = W*in
   wire signed [9:0] m305_13;
   assign m305_13 =10'b0;

   // m305_14 = W*in
   wire signed [9:0] m305_14;
   assign m305_14 =10'b0;

   // m305_15 = W*in
   wire signed [9:0] m305_15;
   assign m305_15 =10'b0;

   // m305_16 = W*in
   wire signed [9:0] m305_16;
   assign m305_16 =10'b0;

   // m305_17 = W*in
   wire signed [9:0] m305_17;
   assign m305_17 =10'b0;

   // m305_18 = W*in
   wire signed [9:0] m305_18;
   assign m305_18 =10'b0;

   // m305_19 = W*in
   wire signed [9:0] m305_19;
   assign m305_19 =10'b0;

   // m305_20 = W*in
   wire signed [9:0] m305_20;
   assign m305_20 =10'b0;

   // m305_21 = W*in
   wire signed [9:0] m305_21;
   assign m305_21 =10'b0;

   // m305_22 = W*in
   wire signed [9:0] m305_22;
   assign m305_22 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_23 = W*in
   wire signed [9:0] m305_23;
   assign m305_23 =10'b0;

   // m305_24 = W*in
   wire signed [9:0] m305_24;
   assign m305_24 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_25 = W*in
   wire signed [9:0] m305_25;
   assign m305_25 =10'b0;

   // m305_26 = W*in
   wire signed [9:0] m305_26;
   assign m305_26 =10'b0;

   // m305_27 = W*in
   wire signed [9:0] m305_27;
   assign m305_27 =10'b0;

   // m305_28 = W*in
   wire signed [9:0] m305_28;
   assign m305_28 =10'b0;

   // m305_29 = W*in
   wire signed [9:0] m305_29;
   assign m305_29 =10'b0;

   // m305_30 = W*in
   wire signed [9:0] m305_30;
   assign m305_30 =10'b0;

   // m305_31 = W*in
   wire signed [9:0] m305_31;
   assign m305_31 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_32 = W*in
   wire signed [9:0] m305_32;
   assign m305_32 =10'b0;

   // m305_33 = W*in
   wire signed [9:0] m305_33;
   assign m305_33 =10'b0;

   // m305_34 = W*in
   wire signed [9:0] m305_34;
   assign m305_34 =10'b0;

   // m305_35 = W*in
   wire signed [9:0] m305_35;
   assign m305_35 =10'b0;

   // m305_36 = W*in
   wire signed [9:0] m305_36;
   assign m305_36 =10'b0;

   // m305_37 = W*in
   wire signed [9:0] m305_37;
   assign m305_37 =10'b0;

   // m305_38 = W*in
   wire signed [9:0] m305_38;
   assign m305_38 =10'b0;

   // m305_39 = W*in
   wire signed [9:0] m305_39;
   assign m305_39 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_40 = W*in
   wire signed [9:0] m305_40;
   assign m305_40 =10'b0;

   // m305_41 = W*in
   wire signed [9:0] m305_41;
   assign m305_41 =10'b0;

   // m305_42 = W*in
   wire signed [9:0] m305_42;
   assign m305_42 =10'b0;

   // m305_43 = W*in
   wire signed [9:0] m305_43;
   assign m305_43 =10'b0;

   // m305_44 = W*in
   wire signed [9:0] m305_44;
   assign m305_44 =10'b0;

   // m305_45 = W*in
   wire signed [9:0] m305_45;
   assign m305_45 =10'b0;

   // m305_46 = W*in
   wire signed [9:0] m305_46;
   assign m305_46 =10'b0;

   // m305_47 = W*in
   wire signed [9:0] m305_47;
   assign m305_47 =10'b0;

   // m305_48 = W*in
   wire signed [9:0] m305_48;
   assign m305_48 ={ {4{in305[5]}} , in305[5:0] };

   // m305_49 = W*in
   wire signed [9:0] m305_49;
   assign m305_49 =10'b0;

   // m305_50 = W*in
   wire signed [9:0] m305_50;
   assign m305_50 =10'b0;

   // m305_51 = W*in
   wire signed [9:0] m305_51;
   assign m305_51 =10'b0;

   // m305_52 = W*in
   wire signed [9:0] m305_52;
   assign m305_52 =10'b0;

   // m305_53 = W*in
   wire signed [9:0] m305_53;
   assign m305_53 =10'b0;

   // m305_54 = W*in
   wire signed [9:0] m305_54;
   assign m305_54 =10'b0;

   // m305_55 = W*in
   wire signed [9:0] m305_55;
   assign m305_55 =10'b0;

   // m305_56 = W*in
   wire signed [9:0] m305_56;
   assign m305_56 =10'b0;

   // m305_57 = W*in
   wire signed [9:0] m305_57;
   assign m305_57 =10'b0;

   // m305_58 = W*in
   wire signed [9:0] m305_58;
   assign m305_58 =10'b0;

   // m305_59 = W*in
   wire signed [9:0] m305_59;
   assign m305_59 =10'b0;

   // m305_60 = W*in
   wire signed [9:0] m305_60;
   assign m305_60 ={ {4{in305[5]}} , in305[5:0] };

   // m305_61 = W*in
   wire signed [9:0] m305_61;
   assign m305_61 =10'b0;

   // m305_62 = W*in
   wire signed [9:0] m305_62;
   assign m305_62 =10'b0;

   // m305_63 = W*in
   wire signed [9:0] m305_63;
   assign m305_63 =10'b0;

   // m305_64 = W*in
   wire signed [9:0] m305_64;
   assign m305_64 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_65 = W*in
   wire signed [9:0] m305_65;
   assign m305_65 =10'b0;

   // m305_66 = W*in
   wire signed [9:0] m305_66;
   assign m305_66 =10'b0;

   // m305_67 = W*in
   wire signed [9:0] m305_67;
   assign m305_67 =10'b0;

   // m305_68 = W*in
   wire signed [9:0] m305_68;
   assign m305_68 =10'b0;

   // m305_69 = W*in
   wire signed [9:0] m305_69;
   assign m305_69 ={ {4{in305[5]}} , in305[5:0] };

   // m305_70 = W*in
   wire signed [9:0] m305_70;
   assign m305_70 ={ {5{in305[5]}} , in305[5:1] };

   // m305_71 = W*in
   wire signed [9:0] m305_71;
   assign m305_71 ={ {5{in305[5]}} , in305[5:1] };

   // m305_72 = W*in
   wire signed [9:0] m305_72;
   assign m305_72 =10'b0;

   // m305_73 = W*in
   wire signed [9:0] m305_73;
   assign m305_73 ={ {5{neg305[5]}} , neg305[5:1] };

   // m305_74 = W*in
   wire signed [9:0] m305_74;
   assign m305_74 =10'b0;

   // m305_75 = W*in
   wire signed [9:0] m305_75;
   assign m305_75 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_76 = W*in
   wire signed [9:0] m305_76;
   assign m305_76 ={ {4{in305[5]}} , in305[5:0] };

   // m305_77 = W*in
   wire signed [9:0] m305_77;
   assign m305_77 =10'b0;

   // m305_78 = W*in
   wire signed [9:0] m305_78;
   assign m305_78 =10'b0;

   // m305_79 = W*in
   wire signed [9:0] m305_79;
   assign m305_79 =10'b0;

   // m305_80 = W*in
   wire signed [9:0] m305_80;
   assign m305_80 =10'b0;

   // m305_81 = W*in
   wire signed [9:0] m305_81;
   assign m305_81 ={ {5{neg305[5]}} , neg305[5:1] };

   // m305_82 = W*in
   wire signed [9:0] m305_82;
   assign m305_82 =10'b0;

   // m305_83 = W*in
   wire signed [9:0] m305_83;
   assign m305_83 =10'b0;

   // m305_84 = W*in
   wire signed [9:0] m305_84;
   assign m305_84 =10'b0;

   // m305_85 = W*in
   wire signed [9:0] m305_85;
   assign m305_85 =10'b0;

   // m305_86 = W*in
   wire signed [9:0] m305_86;
   assign m305_86 =10'b0;

   // m305_87 = W*in
   wire signed [9:0] m305_87;
   assign m305_87 ={ {4{in305[5]}} , in305[5:0] };

   // m305_88 = W*in
   wire signed [9:0] m305_88;
   assign m305_88 =10'b0;

   // m305_89 = W*in
   wire signed [9:0] m305_89;
   assign m305_89 =10'b0;

   // m305_90 = W*in
   wire signed [9:0] m305_90;
   assign m305_90 =10'b0;

   // m305_91 = W*in
   wire signed [9:0] m305_91;
   assign m305_91 =10'b0;

   // m305_92 = W*in
   wire signed [9:0] m305_92;
   assign m305_92 ={ {4{in305[5]}} , in305[5:0] };

   // m305_93 = W*in
   wire signed [9:0] m305_93;
   assign m305_93 =10'b0;

   // m305_94 = W*in
   wire signed [9:0] m305_94;
   assign m305_94 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_95 = W*in
   wire signed [9:0] m305_95;
   assign m305_95 =10'b0;

   // m305_96 = W*in
   wire signed [9:0] m305_96;
   assign m305_96 =10'b0;

   // m305_97 = W*in
   wire signed [9:0] m305_97;
   assign m305_97 =10'b0;

   // m305_98 = W*in
   wire signed [9:0] m305_98;
   assign m305_98 ={ {4{neg305[5]}} , neg305[5:0] };

   // m305_99 = W*in
   wire signed [9:0] m305_99;
   assign m305_99 =10'b0;

   // m305_100 = W*in
   wire signed [9:0] m305_100;
   assign m305_100 =10'b0;

   // m305_101 = W*in
   wire signed [9:0] m305_101;
   assign m305_101 =10'b0;

   // m305_102 = W*in
   wire signed [9:0] m305_102;
   assign m305_102 =10'b0;

   // m305_103 = W*in
   wire signed [9:0] m305_103;
   assign m305_103 =10'b0;

   // m305_104 = W*in
   wire signed [9:0] m305_104;
   assign m305_104 =10'b0;

   // m305_105 = W*in
   wire signed [9:0] m305_105;
   assign m305_105 =10'b0;

   // m305_106 = W*in
   wire signed [9:0] m305_106;
   assign m305_106 =10'b0;

   // m305_107 = W*in
   wire signed [9:0] m305_107;
   assign m305_107 =10'b0;

   // m305_108 = W*in
   wire signed [9:0] m305_108;
   assign m305_108 =10'b0;

   // m305_109 = W*in
   wire signed [9:0] m305_109;
   assign m305_109 =10'b0;

   // m305_110 = W*in
   wire signed [9:0] m305_110;
   assign m305_110 =10'b0;

   // m305_111 = W*in
   wire signed [9:0] m305_111;
   assign m305_111 =10'b0;

   // m305_112 = W*in
   wire signed [9:0] m305_112;
   assign m305_112 =10'b0;

   // m305_113 = W*in
   wire signed [9:0] m305_113;
   assign m305_113 ={ {4{in305[5]}} , in305[5:0] };

   // m305_114 = W*in
   wire signed [9:0] m305_114;
   assign m305_114 =10'b0;

   // m305_115 = W*in
   wire signed [9:0] m305_115;
   assign m305_115 =10'b0;

   // m305_116 = W*in
   wire signed [9:0] m305_116;
   assign m305_116 =10'b0;

   // m305_117 = W*in
   wire signed [9:0] m305_117;
   assign m305_117 =10'b0;

   // m306_1 = W*in
   wire signed [9:0] m306_1;
   assign m306_1 =10'b0;

   // m306_2 = W*in
   wire signed [9:0] m306_2;
   assign m306_2 =10'b0;

   // m306_3 = W*in
   wire signed [9:0] m306_3;
   assign m306_3 =10'b0;

   // m306_4 = W*in
   wire signed [9:0] m306_4;
   assign m306_4 =10'b0;

   // m306_5 = W*in
   wire signed [9:0] m306_5;
   assign m306_5 =10'b0;

   // m306_6 = W*in
   wire signed [9:0] m306_6;
   assign m306_6 =10'b0;

   // m306_7 = W*in
   wire signed [9:0] m306_7;
   assign m306_7 =10'b0;

   // m306_8 = W*in
   wire signed [9:0] m306_8;
   assign m306_8 =10'b0;

   // m306_9 = W*in
   wire signed [9:0] m306_9;
   assign m306_9 =10'b0;

   // m306_10 = W*in
   wire signed [9:0] m306_10;
   assign m306_10 =10'b0;

   // m306_11 = W*in
   wire signed [9:0] m306_11;
   assign m306_11 =10'b0;

   // m306_12 = W*in
   wire signed [9:0] m306_12;
   assign m306_12 =10'b0;

   // m306_13 = W*in
   wire signed [9:0] m306_13;
   assign m306_13 =10'b0;

   // m306_14 = W*in
   wire signed [9:0] m306_14;
   assign m306_14 =10'b0;

   // m306_15 = W*in
   wire signed [9:0] m306_15;
   assign m306_15 =10'b0;

   // m306_16 = W*in
   wire signed [9:0] m306_16;
   assign m306_16 ={ {5{in306[5]}} , in306[5:1] };

   // m306_17 = W*in
   wire signed [9:0] m306_17;
   assign m306_17 =10'b0;

   // m306_18 = W*in
   wire signed [9:0] m306_18;
   assign m306_18 =10'b0;

   // m306_19 = W*in
   wire signed [9:0] m306_19;
   assign m306_19 ={ {5{neg306[5]}} , neg306[5:1] };

   // m306_20 = W*in
   wire signed [9:0] m306_20;
   assign m306_20 =10'b0;

   // m306_21 = W*in
   wire signed [9:0] m306_21;
   assign m306_21 =10'b0;

   // m306_22 = W*in
   wire signed [9:0] m306_22;
   assign m306_22 ={ {4{neg306[5]}} , neg306[5:0] };

   // m306_23 = W*in
   wire signed [9:0] m306_23;
   assign m306_23 =10'b0;

   // m306_24 = W*in
   wire signed [9:0] m306_24;
   assign m306_24 =10'b0;

   // m306_25 = W*in
   wire signed [9:0] m306_25;
   assign m306_25 ={ {5{neg306[5]}} , neg306[5:1] };

   // m306_26 = W*in
   wire signed [9:0] m306_26;
   assign m306_26 =10'b0;

   // m306_27 = W*in
   wire signed [9:0] m306_27;
   assign m306_27 ={ {4{neg306[5]}} , neg306[5:0] };

   // m306_28 = W*in
   wire signed [9:0] m306_28;
   assign m306_28 =10'b0;

   // m306_29 = W*in
   wire signed [9:0] m306_29;
   assign m306_29 =10'b0;

   // m306_30 = W*in
   wire signed [9:0] m306_30;
   assign m306_30 =10'b0;

   // m306_31 = W*in
   wire signed [9:0] m306_31;
   assign m306_31 =10'b0;

   // m306_32 = W*in
   wire signed [9:0] m306_32;
   assign m306_32 =10'b0;

   // m306_33 = W*in
   wire signed [9:0] m306_33;
   assign m306_33 =10'b0;

   // m306_34 = W*in
   wire signed [9:0] m306_34;
   assign m306_34 =10'b0;

   // m306_35 = W*in
   wire signed [9:0] m306_35;
   assign m306_35 =10'b0;

   // m306_36 = W*in
   wire signed [9:0] m306_36;
   assign m306_36 =10'b0;

   // m306_37 = W*in
   wire signed [9:0] m306_37;
   assign m306_37 ={ {4{in306[5]}} , in306[5:0] };

   // m306_38 = W*in
   wire signed [9:0] m306_38;
   assign m306_38 =10'b0;

   // m306_39 = W*in
   wire signed [9:0] m306_39;
   assign m306_39 =10'b0;

   // m306_40 = W*in
   wire signed [9:0] m306_40;
   assign m306_40 =10'b0;

   // m306_41 = W*in
   wire signed [9:0] m306_41;
   assign m306_41 =10'b0;

   // m306_42 = W*in
   wire signed [9:0] m306_42;
   assign m306_42 =10'b0;

   // m306_43 = W*in
   wire signed [9:0] m306_43;
   assign m306_43 =10'b0;

   // m306_44 = W*in
   wire signed [9:0] m306_44;
   assign m306_44 =10'b0;

   // m306_45 = W*in
   wire signed [9:0] m306_45;
   assign m306_45 =10'b0;

   // m306_46 = W*in
   wire signed [9:0] m306_46;
   assign m306_46 =10'b0;

   // m306_47 = W*in
   wire signed [9:0] m306_47;
   assign m306_47 =10'b0;

   // m306_48 = W*in
   wire signed [9:0] m306_48;
   assign m306_48 =10'b0;

   // m306_49 = W*in
   wire signed [9:0] m306_49;
   assign m306_49 =10'b0;

   // m306_50 = W*in
   wire signed [9:0] m306_50;
   assign m306_50 =10'b0;

   // m306_51 = W*in
   wire signed [9:0] m306_51;
   assign m306_51 ={ {4{in306[5]}} , in306[5:0] };

   // m306_52 = W*in
   wire signed [9:0] m306_52;
   assign m306_52 =10'b0;

   // m306_53 = W*in
   wire signed [9:0] m306_53;
   assign m306_53 =10'b0;

   // m306_54 = W*in
   wire signed [9:0] m306_54;
   assign m306_54 =10'b0;

   // m306_55 = W*in
   wire signed [9:0] m306_55;
   assign m306_55 =10'b0;

   // m306_56 = W*in
   wire signed [9:0] m306_56;
   assign m306_56 ={ {4{in306[5]}} , in306[5:0] };

   // m306_57 = W*in
   wire signed [9:0] m306_57;
   assign m306_57 =10'b0;

   // m306_58 = W*in
   wire signed [9:0] m306_58;
   assign m306_58 =10'b0;

   // m306_59 = W*in
   wire signed [9:0] m306_59;
   assign m306_59 ={ {4{neg306[5]}} , neg306[5:0] };

   // m306_60 = W*in
   wire signed [9:0] m306_60;
   assign m306_60 =10'b0;

   // m306_61 = W*in
   wire signed [9:0] m306_61;
   assign m306_61 ={ {4{in306[5]}} , in306[5:0] };

   // m306_62 = W*in
   wire signed [9:0] m306_62;
   assign m306_62 =10'b0;

   // m306_63 = W*in
   wire signed [9:0] m306_63;
   assign m306_63 =10'b0;

   // m306_64 = W*in
   wire signed [9:0] m306_64;
   assign m306_64 =10'b0;

   // m306_65 = W*in
   wire signed [9:0] m306_65;
   assign m306_65 =10'b0;

   // m306_66 = W*in
   wire signed [9:0] m306_66;
   assign m306_66 =10'b0;

   // m306_67 = W*in
   wire signed [9:0] m306_67;
   assign m306_67 =10'b0;

   // m306_68 = W*in
   wire signed [9:0] m306_68;
   assign m306_68 =10'b0;

   // m306_69 = W*in
   wire signed [9:0] m306_69;
   assign m306_69 =10'b0;

   // m306_70 = W*in
   wire signed [9:0] m306_70;
   assign m306_70 =10'b0;

   // m306_71 = W*in
   wire signed [9:0] m306_71;
   assign m306_71 =10'b0;

   // m306_72 = W*in
   wire signed [9:0] m306_72;
   assign m306_72 =10'b0;

   // m306_73 = W*in
   wire signed [9:0] m306_73;
   assign m306_73 =10'b0;

   // m306_74 = W*in
   wire signed [9:0] m306_74;
   assign m306_74 =10'b0;

   // m306_75 = W*in
   wire signed [9:0] m306_75;
   assign m306_75 =10'b0;

   // m306_76 = W*in
   wire signed [9:0] m306_76;
   assign m306_76 =10'b0;

   // m306_77 = W*in
   wire signed [9:0] m306_77;
   assign m306_77 =10'b0;

   // m306_78 = W*in
   wire signed [9:0] m306_78;
   assign m306_78 =10'b0;

   // m306_79 = W*in
   wire signed [9:0] m306_79;
   assign m306_79 =10'b0;

   // m306_80 = W*in
   wire signed [9:0] m306_80;
   assign m306_80 =10'b0;

   // m306_81 = W*in
   wire signed [9:0] m306_81;
   assign m306_81 ={ {5{neg306[5]}} , neg306[5:1] };

   // m306_82 = W*in
   wire signed [9:0] m306_82;
   assign m306_82 =10'b0;

   // m306_83 = W*in
   wire signed [9:0] m306_83;
   assign m306_83 ={ {5{in306[5]}} , in306[5:1] };

   // m306_84 = W*in
   wire signed [9:0] m306_84;
   assign m306_84 =10'b0;

   // m306_85 = W*in
   wire signed [9:0] m306_85;
   assign m306_85 =10'b0;

   // m306_86 = W*in
   wire signed [9:0] m306_86;
   assign m306_86 =10'b0;

   // m306_87 = W*in
   wire signed [9:0] m306_87;
   assign m306_87 =10'b0;

   // m306_88 = W*in
   wire signed [9:0] m306_88;
   assign m306_88 =10'b0;

   // m306_89 = W*in
   wire signed [9:0] m306_89;
   assign m306_89 =10'b0;

   // m306_90 = W*in
   wire signed [9:0] m306_90;
   assign m306_90 =10'b0;

   // m306_91 = W*in
   wire signed [9:0] m306_91;
   assign m306_91 =10'b0;

   // m306_92 = W*in
   wire signed [9:0] m306_92;
   assign m306_92 =10'b0;

   // m306_93 = W*in
   wire signed [9:0] m306_93;
   assign m306_93 =10'b0;

   // m306_94 = W*in
   wire signed [9:0] m306_94;
   assign m306_94 =10'b0;

   // m306_95 = W*in
   wire signed [9:0] m306_95;
   assign m306_95 =10'b0;

   // m306_96 = W*in
   wire signed [9:0] m306_96;
   assign m306_96 =10'b0;

   // m306_97 = W*in
   wire signed [9:0] m306_97;
   assign m306_97 =10'b0;

   // m306_98 = W*in
   wire signed [9:0] m306_98;
   assign m306_98 =10'b0;

   // m306_99 = W*in
   wire signed [9:0] m306_99;
   assign m306_99 =10'b0;

   // m306_100 = W*in
   wire signed [9:0] m306_100;
   assign m306_100 =10'b0;

   // m306_101 = W*in
   wire signed [9:0] m306_101;
   assign m306_101 =10'b0;

   // m306_102 = W*in
   wire signed [9:0] m306_102;
   assign m306_102 =10'b0;

   // m306_103 = W*in
   wire signed [9:0] m306_103;
   assign m306_103 =10'b0;

   // m306_104 = W*in
   wire signed [9:0] m306_104;
   assign m306_104 =10'b0;

   // m306_105 = W*in
   wire signed [9:0] m306_105;
   assign m306_105 =10'b0;

   // m306_106 = W*in
   wire signed [9:0] m306_106;
   assign m306_106 =10'b0;

   // m306_107 = W*in
   wire signed [9:0] m306_107;
   assign m306_107 =10'b0;

   // m306_108 = W*in
   wire signed [9:0] m306_108;
   assign m306_108 =10'b0;

   // m306_109 = W*in
   wire signed [9:0] m306_109;
   assign m306_109 =10'b0;

   // m306_110 = W*in
   wire signed [9:0] m306_110;
   assign m306_110 =10'b0;

   // m306_111 = W*in
   wire signed [9:0] m306_111;
   assign m306_111 =10'b0;

   // m306_112 = W*in
   wire signed [9:0] m306_112;
   assign m306_112 =10'b0;

   // m306_113 = W*in
   wire signed [9:0] m306_113;
   assign m306_113 =10'b0;

   // m306_114 = W*in
   wire signed [9:0] m306_114;
   assign m306_114 ={ {5{neg306[5]}} , neg306[5:1] };

   // m306_115 = W*in
   wire signed [9:0] m306_115;
   assign m306_115 ={ {5{neg306[5]}} , neg306[5:1] };

   // m306_116 = W*in
   wire signed [9:0] m306_116;
   assign m306_116 =10'b0;

   // m306_117 = W*in
   wire signed [9:0] m306_117;
   assign m306_117 =10'b0;

   // m307_1 = W*in
   wire signed [9:0] m307_1;
   assign m307_1 =10'b0;

   // m307_2 = W*in
   wire signed [9:0] m307_2;
   assign m307_2 =10'b0;

   // m307_3 = W*in
   wire signed [9:0] m307_3;
   assign m307_3 =10'b0;

   // m307_4 = W*in
   wire signed [9:0] m307_4;
   assign m307_4 =10'b0;

   // m307_5 = W*in
   wire signed [9:0] m307_5;
   assign m307_5 =10'b0;

   // m307_6 = W*in
   wire signed [9:0] m307_6;
   assign m307_6 =10'b0;

   // m307_7 = W*in
   wire signed [9:0] m307_7;
   assign m307_7 =10'b0;

   // m307_8 = W*in
   wire signed [9:0] m307_8;
   assign m307_8 =10'b0;

   // m307_9 = W*in
   wire signed [9:0] m307_9;
   assign m307_9 =10'b0;

   // m307_10 = W*in
   wire signed [9:0] m307_10;
   assign m307_10 =10'b0;

   // m307_11 = W*in
   wire signed [9:0] m307_11;
   assign m307_11 =10'b0;

   // m307_12 = W*in
   wire signed [9:0] m307_12;
   assign m307_12 =10'b0;

   // m307_13 = W*in
   wire signed [9:0] m307_13;
   assign m307_13 =10'b0;

   // m307_14 = W*in
   wire signed [9:0] m307_14;
   assign m307_14 =10'b0;

   // m307_15 = W*in
   wire signed [9:0] m307_15;
   assign m307_15 =10'b0;

   // m307_16 = W*in
   wire signed [9:0] m307_16;
   assign m307_16 =10'b0;

   // m307_17 = W*in
   wire signed [9:0] m307_17;
   assign m307_17 =10'b0;

   // m307_18 = W*in
   wire signed [9:0] m307_18;
   assign m307_18 =10'b0;

   // m307_19 = W*in
   wire signed [9:0] m307_19;
   assign m307_19 ={ {5{neg307[5]}} , neg307[5:1] };

   // m307_20 = W*in
   wire signed [9:0] m307_20;
   assign m307_20 =10'b0;

   // m307_21 = W*in
   wire signed [9:0] m307_21;
   assign m307_21 =10'b0;

   // m307_22 = W*in
   wire signed [9:0] m307_22;
   assign m307_22 =10'b0;

   // m307_23 = W*in
   wire signed [9:0] m307_23;
   assign m307_23 =10'b0;

   // m307_24 = W*in
   wire signed [9:0] m307_24;
   assign m307_24 =10'b0;

   // m307_25 = W*in
   wire signed [9:0] m307_25;
   assign m307_25 ={ {5{neg307[5]}} , neg307[5:1] };

   // m307_26 = W*in
   wire signed [9:0] m307_26;
   assign m307_26 =10'b0;

   // m307_27 = W*in
   wire signed [9:0] m307_27;
   assign m307_27 ={ {5{in307[5]}} , in307[5:1] };

   // m307_28 = W*in
   wire signed [9:0] m307_28;
   assign m307_28 =10'b0;

   // m307_29 = W*in
   wire signed [9:0] m307_29;
   assign m307_29 =10'b0;

   // m307_30 = W*in
   wire signed [9:0] m307_30;
   assign m307_30 =10'b0;

   // m307_31 = W*in
   wire signed [9:0] m307_31;
   assign m307_31 =10'b0;

   // m307_32 = W*in
   wire signed [9:0] m307_32;
   assign m307_32 =10'b0;

   // m307_33 = W*in
   wire signed [9:0] m307_33;
   assign m307_33 =10'b0;

   // m307_34 = W*in
   wire signed [9:0] m307_34;
   assign m307_34 =10'b0;

   // m307_35 = W*in
   wire signed [9:0] m307_35;
   assign m307_35 ={ {4{in307[5]}} , in307[5:0] };

   // m307_36 = W*in
   wire signed [9:0] m307_36;
   assign m307_36 =10'b0;

   // m307_37 = W*in
   wire signed [9:0] m307_37;
   assign m307_37 =10'b0;

   // m307_38 = W*in
   wire signed [9:0] m307_38;
   assign m307_38 =10'b0;

   // m307_39 = W*in
   wire signed [9:0] m307_39;
   assign m307_39 =10'b0;

   // m307_40 = W*in
   wire signed [9:0] m307_40;
   assign m307_40 =10'b0;

   // m307_41 = W*in
   wire signed [9:0] m307_41;
   assign m307_41 =10'b0;

   // m307_42 = W*in
   wire signed [9:0] m307_42;
   assign m307_42 =10'b0;

   // m307_43 = W*in
   wire signed [9:0] m307_43;
   assign m307_43 =10'b0;

   // m307_44 = W*in
   wire signed [9:0] m307_44;
   assign m307_44 =10'b0;

   // m307_45 = W*in
   wire signed [9:0] m307_45;
   assign m307_45 =10'b0;

   // m307_46 = W*in
   wire signed [9:0] m307_46;
   assign m307_46 =10'b0;

   // m307_47 = W*in
   wire signed [9:0] m307_47;
   assign m307_47 =10'b0;

   // m307_48 = W*in
   wire signed [9:0] m307_48;
   assign m307_48 =10'b0;

   // m307_49 = W*in
   wire signed [9:0] m307_49;
   assign m307_49 =10'b0;

   // m307_50 = W*in
   wire signed [9:0] m307_50;
   assign m307_50 =10'b0;

   // m307_51 = W*in
   wire signed [9:0] m307_51;
   assign m307_51 =10'b0;

   // m307_52 = W*in
   wire signed [9:0] m307_52;
   assign m307_52 =10'b0;

   // m307_53 = W*in
   wire signed [9:0] m307_53;
   assign m307_53 =10'b0;

   // m307_54 = W*in
   wire signed [9:0] m307_54;
   assign m307_54 =10'b0;

   // m307_55 = W*in
   wire signed [9:0] m307_55;
   assign m307_55 =10'b0;

   // m307_56 = W*in
   wire signed [9:0] m307_56;
   assign m307_56 =10'b0;

   // m307_57 = W*in
   wire signed [9:0] m307_57;
   assign m307_57 =10'b0;

   // m307_58 = W*in
   wire signed [9:0] m307_58;
   assign m307_58 =10'b0;

   // m307_59 = W*in
   wire signed [9:0] m307_59;
   assign m307_59 =10'b0;

   // m307_60 = W*in
   wire signed [9:0] m307_60;
   assign m307_60 =10'b0;

   // m307_61 = W*in
   wire signed [9:0] m307_61;
   assign m307_61 =10'b0;

   // m307_62 = W*in
   wire signed [9:0] m307_62;
   assign m307_62 =10'b0;

   // m307_63 = W*in
   wire signed [9:0] m307_63;
   assign m307_63 =10'b0;

   // m307_64 = W*in
   wire signed [9:0] m307_64;
   assign m307_64 ={ {5{in307[5]}} , in307[5:1] };

   // m307_65 = W*in
   wire signed [9:0] m307_65;
   assign m307_65 ={ {5{neg307[5]}} , neg307[5:1] };

   // m307_66 = W*in
   wire signed [9:0] m307_66;
   assign m307_66 =10'b0;

   // m307_67 = W*in
   wire signed [9:0] m307_67;
   assign m307_67 ={ {4{neg307[5]}} , neg307[5:0] };

   // m307_68 = W*in
   wire signed [9:0] m307_68;
   assign m307_68 =10'b0;

   // m307_69 = W*in
   wire signed [9:0] m307_69;
   assign m307_69 ={ {5{neg307[5]}} , neg307[5:1] };

   // m307_70 = W*in
   wire signed [9:0] m307_70;
   assign m307_70 ={ {5{neg307[5]}} , neg307[5:1] };

   // m307_71 = W*in
   wire signed [9:0] m307_71;
   assign m307_71 =10'b0;

   // m307_72 = W*in
   wire signed [9:0] m307_72;
   assign m307_72 =10'b0;

   // m307_73 = W*in
   wire signed [9:0] m307_73;
   assign m307_73 =10'b0;

   // m307_74 = W*in
   wire signed [9:0] m307_74;
   assign m307_74 =10'b0;

   // m307_75 = W*in
   wire signed [9:0] m307_75;
   assign m307_75 =10'b0;

   // m307_76 = W*in
   wire signed [9:0] m307_76;
   assign m307_76 =10'b0;

   // m307_77 = W*in
   wire signed [9:0] m307_77;
   assign m307_77 =10'b0;

   // m307_78 = W*in
   wire signed [9:0] m307_78;
   assign m307_78 =10'b0;

   // m307_79 = W*in
   wire signed [9:0] m307_79;
   assign m307_79 =10'b0;

   // m307_80 = W*in
   wire signed [9:0] m307_80;
   assign m307_80 =10'b0;

   // m307_81 = W*in
   wire signed [9:0] m307_81;
   assign m307_81 =10'b0;

   // m307_82 = W*in
   wire signed [9:0] m307_82;
   assign m307_82 =10'b0;

   // m307_83 = W*in
   wire signed [9:0] m307_83;
   assign m307_83 ={ {5{in307[5]}} , in307[5:1] };

   // m307_84 = W*in
   wire signed [9:0] m307_84;
   assign m307_84 =10'b0;

   // m307_85 = W*in
   wire signed [9:0] m307_85;
   assign m307_85 =10'b0;

   // m307_86 = W*in
   wire signed [9:0] m307_86;
   assign m307_86 =10'b0;

   // m307_87 = W*in
   wire signed [9:0] m307_87;
   assign m307_87 =10'b0;

   // m307_88 = W*in
   wire signed [9:0] m307_88;
   assign m307_88 =10'b0;

   // m307_89 = W*in
   wire signed [9:0] m307_89;
   assign m307_89 =10'b0;

   // m307_90 = W*in
   wire signed [9:0] m307_90;
   assign m307_90 =10'b0;

   // m307_91 = W*in
   wire signed [9:0] m307_91;
   assign m307_91 =10'b0;

   // m307_92 = W*in
   wire signed [9:0] m307_92;
   assign m307_92 =10'b0;

   // m307_93 = W*in
   wire signed [9:0] m307_93;
   assign m307_93 =10'b0;

   // m307_94 = W*in
   wire signed [9:0] m307_94;
   assign m307_94 =10'b0;

   // m307_95 = W*in
   wire signed [9:0] m307_95;
   assign m307_95 =10'b0;

   // m307_96 = W*in
   wire signed [9:0] m307_96;
   assign m307_96 =10'b0;

   // m307_97 = W*in
   wire signed [9:0] m307_97;
   assign m307_97 =10'b0;

   // m307_98 = W*in
   wire signed [9:0] m307_98;
   assign m307_98 =10'b0;

   // m307_99 = W*in
   wire signed [9:0] m307_99;
   assign m307_99 =10'b0;

   // m307_100 = W*in
   wire signed [9:0] m307_100;
   assign m307_100 =10'b0;

   // m307_101 = W*in
   wire signed [9:0] m307_101;
   assign m307_101 =10'b0;

   // m307_102 = W*in
   wire signed [9:0] m307_102;
   assign m307_102 =10'b0;

   // m307_103 = W*in
   wire signed [9:0] m307_103;
   assign m307_103 =10'b0;

   // m307_104 = W*in
   wire signed [9:0] m307_104;
   assign m307_104 =10'b0;

   // m307_105 = W*in
   wire signed [9:0] m307_105;
   assign m307_105 =10'b0;

   // m307_106 = W*in
   wire signed [9:0] m307_106;
   assign m307_106 =10'b0;

   // m307_107 = W*in
   wire signed [9:0] m307_107;
   assign m307_107 =10'b0;

   // m307_108 = W*in
   wire signed [9:0] m307_108;
   assign m307_108 =10'b0;

   // m307_109 = W*in
   wire signed [9:0] m307_109;
   assign m307_109 =10'b0;

   // m307_110 = W*in
   wire signed [9:0] m307_110;
   assign m307_110 =10'b0;

   // m307_111 = W*in
   wire signed [9:0] m307_111;
   assign m307_111 =10'b0;

   // m307_112 = W*in
   wire signed [9:0] m307_112;
   assign m307_112 =10'b0;

   // m307_113 = W*in
   wire signed [9:0] m307_113;
   assign m307_113 =10'b0;

   // m307_114 = W*in
   wire signed [9:0] m307_114;
   assign m307_114 =10'b0;

   // m307_115 = W*in
   wire signed [9:0] m307_115;
   assign m307_115 ={ {5{in307[5]}} , in307[5:1] };

   // m307_116 = W*in
   wire signed [9:0] m307_116;
   assign m307_116 =10'b0;

   // m307_117 = W*in
   wire signed [9:0] m307_117;
   assign m307_117 ={ {4{in307[5]}} , in307[5:0] };

   // m308_1 = W*in
   wire signed [9:0] m308_1;
   assign m308_1 =10'b0;

   // m308_2 = W*in
   wire signed [9:0] m308_2;
   assign m308_2 =10'b0;

   // m308_3 = W*in
   wire signed [9:0] m308_3;
   assign m308_3 =10'b0;

   // m308_4 = W*in
   wire signed [9:0] m308_4;
   assign m308_4 =10'b0;

   // m308_5 = W*in
   wire signed [9:0] m308_5;
   assign m308_5 =10'b0;

   // m308_6 = W*in
   wire signed [9:0] m308_6;
   assign m308_6 =10'b0;

   // m308_7 = W*in
   wire signed [9:0] m308_7;
   assign m308_7 =10'b0;

   // m308_8 = W*in
   wire signed [9:0] m308_8;
   assign m308_8 =10'b0;

   // m308_9 = W*in
   wire signed [9:0] m308_9;
   assign m308_9 =10'b0;

   // m308_10 = W*in
   wire signed [9:0] m308_10;
   assign m308_10 =10'b0;

   // m308_11 = W*in
   wire signed [9:0] m308_11;
   assign m308_11 =10'b0;

   // m308_12 = W*in
   wire signed [9:0] m308_12;
   assign m308_12 =10'b0;

   // m308_13 = W*in
   wire signed [9:0] m308_13;
   assign m308_13 =10'b0;

   // m308_14 = W*in
   wire signed [9:0] m308_14;
   assign m308_14 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_15 = W*in
   wire signed [9:0] m308_15;
   assign m308_15 =10'b0;

   // m308_16 = W*in
   wire signed [9:0] m308_16;
   assign m308_16 =10'b0;

   // m308_17 = W*in
   wire signed [9:0] m308_17;
   assign m308_17 ={ {5{in308[5]}} , in308[5:1] };

   // m308_18 = W*in
   wire signed [9:0] m308_18;
   assign m308_18 ={ {5{neg308[5]}} , neg308[5:1] };

   // m308_19 = W*in
   wire signed [9:0] m308_19;
   assign m308_19 =10'b0;

   // m308_20 = W*in
   wire signed [9:0] m308_20;
   assign m308_20 ={ {5{in308[5]}} , in308[5:1] };

   // m308_21 = W*in
   wire signed [9:0] m308_21;
   assign m308_21 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_22 = W*in
   wire signed [9:0] m308_22;
   assign m308_22 =10'b0;

   // m308_23 = W*in
   wire signed [9:0] m308_23;
   assign m308_23 =10'b0;

   // m308_24 = W*in
   wire signed [9:0] m308_24;
   assign m308_24 =10'b0;

   // m308_25 = W*in
   wire signed [9:0] m308_25;
   assign m308_25 ={ {5{in308[5]}} , in308[5:1] };

   // m308_26 = W*in
   wire signed [9:0] m308_26;
   assign m308_26 ={ {5{neg308[5]}} , neg308[5:1] };

   // m308_27 = W*in
   wire signed [9:0] m308_27;
   assign m308_27 ={ {4{in308[5]}} , in308[5:0] };

   // m308_28 = W*in
   wire signed [9:0] m308_28;
   assign m308_28 ={ {4{in308[5]}} , in308[5:0] };

   // m308_29 = W*in
   wire signed [9:0] m308_29;
   assign m308_29 =10'b0;

   // m308_30 = W*in
   wire signed [9:0] m308_30;
   assign m308_30 =10'b0;

   // m308_31 = W*in
   wire signed [9:0] m308_31;
   assign m308_31 =10'b0;

   // m308_32 = W*in
   wire signed [9:0] m308_32;
   assign m308_32 =10'b0;

   // m308_33 = W*in
   wire signed [9:0] m308_33;
   assign m308_33 =10'b0;

   // m308_34 = W*in
   wire signed [9:0] m308_34;
   assign m308_34 =10'b0;

   // m308_35 = W*in
   wire signed [9:0] m308_35;
   assign m308_35 ={ {5{in308[5]}} , in308[5:1] };

   // m308_36 = W*in
   wire signed [9:0] m308_36;
   assign m308_36 =10'b0;

   // m308_37 = W*in
   wire signed [9:0] m308_37;
   assign m308_37 =10'b0;

   // m308_38 = W*in
   wire signed [9:0] m308_38;
   assign m308_38 =10'b0;

   // m308_39 = W*in
   wire signed [9:0] m308_39;
   assign m308_39 =10'b0;

   // m308_40 = W*in
   wire signed [9:0] m308_40;
   assign m308_40 =10'b0;

   // m308_41 = W*in
   wire signed [9:0] m308_41;
   assign m308_41 =10'b0;

   // m308_42 = W*in
   wire signed [9:0] m308_42;
   assign m308_42 =10'b0;

   // m308_43 = W*in
   wire signed [9:0] m308_43;
   assign m308_43 =10'b0;

   // m308_44 = W*in
   wire signed [9:0] m308_44;
   assign m308_44 =10'b0;

   // m308_45 = W*in
   wire signed [9:0] m308_45;
   assign m308_45 =10'b0;

   // m308_46 = W*in
   wire signed [9:0] m308_46;
   assign m308_46 =10'b0;

   // m308_47 = W*in
   wire signed [9:0] m308_47;
   assign m308_47 =10'b0;

   // m308_48 = W*in
   wire signed [9:0] m308_48;
   assign m308_48 =10'b0;

   // m308_49 = W*in
   wire signed [9:0] m308_49;
   assign m308_49 =10'b0;

   // m308_50 = W*in
   wire signed [9:0] m308_50;
   assign m308_50 =10'b0;

   // m308_51 = W*in
   wire signed [9:0] m308_51;
   assign m308_51 =10'b0;

   // m308_52 = W*in
   wire signed [9:0] m308_52;
   assign m308_52 =10'b0;

   // m308_53 = W*in
   wire signed [9:0] m308_53;
   assign m308_53 =10'b0;

   // m308_54 = W*in
   wire signed [9:0] m308_54;
   assign m308_54 =10'b0;

   // m308_55 = W*in
   wire signed [9:0] m308_55;
   assign m308_55 =10'b0;

   // m308_56 = W*in
   wire signed [9:0] m308_56;
   assign m308_56 =10'b0;

   // m308_57 = W*in
   wire signed [9:0] m308_57;
   assign m308_57 =10'b0;

   // m308_58 = W*in
   wire signed [9:0] m308_58;
   assign m308_58 =10'b0;

   // m308_59 = W*in
   wire signed [9:0] m308_59;
   assign m308_59 ={ {4{in308[5]}} , in308[5:0] };

   // m308_60 = W*in
   wire signed [9:0] m308_60;
   assign m308_60 ={ {4{in308[5]}} , in308[5:0] };

   // m308_61 = W*in
   wire signed [9:0] m308_61;
   assign m308_61 ={ {4{in308[5]}} , in308[5:0] };

   // m308_62 = W*in
   wire signed [9:0] m308_62;
   assign m308_62 =10'b0;

   // m308_63 = W*in
   wire signed [9:0] m308_63;
   assign m308_63 =10'b0;

   // m308_64 = W*in
   wire signed [9:0] m308_64;
   assign m308_64 ={ {5{neg308[5]}} , neg308[5:1] };

   // m308_65 = W*in
   wire signed [9:0] m308_65;
   assign m308_65 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_66 = W*in
   wire signed [9:0] m308_66;
   assign m308_66 =10'b0;

   // m308_67 = W*in
   wire signed [9:0] m308_67;
   assign m308_67 =10'b0;

   // m308_68 = W*in
   wire signed [9:0] m308_68;
   assign m308_68 =10'b0;

   // m308_69 = W*in
   wire signed [9:0] m308_69;
   assign m308_69 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_70 = W*in
   wire signed [9:0] m308_70;
   assign m308_70 ={ {5{neg308[5]}} , neg308[5:1] };

   // m308_71 = W*in
   wire signed [9:0] m308_71;
   assign m308_71 ={ {5{in308[5]}} , in308[5:1] };

   // m308_72 = W*in
   wire signed [9:0] m308_72;
   assign m308_72 =10'b0;

   // m308_73 = W*in
   wire signed [9:0] m308_73;
   assign m308_73 =10'b0;

   // m308_74 = W*in
   wire signed [9:0] m308_74;
   assign m308_74 =10'b0;

   // m308_75 = W*in
   wire signed [9:0] m308_75;
   assign m308_75 =10'b0;

   // m308_76 = W*in
   wire signed [9:0] m308_76;
   assign m308_76 =10'b0;

   // m308_77 = W*in
   wire signed [9:0] m308_77;
   assign m308_77 =10'b0;

   // m308_78 = W*in
   wire signed [9:0] m308_78;
   assign m308_78 =10'b0;

   // m308_79 = W*in
   wire signed [9:0] m308_79;
   assign m308_79 =10'b0;

   // m308_80 = W*in
   wire signed [9:0] m308_80;
   assign m308_80 =10'b0;

   // m308_81 = W*in
   wire signed [9:0] m308_81;
   assign m308_81 ={ {5{neg308[5]}} , neg308[5:1] };

   // m308_82 = W*in
   wire signed [9:0] m308_82;
   assign m308_82 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_83 = W*in
   wire signed [9:0] m308_83;
   assign m308_83 ={ {5{in308[5]}} , in308[5:1] };

   // m308_84 = W*in
   wire signed [9:0] m308_84;
   assign m308_84 =10'b0;

   // m308_85 = W*in
   wire signed [9:0] m308_85;
   assign m308_85 =10'b0;

   // m308_86 = W*in
   wire signed [9:0] m308_86;
   assign m308_86 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_87 = W*in
   wire signed [9:0] m308_87;
   assign m308_87 =10'b0;

   // m308_88 = W*in
   wire signed [9:0] m308_88;
   assign m308_88 =10'b0;

   // m308_89 = W*in
   wire signed [9:0] m308_89;
   assign m308_89 =10'b0;

   // m308_90 = W*in
   wire signed [9:0] m308_90;
   assign m308_90 =10'b0;

   // m308_91 = W*in
   wire signed [9:0] m308_91;
   assign m308_91 =10'b0;

   // m308_92 = W*in
   wire signed [9:0] m308_92;
   assign m308_92 =10'b0;

   // m308_93 = W*in
   wire signed [9:0] m308_93;
   assign m308_93 ={ {4{neg308[5]}} , neg308[5:0] };

   // m308_94 = W*in
   wire signed [9:0] m308_94;
   assign m308_94 =10'b0;

   // m308_95 = W*in
   wire signed [9:0] m308_95;
   assign m308_95 =10'b0;

   // m308_96 = W*in
   wire signed [9:0] m308_96;
   assign m308_96 =10'b0;

   // m308_97 = W*in
   wire signed [9:0] m308_97;
   assign m308_97 =10'b0;

   // m308_98 = W*in
   wire signed [9:0] m308_98;
   assign m308_98 =10'b0;

   // m308_99 = W*in
   wire signed [9:0] m308_99;
   assign m308_99 =10'b0;

   // m308_100 = W*in
   wire signed [9:0] m308_100;
   assign m308_100 =10'b0;

   // m308_101 = W*in
   wire signed [9:0] m308_101;
   assign m308_101 =10'b0;

   // m308_102 = W*in
   wire signed [9:0] m308_102;
   assign m308_102 =10'b0;

   // m308_103 = W*in
   wire signed [9:0] m308_103;
   assign m308_103 =10'b0;

   // m308_104 = W*in
   wire signed [9:0] m308_104;
   assign m308_104 =10'b0;

   // m308_105 = W*in
   wire signed [9:0] m308_105;
   assign m308_105 =10'b0;

   // m308_106 = W*in
   wire signed [9:0] m308_106;
   assign m308_106 =10'b0;

   // m308_107 = W*in
   wire signed [9:0] m308_107;
   assign m308_107 ={ {4{in308[5]}} , in308[5:0] };

   // m308_108 = W*in
   wire signed [9:0] m308_108;
   assign m308_108 =10'b0;

   // m308_109 = W*in
   wire signed [9:0] m308_109;
   assign m308_109 =10'b0;

   // m308_110 = W*in
   wire signed [9:0] m308_110;
   assign m308_110 =10'b0;

   // m308_111 = W*in
   wire signed [9:0] m308_111;
   assign m308_111 =10'b0;

   // m308_112 = W*in
   wire signed [9:0] m308_112;
   assign m308_112 =10'b0;

   // m308_113 = W*in
   wire signed [9:0] m308_113;
   assign m308_113 =10'b0;

   // m308_114 = W*in
   wire signed [9:0] m308_114;
   assign m308_114 =10'b0;

   // m308_115 = W*in
   wire signed [9:0] m308_115;
   assign m308_115 ={ {5{in308[5]}} , in308[5:1] };

   // m308_116 = W*in
   wire signed [9:0] m308_116;
   assign m308_116 =10'b0;

   // m308_117 = W*in
   wire signed [9:0] m308_117;
   assign m308_117 ={ {4{in308[5]}} , in308[5:0] };

   // m309_1 = W*in
   wire signed [9:0] m309_1;
   assign m309_1 =10'b0;

   // m309_2 = W*in
   wire signed [9:0] m309_2;
   assign m309_2 =10'b0;

   // m309_3 = W*in
   wire signed [9:0] m309_3;
   assign m309_3 =10'b0;

   // m309_4 = W*in
   wire signed [9:0] m309_4;
   assign m309_4 =10'b0;

   // m309_5 = W*in
   wire signed [9:0] m309_5;
   assign m309_5 =10'b0;

   // m309_6 = W*in
   wire signed [9:0] m309_6;
   assign m309_6 =10'b0;

   // m309_7 = W*in
   wire signed [9:0] m309_7;
   assign m309_7 =10'b0;

   // m309_8 = W*in
   wire signed [9:0] m309_8;
   assign m309_8 =10'b0;

   // m309_9 = W*in
   wire signed [9:0] m309_9;
   assign m309_9 =10'b0;

   // m309_10 = W*in
   wire signed [9:0] m309_10;
   assign m309_10 =10'b0;

   // m309_11 = W*in
   wire signed [9:0] m309_11;
   assign m309_11 =10'b0;

   // m309_12 = W*in
   wire signed [9:0] m309_12;
   assign m309_12 =10'b0;

   // m309_13 = W*in
   wire signed [9:0] m309_13;
   assign m309_13 =10'b0;

   // m309_14 = W*in
   wire signed [9:0] m309_14;
   assign m309_14 =10'b0;

   // m309_15 = W*in
   wire signed [9:0] m309_15;
   assign m309_15 =10'b0;

   // m309_16 = W*in
   wire signed [9:0] m309_16;
   assign m309_16 =10'b0;

   // m309_17 = W*in
   wire signed [9:0] m309_17;
   assign m309_17 =10'b0;

   // m309_18 = W*in
   wire signed [9:0] m309_18;
   assign m309_18 =10'b0;

   // m309_19 = W*in
   wire signed [9:0] m309_19;
   assign m309_19 ={ {5{neg309[5]}} , neg309[5:1] };

   // m309_20 = W*in
   wire signed [9:0] m309_20;
   assign m309_20 =10'b0;

   // m309_21 = W*in
   wire signed [9:0] m309_21;
   assign m309_21 =10'b0;

   // m309_22 = W*in
   wire signed [9:0] m309_22;
   assign m309_22 =10'b0;

   // m309_23 = W*in
   wire signed [9:0] m309_23;
   assign m309_23 =10'b0;

   // m309_24 = W*in
   wire signed [9:0] m309_24;
   assign m309_24 =10'b0;

   // m309_25 = W*in
   wire signed [9:0] m309_25;
   assign m309_25 =10'b0;

   // m309_26 = W*in
   wire signed [9:0] m309_26;
   assign m309_26 =10'b0;

   // m309_27 = W*in
   wire signed [9:0] m309_27;
   assign m309_27 =10'b0;

   // m309_28 = W*in
   wire signed [9:0] m309_28;
   assign m309_28 =10'b0;

   // m309_29 = W*in
   wire signed [9:0] m309_29;
   assign m309_29 =10'b0;

   // m309_30 = W*in
   wire signed [9:0] m309_30;
   assign m309_30 ={ {5{neg309[5]}} , neg309[5:1] };

   // m309_31 = W*in
   wire signed [9:0] m309_31;
   assign m309_31 =10'b0;

   // m309_32 = W*in
   wire signed [9:0] m309_32;
   assign m309_32 =10'b0;

   // m309_33 = W*in
   wire signed [9:0] m309_33;
   assign m309_33 =10'b0;

   // m309_34 = W*in
   wire signed [9:0] m309_34;
   assign m309_34 ={ {5{in309[5]}} , in309[5:1] };

   // m309_35 = W*in
   wire signed [9:0] m309_35;
   assign m309_35 =10'b0;

   // m309_36 = W*in
   wire signed [9:0] m309_36;
   assign m309_36 =10'b0;

   // m309_37 = W*in
   wire signed [9:0] m309_37;
   assign m309_37 =10'b0;

   // m309_38 = W*in
   wire signed [9:0] m309_38;
   assign m309_38 =10'b0;

   // m309_39 = W*in
   wire signed [9:0] m309_39;
   assign m309_39 =10'b0;

   // m309_40 = W*in
   wire signed [9:0] m309_40;
   assign m309_40 =10'b0;

   // m309_41 = W*in
   wire signed [9:0] m309_41;
   assign m309_41 =10'b0;

   // m309_42 = W*in
   wire signed [9:0] m309_42;
   assign m309_42 =10'b0;

   // m309_43 = W*in
   wire signed [9:0] m309_43;
   assign m309_43 =10'b0;

   // m309_44 = W*in
   wire signed [9:0] m309_44;
   assign m309_44 =10'b0;

   // m309_45 = W*in
   wire signed [9:0] m309_45;
   assign m309_45 =10'b0;

   // m309_46 = W*in
   wire signed [9:0] m309_46;
   assign m309_46 =10'b0;

   // m309_47 = W*in
   wire signed [9:0] m309_47;
   assign m309_47 =10'b0;

   // m309_48 = W*in
   wire signed [9:0] m309_48;
   assign m309_48 =10'b0;

   // m309_49 = W*in
   wire signed [9:0] m309_49;
   assign m309_49 =10'b0;

   // m309_50 = W*in
   wire signed [9:0] m309_50;
   assign m309_50 =10'b0;

   // m309_51 = W*in
   wire signed [9:0] m309_51;
   assign m309_51 =10'b0;

   // m309_52 = W*in
   wire signed [9:0] m309_52;
   assign m309_52 =10'b0;

   // m309_53 = W*in
   wire signed [9:0] m309_53;
   assign m309_53 =10'b0;

   // m309_54 = W*in
   wire signed [9:0] m309_54;
   assign m309_54 =10'b0;

   // m309_55 = W*in
   wire signed [9:0] m309_55;
   assign m309_55 =10'b0;

   // m309_56 = W*in
   wire signed [9:0] m309_56;
   assign m309_56 =10'b0;

   // m309_57 = W*in
   wire signed [9:0] m309_57;
   assign m309_57 =10'b0;

   // m309_58 = W*in
   wire signed [9:0] m309_58;
   assign m309_58 =10'b0;

   // m309_59 = W*in
   wire signed [9:0] m309_59;
   assign m309_59 =10'b0;

   // m309_60 = W*in
   wire signed [9:0] m309_60;
   assign m309_60 =10'b0;

   // m309_61 = W*in
   wire signed [9:0] m309_61;
   assign m309_61 =10'b0;

   // m309_62 = W*in
   wire signed [9:0] m309_62;
   assign m309_62 =10'b0;

   // m309_63 = W*in
   wire signed [9:0] m309_63;
   assign m309_63 =10'b0;

   // m309_64 = W*in
   wire signed [9:0] m309_64;
   assign m309_64 ={ {5{in309[5]}} , in309[5:1] };

   // m309_65 = W*in
   wire signed [9:0] m309_65;
   assign m309_65 =10'b0;

   // m309_66 = W*in
   wire signed [9:0] m309_66;
   assign m309_66 =10'b0;

   // m309_67 = W*in
   wire signed [9:0] m309_67;
   assign m309_67 =10'b0;

   // m309_68 = W*in
   wire signed [9:0] m309_68;
   assign m309_68 =10'b0;

   // m309_69 = W*in
   wire signed [9:0] m309_69;
   assign m309_69 =10'b0;

   // m309_70 = W*in
   wire signed [9:0] m309_70;
   assign m309_70 =10'b0;

   // m309_71 = W*in
   wire signed [9:0] m309_71;
   assign m309_71 =10'b0;

   // m309_72 = W*in
   wire signed [9:0] m309_72;
   assign m309_72 =10'b0;

   // m309_73 = W*in
   wire signed [9:0] m309_73;
   assign m309_73 =10'b0;

   // m309_74 = W*in
   wire signed [9:0] m309_74;
   assign m309_74 =10'b0;

   // m309_75 = W*in
   wire signed [9:0] m309_75;
   assign m309_75 =10'b0;

   // m309_76 = W*in
   wire signed [9:0] m309_76;
   assign m309_76 =10'b0;

   // m309_77 = W*in
   wire signed [9:0] m309_77;
   assign m309_77 =10'b0;

   // m309_78 = W*in
   wire signed [9:0] m309_78;
   assign m309_78 =10'b0;

   // m309_79 = W*in
   wire signed [9:0] m309_79;
   assign m309_79 =10'b0;

   // m309_80 = W*in
   wire signed [9:0] m309_80;
   assign m309_80 =10'b0;

   // m309_81 = W*in
   wire signed [9:0] m309_81;
   assign m309_81 =10'b0;

   // m309_82 = W*in
   wire signed [9:0] m309_82;
   assign m309_82 =10'b0;

   // m309_83 = W*in
   wire signed [9:0] m309_83;
   assign m309_83 =10'b0;

   // m309_84 = W*in
   wire signed [9:0] m309_84;
   assign m309_84 =10'b0;

   // m309_85 = W*in
   wire signed [9:0] m309_85;
   assign m309_85 ={ {5{neg309[5]}} , neg309[5:1] };

   // m309_86 = W*in
   wire signed [9:0] m309_86;
   assign m309_86 =10'b0;

   // m309_87 = W*in
   wire signed [9:0] m309_87;
   assign m309_87 =10'b0;

   // m309_88 = W*in
   wire signed [9:0] m309_88;
   assign m309_88 =10'b0;

   // m309_89 = W*in
   wire signed [9:0] m309_89;
   assign m309_89 =10'b0;

   // m309_90 = W*in
   wire signed [9:0] m309_90;
   assign m309_90 =10'b0;

   // m309_91 = W*in
   wire signed [9:0] m309_91;
   assign m309_91 =10'b0;

   // m309_92 = W*in
   wire signed [9:0] m309_92;
   assign m309_92 =10'b0;

   // m309_93 = W*in
   wire signed [9:0] m309_93;
   assign m309_93 =10'b0;

   // m309_94 = W*in
   wire signed [9:0] m309_94;
   assign m309_94 =10'b0;

   // m309_95 = W*in
   wire signed [9:0] m309_95;
   assign m309_95 =10'b0;

   // m309_96 = W*in
   wire signed [9:0] m309_96;
   assign m309_96 =10'b0;

   // m309_97 = W*in
   wire signed [9:0] m309_97;
   assign m309_97 =10'b0;

   // m309_98 = W*in
   wire signed [9:0] m309_98;
   assign m309_98 =10'b0;

   // m309_99 = W*in
   wire signed [9:0] m309_99;
   assign m309_99 ={ {4{in309[5]}} , in309[5:0] };

   // m309_100 = W*in
   wire signed [9:0] m309_100;
   assign m309_100 =10'b0;

   // m309_101 = W*in
   wire signed [9:0] m309_101;
   assign m309_101 =10'b0;

   // m309_102 = W*in
   wire signed [9:0] m309_102;
   assign m309_102 =10'b0;

   // m309_103 = W*in
   wire signed [9:0] m309_103;
   assign m309_103 =10'b0;

   // m309_104 = W*in
   wire signed [9:0] m309_104;
   assign m309_104 =10'b0;

   // m309_105 = W*in
   wire signed [9:0] m309_105;
   assign m309_105 =10'b0;

   // m309_106 = W*in
   wire signed [9:0] m309_106;
   assign m309_106 =10'b0;

   // m309_107 = W*in
   wire signed [9:0] m309_107;
   assign m309_107 =10'b0;

   // m309_108 = W*in
   wire signed [9:0] m309_108;
   assign m309_108 =10'b0;

   // m309_109 = W*in
   wire signed [9:0] m309_109;
   assign m309_109 =10'b0;

   // m309_110 = W*in
   wire signed [9:0] m309_110;
   assign m309_110 =10'b0;

   // m309_111 = W*in
   wire signed [9:0] m309_111;
   assign m309_111 =10'b0;

   // m309_112 = W*in
   wire signed [9:0] m309_112;
   assign m309_112 =10'b0;

   // m309_113 = W*in
   wire signed [9:0] m309_113;
   assign m309_113 =10'b0;

   // m309_114 = W*in
   wire signed [9:0] m309_114;
   assign m309_114 =10'b0;

   // m309_115 = W*in
   wire signed [9:0] m309_115;
   assign m309_115 =10'b0;

   // m309_116 = W*in
   wire signed [9:0] m309_116;
   assign m309_116 =10'b0;

   // m309_117 = W*in
   wire signed [9:0] m309_117;
   assign m309_117 =10'b0;

   // m310_1 = W*in
   wire signed [9:0] m310_1;
   assign m310_1 =10'b0;

   // m310_2 = W*in
   wire signed [9:0] m310_2;
   assign m310_2 =10'b0;

   // m310_3 = W*in
   wire signed [9:0] m310_3;
   assign m310_3 =10'b0;

   // m310_4 = W*in
   wire signed [9:0] m310_4;
   assign m310_4 =10'b0;

   // m310_5 = W*in
   wire signed [9:0] m310_5;
   assign m310_5 =10'b0;

   // m310_6 = W*in
   wire signed [9:0] m310_6;
   assign m310_6 =10'b0;

   // m310_7 = W*in
   wire signed [9:0] m310_7;
   assign m310_7 =10'b0;

   // m310_8 = W*in
   wire signed [9:0] m310_8;
   assign m310_8 =10'b0;

   // m310_9 = W*in
   wire signed [9:0] m310_9;
   assign m310_9 =10'b0;

   // m310_10 = W*in
   wire signed [9:0] m310_10;
   assign m310_10 =10'b0;

   // m310_11 = W*in
   wire signed [9:0] m310_11;
   assign m310_11 =10'b0;

   // m310_12 = W*in
   wire signed [9:0] m310_12;
   assign m310_12 =10'b0;

   // m310_13 = W*in
   wire signed [9:0] m310_13;
   assign m310_13 =10'b0;

   // m310_14 = W*in
   wire signed [9:0] m310_14;
   assign m310_14 =10'b0;

   // m310_15 = W*in
   wire signed [9:0] m310_15;
   assign m310_15 =10'b0;

   // m310_16 = W*in
   wire signed [9:0] m310_16;
   assign m310_16 ={ {5{neg310[5]}} , neg310[5:1] };

   // m310_17 = W*in
   wire signed [9:0] m310_17;
   assign m310_17 =10'b0;

   // m310_18 = W*in
   wire signed [9:0] m310_18;
   assign m310_18 =10'b0;

   // m310_19 = W*in
   wire signed [9:0] m310_19;
   assign m310_19 =10'b0;

   // m310_20 = W*in
   wire signed [9:0] m310_20;
   assign m310_20 ={ {5{in310[5]}} , in310[5:1] };

   // m310_21 = W*in
   wire signed [9:0] m310_21;
   assign m310_21 ={ {5{in310[5]}} , in310[5:1] };

   // m310_22 = W*in
   wire signed [9:0] m310_22;
   assign m310_22 =10'b0;

   // m310_23 = W*in
   wire signed [9:0] m310_23;
   assign m310_23 =10'b0;

   // m310_24 = W*in
   wire signed [9:0] m310_24;
   assign m310_24 =10'b0;

   // m310_25 = W*in
   wire signed [9:0] m310_25;
   assign m310_25 ={ {5{neg310[5]}} , neg310[5:1] };

   // m310_26 = W*in
   wire signed [9:0] m310_26;
   assign m310_26 =10'b0;

   // m310_27 = W*in
   wire signed [9:0] m310_27;
   assign m310_27 ={ {5{neg310[5]}} , neg310[5:1] };

   // m310_28 = W*in
   wire signed [9:0] m310_28;
   assign m310_28 =10'b0;

   // m310_29 = W*in
   wire signed [9:0] m310_29;
   assign m310_29 =10'b0;

   // m310_30 = W*in
   wire signed [9:0] m310_30;
   assign m310_30 =10'b0;

   // m310_31 = W*in
   wire signed [9:0] m310_31;
   assign m310_31 =10'b0;

   // m310_32 = W*in
   wire signed [9:0] m310_32;
   assign m310_32 =10'b0;

   // m310_33 = W*in
   wire signed [9:0] m310_33;
   assign m310_33 =10'b0;

   // m310_34 = W*in
   wire signed [9:0] m310_34;
   assign m310_34 ={ {5{in310[5]}} , in310[5:1] };

   // m310_35 = W*in
   wire signed [9:0] m310_35;
   assign m310_35 =10'b0;

   // m310_36 = W*in
   wire signed [9:0] m310_36;
   assign m310_36 =10'b0;

   // m310_37 = W*in
   wire signed [9:0] m310_37;
   assign m310_37 =10'b0;

   // m310_38 = W*in
   wire signed [9:0] m310_38;
   assign m310_38 =10'b0;

   // m310_39 = W*in
   wire signed [9:0] m310_39;
   assign m310_39 =10'b0;

   // m310_40 = W*in
   wire signed [9:0] m310_40;
   assign m310_40 =10'b0;

   // m310_41 = W*in
   wire signed [9:0] m310_41;
   assign m310_41 ={ {4{in310[5]}} , in310[5:0] };

   // m310_42 = W*in
   wire signed [9:0] m310_42;
   assign m310_42 =10'b0;

   // m310_43 = W*in
   wire signed [9:0] m310_43;
   assign m310_43 =10'b0;

   // m310_44 = W*in
   wire signed [9:0] m310_44;
   assign m310_44 =10'b0;

   // m310_45 = W*in
   wire signed [9:0] m310_45;
   assign m310_45 ={ {4{neg310[5]}} , neg310[5:0] };

   // m310_46 = W*in
   wire signed [9:0] m310_46;
   assign m310_46 =10'b0;

   // m310_47 = W*in
   wire signed [9:0] m310_47;
   assign m310_47 =10'b0;

   // m310_48 = W*in
   wire signed [9:0] m310_48;
   assign m310_48 =10'b0;

   // m310_49 = W*in
   wire signed [9:0] m310_49;
   assign m310_49 =10'b0;

   // m310_50 = W*in
   wire signed [9:0] m310_50;
   assign m310_50 =10'b0;

   // m310_51 = W*in
   wire signed [9:0] m310_51;
   assign m310_51 =10'b0;

   // m310_52 = W*in
   wire signed [9:0] m310_52;
   assign m310_52 =10'b0;

   // m310_53 = W*in
   wire signed [9:0] m310_53;
   assign m310_53 =10'b0;

   // m310_54 = W*in
   wire signed [9:0] m310_54;
   assign m310_54 =10'b0;

   // m310_55 = W*in
   wire signed [9:0] m310_55;
   assign m310_55 =10'b0;

   // m310_56 = W*in
   wire signed [9:0] m310_56;
   assign m310_56 =10'b0;

   // m310_57 = W*in
   wire signed [9:0] m310_57;
   assign m310_57 =10'b0;

   // m310_58 = W*in
   wire signed [9:0] m310_58;
   assign m310_58 =10'b0;

   // m310_59 = W*in
   wire signed [9:0] m310_59;
   assign m310_59 =10'b0;

   // m310_60 = W*in
   wire signed [9:0] m310_60;
   assign m310_60 =10'b0;

   // m310_61 = W*in
   wire signed [9:0] m310_61;
   assign m310_61 =10'b0;

   // m310_62 = W*in
   wire signed [9:0] m310_62;
   assign m310_62 =10'b0;

   // m310_63 = W*in
   wire signed [9:0] m310_63;
   assign m310_63 =10'b0;

   // m310_64 = W*in
   wire signed [9:0] m310_64;
   assign m310_64 =10'b0;

   // m310_65 = W*in
   wire signed [9:0] m310_65;
   assign m310_65 ={ {5{in310[5]}} , in310[5:1] };

   // m310_66 = W*in
   wire signed [9:0] m310_66;
   assign m310_66 ={ {5{in310[5]}} , in310[5:1] };

   // m310_67 = W*in
   wire signed [9:0] m310_67;
   assign m310_67 =10'b0;

   // m310_68 = W*in
   wire signed [9:0] m310_68;
   assign m310_68 =10'b0;

   // m310_69 = W*in
   wire signed [9:0] m310_69;
   assign m310_69 ={ {5{in310[5]}} , in310[5:1] };

   // m310_70 = W*in
   wire signed [9:0] m310_70;
   assign m310_70 ={ {5{in310[5]}} , in310[5:1] };

   // m310_71 = W*in
   wire signed [9:0] m310_71;
   assign m310_71 =10'b0;

   // m310_72 = W*in
   wire signed [9:0] m310_72;
   assign m310_72 ={ {5{in310[5]}} , in310[5:1] };

   // m310_73 = W*in
   wire signed [9:0] m310_73;
   assign m310_73 =10'b0;

   // m310_74 = W*in
   wire signed [9:0] m310_74;
   assign m310_74 ={ {5{in310[5]}} , in310[5:1] };

   // m310_75 = W*in
   wire signed [9:0] m310_75;
   assign m310_75 =10'b0;

   // m310_76 = W*in
   wire signed [9:0] m310_76;
   assign m310_76 =10'b0;

   // m310_77 = W*in
   wire signed [9:0] m310_77;
   assign m310_77 =10'b0;

   // m310_78 = W*in
   wire signed [9:0] m310_78;
   assign m310_78 =10'b0;

   // m310_79 = W*in
   wire signed [9:0] m310_79;
   assign m310_79 =10'b0;

   // m310_80 = W*in
   wire signed [9:0] m310_80;
   assign m310_80 ={ {5{neg310[5]}} , neg310[5:1] };

   // m310_81 = W*in
   wire signed [9:0] m310_81;
   assign m310_81 =10'b0;

   // m310_82 = W*in
   wire signed [9:0] m310_82;
   assign m310_82 =10'b0;

   // m310_83 = W*in
   wire signed [9:0] m310_83;
   assign m310_83 =10'b0;

   // m310_84 = W*in
   wire signed [9:0] m310_84;
   assign m310_84 =10'b0;

   // m310_85 = W*in
   wire signed [9:0] m310_85;
   assign m310_85 =10'b0;

   // m310_86 = W*in
   wire signed [9:0] m310_86;
   assign m310_86 =10'b0;

   // m310_87 = W*in
   wire signed [9:0] m310_87;
   assign m310_87 =10'b0;

   // m310_88 = W*in
   wire signed [9:0] m310_88;
   assign m310_88 =10'b0;

   // m310_89 = W*in
   wire signed [9:0] m310_89;
   assign m310_89 =10'b0;

   // m310_90 = W*in
   wire signed [9:0] m310_90;
   assign m310_90 =10'b0;

   // m310_91 = W*in
   wire signed [9:0] m310_91;
   assign m310_91 =10'b0;

   // m310_92 = W*in
   wire signed [9:0] m310_92;
   assign m310_92 =10'b0;

   // m310_93 = W*in
   wire signed [9:0] m310_93;
   assign m310_93 =10'b0;

   // m310_94 = W*in
   wire signed [9:0] m310_94;
   assign m310_94 =10'b0;

   // m310_95 = W*in
   wire signed [9:0] m310_95;
   assign m310_95 =10'b0;

   // m310_96 = W*in
   wire signed [9:0] m310_96;
   assign m310_96 =10'b0;

   // m310_97 = W*in
   wire signed [9:0] m310_97;
   assign m310_97 =10'b0;

   // m310_98 = W*in
   wire signed [9:0] m310_98;
   assign m310_98 =10'b0;

   // m310_99 = W*in
   wire signed [9:0] m310_99;
   assign m310_99 =10'b0;

   // m310_100 = W*in
   wire signed [9:0] m310_100;
   assign m310_100 =10'b0;

   // m310_101 = W*in
   wire signed [9:0] m310_101;
   assign m310_101 =10'b0;

   // m310_102 = W*in
   wire signed [9:0] m310_102;
   assign m310_102 =10'b0;

   // m310_103 = W*in
   wire signed [9:0] m310_103;
   assign m310_103 =10'b0;

   // m310_104 = W*in
   wire signed [9:0] m310_104;
   assign m310_104 =10'b0;

   // m310_105 = W*in
   wire signed [9:0] m310_105;
   assign m310_105 =10'b0;

   // m310_106 = W*in
   wire signed [9:0] m310_106;
   assign m310_106 =10'b0;

   // m310_107 = W*in
   wire signed [9:0] m310_107;
   assign m310_107 =10'b0;

   // m310_108 = W*in
   wire signed [9:0] m310_108;
   assign m310_108 ={ {4{in310[5]}} , in310[5:0] };

   // m310_109 = W*in
   wire signed [9:0] m310_109;
   assign m310_109 ={ {4{in310[5]}} , in310[5:0] };

   // m310_110 = W*in
   wire signed [9:0] m310_110;
   assign m310_110 =10'b0;

   // m310_111 = W*in
   wire signed [9:0] m310_111;
   assign m310_111 =10'b0;

   // m310_112 = W*in
   wire signed [9:0] m310_112;
   assign m310_112 =10'b0;

   // m310_113 = W*in
   wire signed [9:0] m310_113;
   assign m310_113 =10'b0;

   // m310_114 = W*in
   wire signed [9:0] m310_114;
   assign m310_114 ={ {5{in310[5]}} , in310[5:1] };

   // m310_115 = W*in
   wire signed [9:0] m310_115;
   assign m310_115 =10'b0;

   // m310_116 = W*in
   wire signed [9:0] m310_116;
   assign m310_116 =10'b0;

   // m310_117 = W*in
   wire signed [9:0] m310_117;
   assign m310_117 =10'b0;

   // m311_1 = W*in
   wire signed [9:0] m311_1;
   assign m311_1 =10'b0;

   // m311_2 = W*in
   wire signed [9:0] m311_2;
   assign m311_2 =10'b0;

   // m311_3 = W*in
   wire signed [9:0] m311_3;
   assign m311_3 =10'b0;

   // m311_4 = W*in
   wire signed [9:0] m311_4;
   assign m311_4 =10'b0;

   // m311_5 = W*in
   wire signed [9:0] m311_5;
   assign m311_5 =10'b0;

   // m311_6 = W*in
   wire signed [9:0] m311_6;
   assign m311_6 =10'b0;

   // m311_7 = W*in
   wire signed [9:0] m311_7;
   assign m311_7 =10'b0;

   // m311_8 = W*in
   wire signed [9:0] m311_8;
   assign m311_8 =10'b0;

   // m311_9 = W*in
   wire signed [9:0] m311_9;
   assign m311_9 =10'b0;

   // m311_10 = W*in
   wire signed [9:0] m311_10;
   assign m311_10 =10'b0;

   // m311_11 = W*in
   wire signed [9:0] m311_11;
   assign m311_11 =10'b0;

   // m311_12 = W*in
   wire signed [9:0] m311_12;
   assign m311_12 =10'b0;

   // m311_13 = W*in
   wire signed [9:0] m311_13;
   assign m311_13 =10'b0;

   // m311_14 = W*in
   wire signed [9:0] m311_14;
   assign m311_14 =10'b0;

   // m311_15 = W*in
   wire signed [9:0] m311_15;
   assign m311_15 =10'b0;

   // m311_16 = W*in
   wire signed [9:0] m311_16;
   assign m311_16 ={ {5{in311[5]}} , in311[5:1] };

   // m311_17 = W*in
   wire signed [9:0] m311_17;
   assign m311_17 ={ {4{in311[5]}} , in311[5:0] };

   // m311_18 = W*in
   wire signed [9:0] m311_18;
   assign m311_18 ={ {5{neg311[5]}} , neg311[5:1] };

   // m311_19 = W*in
   wire signed [9:0] m311_19;
   assign m311_19 ={ {5{neg311[5]}} , neg311[5:1] };

   // m311_20 = W*in
   wire signed [9:0] m311_20;
   assign m311_20 ={ {5{in311[5]}} , in311[5:1] };

   // m311_21 = W*in
   wire signed [9:0] m311_21;
   assign m311_21 =10'b0;

   // m311_22 = W*in
   wire signed [9:0] m311_22;
   assign m311_22 =10'b0;

   // m311_23 = W*in
   wire signed [9:0] m311_23;
   assign m311_23 =10'b0;

   // m311_24 = W*in
   wire signed [9:0] m311_24;
   assign m311_24 =10'b0;

   // m311_25 = W*in
   wire signed [9:0] m311_25;
   assign m311_25 =10'b0;

   // m311_26 = W*in
   wire signed [9:0] m311_26;
   assign m311_26 ={ {5{neg311[5]}} , neg311[5:1] };

   // m311_27 = W*in
   wire signed [9:0] m311_27;
   assign m311_27 =10'b0;

   // m311_28 = W*in
   wire signed [9:0] m311_28;
   assign m311_28 =10'b0;

   // m311_29 = W*in
   wire signed [9:0] m311_29;
   assign m311_29 =10'b0;

   // m311_30 = W*in
   wire signed [9:0] m311_30;
   assign m311_30 ={ {5{in311[5]}} , in311[5:1] };

   // m311_31 = W*in
   wire signed [9:0] m311_31;
   assign m311_31 =10'b0;

   // m311_32 = W*in
   wire signed [9:0] m311_32;
   assign m311_32 =10'b0;

   // m311_33 = W*in
   wire signed [9:0] m311_33;
   assign m311_33 =10'b0;

   // m311_34 = W*in
   wire signed [9:0] m311_34;
   assign m311_34 =10'b0;

   // m311_35 = W*in
   wire signed [9:0] m311_35;
   assign m311_35 ={ {5{in311[5]}} , in311[5:1] };

   // m311_36 = W*in
   wire signed [9:0] m311_36;
   assign m311_36 =10'b0;

   // m311_37 = W*in
   wire signed [9:0] m311_37;
   assign m311_37 =10'b0;

   // m311_38 = W*in
   wire signed [9:0] m311_38;
   assign m311_38 =10'b0;

   // m311_39 = W*in
   wire signed [9:0] m311_39;
   assign m311_39 =10'b0;

   // m311_40 = W*in
   wire signed [9:0] m311_40;
   assign m311_40 =10'b0;

   // m311_41 = W*in
   wire signed [9:0] m311_41;
   assign m311_41 ={ {4{in311[5]}} , in311[5:0] };

   // m311_42 = W*in
   wire signed [9:0] m311_42;
   assign m311_42 =10'b0;

   // m311_43 = W*in
   wire signed [9:0] m311_43;
   assign m311_43 =10'b0;

   // m311_44 = W*in
   wire signed [9:0] m311_44;
   assign m311_44 =10'b0;

   // m311_45 = W*in
   wire signed [9:0] m311_45;
   assign m311_45 =10'b0;

   // m311_46 = W*in
   wire signed [9:0] m311_46;
   assign m311_46 =10'b0;

   // m311_47 = W*in
   wire signed [9:0] m311_47;
   assign m311_47 =10'b0;

   // m311_48 = W*in
   wire signed [9:0] m311_48;
   assign m311_48 =10'b0;

   // m311_49 = W*in
   wire signed [9:0] m311_49;
   assign m311_49 =10'b0;

   // m311_50 = W*in
   wire signed [9:0] m311_50;
   assign m311_50 =10'b0;

   // m311_51 = W*in
   wire signed [9:0] m311_51;
   assign m311_51 =10'b0;

   // m311_52 = W*in
   wire signed [9:0] m311_52;
   assign m311_52 =10'b0;

   // m311_53 = W*in
   wire signed [9:0] m311_53;
   assign m311_53 =10'b0;

   // m311_54 = W*in
   wire signed [9:0] m311_54;
   assign m311_54 =10'b0;

   // m311_55 = W*in
   wire signed [9:0] m311_55;
   assign m311_55 =10'b0;

   // m311_56 = W*in
   wire signed [9:0] m311_56;
   assign m311_56 =10'b0;

   // m311_57 = W*in
   wire signed [9:0] m311_57;
   assign m311_57 =10'b0;

   // m311_58 = W*in
   wire signed [9:0] m311_58;
   assign m311_58 =10'b0;

   // m311_59 = W*in
   wire signed [9:0] m311_59;
   assign m311_59 =10'b0;

   // m311_60 = W*in
   wire signed [9:0] m311_60;
   assign m311_60 =10'b0;

   // m311_61 = W*in
   wire signed [9:0] m311_61;
   assign m311_61 =10'b0;

   // m311_62 = W*in
   wire signed [9:0] m311_62;
   assign m311_62 =10'b0;

   // m311_63 = W*in
   wire signed [9:0] m311_63;
   assign m311_63 =10'b0;

   // m311_64 = W*in
   wire signed [9:0] m311_64;
   assign m311_64 =10'b0;

   // m311_65 = W*in
   wire signed [9:0] m311_65;
   assign m311_65 =10'b0;

   // m311_66 = W*in
   wire signed [9:0] m311_66;
   assign m311_66 =10'b0;

   // m311_67 = W*in
   wire signed [9:0] m311_67;
   assign m311_67 =10'b0;

   // m311_68 = W*in
   wire signed [9:0] m311_68;
   assign m311_68 =10'b0;

   // m311_69 = W*in
   wire signed [9:0] m311_69;
   assign m311_69 =10'b0;

   // m311_70 = W*in
   wire signed [9:0] m311_70;
   assign m311_70 ={ {5{neg311[5]}} , neg311[5:1] };

   // m311_71 = W*in
   wire signed [9:0] m311_71;
   assign m311_71 =10'b0;

   // m311_72 = W*in
   wire signed [9:0] m311_72;
   assign m311_72 ={ {5{neg311[5]}} , neg311[5:1] };

   // m311_73 = W*in
   wire signed [9:0] m311_73;
   assign m311_73 =10'b0;

   // m311_74 = W*in
   wire signed [9:0] m311_74;
   assign m311_74 =10'b0;

   // m311_75 = W*in
   wire signed [9:0] m311_75;
   assign m311_75 =10'b0;

   // m311_76 = W*in
   wire signed [9:0] m311_76;
   assign m311_76 =10'b0;

   // m311_77 = W*in
   wire signed [9:0] m311_77;
   assign m311_77 =10'b0;

   // m311_78 = W*in
   wire signed [9:0] m311_78;
   assign m311_78 =10'b0;

   // m311_79 = W*in
   wire signed [9:0] m311_79;
   assign m311_79 =10'b0;

   // m311_80 = W*in
   wire signed [9:0] m311_80;
   assign m311_80 ={ {5{in311[5]}} , in311[5:1] };

   // m311_81 = W*in
   wire signed [9:0] m311_81;
   assign m311_81 =10'b0;

   // m311_82 = W*in
   wire signed [9:0] m311_82;
   assign m311_82 =10'b0;

   // m311_83 = W*in
   wire signed [9:0] m311_83;
   assign m311_83 ={ {5{in311[5]}} , in311[5:1] };

   // m311_84 = W*in
   wire signed [9:0] m311_84;
   assign m311_84 =10'b0;

   // m311_85 = W*in
   wire signed [9:0] m311_85;
   assign m311_85 =10'b0;

   // m311_86 = W*in
   wire signed [9:0] m311_86;
   assign m311_86 =10'b0;

   // m311_87 = W*in
   wire signed [9:0] m311_87;
   assign m311_87 =10'b0;

   // m311_88 = W*in
   wire signed [9:0] m311_88;
   assign m311_88 =10'b0;

   // m311_89 = W*in
   wire signed [9:0] m311_89;
   assign m311_89 =10'b0;

   // m311_90 = W*in
   wire signed [9:0] m311_90;
   assign m311_90 =10'b0;

   // m311_91 = W*in
   wire signed [9:0] m311_91;
   assign m311_91 =10'b0;

   // m311_92 = W*in
   wire signed [9:0] m311_92;
   assign m311_92 =10'b0;

   // m311_93 = W*in
   wire signed [9:0] m311_93;
   assign m311_93 =10'b0;

   // m311_94 = W*in
   wire signed [9:0] m311_94;
   assign m311_94 =10'b0;

   // m311_95 = W*in
   wire signed [9:0] m311_95;
   assign m311_95 =10'b0;

   // m311_96 = W*in
   wire signed [9:0] m311_96;
   assign m311_96 =10'b0;

   // m311_97 = W*in
   wire signed [9:0] m311_97;
   assign m311_97 =10'b0;

   // m311_98 = W*in
   wire signed [9:0] m311_98;
   assign m311_98 =10'b0;

   // m311_99 = W*in
   wire signed [9:0] m311_99;
   assign m311_99 =10'b0;

   // m311_100 = W*in
   wire signed [9:0] m311_100;
   assign m311_100 =10'b0;

   // m311_101 = W*in
   wire signed [9:0] m311_101;
   assign m311_101 =10'b0;

   // m311_102 = W*in
   wire signed [9:0] m311_102;
   assign m311_102 =10'b0;

   // m311_103 = W*in
   wire signed [9:0] m311_103;
   assign m311_103 =10'b0;

   // m311_104 = W*in
   wire signed [9:0] m311_104;
   assign m311_104 =10'b0;

   // m311_105 = W*in
   wire signed [9:0] m311_105;
   assign m311_105 =10'b0;

   // m311_106 = W*in
   wire signed [9:0] m311_106;
   assign m311_106 =10'b0;

   // m311_107 = W*in
   wire signed [9:0] m311_107;
   assign m311_107 =10'b0;

   // m311_108 = W*in
   wire signed [9:0] m311_108;
   assign m311_108 ={ {4{in311[5]}} , in311[5:0] };

   // m311_109 = W*in
   wire signed [9:0] m311_109;
   assign m311_109 ={ {4{in311[5]}} , in311[5:0] };

   // m311_110 = W*in
   wire signed [9:0] m311_110;
   assign m311_110 =10'b0;

   // m311_111 = W*in
   wire signed [9:0] m311_111;
   assign m311_111 =10'b0;

   // m311_112 = W*in
   wire signed [9:0] m311_112;
   assign m311_112 =10'b0;

   // m311_113 = W*in
   wire signed [9:0] m311_113;
   assign m311_113 =10'b0;

   // m311_114 = W*in
   wire signed [9:0] m311_114;
   assign m311_114 =10'b0;

   // m311_115 = W*in
   wire signed [9:0] m311_115;
   assign m311_115 ={ {5{in311[5]}} , in311[5:1] };

   // m311_116 = W*in
   wire signed [9:0] m311_116;
   assign m311_116 ={ {4{in311[5]}} , in311[5:0] };

   // m311_117 = W*in
   wire signed [9:0] m311_117;
   assign m311_117 =10'b0;

   // m312_1 = W*in
   wire signed [9:0] m312_1;
   assign m312_1 =10'b0;

   // m312_2 = W*in
   wire signed [9:0] m312_2;
   assign m312_2 =10'b0;

   // m312_3 = W*in
   wire signed [9:0] m312_3;
   assign m312_3 =10'b0;

   // m312_4 = W*in
   wire signed [9:0] m312_4;
   assign m312_4 =10'b0;

   // m312_5 = W*in
   wire signed [9:0] m312_5;
   assign m312_5 =10'b0;

   // m312_6 = W*in
   wire signed [9:0] m312_6;
   assign m312_6 =10'b0;

   // m312_7 = W*in
   wire signed [9:0] m312_7;
   assign m312_7 =10'b0;

   // m312_8 = W*in
   wire signed [9:0] m312_8;
   assign m312_8 ={ {4{in312[5]}} , in312[5:0] };

   // m312_9 = W*in
   wire signed [9:0] m312_9;
   assign m312_9 =10'b0;

   // m312_10 = W*in
   wire signed [9:0] m312_10;
   assign m312_10 =10'b0;

   // m312_11 = W*in
   wire signed [9:0] m312_11;
   assign m312_11 =10'b0;

   // m312_12 = W*in
   wire signed [9:0] m312_12;
   assign m312_12 =10'b0;

   // m312_13 = W*in
   wire signed [9:0] m312_13;
   assign m312_13 =10'b0;

   // m312_14 = W*in
   wire signed [9:0] m312_14;
   assign m312_14 =10'b0;

   // m312_15 = W*in
   wire signed [9:0] m312_15;
   assign m312_15 =10'b0;

   // m312_16 = W*in
   wire signed [9:0] m312_16;
   assign m312_16 ={ {5{in312[5]}} , in312[5:1] };

   // m312_17 = W*in
   wire signed [9:0] m312_17;
   assign m312_17 =10'b0;

   // m312_18 = W*in
   wire signed [9:0] m312_18;
   assign m312_18 ={ {5{neg312[5]}} , neg312[5:1] };

   // m312_19 = W*in
   wire signed [9:0] m312_19;
   assign m312_19 =10'b0;

   // m312_20 = W*in
   wire signed [9:0] m312_20;
   assign m312_20 ={ {5{in312[5]}} , in312[5:1] };

   // m312_21 = W*in
   wire signed [9:0] m312_21;
   assign m312_21 =10'b0;

   // m312_22 = W*in
   wire signed [9:0] m312_22;
   assign m312_22 =10'b0;

   // m312_23 = W*in
   wire signed [9:0] m312_23;
   assign m312_23 =10'b0;

   // m312_24 = W*in
   wire signed [9:0] m312_24;
   assign m312_24 =10'b0;

   // m312_25 = W*in
   wire signed [9:0] m312_25;
   assign m312_25 =10'b0;

   // m312_26 = W*in
   wire signed [9:0] m312_26;
   assign m312_26 ={ {4{neg312[5]}} , neg312[5:0] };

   // m312_27 = W*in
   wire signed [9:0] m312_27;
   assign m312_27 ={ {5{neg312[5]}} , neg312[5:1] };

   // m312_28 = W*in
   wire signed [9:0] m312_28;
   assign m312_28 =10'b0;

   // m312_29 = W*in
   wire signed [9:0] m312_29;
   assign m312_29 =10'b0;

   // m312_30 = W*in
   wire signed [9:0] m312_30;
   assign m312_30 ={ {4{in312[5]}} , in312[5:0] };

   // m312_31 = W*in
   wire signed [9:0] m312_31;
   assign m312_31 ={ {4{in312[5]}} , in312[5:0] };

   // m312_32 = W*in
   wire signed [9:0] m312_32;
   assign m312_32 =10'b0;

   // m312_33 = W*in
   wire signed [9:0] m312_33;
   assign m312_33 ={ {4{neg312[5]}} , neg312[5:0] };

   // m312_34 = W*in
   wire signed [9:0] m312_34;
   assign m312_34 =10'b0;

   // m312_35 = W*in
   wire signed [9:0] m312_35;
   assign m312_35 ={ {5{in312[5]}} , in312[5:1] };

   // m312_36 = W*in
   wire signed [9:0] m312_36;
   assign m312_36 =10'b0;

   // m312_37 = W*in
   wire signed [9:0] m312_37;
   assign m312_37 =10'b0;

   // m312_38 = W*in
   wire signed [9:0] m312_38;
   assign m312_38 =10'b0;

   // m312_39 = W*in
   wire signed [9:0] m312_39;
   assign m312_39 =10'b0;

   // m312_40 = W*in
   wire signed [9:0] m312_40;
   assign m312_40 =10'b0;

   // m312_41 = W*in
   wire signed [9:0] m312_41;
   assign m312_41 ={ {4{in312[5]}} , in312[5:0] };

   // m312_42 = W*in
   wire signed [9:0] m312_42;
   assign m312_42 =10'b0;

   // m312_43 = W*in
   wire signed [9:0] m312_43;
   assign m312_43 ={ {4{neg312[5]}} , neg312[5:0] };

   // m312_44 = W*in
   wire signed [9:0] m312_44;
   assign m312_44 =10'b0;

   // m312_45 = W*in
   wire signed [9:0] m312_45;
   assign m312_45 =10'b0;

   // m312_46 = W*in
   wire signed [9:0] m312_46;
   assign m312_46 =10'b0;

   // m312_47 = W*in
   wire signed [9:0] m312_47;
   assign m312_47 =10'b0;

   // m312_48 = W*in
   wire signed [9:0] m312_48;
   assign m312_48 =10'b0;

   // m312_49 = W*in
   wire signed [9:0] m312_49;
   assign m312_49 =10'b0;

   // m312_50 = W*in
   wire signed [9:0] m312_50;
   assign m312_50 =10'b0;

   // m312_51 = W*in
   wire signed [9:0] m312_51;
   assign m312_51 =10'b0;

   // m312_52 = W*in
   wire signed [9:0] m312_52;
   assign m312_52 =10'b0;

   // m312_53 = W*in
   wire signed [9:0] m312_53;
   assign m312_53 =10'b0;

   // m312_54 = W*in
   wire signed [9:0] m312_54;
   assign m312_54 =10'b0;

   // m312_55 = W*in
   wire signed [9:0] m312_55;
   assign m312_55 =10'b0;

   // m312_56 = W*in
   wire signed [9:0] m312_56;
   assign m312_56 =10'b0;

   // m312_57 = W*in
   wire signed [9:0] m312_57;
   assign m312_57 =10'b0;

   // m312_58 = W*in
   wire signed [9:0] m312_58;
   assign m312_58 =10'b0;

   // m312_59 = W*in
   wire signed [9:0] m312_59;
   assign m312_59 =10'b0;

   // m312_60 = W*in
   wire signed [9:0] m312_60;
   assign m312_60 =10'b0;

   // m312_61 = W*in
   wire signed [9:0] m312_61;
   assign m312_61 =10'b0;

   // m312_62 = W*in
   wire signed [9:0] m312_62;
   assign m312_62 =10'b0;

   // m312_63 = W*in
   wire signed [9:0] m312_63;
   assign m312_63 =10'b0;

   // m312_64 = W*in
   wire signed [9:0] m312_64;
   assign m312_64 =10'b0;

   // m312_65 = W*in
   wire signed [9:0] m312_65;
   assign m312_65 =10'b0;

   // m312_66 = W*in
   wire signed [9:0] m312_66;
   assign m312_66 =10'b0;

   // m312_67 = W*in
   wire signed [9:0] m312_67;
   assign m312_67 =10'b0;

   // m312_68 = W*in
   wire signed [9:0] m312_68;
   assign m312_68 =10'b0;

   // m312_69 = W*in
   wire signed [9:0] m312_69;
   assign m312_69 ={ {5{neg312[5]}} , neg312[5:1] };

   // m312_70 = W*in
   wire signed [9:0] m312_70;
   assign m312_70 =10'b0;

   // m312_71 = W*in
   wire signed [9:0] m312_71;
   assign m312_71 =10'b0;

   // m312_72 = W*in
   wire signed [9:0] m312_72;
   assign m312_72 ={ {5{neg312[5]}} , neg312[5:1] };

   // m312_73 = W*in
   wire signed [9:0] m312_73;
   assign m312_73 =10'b0;

   // m312_74 = W*in
   wire signed [9:0] m312_74;
   assign m312_74 =10'b0;

   // m312_75 = W*in
   wire signed [9:0] m312_75;
   assign m312_75 =10'b0;

   // m312_76 = W*in
   wire signed [9:0] m312_76;
   assign m312_76 =10'b0;

   // m312_77 = W*in
   wire signed [9:0] m312_77;
   assign m312_77 =10'b0;

   // m312_78 = W*in
   wire signed [9:0] m312_78;
   assign m312_78 ={ {4{neg312[5]}} , neg312[5:0] };

   // m312_79 = W*in
   wire signed [9:0] m312_79;
   assign m312_79 ={ {4{in312[5]}} , in312[5:0] };

   // m312_80 = W*in
   wire signed [9:0] m312_80;
   assign m312_80 ={ {4{in312[5]}} , in312[5:0] };

   // m312_81 = W*in
   wire signed [9:0] m312_81;
   assign m312_81 ={ {5{in312[5]}} , in312[5:1] };

   // m312_82 = W*in
   wire signed [9:0] m312_82;
   assign m312_82 =10'b0;

   // m312_83 = W*in
   wire signed [9:0] m312_83;
   assign m312_83 =10'b0;

   // m312_84 = W*in
   wire signed [9:0] m312_84;
   assign m312_84 ={ {5{neg312[5]}} , neg312[5:1] };

   // m312_85 = W*in
   wire signed [9:0] m312_85;
   assign m312_85 =10'b0;

   // m312_86 = W*in
   wire signed [9:0] m312_86;
   assign m312_86 =10'b0;

   // m312_87 = W*in
   wire signed [9:0] m312_87;
   assign m312_87 =10'b0;

   // m312_88 = W*in
   wire signed [9:0] m312_88;
   assign m312_88 =10'b0;

   // m312_89 = W*in
   wire signed [9:0] m312_89;
   assign m312_89 =10'b0;

   // m312_90 = W*in
   wire signed [9:0] m312_90;
   assign m312_90 =10'b0;

   // m312_91 = W*in
   wire signed [9:0] m312_91;
   assign m312_91 =10'b0;

   // m312_92 = W*in
   wire signed [9:0] m312_92;
   assign m312_92 =10'b0;

   // m312_93 = W*in
   wire signed [9:0] m312_93;
   assign m312_93 =10'b0;

   // m312_94 = W*in
   wire signed [9:0] m312_94;
   assign m312_94 =10'b0;

   // m312_95 = W*in
   wire signed [9:0] m312_95;
   assign m312_95 =10'b0;

   // m312_96 = W*in
   wire signed [9:0] m312_96;
   assign m312_96 =10'b0;

   // m312_97 = W*in
   wire signed [9:0] m312_97;
   assign m312_97 =10'b0;

   // m312_98 = W*in
   wire signed [9:0] m312_98;
   assign m312_98 ={ {4{in312[5]}} , in312[5:0] };

   // m312_99 = W*in
   wire signed [9:0] m312_99;
   assign m312_99 =10'b0;

   // m312_100 = W*in
   wire signed [9:0] m312_100;
   assign m312_100 =10'b0;

   // m312_101 = W*in
   wire signed [9:0] m312_101;
   assign m312_101 =10'b0;

   // m312_102 = W*in
   wire signed [9:0] m312_102;
   assign m312_102 =10'b0;

   // m312_103 = W*in
   wire signed [9:0] m312_103;
   assign m312_103 =10'b0;

   // m312_104 = W*in
   wire signed [9:0] m312_104;
   assign m312_104 =10'b0;

   // m312_105 = W*in
   wire signed [9:0] m312_105;
   assign m312_105 =10'b0;

   // m312_106 = W*in
   wire signed [9:0] m312_106;
   assign m312_106 =10'b0;

   // m312_107 = W*in
   wire signed [9:0] m312_107;
   assign m312_107 =10'b0;

   // m312_108 = W*in
   wire signed [9:0] m312_108;
   assign m312_108 ={ {4{in312[5]}} , in312[5:0] };

   // m312_109 = W*in
   wire signed [9:0] m312_109;
   assign m312_109 ={ {5{in312[5]}} , in312[5:1] };

   // m312_110 = W*in
   wire signed [9:0] m312_110;
   assign m312_110 =10'b0;

   // m312_111 = W*in
   wire signed [9:0] m312_111;
   assign m312_111 =10'b0;

   // m312_112 = W*in
   wire signed [9:0] m312_112;
   assign m312_112 =10'b0;

   // m312_113 = W*in
   wire signed [9:0] m312_113;
   assign m312_113 =10'b0;

   // m312_114 = W*in
   wire signed [9:0] m312_114;
   assign m312_114 =10'b0;

   // m312_115 = W*in
   wire signed [9:0] m312_115;
   assign m312_115 ={ {5{in312[5]}} , in312[5:1] };

   // m312_116 = W*in
   wire signed [9:0] m312_116;
   assign m312_116 ={ {4{in312[5]}} , in312[5:0] };

   // m312_117 = W*in
   wire signed [9:0] m312_117;
   assign m312_117 =10'b0;

   // m313_1 = W*in
   wire signed [9:0] m313_1;
   assign m313_1 =10'b0;

   // m313_2 = W*in
   wire signed [9:0] m313_2;
   assign m313_2 =10'b0;

   // m313_3 = W*in
   wire signed [9:0] m313_3;
   assign m313_3 =10'b0;

   // m313_4 = W*in
   wire signed [9:0] m313_4;
   assign m313_4 =10'b0;

   // m313_5 = W*in
   wire signed [9:0] m313_5;
   assign m313_5 =10'b0;

   // m313_6 = W*in
   wire signed [9:0] m313_6;
   assign m313_6 =10'b0;

   // m313_7 = W*in
   wire signed [9:0] m313_7;
   assign m313_7 =10'b0;

   // m313_8 = W*in
   wire signed [9:0] m313_8;
   assign m313_8 =10'b0;

   // m313_9 = W*in
   wire signed [9:0] m313_9;
   assign m313_9 =10'b0;

   // m313_10 = W*in
   wire signed [9:0] m313_10;
   assign m313_10 =10'b0;

   // m313_11 = W*in
   wire signed [9:0] m313_11;
   assign m313_11 =10'b0;

   // m313_12 = W*in
   wire signed [9:0] m313_12;
   assign m313_12 =10'b0;

   // m313_13 = W*in
   wire signed [9:0] m313_13;
   assign m313_13 =10'b0;

   // m313_14 = W*in
   wire signed [9:0] m313_14;
   assign m313_14 =10'b0;

   // m313_15 = W*in
   wire signed [9:0] m313_15;
   assign m313_15 =10'b0;

   // m313_16 = W*in
   wire signed [9:0] m313_16;
   assign m313_16 =10'b0;

   // m313_17 = W*in
   wire signed [9:0] m313_17;
   assign m313_17 =10'b0;

   // m313_18 = W*in
   wire signed [9:0] m313_18;
   assign m313_18 ={ {5{neg313[5]}} , neg313[5:1] };

   // m313_19 = W*in
   wire signed [9:0] m313_19;
   assign m313_19 =10'b0;

   // m313_20 = W*in
   wire signed [9:0] m313_20;
   assign m313_20 ={ {5{in313[5]}} , in313[5:1] };

   // m313_21 = W*in
   wire signed [9:0] m313_21;
   assign m313_21 =10'b0;

   // m313_22 = W*in
   wire signed [9:0] m313_22;
   assign m313_22 =10'b0;

   // m313_23 = W*in
   wire signed [9:0] m313_23;
   assign m313_23 =10'b0;

   // m313_24 = W*in
   wire signed [9:0] m313_24;
   assign m313_24 =10'b0;

   // m313_25 = W*in
   wire signed [9:0] m313_25;
   assign m313_25 =10'b0;

   // m313_26 = W*in
   wire signed [9:0] m313_26;
   assign m313_26 ={ {5{neg313[5]}} , neg313[5:1] };

   // m313_27 = W*in
   wire signed [9:0] m313_27;
   assign m313_27 =10'b0;

   // m313_28 = W*in
   wire signed [9:0] m313_28;
   assign m313_28 =10'b0;

   // m313_29 = W*in
   wire signed [9:0] m313_29;
   assign m313_29 =10'b0;

   // m313_30 = W*in
   wire signed [9:0] m313_30;
   assign m313_30 ={ {5{in313[5]}} , in313[5:1] };

   // m313_31 = W*in
   wire signed [9:0] m313_31;
   assign m313_31 =10'b0;

   // m313_32 = W*in
   wire signed [9:0] m313_32;
   assign m313_32 =10'b0;

   // m313_33 = W*in
   wire signed [9:0] m313_33;
   assign m313_33 =10'b0;

   // m313_34 = W*in
   wire signed [9:0] m313_34;
   assign m313_34 =10'b0;

   // m313_35 = W*in
   wire signed [9:0] m313_35;
   assign m313_35 =10'b0;

   // m313_36 = W*in
   wire signed [9:0] m313_36;
   assign m313_36 =10'b0;

   // m313_37 = W*in
   wire signed [9:0] m313_37;
   assign m313_37 =10'b0;

   // m313_38 = W*in
   wire signed [9:0] m313_38;
   assign m313_38 =10'b0;

   // m313_39 = W*in
   wire signed [9:0] m313_39;
   assign m313_39 =10'b0;

   // m313_40 = W*in
   wire signed [9:0] m313_40;
   assign m313_40 =10'b0;

   // m313_41 = W*in
   wire signed [9:0] m313_41;
   assign m313_41 =10'b0;

   // m313_42 = W*in
   wire signed [9:0] m313_42;
   assign m313_42 =10'b0;

   // m313_43 = W*in
   wire signed [9:0] m313_43;
   assign m313_43 =10'b0;

   // m313_44 = W*in
   wire signed [9:0] m313_44;
   assign m313_44 =10'b0;

   // m313_45 = W*in
   wire signed [9:0] m313_45;
   assign m313_45 =10'b0;

   // m313_46 = W*in
   wire signed [9:0] m313_46;
   assign m313_46 =10'b0;

   // m313_47 = W*in
   wire signed [9:0] m313_47;
   assign m313_47 =10'b0;

   // m313_48 = W*in
   wire signed [9:0] m313_48;
   assign m313_48 =10'b0;

   // m313_49 = W*in
   wire signed [9:0] m313_49;
   assign m313_49 =10'b0;

   // m313_50 = W*in
   wire signed [9:0] m313_50;
   assign m313_50 =10'b0;

   // m313_51 = W*in
   wire signed [9:0] m313_51;
   assign m313_51 =10'b0;

   // m313_52 = W*in
   wire signed [9:0] m313_52;
   assign m313_52 =10'b0;

   // m313_53 = W*in
   wire signed [9:0] m313_53;
   assign m313_53 =10'b0;

   // m313_54 = W*in
   wire signed [9:0] m313_54;
   assign m313_54 =10'b0;

   // m313_55 = W*in
   wire signed [9:0] m313_55;
   assign m313_55 =10'b0;

   // m313_56 = W*in
   wire signed [9:0] m313_56;
   assign m313_56 =10'b0;

   // m313_57 = W*in
   wire signed [9:0] m313_57;
   assign m313_57 =10'b0;

   // m313_58 = W*in
   wire signed [9:0] m313_58;
   assign m313_58 =10'b0;

   // m313_59 = W*in
   wire signed [9:0] m313_59;
   assign m313_59 =10'b0;

   // m313_60 = W*in
   wire signed [9:0] m313_60;
   assign m313_60 =10'b0;

   // m313_61 = W*in
   wire signed [9:0] m313_61;
   assign m313_61 =10'b0;

   // m313_62 = W*in
   wire signed [9:0] m313_62;
   assign m313_62 =10'b0;

   // m313_63 = W*in
   wire signed [9:0] m313_63;
   assign m313_63 =10'b0;

   // m313_64 = W*in
   wire signed [9:0] m313_64;
   assign m313_64 =10'b0;

   // m313_65 = W*in
   wire signed [9:0] m313_65;
   assign m313_65 =10'b0;

   // m313_66 = W*in
   wire signed [9:0] m313_66;
   assign m313_66 =10'b0;

   // m313_67 = W*in
   wire signed [9:0] m313_67;
   assign m313_67 =10'b0;

   // m313_68 = W*in
   wire signed [9:0] m313_68;
   assign m313_68 =10'b0;

   // m313_69 = W*in
   wire signed [9:0] m313_69;
   assign m313_69 =10'b0;

   // m313_70 = W*in
   wire signed [9:0] m313_70;
   assign m313_70 =10'b0;

   // m313_71 = W*in
   wire signed [9:0] m313_71;
   assign m313_71 =10'b0;

   // m313_72 = W*in
   wire signed [9:0] m313_72;
   assign m313_72 =10'b0;

   // m313_73 = W*in
   wire signed [9:0] m313_73;
   assign m313_73 =10'b0;

   // m313_74 = W*in
   wire signed [9:0] m313_74;
   assign m313_74 =10'b0;

   // m313_75 = W*in
   wire signed [9:0] m313_75;
   assign m313_75 =10'b0;

   // m313_76 = W*in
   wire signed [9:0] m313_76;
   assign m313_76 =10'b0;

   // m313_77 = W*in
   wire signed [9:0] m313_77;
   assign m313_77 =10'b0;

   // m313_78 = W*in
   wire signed [9:0] m313_78;
   assign m313_78 =10'b0;

   // m313_79 = W*in
   wire signed [9:0] m313_79;
   assign m313_79 =10'b0;

   // m313_80 = W*in
   wire signed [9:0] m313_80;
   assign m313_80 ={ {5{in313[5]}} , in313[5:1] };

   // m313_81 = W*in
   wire signed [9:0] m313_81;
   assign m313_81 =10'b0;

   // m313_82 = W*in
   wire signed [9:0] m313_82;
   assign m313_82 =10'b0;

   // m313_83 = W*in
   wire signed [9:0] m313_83;
   assign m313_83 ={ {5{in313[5]}} , in313[5:1] };

   // m313_84 = W*in
   wire signed [9:0] m313_84;
   assign m313_84 =10'b0;

   // m313_85 = W*in
   wire signed [9:0] m313_85;
   assign m313_85 =10'b0;

   // m313_86 = W*in
   wire signed [9:0] m313_86;
   assign m313_86 =10'b0;

   // m313_87 = W*in
   wire signed [9:0] m313_87;
   assign m313_87 =10'b0;

   // m313_88 = W*in
   wire signed [9:0] m313_88;
   assign m313_88 =10'b0;

   // m313_89 = W*in
   wire signed [9:0] m313_89;
   assign m313_89 =10'b0;

   // m313_90 = W*in
   wire signed [9:0] m313_90;
   assign m313_90 =10'b0;

   // m313_91 = W*in
   wire signed [9:0] m313_91;
   assign m313_91 =10'b0;

   // m313_92 = W*in
   wire signed [9:0] m313_92;
   assign m313_92 =10'b0;

   // m313_93 = W*in
   wire signed [9:0] m313_93;
   assign m313_93 =10'b0;

   // m313_94 = W*in
   wire signed [9:0] m313_94;
   assign m313_94 =10'b0;

   // m313_95 = W*in
   wire signed [9:0] m313_95;
   assign m313_95 =10'b0;

   // m313_96 = W*in
   wire signed [9:0] m313_96;
   assign m313_96 =10'b0;

   // m313_97 = W*in
   wire signed [9:0] m313_97;
   assign m313_97 =10'b0;

   // m313_98 = W*in
   wire signed [9:0] m313_98;
   assign m313_98 =10'b0;

   // m313_99 = W*in
   wire signed [9:0] m313_99;
   assign m313_99 =10'b0;

   // m313_100 = W*in
   wire signed [9:0] m313_100;
   assign m313_100 =10'b0;

   // m313_101 = W*in
   wire signed [9:0] m313_101;
   assign m313_101 =10'b0;

   // m313_102 = W*in
   wire signed [9:0] m313_102;
   assign m313_102 =10'b0;

   // m313_103 = W*in
   wire signed [9:0] m313_103;
   assign m313_103 =10'b0;

   // m313_104 = W*in
   wire signed [9:0] m313_104;
   assign m313_104 =10'b0;

   // m313_105 = W*in
   wire signed [9:0] m313_105;
   assign m313_105 =10'b0;

   // m313_106 = W*in
   wire signed [9:0] m313_106;
   assign m313_106 =10'b0;

   // m313_107 = W*in
   wire signed [9:0] m313_107;
   assign m313_107 =10'b0;

   // m313_108 = W*in
   wire signed [9:0] m313_108;
   assign m313_108 =10'b0;

   // m313_109 = W*in
   wire signed [9:0] m313_109;
   assign m313_109 =10'b0;

   // m313_110 = W*in
   wire signed [9:0] m313_110;
   assign m313_110 =10'b0;

   // m313_111 = W*in
   wire signed [9:0] m313_111;
   assign m313_111 =10'b0;

   // m313_112 = W*in
   wire signed [9:0] m313_112;
   assign m313_112 =10'b0;

   // m313_113 = W*in
   wire signed [9:0] m313_113;
   assign m313_113 =10'b0;

   // m313_114 = W*in
   wire signed [9:0] m313_114;
   assign m313_114 =10'b0;

   // m313_115 = W*in
   wire signed [9:0] m313_115;
   assign m313_115 =10'b0;

   // m313_116 = W*in
   wire signed [9:0] m313_116;
   assign m313_116 =10'b0;

   // m313_117 = W*in
   wire signed [9:0] m313_117;
   assign m313_117 =10'b0;

   // m314_1 = W*in
   wire signed [9:0] m314_1;
   assign m314_1 =10'b0;

   // m314_2 = W*in
   wire signed [9:0] m314_2;
   assign m314_2 =10'b0;

   // m314_3 = W*in
   wire signed [9:0] m314_3;
   assign m314_3 =10'b0;

   // m314_4 = W*in
   wire signed [9:0] m314_4;
   assign m314_4 =10'b0;

   // m314_5 = W*in
   wire signed [9:0] m314_5;
   assign m314_5 =10'b0;

   // m314_6 = W*in
   wire signed [9:0] m314_6;
   assign m314_6 =10'b0;

   // m314_7 = W*in
   wire signed [9:0] m314_7;
   assign m314_7 =10'b0;

   // m314_8 = W*in
   wire signed [9:0] m314_8;
   assign m314_8 =10'b0;

   // m314_9 = W*in
   wire signed [9:0] m314_9;
   assign m314_9 =10'b0;

   // m314_10 = W*in
   wire signed [9:0] m314_10;
   assign m314_10 =10'b0;

   // m314_11 = W*in
   wire signed [9:0] m314_11;
   assign m314_11 =10'b0;

   // m314_12 = W*in
   wire signed [9:0] m314_12;
   assign m314_12 =10'b0;

   // m314_13 = W*in
   wire signed [9:0] m314_13;
   assign m314_13 =10'b0;

   // m314_14 = W*in
   wire signed [9:0] m314_14;
   assign m314_14 =10'b0;

   // m314_15 = W*in
   wire signed [9:0] m314_15;
   assign m314_15 =10'b0;

   // m314_16 = W*in
   wire signed [9:0] m314_16;
   assign m314_16 =10'b0;

   // m314_17 = W*in
   wire signed [9:0] m314_17;
   assign m314_17 =10'b0;

   // m314_18 = W*in
   wire signed [9:0] m314_18;
   assign m314_18 =10'b0;

   // m314_19 = W*in
   wire signed [9:0] m314_19;
   assign m314_19 ={ {5{in314[5]}} , in314[5:1] };

   // m314_20 = W*in
   wire signed [9:0] m314_20;
   assign m314_20 ={ {5{in314[5]}} , in314[5:1] };

   // m314_21 = W*in
   wire signed [9:0] m314_21;
   assign m314_21 =10'b0;

   // m314_22 = W*in
   wire signed [9:0] m314_22;
   assign m314_22 =10'b0;

   // m314_23 = W*in
   wire signed [9:0] m314_23;
   assign m314_23 =10'b0;

   // m314_24 = W*in
   wire signed [9:0] m314_24;
   assign m314_24 =10'b0;

   // m314_25 = W*in
   wire signed [9:0] m314_25;
   assign m314_25 =10'b0;

   // m314_26 = W*in
   wire signed [9:0] m314_26;
   assign m314_26 ={ {5{neg314[5]}} , neg314[5:1] };

   // m314_27 = W*in
   wire signed [9:0] m314_27;
   assign m314_27 ={ {5{in314[5]}} , in314[5:1] };

   // m314_28 = W*in
   wire signed [9:0] m314_28;
   assign m314_28 =10'b0;

   // m314_29 = W*in
   wire signed [9:0] m314_29;
   assign m314_29 =10'b0;

   // m314_30 = W*in
   wire signed [9:0] m314_30;
   assign m314_30 ={ {5{in314[5]}} , in314[5:1] };

   // m314_31 = W*in
   wire signed [9:0] m314_31;
   assign m314_31 =10'b0;

   // m314_32 = W*in
   wire signed [9:0] m314_32;
   assign m314_32 =10'b0;

   // m314_33 = W*in
   wire signed [9:0] m314_33;
   assign m314_33 =10'b0;

   // m314_34 = W*in
   wire signed [9:0] m314_34;
   assign m314_34 =10'b0;

   // m314_35 = W*in
   wire signed [9:0] m314_35;
   assign m314_35 ={ {5{in314[5]}} , in314[5:1] };

   // m314_36 = W*in
   wire signed [9:0] m314_36;
   assign m314_36 =10'b0;

   // m314_37 = W*in
   wire signed [9:0] m314_37;
   assign m314_37 =10'b0;

   // m314_38 = W*in
   wire signed [9:0] m314_38;
   assign m314_38 =10'b0;

   // m314_39 = W*in
   wire signed [9:0] m314_39;
   assign m314_39 =10'b0;

   // m314_40 = W*in
   wire signed [9:0] m314_40;
   assign m314_40 =10'b0;

   // m314_41 = W*in
   wire signed [9:0] m314_41;
   assign m314_41 =10'b0;

   // m314_42 = W*in
   wire signed [9:0] m314_42;
   assign m314_42 =10'b0;

   // m314_43 = W*in
   wire signed [9:0] m314_43;
   assign m314_43 =10'b0;

   // m314_44 = W*in
   wire signed [9:0] m314_44;
   assign m314_44 =10'b0;

   // m314_45 = W*in
   wire signed [9:0] m314_45;
   assign m314_45 =10'b0;

   // m314_46 = W*in
   wire signed [9:0] m314_46;
   assign m314_46 =10'b0;

   // m314_47 = W*in
   wire signed [9:0] m314_47;
   assign m314_47 =10'b0;

   // m314_48 = W*in
   wire signed [9:0] m314_48;
   assign m314_48 =10'b0;

   // m314_49 = W*in
   wire signed [9:0] m314_49;
   assign m314_49 =10'b0;

   // m314_50 = W*in
   wire signed [9:0] m314_50;
   assign m314_50 =10'b0;

   // m314_51 = W*in
   wire signed [9:0] m314_51;
   assign m314_51 =10'b0;

   // m314_52 = W*in
   wire signed [9:0] m314_52;
   assign m314_52 =10'b0;

   // m314_53 = W*in
   wire signed [9:0] m314_53;
   assign m314_53 =10'b0;

   // m314_54 = W*in
   wire signed [9:0] m314_54;
   assign m314_54 =10'b0;

   // m314_55 = W*in
   wire signed [9:0] m314_55;
   assign m314_55 =10'b0;

   // m314_56 = W*in
   wire signed [9:0] m314_56;
   assign m314_56 =10'b0;

   // m314_57 = W*in
   wire signed [9:0] m314_57;
   assign m314_57 =10'b0;

   // m314_58 = W*in
   wire signed [9:0] m314_58;
   assign m314_58 =10'b0;

   // m314_59 = W*in
   wire signed [9:0] m314_59;
   assign m314_59 =10'b0;

   // m314_60 = W*in
   wire signed [9:0] m314_60;
   assign m314_60 =10'b0;

   // m314_61 = W*in
   wire signed [9:0] m314_61;
   assign m314_61 =10'b0;

   // m314_62 = W*in
   wire signed [9:0] m314_62;
   assign m314_62 =10'b0;

   // m314_63 = W*in
   wire signed [9:0] m314_63;
   assign m314_63 =10'b0;

   // m314_64 = W*in
   wire signed [9:0] m314_64;
   assign m314_64 =10'b0;

   // m314_65 = W*in
   wire signed [9:0] m314_65;
   assign m314_65 =10'b0;

   // m314_66 = W*in
   wire signed [9:0] m314_66;
   assign m314_66 =10'b0;

   // m314_67 = W*in
   wire signed [9:0] m314_67;
   assign m314_67 =10'b0;

   // m314_68 = W*in
   wire signed [9:0] m314_68;
   assign m314_68 =10'b0;

   // m314_69 = W*in
   wire signed [9:0] m314_69;
   assign m314_69 =10'b0;

   // m314_70 = W*in
   wire signed [9:0] m314_70;
   assign m314_70 =10'b0;

   // m314_71 = W*in
   wire signed [9:0] m314_71;
   assign m314_71 =10'b0;

   // m314_72 = W*in
   wire signed [9:0] m314_72;
   assign m314_72 =10'b0;

   // m314_73 = W*in
   wire signed [9:0] m314_73;
   assign m314_73 =10'b0;

   // m314_74 = W*in
   wire signed [9:0] m314_74;
   assign m314_74 =10'b0;

   // m314_75 = W*in
   wire signed [9:0] m314_75;
   assign m314_75 =10'b0;

   // m314_76 = W*in
   wire signed [9:0] m314_76;
   assign m314_76 =10'b0;

   // m314_77 = W*in
   wire signed [9:0] m314_77;
   assign m314_77 =10'b0;

   // m314_78 = W*in
   wire signed [9:0] m314_78;
   assign m314_78 =10'b0;

   // m314_79 = W*in
   wire signed [9:0] m314_79;
   assign m314_79 =10'b0;

   // m314_80 = W*in
   wire signed [9:0] m314_80;
   assign m314_80 =10'b0;

   // m314_81 = W*in
   wire signed [9:0] m314_81;
   assign m314_81 =10'b0;

   // m314_82 = W*in
   wire signed [9:0] m314_82;
   assign m314_82 =10'b0;

   // m314_83 = W*in
   wire signed [9:0] m314_83;
   assign m314_83 =10'b0;

   // m314_84 = W*in
   wire signed [9:0] m314_84;
   assign m314_84 =10'b0;

   // m314_85 = W*in
   wire signed [9:0] m314_85;
   assign m314_85 =10'b0;

   // m314_86 = W*in
   wire signed [9:0] m314_86;
   assign m314_86 =10'b0;

   // m314_87 = W*in
   wire signed [9:0] m314_87;
   assign m314_87 =10'b0;

   // m314_88 = W*in
   wire signed [9:0] m314_88;
   assign m314_88 =10'b0;

   // m314_89 = W*in
   wire signed [9:0] m314_89;
   assign m314_89 =10'b0;

   // m314_90 = W*in
   wire signed [9:0] m314_90;
   assign m314_90 =10'b0;

   // m314_91 = W*in
   wire signed [9:0] m314_91;
   assign m314_91 =10'b0;

   // m314_92 = W*in
   wire signed [9:0] m314_92;
   assign m314_92 =10'b0;

   // m314_93 = W*in
   wire signed [9:0] m314_93;
   assign m314_93 =10'b0;

   // m314_94 = W*in
   wire signed [9:0] m314_94;
   assign m314_94 =10'b0;

   // m314_95 = W*in
   wire signed [9:0] m314_95;
   assign m314_95 =10'b0;

   // m314_96 = W*in
   wire signed [9:0] m314_96;
   assign m314_96 =10'b0;

   // m314_97 = W*in
   wire signed [9:0] m314_97;
   assign m314_97 =10'b0;

   // m314_98 = W*in
   wire signed [9:0] m314_98;
   assign m314_98 =10'b0;

   // m314_99 = W*in
   wire signed [9:0] m314_99;
   assign m314_99 =10'b0;

   // m314_100 = W*in
   wire signed [9:0] m314_100;
   assign m314_100 =10'b0;

   // m314_101 = W*in
   wire signed [9:0] m314_101;
   assign m314_101 =10'b0;

   // m314_102 = W*in
   wire signed [9:0] m314_102;
   assign m314_102 =10'b0;

   // m314_103 = W*in
   wire signed [9:0] m314_103;
   assign m314_103 =10'b0;

   // m314_104 = W*in
   wire signed [9:0] m314_104;
   assign m314_104 =10'b0;

   // m314_105 = W*in
   wire signed [9:0] m314_105;
   assign m314_105 =10'b0;

   // m314_106 = W*in
   wire signed [9:0] m314_106;
   assign m314_106 =10'b0;

   // m314_107 = W*in
   wire signed [9:0] m314_107;
   assign m314_107 =10'b0;

   // m314_108 = W*in
   wire signed [9:0] m314_108;
   assign m314_108 ={ {5{in314[5]}} , in314[5:1] };

   // m314_109 = W*in
   wire signed [9:0] m314_109;
   assign m314_109 =10'b0;

   // m314_110 = W*in
   wire signed [9:0] m314_110;
   assign m314_110 =10'b0;

   // m314_111 = W*in
   wire signed [9:0] m314_111;
   assign m314_111 =10'b0;

   // m314_112 = W*in
   wire signed [9:0] m314_112;
   assign m314_112 =10'b0;

   // m314_113 = W*in
   wire signed [9:0] m314_113;
   assign m314_113 =10'b0;

   // m314_114 = W*in
   wire signed [9:0] m314_114;
   assign m314_114 =10'b0;

   // m314_115 = W*in
   wire signed [9:0] m314_115;
   assign m314_115 =10'b0;

   // m314_116 = W*in
   wire signed [9:0] m314_116;
   assign m314_116 =10'b0;

   // m314_117 = W*in
   wire signed [9:0] m314_117;
   assign m314_117 =10'b0;

   // m315_1 = W*in
   wire signed [9:0] m315_1;
   assign m315_1 =10'b0;

   // m315_2 = W*in
   wire signed [9:0] m315_2;
   assign m315_2 =10'b0;

   // m315_3 = W*in
   wire signed [9:0] m315_3;
   assign m315_3 =10'b0;

   // m315_4 = W*in
   wire signed [9:0] m315_4;
   assign m315_4 =10'b0;

   // m315_5 = W*in
   wire signed [9:0] m315_5;
   assign m315_5 =10'b0;

   // m315_6 = W*in
   wire signed [9:0] m315_6;
   assign m315_6 =10'b0;

   // m315_7 = W*in
   wire signed [9:0] m315_7;
   assign m315_7 =10'b0;

   // m315_8 = W*in
   wire signed [9:0] m315_8;
   assign m315_8 =10'b0;

   // m315_9 = W*in
   wire signed [9:0] m315_9;
   assign m315_9 =10'b0;

   // m315_10 = W*in
   wire signed [9:0] m315_10;
   assign m315_10 =10'b0;

   // m315_11 = W*in
   wire signed [9:0] m315_11;
   assign m315_11 =10'b0;

   // m315_12 = W*in
   wire signed [9:0] m315_12;
   assign m315_12 =10'b0;

   // m315_13 = W*in
   wire signed [9:0] m315_13;
   assign m315_13 =10'b0;

   // m315_14 = W*in
   wire signed [9:0] m315_14;
   assign m315_14 =10'b0;

   // m315_15 = W*in
   wire signed [9:0] m315_15;
   assign m315_15 =10'b0;

   // m315_16 = W*in
   wire signed [9:0] m315_16;
   assign m315_16 =10'b0;

   // m315_17 = W*in
   wire signed [9:0] m315_17;
   assign m315_17 ={ {5{in315[5]}} , in315[5:1] };

   // m315_18 = W*in
   wire signed [9:0] m315_18;
   assign m315_18 ={ {5{neg315[5]}} , neg315[5:1] };

   // m315_19 = W*in
   wire signed [9:0] m315_19;
   assign m315_19 =10'b0;

   // m315_20 = W*in
   wire signed [9:0] m315_20;
   assign m315_20 ={ {4{in315[5]}} , in315[5:0] };

   // m315_21 = W*in
   wire signed [9:0] m315_21;
   assign m315_21 =10'b0;

   // m315_22 = W*in
   wire signed [9:0] m315_22;
   assign m315_22 =10'b0;

   // m315_23 = W*in
   wire signed [9:0] m315_23;
   assign m315_23 =10'b0;

   // m315_24 = W*in
   wire signed [9:0] m315_24;
   assign m315_24 =10'b0;

   // m315_25 = W*in
   wire signed [9:0] m315_25;
   assign m315_25 ={ {5{neg315[5]}} , neg315[5:1] };

   // m315_26 = W*in
   wire signed [9:0] m315_26;
   assign m315_26 =10'b0;

   // m315_27 = W*in
   wire signed [9:0] m315_27;
   assign m315_27 ={ {5{in315[5]}} , in315[5:1] };

   // m315_28 = W*in
   wire signed [9:0] m315_28;
   assign m315_28 =10'b0;

   // m315_29 = W*in
   wire signed [9:0] m315_29;
   assign m315_29 =10'b0;

   // m315_30 = W*in
   wire signed [9:0] m315_30;
   assign m315_30 =10'b0;

   // m315_31 = W*in
   wire signed [9:0] m315_31;
   assign m315_31 =10'b0;

   // m315_32 = W*in
   wire signed [9:0] m315_32;
   assign m315_32 =10'b0;

   // m315_33 = W*in
   wire signed [9:0] m315_33;
   assign m315_33 =10'b0;

   // m315_34 = W*in
   wire signed [9:0] m315_34;
   assign m315_34 =10'b0;

   // m315_35 = W*in
   wire signed [9:0] m315_35;
   assign m315_35 =10'b0;

   // m315_36 = W*in
   wire signed [9:0] m315_36;
   assign m315_36 =10'b0;

   // m315_37 = W*in
   wire signed [9:0] m315_37;
   assign m315_37 =10'b0;

   // m315_38 = W*in
   wire signed [9:0] m315_38;
   assign m315_38 =10'b0;

   // m315_39 = W*in
   wire signed [9:0] m315_39;
   assign m315_39 =10'b0;

   // m315_40 = W*in
   wire signed [9:0] m315_40;
   assign m315_40 =10'b0;

   // m315_41 = W*in
   wire signed [9:0] m315_41;
   assign m315_41 ={ {4{in315[5]}} , in315[5:0] };

   // m315_42 = W*in
   wire signed [9:0] m315_42;
   assign m315_42 =10'b0;

   // m315_43 = W*in
   wire signed [9:0] m315_43;
   assign m315_43 =10'b0;

   // m315_44 = W*in
   wire signed [9:0] m315_44;
   assign m315_44 =10'b0;

   // m315_45 = W*in
   wire signed [9:0] m315_45;
   assign m315_45 =10'b0;

   // m315_46 = W*in
   wire signed [9:0] m315_46;
   assign m315_46 =10'b0;

   // m315_47 = W*in
   wire signed [9:0] m315_47;
   assign m315_47 =10'b0;

   // m315_48 = W*in
   wire signed [9:0] m315_48;
   assign m315_48 =10'b0;

   // m315_49 = W*in
   wire signed [9:0] m315_49;
   assign m315_49 =10'b0;

   // m315_50 = W*in
   wire signed [9:0] m315_50;
   assign m315_50 =10'b0;

   // m315_51 = W*in
   wire signed [9:0] m315_51;
   assign m315_51 =10'b0;

   // m315_52 = W*in
   wire signed [9:0] m315_52;
   assign m315_52 =10'b0;

   // m315_53 = W*in
   wire signed [9:0] m315_53;
   assign m315_53 =10'b0;

   // m315_54 = W*in
   wire signed [9:0] m315_54;
   assign m315_54 =10'b0;

   // m315_55 = W*in
   wire signed [9:0] m315_55;
   assign m315_55 =10'b0;

   // m315_56 = W*in
   wire signed [9:0] m315_56;
   assign m315_56 =10'b0;

   // m315_57 = W*in
   wire signed [9:0] m315_57;
   assign m315_57 =10'b0;

   // m315_58 = W*in
   wire signed [9:0] m315_58;
   assign m315_58 =10'b0;

   // m315_59 = W*in
   wire signed [9:0] m315_59;
   assign m315_59 =10'b0;

   // m315_60 = W*in
   wire signed [9:0] m315_60;
   assign m315_60 =10'b0;

   // m315_61 = W*in
   wire signed [9:0] m315_61;
   assign m315_61 =10'b0;

   // m315_62 = W*in
   wire signed [9:0] m315_62;
   assign m315_62 =10'b0;

   // m315_63 = W*in
   wire signed [9:0] m315_63;
   assign m315_63 =10'b0;

   // m315_64 = W*in
   wire signed [9:0] m315_64;
   assign m315_64 ={ {5{neg315[5]}} , neg315[5:1] };

   // m315_65 = W*in
   wire signed [9:0] m315_65;
   assign m315_65 =10'b0;

   // m315_66 = W*in
   wire signed [9:0] m315_66;
   assign m315_66 =10'b0;

   // m315_67 = W*in
   wire signed [9:0] m315_67;
   assign m315_67 =10'b0;

   // m315_68 = W*in
   wire signed [9:0] m315_68;
   assign m315_68 =10'b0;

   // m315_69 = W*in
   wire signed [9:0] m315_69;
   assign m315_69 =10'b0;

   // m315_70 = W*in
   wire signed [9:0] m315_70;
   assign m315_70 =10'b0;

   // m315_71 = W*in
   wire signed [9:0] m315_71;
   assign m315_71 =10'b0;

   // m315_72 = W*in
   wire signed [9:0] m315_72;
   assign m315_72 =10'b0;

   // m315_73 = W*in
   wire signed [9:0] m315_73;
   assign m315_73 ={ {5{neg315[5]}} , neg315[5:1] };

   // m315_74 = W*in
   wire signed [9:0] m315_74;
   assign m315_74 =10'b0;

   // m315_75 = W*in
   wire signed [9:0] m315_75;
   assign m315_75 =10'b0;

   // m315_76 = W*in
   wire signed [9:0] m315_76;
   assign m315_76 =10'b0;

   // m315_77 = W*in
   wire signed [9:0] m315_77;
   assign m315_77 ={ {4{neg315[5]}} , neg315[5:0] };

   // m315_78 = W*in
   wire signed [9:0] m315_78;
   assign m315_78 =10'b0;

   // m315_79 = W*in
   wire signed [9:0] m315_79;
   assign m315_79 =10'b0;

   // m315_80 = W*in
   wire signed [9:0] m315_80;
   assign m315_80 =10'b0;

   // m315_81 = W*in
   wire signed [9:0] m315_81;
   assign m315_81 =10'b0;

   // m315_82 = W*in
   wire signed [9:0] m315_82;
   assign m315_82 =10'b0;

   // m315_83 = W*in
   wire signed [9:0] m315_83;
   assign m315_83 =10'b0;

   // m315_84 = W*in
   wire signed [9:0] m315_84;
   assign m315_84 =10'b0;

   // m315_85 = W*in
   wire signed [9:0] m315_85;
   assign m315_85 ={ {4{in315[5]}} , in315[5:0] };

   // m315_86 = W*in
   wire signed [9:0] m315_86;
   assign m315_86 =10'b0;

   // m315_87 = W*in
   wire signed [9:0] m315_87;
   assign m315_87 =10'b0;

   // m315_88 = W*in
   wire signed [9:0] m315_88;
   assign m315_88 =10'b0;

   // m315_89 = W*in
   wire signed [9:0] m315_89;
   assign m315_89 ={ {4{in315[5]}} , in315[5:0] };

   // m315_90 = W*in
   wire signed [9:0] m315_90;
   assign m315_90 =10'b0;

   // m315_91 = W*in
   wire signed [9:0] m315_91;
   assign m315_91 =10'b0;

   // m315_92 = W*in
   wire signed [9:0] m315_92;
   assign m315_92 =10'b0;

   // m315_93 = W*in
   wire signed [9:0] m315_93;
   assign m315_93 =10'b0;

   // m315_94 = W*in
   wire signed [9:0] m315_94;
   assign m315_94 =10'b0;

   // m315_95 = W*in
   wire signed [9:0] m315_95;
   assign m315_95 =10'b0;

   // m315_96 = W*in
   wire signed [9:0] m315_96;
   assign m315_96 =10'b0;

   // m315_97 = W*in
   wire signed [9:0] m315_97;
   assign m315_97 ={ {4{neg315[5]}} , neg315[5:0] };

   // m315_98 = W*in
   wire signed [9:0] m315_98;
   assign m315_98 =10'b0;

   // m315_99 = W*in
   wire signed [9:0] m315_99;
   assign m315_99 =10'b0;

   // m315_100 = W*in
   wire signed [9:0] m315_100;
   assign m315_100 =10'b0;

   // m315_101 = W*in
   wire signed [9:0] m315_101;
   assign m315_101 =10'b0;

   // m315_102 = W*in
   wire signed [9:0] m315_102;
   assign m315_102 =10'b0;

   // m315_103 = W*in
   wire signed [9:0] m315_103;
   assign m315_103 =10'b0;

   // m315_104 = W*in
   wire signed [9:0] m315_104;
   assign m315_104 =10'b0;

   // m315_105 = W*in
   wire signed [9:0] m315_105;
   assign m315_105 =10'b0;

   // m315_106 = W*in
   wire signed [9:0] m315_106;
   assign m315_106 =10'b0;

   // m315_107 = W*in
   wire signed [9:0] m315_107;
   assign m315_107 =10'b0;

   // m315_108 = W*in
   wire signed [9:0] m315_108;
   assign m315_108 ={ {4{in315[5]}} , in315[5:0] };

   // m315_109 = W*in
   wire signed [9:0] m315_109;
   assign m315_109 =10'b0;

   // m315_110 = W*in
   wire signed [9:0] m315_110;
   assign m315_110 =10'b0;

   // m315_111 = W*in
   wire signed [9:0] m315_111;
   assign m315_111 =10'b0;

   // m315_112 = W*in
   wire signed [9:0] m315_112;
   assign m315_112 =10'b0;

   // m315_113 = W*in
   wire signed [9:0] m315_113;
   assign m315_113 =10'b0;

   // m315_114 = W*in
   wire signed [9:0] m315_114;
   assign m315_114 =10'b0;

   // m315_115 = W*in
   wire signed [9:0] m315_115;
   assign m315_115 =10'b0;

   // m315_116 = W*in
   wire signed [9:0] m315_116;
   assign m315_116 =10'b0;

   // m315_117 = W*in
   wire signed [9:0] m315_117;
   assign m315_117 =10'b0;

   // m316_1 = W*in
   wire signed [9:0] m316_1;
   assign m316_1 =10'b0;

   // m316_2 = W*in
   wire signed [9:0] m316_2;
   assign m316_2 =10'b0;

   // m316_3 = W*in
   wire signed [9:0] m316_3;
   assign m316_3 =10'b0;

   // m316_4 = W*in
   wire signed [9:0] m316_4;
   assign m316_4 ={ {4{in316[5]}} , in316[5:0] };

   // m316_5 = W*in
   wire signed [9:0] m316_5;
   assign m316_5 =10'b0;

   // m316_6 = W*in
   wire signed [9:0] m316_6;
   assign m316_6 =10'b0;

   // m316_7 = W*in
   wire signed [9:0] m316_7;
   assign m316_7 =10'b0;

   // m316_8 = W*in
   wire signed [9:0] m316_8;
   assign m316_8 =10'b0;

   // m316_9 = W*in
   wire signed [9:0] m316_9;
   assign m316_9 =10'b0;

   // m316_10 = W*in
   wire signed [9:0] m316_10;
   assign m316_10 =10'b0;

   // m316_11 = W*in
   wire signed [9:0] m316_11;
   assign m316_11 =10'b0;

   // m316_12 = W*in
   wire signed [9:0] m316_12;
   assign m316_12 =10'b0;

   // m316_13 = W*in
   wire signed [9:0] m316_13;
   assign m316_13 =10'b0;

   // m316_14 = W*in
   wire signed [9:0] m316_14;
   assign m316_14 ={ {4{neg316[5]}} , neg316[5:0] };

   // m316_15 = W*in
   wire signed [9:0] m316_15;
   assign m316_15 =10'b0;

   // m316_16 = W*in
   wire signed [9:0] m316_16;
   assign m316_16 ={ {5{in316[5]}} , in316[5:1] };

   // m316_17 = W*in
   wire signed [9:0] m316_17;
   assign m316_17 =10'b0;

   // m316_18 = W*in
   wire signed [9:0] m316_18;
   assign m316_18 ={ {5{neg316[5]}} , neg316[5:1] };

   // m316_19 = W*in
   wire signed [9:0] m316_19;
   assign m316_19 ={ {5{neg316[5]}} , neg316[5:1] };

   // m316_20 = W*in
   wire signed [9:0] m316_20;
   assign m316_20 ={ {4{in316[5]}} , in316[5:0] };

   // m316_21 = W*in
   wire signed [9:0] m316_21;
   assign m316_21 ={ {5{neg316[5]}} , neg316[5:1] };

   // m316_22 = W*in
   wire signed [9:0] m316_22;
   assign m316_22 =10'b0;

   // m316_23 = W*in
   wire signed [9:0] m316_23;
   assign m316_23 =10'b0;

   // m316_24 = W*in
   wire signed [9:0] m316_24;
   assign m316_24 =10'b0;

   // m316_25 = W*in
   wire signed [9:0] m316_25;
   assign m316_25 =10'b0;

   // m316_26 = W*in
   wire signed [9:0] m316_26;
   assign m316_26 =10'b0;

   // m316_27 = W*in
   wire signed [9:0] m316_27;
   assign m316_27 =10'b0;

   // m316_28 = W*in
   wire signed [9:0] m316_28;
   assign m316_28 =10'b0;

   // m316_29 = W*in
   wire signed [9:0] m316_29;
   assign m316_29 =10'b0;

   // m316_30 = W*in
   wire signed [9:0] m316_30;
   assign m316_30 ={ {4{in316[5]}} , in316[5:0] };

   // m316_31 = W*in
   wire signed [9:0] m316_31;
   assign m316_31 =10'b0;

   // m316_32 = W*in
   wire signed [9:0] m316_32;
   assign m316_32 =10'b0;

   // m316_33 = W*in
   wire signed [9:0] m316_33;
   assign m316_33 =10'b0;

   // m316_34 = W*in
   wire signed [9:0] m316_34;
   assign m316_34 ={ {5{neg316[5]}} , neg316[5:1] };

   // m316_35 = W*in
   wire signed [9:0] m316_35;
   assign m316_35 ={ {5{in316[5]}} , in316[5:1] };

   // m316_36 = W*in
   wire signed [9:0] m316_36;
   assign m316_36 =10'b0;

   // m316_37 = W*in
   wire signed [9:0] m316_37;
   assign m316_37 =10'b0;

   // m316_38 = W*in
   wire signed [9:0] m316_38;
   assign m316_38 =10'b0;

   // m316_39 = W*in
   wire signed [9:0] m316_39;
   assign m316_39 =10'b0;

   // m316_40 = W*in
   wire signed [9:0] m316_40;
   assign m316_40 =10'b0;

   // m316_41 = W*in
   wire signed [9:0] m316_41;
   assign m316_41 =10'b0;

   // m316_42 = W*in
   wire signed [9:0] m316_42;
   assign m316_42 =10'b0;

   // m316_43 = W*in
   wire signed [9:0] m316_43;
   assign m316_43 =10'b0;

   // m316_44 = W*in
   wire signed [9:0] m316_44;
   assign m316_44 =10'b0;

   // m316_45 = W*in
   wire signed [9:0] m316_45;
   assign m316_45 =10'b0;

   // m316_46 = W*in
   wire signed [9:0] m316_46;
   assign m316_46 =10'b0;

   // m316_47 = W*in
   wire signed [9:0] m316_47;
   assign m316_47 =10'b0;

   // m316_48 = W*in
   wire signed [9:0] m316_48;
   assign m316_48 =10'b0;

   // m316_49 = W*in
   wire signed [9:0] m316_49;
   assign m316_49 =10'b0;

   // m316_50 = W*in
   wire signed [9:0] m316_50;
   assign m316_50 =10'b0;

   // m316_51 = W*in
   wire signed [9:0] m316_51;
   assign m316_51 =10'b0;

   // m316_52 = W*in
   wire signed [9:0] m316_52;
   assign m316_52 =10'b0;

   // m316_53 = W*in
   wire signed [9:0] m316_53;
   assign m316_53 =10'b0;

   // m316_54 = W*in
   wire signed [9:0] m316_54;
   assign m316_54 =10'b0;

   // m316_55 = W*in
   wire signed [9:0] m316_55;
   assign m316_55 =10'b0;

   // m316_56 = W*in
   wire signed [9:0] m316_56;
   assign m316_56 ={ {4{in316[5]}} , in316[5:0] };

   // m316_57 = W*in
   wire signed [9:0] m316_57;
   assign m316_57 =10'b0;

   // m316_58 = W*in
   wire signed [9:0] m316_58;
   assign m316_58 =10'b0;

   // m316_59 = W*in
   wire signed [9:0] m316_59;
   assign m316_59 =10'b0;

   // m316_60 = W*in
   wire signed [9:0] m316_60;
   assign m316_60 =10'b0;

   // m316_61 = W*in
   wire signed [9:0] m316_61;
   assign m316_61 =10'b0;

   // m316_62 = W*in
   wire signed [9:0] m316_62;
   assign m316_62 =10'b0;

   // m316_63 = W*in
   wire signed [9:0] m316_63;
   assign m316_63 =10'b0;

   // m316_64 = W*in
   wire signed [9:0] m316_64;
   assign m316_64 =10'b0;

   // m316_65 = W*in
   wire signed [9:0] m316_65;
   assign m316_65 =10'b0;

   // m316_66 = W*in
   wire signed [9:0] m316_66;
   assign m316_66 =10'b0;

   // m316_67 = W*in
   wire signed [9:0] m316_67;
   assign m316_67 =10'b0;

   // m316_68 = W*in
   wire signed [9:0] m316_68;
   assign m316_68 =10'b0;

   // m316_69 = W*in
   wire signed [9:0] m316_69;
   assign m316_69 =10'b0;

   // m316_70 = W*in
   wire signed [9:0] m316_70;
   assign m316_70 ={ {4{neg316[5]}} , neg316[5:0] };

   // m316_71 = W*in
   wire signed [9:0] m316_71;
   assign m316_71 =10'b0;

   // m316_72 = W*in
   wire signed [9:0] m316_72;
   assign m316_72 ={ {5{neg316[5]}} , neg316[5:1] };

   // m316_73 = W*in
   wire signed [9:0] m316_73;
   assign m316_73 =10'b0;

   // m316_74 = W*in
   wire signed [9:0] m316_74;
   assign m316_74 =10'b0;

   // m316_75 = W*in
   wire signed [9:0] m316_75;
   assign m316_75 ={ {4{in316[5]}} , in316[5:0] };

   // m316_76 = W*in
   wire signed [9:0] m316_76;
   assign m316_76 =10'b0;

   // m316_77 = W*in
   wire signed [9:0] m316_77;
   assign m316_77 =10'b0;

   // m316_78 = W*in
   wire signed [9:0] m316_78;
   assign m316_78 =10'b0;

   // m316_79 = W*in
   wire signed [9:0] m316_79;
   assign m316_79 =10'b0;

   // m316_80 = W*in
   wire signed [9:0] m316_80;
   assign m316_80 =10'b0;

   // m316_81 = W*in
   wire signed [9:0] m316_81;
   assign m316_81 =10'b0;

   // m316_82 = W*in
   wire signed [9:0] m316_82;
   assign m316_82 =10'b0;

   // m316_83 = W*in
   wire signed [9:0] m316_83;
   assign m316_83 ={ {4{in316[5]}} , in316[5:0] };

   // m316_84 = W*in
   wire signed [9:0] m316_84;
   assign m316_84 ={ {5{neg316[5]}} , neg316[5:1] };

   // m316_85 = W*in
   wire signed [9:0] m316_85;
   assign m316_85 =10'b0;

   // m316_86 = W*in
   wire signed [9:0] m316_86;
   assign m316_86 =10'b0;

   // m316_87 = W*in
   wire signed [9:0] m316_87;
   assign m316_87 =10'b0;

   // m316_88 = W*in
   wire signed [9:0] m316_88;
   assign m316_88 =10'b0;

   // m316_89 = W*in
   wire signed [9:0] m316_89;
   assign m316_89 =10'b0;

   // m316_90 = W*in
   wire signed [9:0] m316_90;
   assign m316_90 =10'b0;

   // m316_91 = W*in
   wire signed [9:0] m316_91;
   assign m316_91 =10'b0;

   // m316_92 = W*in
   wire signed [9:0] m316_92;
   assign m316_92 =10'b0;

   // m316_93 = W*in
   wire signed [9:0] m316_93;
   assign m316_93 =10'b0;

   // m316_94 = W*in
   wire signed [9:0] m316_94;
   assign m316_94 =10'b0;

   // m316_95 = W*in
   wire signed [9:0] m316_95;
   assign m316_95 =10'b0;

   // m316_96 = W*in
   wire signed [9:0] m316_96;
   assign m316_96 =10'b0;

   // m316_97 = W*in
   wire signed [9:0] m316_97;
   assign m316_97 =10'b0;

   // m316_98 = W*in
   wire signed [9:0] m316_98;
   assign m316_98 =10'b0;

   // m316_99 = W*in
   wire signed [9:0] m316_99;
   assign m316_99 =10'b0;

   // m316_100 = W*in
   wire signed [9:0] m316_100;
   assign m316_100 =10'b0;

   // m316_101 = W*in
   wire signed [9:0] m316_101;
   assign m316_101 =10'b0;

   // m316_102 = W*in
   wire signed [9:0] m316_102;
   assign m316_102 =10'b0;

   // m316_103 = W*in
   wire signed [9:0] m316_103;
   assign m316_103 =10'b0;

   // m316_104 = W*in
   wire signed [9:0] m316_104;
   assign m316_104 =10'b0;

   // m316_105 = W*in
   wire signed [9:0] m316_105;
   assign m316_105 =10'b0;

   // m316_106 = W*in
   wire signed [9:0] m316_106;
   assign m316_106 =10'b0;

   // m316_107 = W*in
   wire signed [9:0] m316_107;
   assign m316_107 =10'b0;

   // m316_108 = W*in
   wire signed [9:0] m316_108;
   assign m316_108 ={ {5{in316[5]}} , in316[5:1] };

   // m316_109 = W*in
   wire signed [9:0] m316_109;
   assign m316_109 ={ {5{in316[5]}} , in316[5:1] };

   // m316_110 = W*in
   wire signed [9:0] m316_110;
   assign m316_110 ={ {4{neg316[5]}} , neg316[5:0] };

   // m316_111 = W*in
   wire signed [9:0] m316_111;
   assign m316_111 =10'b0;

   // m316_112 = W*in
   wire signed [9:0] m316_112;
   assign m316_112 =10'b0;

   // m316_113 = W*in
   wire signed [9:0] m316_113;
   assign m316_113 ={ {4{in316[5]}} , in316[5:0] };

   // m316_114 = W*in
   wire signed [9:0] m316_114;
   assign m316_114 =10'b0;

   // m316_115 = W*in
   wire signed [9:0] m316_115;
   assign m316_115 ={ {4{in316[5]}} , in316[5:0] };

   // m316_116 = W*in
   wire signed [9:0] m316_116;
   assign m316_116 =10'b0;

   // m316_117 = W*in
   wire signed [9:0] m316_117;
   assign m316_117 =10'b0;

   // m317_1 = W*in
   wire signed [9:0] m317_1;
   assign m317_1 =10'b0;

   // m317_2 = W*in
   wire signed [9:0] m317_2;
   assign m317_2 =10'b0;

   // m317_3 = W*in
   wire signed [9:0] m317_3;
   assign m317_3 =10'b0;

   // m317_4 = W*in
   wire signed [9:0] m317_4;
   assign m317_4 =10'b0;

   // m317_5 = W*in
   wire signed [9:0] m317_5;
   assign m317_5 =10'b0;

   // m317_6 = W*in
   wire signed [9:0] m317_6;
   assign m317_6 =10'b0;

   // m317_7 = W*in
   wire signed [9:0] m317_7;
   assign m317_7 =10'b0;

   // m317_8 = W*in
   wire signed [9:0] m317_8;
   assign m317_8 =10'b0;

   // m317_9 = W*in
   wire signed [9:0] m317_9;
   assign m317_9 =10'b0;

   // m317_10 = W*in
   wire signed [9:0] m317_10;
   assign m317_10 =10'b0;

   // m317_11 = W*in
   wire signed [9:0] m317_11;
   assign m317_11 =10'b0;

   // m317_12 = W*in
   wire signed [9:0] m317_12;
   assign m317_12 =10'b0;

   // m317_13 = W*in
   wire signed [9:0] m317_13;
   assign m317_13 =10'b0;

   // m317_14 = W*in
   wire signed [9:0] m317_14;
   assign m317_14 =10'b0;

   // m317_15 = W*in
   wire signed [9:0] m317_15;
   assign m317_15 =10'b0;

   // m317_16 = W*in
   wire signed [9:0] m317_16;
   assign m317_16 ={ {5{in317[5]}} , in317[5:1] };

   // m317_17 = W*in
   wire signed [9:0] m317_17;
   assign m317_17 =10'b0;

   // m317_18 = W*in
   wire signed [9:0] m317_18;
   assign m317_18 =10'b0;

   // m317_19 = W*in
   wire signed [9:0] m317_19;
   assign m317_19 =10'b0;

   // m317_20 = W*in
   wire signed [9:0] m317_20;
   assign m317_20 =10'b0;

   // m317_21 = W*in
   wire signed [9:0] m317_21;
   assign m317_21 ={ {5{neg317[5]}} , neg317[5:1] };

   // m317_22 = W*in
   wire signed [9:0] m317_22;
   assign m317_22 =10'b0;

   // m317_23 = W*in
   wire signed [9:0] m317_23;
   assign m317_23 =10'b0;

   // m317_24 = W*in
   wire signed [9:0] m317_24;
   assign m317_24 =10'b0;

   // m317_25 = W*in
   wire signed [9:0] m317_25;
   assign m317_25 =10'b0;

   // m317_26 = W*in
   wire signed [9:0] m317_26;
   assign m317_26 =10'b0;

   // m317_27 = W*in
   wire signed [9:0] m317_27;
   assign m317_27 =10'b0;

   // m317_28 = W*in
   wire signed [9:0] m317_28;
   assign m317_28 =10'b0;

   // m317_29 = W*in
   wire signed [9:0] m317_29;
   assign m317_29 =10'b0;

   // m317_30 = W*in
   wire signed [9:0] m317_30;
   assign m317_30 ={ {4{in317[5]}} , in317[5:0] };

   // m317_31 = W*in
   wire signed [9:0] m317_31;
   assign m317_31 =10'b0;

   // m317_32 = W*in
   wire signed [9:0] m317_32;
   assign m317_32 =10'b0;

   // m317_33 = W*in
   wire signed [9:0] m317_33;
   assign m317_33 =10'b0;

   // m317_34 = W*in
   wire signed [9:0] m317_34;
   assign m317_34 =10'b0;

   // m317_35 = W*in
   wire signed [9:0] m317_35;
   assign m317_35 =10'b0;

   // m317_36 = W*in
   wire signed [9:0] m317_36;
   assign m317_36 =10'b0;

   // m317_37 = W*in
   wire signed [9:0] m317_37;
   assign m317_37 =10'b0;

   // m317_38 = W*in
   wire signed [9:0] m317_38;
   assign m317_38 =10'b0;

   // m317_39 = W*in
   wire signed [9:0] m317_39;
   assign m317_39 =10'b0;

   // m317_40 = W*in
   wire signed [9:0] m317_40;
   assign m317_40 =10'b0;

   // m317_41 = W*in
   wire signed [9:0] m317_41;
   assign m317_41 =10'b0;

   // m317_42 = W*in
   wire signed [9:0] m317_42;
   assign m317_42 =10'b0;

   // m317_43 = W*in
   wire signed [9:0] m317_43;
   assign m317_43 =10'b0;

   // m317_44 = W*in
   wire signed [9:0] m317_44;
   assign m317_44 =10'b0;

   // m317_45 = W*in
   wire signed [9:0] m317_45;
   assign m317_45 =10'b0;

   // m317_46 = W*in
   wire signed [9:0] m317_46;
   assign m317_46 =10'b0;

   // m317_47 = W*in
   wire signed [9:0] m317_47;
   assign m317_47 =10'b0;

   // m317_48 = W*in
   wire signed [9:0] m317_48;
   assign m317_48 =10'b0;

   // m317_49 = W*in
   wire signed [9:0] m317_49;
   assign m317_49 =10'b0;

   // m317_50 = W*in
   wire signed [9:0] m317_50;
   assign m317_50 =10'b0;

   // m317_51 = W*in
   wire signed [9:0] m317_51;
   assign m317_51 =10'b0;

   // m317_52 = W*in
   wire signed [9:0] m317_52;
   assign m317_52 =10'b0;

   // m317_53 = W*in
   wire signed [9:0] m317_53;
   assign m317_53 =10'b0;

   // m317_54 = W*in
   wire signed [9:0] m317_54;
   assign m317_54 =10'b0;

   // m317_55 = W*in
   wire signed [9:0] m317_55;
   assign m317_55 =10'b0;

   // m317_56 = W*in
   wire signed [9:0] m317_56;
   assign m317_56 =10'b0;

   // m317_57 = W*in
   wire signed [9:0] m317_57;
   assign m317_57 =10'b0;

   // m317_58 = W*in
   wire signed [9:0] m317_58;
   assign m317_58 =10'b0;

   // m317_59 = W*in
   wire signed [9:0] m317_59;
   assign m317_59 =10'b0;

   // m317_60 = W*in
   wire signed [9:0] m317_60;
   assign m317_60 =10'b0;

   // m317_61 = W*in
   wire signed [9:0] m317_61;
   assign m317_61 =10'b0;

   // m317_62 = W*in
   wire signed [9:0] m317_62;
   assign m317_62 =10'b0;

   // m317_63 = W*in
   wire signed [9:0] m317_63;
   assign m317_63 =10'b0;

   // m317_64 = W*in
   wire signed [9:0] m317_64;
   assign m317_64 =10'b0;

   // m317_65 = W*in
   wire signed [9:0] m317_65;
   assign m317_65 =10'b0;

   // m317_66 = W*in
   wire signed [9:0] m317_66;
   assign m317_66 =10'b0;

   // m317_67 = W*in
   wire signed [9:0] m317_67;
   assign m317_67 =10'b0;

   // m317_68 = W*in
   wire signed [9:0] m317_68;
   assign m317_68 =10'b0;

   // m317_69 = W*in
   wire signed [9:0] m317_69;
   assign m317_69 =10'b0;

   // m317_70 = W*in
   wire signed [9:0] m317_70;
   assign m317_70 =10'b0;

   // m317_71 = W*in
   wire signed [9:0] m317_71;
   assign m317_71 =10'b0;

   // m317_72 = W*in
   wire signed [9:0] m317_72;
   assign m317_72 =10'b0;

   // m317_73 = W*in
   wire signed [9:0] m317_73;
   assign m317_73 =10'b0;

   // m317_74 = W*in
   wire signed [9:0] m317_74;
   assign m317_74 =10'b0;

   // m317_75 = W*in
   wire signed [9:0] m317_75;
   assign m317_75 ={ {4{in317[5]}} , in317[5:0] };

   // m317_76 = W*in
   wire signed [9:0] m317_76;
   assign m317_76 =10'b0;

   // m317_77 = W*in
   wire signed [9:0] m317_77;
   assign m317_77 =10'b0;

   // m317_78 = W*in
   wire signed [9:0] m317_78;
   assign m317_78 =10'b0;

   // m317_79 = W*in
   wire signed [9:0] m317_79;
   assign m317_79 =10'b0;

   // m317_80 = W*in
   wire signed [9:0] m317_80;
   assign m317_80 =10'b0;

   // m317_81 = W*in
   wire signed [9:0] m317_81;
   assign m317_81 ={ {5{in317[5]}} , in317[5:1] };

   // m317_82 = W*in
   wire signed [9:0] m317_82;
   assign m317_82 =10'b0;

   // m317_83 = W*in
   wire signed [9:0] m317_83;
   assign m317_83 =10'b0;

   // m317_84 = W*in
   wire signed [9:0] m317_84;
   assign m317_84 =10'b0;

   // m317_85 = W*in
   wire signed [9:0] m317_85;
   assign m317_85 =10'b0;

   // m317_86 = W*in
   wire signed [9:0] m317_86;
   assign m317_86 ={ {4{neg317[5]}} , neg317[5:0] };

   // m317_87 = W*in
   wire signed [9:0] m317_87;
   assign m317_87 =10'b0;

   // m317_88 = W*in
   wire signed [9:0] m317_88;
   assign m317_88 =10'b0;

   // m317_89 = W*in
   wire signed [9:0] m317_89;
   assign m317_89 =10'b0;

   // m317_90 = W*in
   wire signed [9:0] m317_90;
   assign m317_90 =10'b0;

   // m317_91 = W*in
   wire signed [9:0] m317_91;
   assign m317_91 =10'b0;

   // m317_92 = W*in
   wire signed [9:0] m317_92;
   assign m317_92 =10'b0;

   // m317_93 = W*in
   wire signed [9:0] m317_93;
   assign m317_93 =10'b0;

   // m317_94 = W*in
   wire signed [9:0] m317_94;
   assign m317_94 =10'b0;

   // m317_95 = W*in
   wire signed [9:0] m317_95;
   assign m317_95 =10'b0;

   // m317_96 = W*in
   wire signed [9:0] m317_96;
   assign m317_96 =10'b0;

   // m317_97 = W*in
   wire signed [9:0] m317_97;
   assign m317_97 =10'b0;

   // m317_98 = W*in
   wire signed [9:0] m317_98;
   assign m317_98 =10'b0;

   // m317_99 = W*in
   wire signed [9:0] m317_99;
   assign m317_99 =10'b0;

   // m317_100 = W*in
   wire signed [9:0] m317_100;
   assign m317_100 =10'b0;

   // m317_101 = W*in
   wire signed [9:0] m317_101;
   assign m317_101 =10'b0;

   // m317_102 = W*in
   wire signed [9:0] m317_102;
   assign m317_102 =10'b0;

   // m317_103 = W*in
   wire signed [9:0] m317_103;
   assign m317_103 =10'b0;

   // m317_104 = W*in
   wire signed [9:0] m317_104;
   assign m317_104 =10'b0;

   // m317_105 = W*in
   wire signed [9:0] m317_105;
   assign m317_105 =10'b0;

   // m317_106 = W*in
   wire signed [9:0] m317_106;
   assign m317_106 =10'b0;

   // m317_107 = W*in
   wire signed [9:0] m317_107;
   assign m317_107 =10'b0;

   // m317_108 = W*in
   wire signed [9:0] m317_108;
   assign m317_108 ={ {4{in317[5]}} , in317[5:0] };

   // m317_109 = W*in
   wire signed [9:0] m317_109;
   assign m317_109 ={ {5{in317[5]}} , in317[5:1] };

   // m317_110 = W*in
   wire signed [9:0] m317_110;
   assign m317_110 =10'b0;

   // m317_111 = W*in
   wire signed [9:0] m317_111;
   assign m317_111 =10'b0;

   // m317_112 = W*in
   wire signed [9:0] m317_112;
   assign m317_112 =10'b0;

   // m317_113 = W*in
   wire signed [9:0] m317_113;
   assign m317_113 =10'b0;

   // m317_114 = W*in
   wire signed [9:0] m317_114;
   assign m317_114 ={ {5{neg317[5]}} , neg317[5:1] };

   // m317_115 = W*in
   wire signed [9:0] m317_115;
   assign m317_115 =10'b0;

   // m317_116 = W*in
   wire signed [9:0] m317_116;
   assign m317_116 =10'b0;

   // m317_117 = W*in
   wire signed [9:0] m317_117;
   assign m317_117 =10'b0;

   // m318_1 = W*in
   wire signed [9:0] m318_1;
   assign m318_1 =10'b0;

   // m318_2 = W*in
   wire signed [9:0] m318_2;
   assign m318_2 =10'b0;

   // m318_3 = W*in
   wire signed [9:0] m318_3;
   assign m318_3 =10'b0;

   // m318_4 = W*in
   wire signed [9:0] m318_4;
   assign m318_4 =10'b0;

   // m318_5 = W*in
   wire signed [9:0] m318_5;
   assign m318_5 =10'b0;

   // m318_6 = W*in
   wire signed [9:0] m318_6;
   assign m318_6 =10'b0;

   // m318_7 = W*in
   wire signed [9:0] m318_7;
   assign m318_7 =10'b0;

   // m318_8 = W*in
   wire signed [9:0] m318_8;
   assign m318_8 =10'b0;

   // m318_9 = W*in
   wire signed [9:0] m318_9;
   assign m318_9 =10'b0;

   // m318_10 = W*in
   wire signed [9:0] m318_10;
   assign m318_10 =10'b0;

   // m318_11 = W*in
   wire signed [9:0] m318_11;
   assign m318_11 =10'b0;

   // m318_12 = W*in
   wire signed [9:0] m318_12;
   assign m318_12 =10'b0;

   // m318_13 = W*in
   wire signed [9:0] m318_13;
   assign m318_13 =10'b0;

   // m318_14 = W*in
   wire signed [9:0] m318_14;
   assign m318_14 =10'b0;

   // m318_15 = W*in
   wire signed [9:0] m318_15;
   assign m318_15 =10'b0;

   // m318_16 = W*in
   wire signed [9:0] m318_16;
   assign m318_16 =10'b0;

   // m318_17 = W*in
   wire signed [9:0] m318_17;
   assign m318_17 =10'b0;

   // m318_18 = W*in
   wire signed [9:0] m318_18;
   assign m318_18 =10'b0;

   // m318_19 = W*in
   wire signed [9:0] m318_19;
   assign m318_19 =10'b0;

   // m318_20 = W*in
   wire signed [9:0] m318_20;
   assign m318_20 =10'b0;

   // m318_21 = W*in
   wire signed [9:0] m318_21;
   assign m318_21 =10'b0;

   // m318_22 = W*in
   wire signed [9:0] m318_22;
   assign m318_22 =10'b0;

   // m318_23 = W*in
   wire signed [9:0] m318_23;
   assign m318_23 =10'b0;

   // m318_24 = W*in
   wire signed [9:0] m318_24;
   assign m318_24 =10'b0;

   // m318_25 = W*in
   wire signed [9:0] m318_25;
   assign m318_25 =10'b0;

   // m318_26 = W*in
   wire signed [9:0] m318_26;
   assign m318_26 =10'b0;

   // m318_27 = W*in
   wire signed [9:0] m318_27;
   assign m318_27 =10'b0;

   // m318_28 = W*in
   wire signed [9:0] m318_28;
   assign m318_28 =10'b0;

   // m318_29 = W*in
   wire signed [9:0] m318_29;
   assign m318_29 =10'b0;

   // m318_30 = W*in
   wire signed [9:0] m318_30;
   assign m318_30 =10'b0;

   // m318_31 = W*in
   wire signed [9:0] m318_31;
   assign m318_31 =10'b0;

   // m318_32 = W*in
   wire signed [9:0] m318_32;
   assign m318_32 =10'b0;

   // m318_33 = W*in
   wire signed [9:0] m318_33;
   assign m318_33 =10'b0;

   // m318_34 = W*in
   wire signed [9:0] m318_34;
   assign m318_34 =10'b0;

   // m318_35 = W*in
   wire signed [9:0] m318_35;
   assign m318_35 =10'b0;

   // m318_36 = W*in
   wire signed [9:0] m318_36;
   assign m318_36 =10'b0;

   // m318_37 = W*in
   wire signed [9:0] m318_37;
   assign m318_37 =10'b0;

   // m318_38 = W*in
   wire signed [9:0] m318_38;
   assign m318_38 =10'b0;

   // m318_39 = W*in
   wire signed [9:0] m318_39;
   assign m318_39 =10'b0;

   // m318_40 = W*in
   wire signed [9:0] m318_40;
   assign m318_40 =10'b0;

   // m318_41 = W*in
   wire signed [9:0] m318_41;
   assign m318_41 =10'b0;

   // m318_42 = W*in
   wire signed [9:0] m318_42;
   assign m318_42 =10'b0;

   // m318_43 = W*in
   wire signed [9:0] m318_43;
   assign m318_43 =10'b0;

   // m318_44 = W*in
   wire signed [9:0] m318_44;
   assign m318_44 =10'b0;

   // m318_45 = W*in
   wire signed [9:0] m318_45;
   assign m318_45 =10'b0;

   // m318_46 = W*in
   wire signed [9:0] m318_46;
   assign m318_46 =10'b0;

   // m318_47 = W*in
   wire signed [9:0] m318_47;
   assign m318_47 =10'b0;

   // m318_48 = W*in
   wire signed [9:0] m318_48;
   assign m318_48 =10'b0;

   // m318_49 = W*in
   wire signed [9:0] m318_49;
   assign m318_49 =10'b0;

   // m318_50 = W*in
   wire signed [9:0] m318_50;
   assign m318_50 =10'b0;

   // m318_51 = W*in
   wire signed [9:0] m318_51;
   assign m318_51 =10'b0;

   // m318_52 = W*in
   wire signed [9:0] m318_52;
   assign m318_52 =10'b0;

   // m318_53 = W*in
   wire signed [9:0] m318_53;
   assign m318_53 =10'b0;

   // m318_54 = W*in
   wire signed [9:0] m318_54;
   assign m318_54 =10'b0;

   // m318_55 = W*in
   wire signed [9:0] m318_55;
   assign m318_55 =10'b0;

   // m318_56 = W*in
   wire signed [9:0] m318_56;
   assign m318_56 =10'b0;

   // m318_57 = W*in
   wire signed [9:0] m318_57;
   assign m318_57 =10'b0;

   // m318_58 = W*in
   wire signed [9:0] m318_58;
   assign m318_58 =10'b0;

   // m318_59 = W*in
   wire signed [9:0] m318_59;
   assign m318_59 =10'b0;

   // m318_60 = W*in
   wire signed [9:0] m318_60;
   assign m318_60 =10'b0;

   // m318_61 = W*in
   wire signed [9:0] m318_61;
   assign m318_61 =10'b0;

   // m318_62 = W*in
   wire signed [9:0] m318_62;
   assign m318_62 =10'b0;

   // m318_63 = W*in
   wire signed [9:0] m318_63;
   assign m318_63 =10'b0;

   // m318_64 = W*in
   wire signed [9:0] m318_64;
   assign m318_64 =10'b0;

   // m318_65 = W*in
   wire signed [9:0] m318_65;
   assign m318_65 =10'b0;

   // m318_66 = W*in
   wire signed [9:0] m318_66;
   assign m318_66 =10'b0;

   // m318_67 = W*in
   wire signed [9:0] m318_67;
   assign m318_67 =10'b0;

   // m318_68 = W*in
   wire signed [9:0] m318_68;
   assign m318_68 =10'b0;

   // m318_69 = W*in
   wire signed [9:0] m318_69;
   assign m318_69 =10'b0;

   // m318_70 = W*in
   wire signed [9:0] m318_70;
   assign m318_70 =10'b0;

   // m318_71 = W*in
   wire signed [9:0] m318_71;
   assign m318_71 =10'b0;

   // m318_72 = W*in
   wire signed [9:0] m318_72;
   assign m318_72 =10'b0;

   // m318_73 = W*in
   wire signed [9:0] m318_73;
   assign m318_73 =10'b0;

   // m318_74 = W*in
   wire signed [9:0] m318_74;
   assign m318_74 =10'b0;

   // m318_75 = W*in
   wire signed [9:0] m318_75;
   assign m318_75 =10'b0;

   // m318_76 = W*in
   wire signed [9:0] m318_76;
   assign m318_76 =10'b0;

   // m318_77 = W*in
   wire signed [9:0] m318_77;
   assign m318_77 =10'b0;

   // m318_78 = W*in
   wire signed [9:0] m318_78;
   assign m318_78 =10'b0;

   // m318_79 = W*in
   wire signed [9:0] m318_79;
   assign m318_79 =10'b0;

   // m318_80 = W*in
   wire signed [9:0] m318_80;
   assign m318_80 =10'b0;

   // m318_81 = W*in
   wire signed [9:0] m318_81;
   assign m318_81 =10'b0;

   // m318_82 = W*in
   wire signed [9:0] m318_82;
   assign m318_82 =10'b0;

   // m318_83 = W*in
   wire signed [9:0] m318_83;
   assign m318_83 ={ {5{in318[5]}} , in318[5:1] };

   // m318_84 = W*in
   wire signed [9:0] m318_84;
   assign m318_84 ={ {5{neg318[5]}} , neg318[5:1] };

   // m318_85 = W*in
   wire signed [9:0] m318_85;
   assign m318_85 =10'b0;

   // m318_86 = W*in
   wire signed [9:0] m318_86;
   assign m318_86 =10'b0;

   // m318_87 = W*in
   wire signed [9:0] m318_87;
   assign m318_87 =10'b0;

   // m318_88 = W*in
   wire signed [9:0] m318_88;
   assign m318_88 =10'b0;

   // m318_89 = W*in
   wire signed [9:0] m318_89;
   assign m318_89 =10'b0;

   // m318_90 = W*in
   wire signed [9:0] m318_90;
   assign m318_90 =10'b0;

   // m318_91 = W*in
   wire signed [9:0] m318_91;
   assign m318_91 =10'b0;

   // m318_92 = W*in
   wire signed [9:0] m318_92;
   assign m318_92 =10'b0;

   // m318_93 = W*in
   wire signed [9:0] m318_93;
   assign m318_93 =10'b0;

   // m318_94 = W*in
   wire signed [9:0] m318_94;
   assign m318_94 =10'b0;

   // m318_95 = W*in
   wire signed [9:0] m318_95;
   assign m318_95 =10'b0;

   // m318_96 = W*in
   wire signed [9:0] m318_96;
   assign m318_96 =10'b0;

   // m318_97 = W*in
   wire signed [9:0] m318_97;
   assign m318_97 =10'b0;

   // m318_98 = W*in
   wire signed [9:0] m318_98;
   assign m318_98 =10'b0;

   // m318_99 = W*in
   wire signed [9:0] m318_99;
   assign m318_99 =10'b0;

   // m318_100 = W*in
   wire signed [9:0] m318_100;
   assign m318_100 =10'b0;

   // m318_101 = W*in
   wire signed [9:0] m318_101;
   assign m318_101 =10'b0;

   // m318_102 = W*in
   wire signed [9:0] m318_102;
   assign m318_102 =10'b0;

   // m318_103 = W*in
   wire signed [9:0] m318_103;
   assign m318_103 =10'b0;

   // m318_104 = W*in
   wire signed [9:0] m318_104;
   assign m318_104 =10'b0;

   // m318_105 = W*in
   wire signed [9:0] m318_105;
   assign m318_105 =10'b0;

   // m318_106 = W*in
   wire signed [9:0] m318_106;
   assign m318_106 =10'b0;

   // m318_107 = W*in
   wire signed [9:0] m318_107;
   assign m318_107 =10'b0;

   // m318_108 = W*in
   wire signed [9:0] m318_108;
   assign m318_108 =10'b0;

   // m318_109 = W*in
   wire signed [9:0] m318_109;
   assign m318_109 =10'b0;

   // m318_110 = W*in
   wire signed [9:0] m318_110;
   assign m318_110 =10'b0;

   // m318_111 = W*in
   wire signed [9:0] m318_111;
   assign m318_111 =10'b0;

   // m318_112 = W*in
   wire signed [9:0] m318_112;
   assign m318_112 =10'b0;

   // m318_113 = W*in
   wire signed [9:0] m318_113;
   assign m318_113 =10'b0;

   // m318_114 = W*in
   wire signed [9:0] m318_114;
   assign m318_114 =10'b0;

   // m318_115 = W*in
   wire signed [9:0] m318_115;
   assign m318_115 =10'b0;

   // m318_116 = W*in
   wire signed [9:0] m318_116;
   assign m318_116 =10'b0;

   // m318_117 = W*in
   wire signed [9:0] m318_117;
   assign m318_117 =10'b0;

   // m319_1 = W*in
   wire signed [9:0] m319_1;
   assign m319_1 =10'b0;

   // m319_2 = W*in
   wire signed [9:0] m319_2;
   assign m319_2 =10'b0;

   // m319_3 = W*in
   wire signed [9:0] m319_3;
   assign m319_3 =10'b0;

   // m319_4 = W*in
   wire signed [9:0] m319_4;
   assign m319_4 =10'b0;

   // m319_5 = W*in
   wire signed [9:0] m319_5;
   assign m319_5 =10'b0;

   // m319_6 = W*in
   wire signed [9:0] m319_6;
   assign m319_6 =10'b0;

   // m319_7 = W*in
   wire signed [9:0] m319_7;
   assign m319_7 =10'b0;

   // m319_8 = W*in
   wire signed [9:0] m319_8;
   assign m319_8 =10'b0;

   // m319_9 = W*in
   wire signed [9:0] m319_9;
   assign m319_9 =10'b0;

   // m319_10 = W*in
   wire signed [9:0] m319_10;
   assign m319_10 ={ {4{neg319[5]}} , neg319[5:0] };

   // m319_11 = W*in
   wire signed [9:0] m319_11;
   assign m319_11 =10'b0;

   // m319_12 = W*in
   wire signed [9:0] m319_12;
   assign m319_12 =10'b0;

   // m319_13 = W*in
   wire signed [9:0] m319_13;
   assign m319_13 =10'b0;

   // m319_14 = W*in
   wire signed [9:0] m319_14;
   assign m319_14 =10'b0;

   // m319_15 = W*in
   wire signed [9:0] m319_15;
   assign m319_15 =10'b0;

   // m319_16 = W*in
   wire signed [9:0] m319_16;
   assign m319_16 =10'b0;

   // m319_17 = W*in
   wire signed [9:0] m319_17;
   assign m319_17 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_18 = W*in
   wire signed [9:0] m319_18;
   assign m319_18 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_19 = W*in
   wire signed [9:0] m319_19;
   assign m319_19 =10'b0;

   // m319_20 = W*in
   wire signed [9:0] m319_20;
   assign m319_20 ={ {5{in319[5]}} , in319[5:1] };

   // m319_21 = W*in
   wire signed [9:0] m319_21;
   assign m319_21 ={ {4{neg319[5]}} , neg319[5:0] };

   // m319_22 = W*in
   wire signed [9:0] m319_22;
   assign m319_22 =10'b0;

   // m319_23 = W*in
   wire signed [9:0] m319_23;
   assign m319_23 =10'b0;

   // m319_24 = W*in
   wire signed [9:0] m319_24;
   assign m319_24 =10'b0;

   // m319_25 = W*in
   wire signed [9:0] m319_25;
   assign m319_25 =10'b0;

   // m319_26 = W*in
   wire signed [9:0] m319_26;
   assign m319_26 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_27 = W*in
   wire signed [9:0] m319_27;
   assign m319_27 =10'b0;

   // m319_28 = W*in
   wire signed [9:0] m319_28;
   assign m319_28 =10'b0;

   // m319_29 = W*in
   wire signed [9:0] m319_29;
   assign m319_29 =10'b0;

   // m319_30 = W*in
   wire signed [9:0] m319_30;
   assign m319_30 =10'b0;

   // m319_31 = W*in
   wire signed [9:0] m319_31;
   assign m319_31 =10'b0;

   // m319_32 = W*in
   wire signed [9:0] m319_32;
   assign m319_32 =10'b0;

   // m319_33 = W*in
   wire signed [9:0] m319_33;
   assign m319_33 =10'b0;

   // m319_34 = W*in
   wire signed [9:0] m319_34;
   assign m319_34 =10'b0;

   // m319_35 = W*in
   wire signed [9:0] m319_35;
   assign m319_35 ={ {5{in319[5]}} , in319[5:1] };

   // m319_36 = W*in
   wire signed [9:0] m319_36;
   assign m319_36 =10'b0;

   // m319_37 = W*in
   wire signed [9:0] m319_37;
   assign m319_37 =10'b0;

   // m319_38 = W*in
   wire signed [9:0] m319_38;
   assign m319_38 =10'b0;

   // m319_39 = W*in
   wire signed [9:0] m319_39;
   assign m319_39 =10'b0;

   // m319_40 = W*in
   wire signed [9:0] m319_40;
   assign m319_40 =10'b0;

   // m319_41 = W*in
   wire signed [9:0] m319_41;
   assign m319_41 =10'b0;

   // m319_42 = W*in
   wire signed [9:0] m319_42;
   assign m319_42 =10'b0;

   // m319_43 = W*in
   wire signed [9:0] m319_43;
   assign m319_43 =10'b0;

   // m319_44 = W*in
   wire signed [9:0] m319_44;
   assign m319_44 =10'b0;

   // m319_45 = W*in
   wire signed [9:0] m319_45;
   assign m319_45 =10'b0;

   // m319_46 = W*in
   wire signed [9:0] m319_46;
   assign m319_46 =10'b0;

   // m319_47 = W*in
   wire signed [9:0] m319_47;
   assign m319_47 =10'b0;

   // m319_48 = W*in
   wire signed [9:0] m319_48;
   assign m319_48 =10'b0;

   // m319_49 = W*in
   wire signed [9:0] m319_49;
   assign m319_49 =10'b0;

   // m319_50 = W*in
   wire signed [9:0] m319_50;
   assign m319_50 =10'b0;

   // m319_51 = W*in
   wire signed [9:0] m319_51;
   assign m319_51 =10'b0;

   // m319_52 = W*in
   wire signed [9:0] m319_52;
   assign m319_52 =10'b0;

   // m319_53 = W*in
   wire signed [9:0] m319_53;
   assign m319_53 =10'b0;

   // m319_54 = W*in
   wire signed [9:0] m319_54;
   assign m319_54 =10'b0;

   // m319_55 = W*in
   wire signed [9:0] m319_55;
   assign m319_55 =10'b0;

   // m319_56 = W*in
   wire signed [9:0] m319_56;
   assign m319_56 =10'b0;

   // m319_57 = W*in
   wire signed [9:0] m319_57;
   assign m319_57 =10'b0;

   // m319_58 = W*in
   wire signed [9:0] m319_58;
   assign m319_58 =10'b0;

   // m319_59 = W*in
   wire signed [9:0] m319_59;
   assign m319_59 =10'b0;

   // m319_60 = W*in
   wire signed [9:0] m319_60;
   assign m319_60 =10'b0;

   // m319_61 = W*in
   wire signed [9:0] m319_61;
   assign m319_61 ={ {4{in319[5]}} , in319[5:0] };

   // m319_62 = W*in
   wire signed [9:0] m319_62;
   assign m319_62 =10'b0;

   // m319_63 = W*in
   wire signed [9:0] m319_63;
   assign m319_63 =10'b0;

   // m319_64 = W*in
   wire signed [9:0] m319_64;
   assign m319_64 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_65 = W*in
   wire signed [9:0] m319_65;
   assign m319_65 =10'b0;

   // m319_66 = W*in
   wire signed [9:0] m319_66;
   assign m319_66 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_67 = W*in
   wire signed [9:0] m319_67;
   assign m319_67 =10'b0;

   // m319_68 = W*in
   wire signed [9:0] m319_68;
   assign m319_68 =10'b0;

   // m319_69 = W*in
   wire signed [9:0] m319_69;
   assign m319_69 =10'b0;

   // m319_70 = W*in
   wire signed [9:0] m319_70;
   assign m319_70 ={ {4{neg319[5]}} , neg319[5:0] };

   // m319_71 = W*in
   wire signed [9:0] m319_71;
   assign m319_71 =10'b0;

   // m319_72 = W*in
   wire signed [9:0] m319_72;
   assign m319_72 =10'b0;

   // m319_73 = W*in
   wire signed [9:0] m319_73;
   assign m319_73 ={ {5{in319[5]}} , in319[5:1] };

   // m319_74 = W*in
   wire signed [9:0] m319_74;
   assign m319_74 =10'b0;

   // m319_75 = W*in
   wire signed [9:0] m319_75;
   assign m319_75 =10'b0;

   // m319_76 = W*in
   wire signed [9:0] m319_76;
   assign m319_76 =10'b0;

   // m319_77 = W*in
   wire signed [9:0] m319_77;
   assign m319_77 =10'b0;

   // m319_78 = W*in
   wire signed [9:0] m319_78;
   assign m319_78 =10'b0;

   // m319_79 = W*in
   wire signed [9:0] m319_79;
   assign m319_79 =10'b0;

   // m319_80 = W*in
   wire signed [9:0] m319_80;
   assign m319_80 ={ {4{in319[5]}} , in319[5:0] };

   // m319_81 = W*in
   wire signed [9:0] m319_81;
   assign m319_81 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_82 = W*in
   wire signed [9:0] m319_82;
   assign m319_82 =10'b0;

   // m319_83 = W*in
   wire signed [9:0] m319_83;
   assign m319_83 =10'b0;

   // m319_84 = W*in
   wire signed [9:0] m319_84;
   assign m319_84 ={ {5{neg319[5]}} , neg319[5:1] };

   // m319_85 = W*in
   wire signed [9:0] m319_85;
   assign m319_85 =10'b0;

   // m319_86 = W*in
   wire signed [9:0] m319_86;
   assign m319_86 =10'b0;

   // m319_87 = W*in
   wire signed [9:0] m319_87;
   assign m319_87 =10'b0;

   // m319_88 = W*in
   wire signed [9:0] m319_88;
   assign m319_88 =10'b0;

   // m319_89 = W*in
   wire signed [9:0] m319_89;
   assign m319_89 =10'b0;

   // m319_90 = W*in
   wire signed [9:0] m319_90;
   assign m319_90 =10'b0;

   // m319_91 = W*in
   wire signed [9:0] m319_91;
   assign m319_91 =10'b0;

   // m319_92 = W*in
   wire signed [9:0] m319_92;
   assign m319_92 =10'b0;

   // m319_93 = W*in
   wire signed [9:0] m319_93;
   assign m319_93 =10'b0;

   // m319_94 = W*in
   wire signed [9:0] m319_94;
   assign m319_94 ={ {4{neg319[5]}} , neg319[5:0] };

   // m319_95 = W*in
   wire signed [9:0] m319_95;
   assign m319_95 =10'b0;

   // m319_96 = W*in
   wire signed [9:0] m319_96;
   assign m319_96 =10'b0;

   // m319_97 = W*in
   wire signed [9:0] m319_97;
   assign m319_97 =10'b0;

   // m319_98 = W*in
   wire signed [9:0] m319_98;
   assign m319_98 =10'b0;

   // m319_99 = W*in
   wire signed [9:0] m319_99;
   assign m319_99 =10'b0;

   // m319_100 = W*in
   wire signed [9:0] m319_100;
   assign m319_100 =10'b0;

   // m319_101 = W*in
   wire signed [9:0] m319_101;
   assign m319_101 =10'b0;

   // m319_102 = W*in
   wire signed [9:0] m319_102;
   assign m319_102 =10'b0;

   // m319_103 = W*in
   wire signed [9:0] m319_103;
   assign m319_103 =10'b0;

   // m319_104 = W*in
   wire signed [9:0] m319_104;
   assign m319_104 =10'b0;

   // m319_105 = W*in
   wire signed [9:0] m319_105;
   assign m319_105 ={ {4{in319[5]}} , in319[5:0] };

   // m319_106 = W*in
   wire signed [9:0] m319_106;
   assign m319_106 =10'b0;

   // m319_107 = W*in
   wire signed [9:0] m319_107;
   assign m319_107 =10'b0;

   // m319_108 = W*in
   wire signed [9:0] m319_108;
   assign m319_108 ={ {5{in319[5]}} , in319[5:1] };

   // m319_109 = W*in
   wire signed [9:0] m319_109;
   assign m319_109 =10'b0;

   // m319_110 = W*in
   wire signed [9:0] m319_110;
   assign m319_110 =10'b0;

   // m319_111 = W*in
   wire signed [9:0] m319_111;
   assign m319_111 =10'b0;

   // m319_112 = W*in
   wire signed [9:0] m319_112;
   assign m319_112 =10'b0;

   // m319_113 = W*in
   wire signed [9:0] m319_113;
   assign m319_113 =10'b0;

   // m319_114 = W*in
   wire signed [9:0] m319_114;
   assign m319_114 =10'b0;

   // m319_115 = W*in
   wire signed [9:0] m319_115;
   assign m319_115 =10'b0;

   // m319_116 = W*in
   wire signed [9:0] m319_116;
   assign m319_116 =10'b0;

   // m319_117 = W*in
   wire signed [9:0] m319_117;
   assign m319_117 =10'b0;

   // m320_1 = W*in
   wire signed [9:0] m320_1;
   assign m320_1 =10'b0;

   // m320_2 = W*in
   wire signed [9:0] m320_2;
   assign m320_2 =10'b0;

   // m320_3 = W*in
   wire signed [9:0] m320_3;
   assign m320_3 ={ {4{in320[5]}} , in320[5:0] };

   // m320_4 = W*in
   wire signed [9:0] m320_4;
   assign m320_4 =10'b0;

   // m320_5 = W*in
   wire signed [9:0] m320_5;
   assign m320_5 =10'b0;

   // m320_6 = W*in
   wire signed [9:0] m320_6;
   assign m320_6 =10'b0;

   // m320_7 = W*in
   wire signed [9:0] m320_7;
   assign m320_7 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_8 = W*in
   wire signed [9:0] m320_8;
   assign m320_8 ={ {4{in320[5]}} , in320[5:0] };

   // m320_9 = W*in
   wire signed [9:0] m320_9;
   assign m320_9 =10'b0;

   // m320_10 = W*in
   wire signed [9:0] m320_10;
   assign m320_10 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_11 = W*in
   wire signed [9:0] m320_11;
   assign m320_11 =10'b0;

   // m320_12 = W*in
   wire signed [9:0] m320_12;
   assign m320_12 ={ {4{in320[5]}} , in320[5:0] };

   // m320_13 = W*in
   wire signed [9:0] m320_13;
   assign m320_13 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_14 = W*in
   wire signed [9:0] m320_14;
   assign m320_14 =10'b0;

   // m320_15 = W*in
   wire signed [9:0] m320_15;
   assign m320_15 ={ {4{in320[5]}} , in320[5:0] };

   // m320_16 = W*in
   wire signed [9:0] m320_16;
   assign m320_16 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_17 = W*in
   wire signed [9:0] m320_17;
   assign m320_17 ={ {5{in320[5]}} , in320[5:1] };

   // m320_18 = W*in
   wire signed [9:0] m320_18;
   assign m320_18 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_19 = W*in
   wire signed [9:0] m320_19;
   assign m320_19 =10'b0;

   // m320_20 = W*in
   wire signed [9:0] m320_20;
   assign m320_20 ={ {5{in320[5]}} , in320[5:1] };

   // m320_21 = W*in
   wire signed [9:0] m320_21;
   assign m320_21 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_22 = W*in
   wire signed [9:0] m320_22;
   assign m320_22 =10'b0;

   // m320_23 = W*in
   wire signed [9:0] m320_23;
   assign m320_23 =10'b0;

   // m320_24 = W*in
   wire signed [9:0] m320_24;
   assign m320_24 ={ {4{in320[5]}} , in320[5:0] };

   // m320_25 = W*in
   wire signed [9:0] m320_25;
   assign m320_25 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_26 = W*in
   wire signed [9:0] m320_26;
   assign m320_26 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_27 = W*in
   wire signed [9:0] m320_27;
   assign m320_27 ={ {4{in320[5]}} , in320[5:0] };

   // m320_28 = W*in
   wire signed [9:0] m320_28;
   assign m320_28 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_29 = W*in
   wire signed [9:0] m320_29;
   assign m320_29 =10'b0;

   // m320_30 = W*in
   wire signed [9:0] m320_30;
   assign m320_30 =10'b0;

   // m320_31 = W*in
   wire signed [9:0] m320_31;
   assign m320_31 ={ {4{in320[5]}} , in320[5:0] };

   // m320_32 = W*in
   wire signed [9:0] m320_32;
   assign m320_32 =10'b0;

   // m320_33 = W*in
   wire signed [9:0] m320_33;
   assign m320_33 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_34 = W*in
   wire signed [9:0] m320_34;
   assign m320_34 ={ {5{in320[5]}} , in320[5:1] };

   // m320_35 = W*in
   wire signed [9:0] m320_35;
   assign m320_35 =10'b0;

   // m320_36 = W*in
   wire signed [9:0] m320_36;
   assign m320_36 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_37 = W*in
   wire signed [9:0] m320_37;
   assign m320_37 =10'b0;

   // m320_38 = W*in
   wire signed [9:0] m320_38;
   assign m320_38 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_39 = W*in
   wire signed [9:0] m320_39;
   assign m320_39 ={ {4{in320[5]}} , in320[5:0] };

   // m320_40 = W*in
   wire signed [9:0] m320_40;
   assign m320_40 =10'b0;

   // m320_41 = W*in
   wire signed [9:0] m320_41;
   assign m320_41 =10'b0;

   // m320_42 = W*in
   wire signed [9:0] m320_42;
   assign m320_42 =10'b0;

   // m320_43 = W*in
   wire signed [9:0] m320_43;
   assign m320_43 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_44 = W*in
   wire signed [9:0] m320_44;
   assign m320_44 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_45 = W*in
   wire signed [9:0] m320_45;
   assign m320_45 =10'b0;

   // m320_46 = W*in
   wire signed [9:0] m320_46;
   assign m320_46 =10'b0;

   // m320_47 = W*in
   wire signed [9:0] m320_47;
   assign m320_47 =10'b0;

   // m320_48 = W*in
   wire signed [9:0] m320_48;
   assign m320_48 =10'b0;

   // m320_49 = W*in
   wire signed [9:0] m320_49;
   assign m320_49 =10'b0;

   // m320_50 = W*in
   wire signed [9:0] m320_50;
   assign m320_50 ={ {4{in320[5]}} , in320[5:0] };

   // m320_51 = W*in
   wire signed [9:0] m320_51;
   assign m320_51 =10'b0;

   // m320_52 = W*in
   wire signed [9:0] m320_52;
   assign m320_52 ={ {4{in320[5]}} , in320[5:0] };

   // m320_53 = W*in
   wire signed [9:0] m320_53;
   assign m320_53 =10'b0;

   // m320_54 = W*in
   wire signed [9:0] m320_54;
   assign m320_54 =10'b0;

   // m320_55 = W*in
   wire signed [9:0] m320_55;
   assign m320_55 =10'b0;

   // m320_56 = W*in
   wire signed [9:0] m320_56;
   assign m320_56 =10'b0;

   // m320_57 = W*in
   wire signed [9:0] m320_57;
   assign m320_57 =10'b0;

   // m320_58 = W*in
   wire signed [9:0] m320_58;
   assign m320_58 =10'b0;

   // m320_59 = W*in
   wire signed [9:0] m320_59;
   assign m320_59 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_60 = W*in
   wire signed [9:0] m320_60;
   assign m320_60 =10'b0;

   // m320_61 = W*in
   wire signed [9:0] m320_61;
   assign m320_61 =10'b0;

   // m320_62 = W*in
   wire signed [9:0] m320_62;
   assign m320_62 =10'b0;

   // m320_63 = W*in
   wire signed [9:0] m320_63;
   assign m320_63 =10'b0;

   // m320_64 = W*in
   wire signed [9:0] m320_64;
   assign m320_64 =10'b0;

   // m320_65 = W*in
   wire signed [9:0] m320_65;
   assign m320_65 ={ {5{in320[5]}} , in320[5:1] };

   // m320_66 = W*in
   wire signed [9:0] m320_66;
   assign m320_66 =10'b0;

   // m320_67 = W*in
   wire signed [9:0] m320_67;
   assign m320_67 =10'b0;

   // m320_68 = W*in
   wire signed [9:0] m320_68;
   assign m320_68 =10'b0;

   // m320_69 = W*in
   wire signed [9:0] m320_69;
   assign m320_69 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_70 = W*in
   wire signed [9:0] m320_70;
   assign m320_70 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_71 = W*in
   wire signed [9:0] m320_71;
   assign m320_71 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_72 = W*in
   wire signed [9:0] m320_72;
   assign m320_72 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_73 = W*in
   wire signed [9:0] m320_73;
   assign m320_73 ={ {4{in320[5]}} , in320[5:0] };

   // m320_74 = W*in
   wire signed [9:0] m320_74;
   assign m320_74 =10'b0;

   // m320_75 = W*in
   wire signed [9:0] m320_75;
   assign m320_75 =10'b0;

   // m320_76 = W*in
   wire signed [9:0] m320_76;
   assign m320_76 =10'b0;

   // m320_77 = W*in
   wire signed [9:0] m320_77;
   assign m320_77 =10'b0;

   // m320_78 = W*in
   wire signed [9:0] m320_78;
   assign m320_78 =10'b0;

   // m320_79 = W*in
   wire signed [9:0] m320_79;
   assign m320_79 =10'b0;

   // m320_80 = W*in
   wire signed [9:0] m320_80;
   assign m320_80 ={ {3{in320[5]}} , in320 , {1{1'b0}} };

   // m320_81 = W*in
   wire signed [9:0] m320_81;
   assign m320_81 =10'b0;

   // m320_82 = W*in
   wire signed [9:0] m320_82;
   assign m320_82 =10'b0;

   // m320_83 = W*in
   wire signed [9:0] m320_83;
   assign m320_83 =10'b0;

   // m320_84 = W*in
   wire signed [9:0] m320_84;
   assign m320_84 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_85 = W*in
   wire signed [9:0] m320_85;
   assign m320_85 ={ {5{neg320[5]}} , neg320[5:1] };

   // m320_86 = W*in
   wire signed [9:0] m320_86;
   assign m320_86 =10'b0;

   // m320_87 = W*in
   wire signed [9:0] m320_87;
   assign m320_87 =10'b0;

   // m320_88 = W*in
   wire signed [9:0] m320_88;
   assign m320_88 ={ {4{in320[5]}} , in320[5:0] };

   // m320_89 = W*in
   wire signed [9:0] m320_89;
   assign m320_89 =10'b0;

   // m320_90 = W*in
   wire signed [9:0] m320_90;
   assign m320_90 =10'b0;

   // m320_91 = W*in
   wire signed [9:0] m320_91;
   assign m320_91 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_92 = W*in
   wire signed [9:0] m320_92;
   assign m320_92 =10'b0;

   // m320_93 = W*in
   wire signed [9:0] m320_93;
   assign m320_93 =10'b0;

   // m320_94 = W*in
   wire signed [9:0] m320_94;
   assign m320_94 =10'b0;

   // m320_95 = W*in
   wire signed [9:0] m320_95;
   assign m320_95 =10'b0;

   // m320_96 = W*in
   wire signed [9:0] m320_96;
   assign m320_96 =10'b0;

   // m320_97 = W*in
   wire signed [9:0] m320_97;
   assign m320_97 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_98 = W*in
   wire signed [9:0] m320_98;
   assign m320_98 ={ {4{in320[5]}} , in320[5:0] };

   // m320_99 = W*in
   wire signed [9:0] m320_99;
   assign m320_99 =10'b0;

   // m320_100 = W*in
   wire signed [9:0] m320_100;
   assign m320_100 =10'b0;

   // m320_101 = W*in
   wire signed [9:0] m320_101;
   assign m320_101 =10'b0;

   // m320_102 = W*in
   wire signed [9:0] m320_102;
   assign m320_102 =10'b0;

   // m320_103 = W*in
   wire signed [9:0] m320_103;
   assign m320_103 =10'b0;

   // m320_104 = W*in
   wire signed [9:0] m320_104;
   assign m320_104 =10'b0;

   // m320_105 = W*in
   wire signed [9:0] m320_105;
   assign m320_105 ={ {3{in320[5]}} , in320 , {1{1'b0}} };

   // m320_106 = W*in
   wire signed [9:0] m320_106;
   assign m320_106 =10'b0;

   // m320_107 = W*in
   wire signed [9:0] m320_107;
   assign m320_107 ={ {4{in320[5]}} , in320[5:0] };

   // m320_108 = W*in
   wire signed [9:0] m320_108;
   assign m320_108 =10'b0;

   // m320_109 = W*in
   wire signed [9:0] m320_109;
   assign m320_109 =10'b0;

   // m320_110 = W*in
   wire signed [9:0] m320_110;
   assign m320_110 =10'b0;

   // m320_111 = W*in
   wire signed [9:0] m320_111;
   assign m320_111 ={ {4{neg320[5]}} , neg320[5:0] };

   // m320_112 = W*in
   wire signed [9:0] m320_112;
   assign m320_112 =10'b0;

   // m320_113 = W*in
   wire signed [9:0] m320_113;
   assign m320_113 =10'b0;

   // m320_114 = W*in
   wire signed [9:0] m320_114;
   assign m320_114 ={ {5{in320[5]}} , in320[5:1] };

   // m320_115 = W*in
   wire signed [9:0] m320_115;
   assign m320_115 =10'b0;

   // m320_116 = W*in
   wire signed [9:0] m320_116;
   assign m320_116 =10'b0;

   // m320_117 = W*in
   wire signed [9:0] m320_117;
   assign m320_117 =10'b0;

   // m321_1 = W*in
   wire signed [9:0] m321_1;
   assign m321_1 =10'b0;

   // m321_2 = W*in
   wire signed [9:0] m321_2;
   assign m321_2 =10'b0;

   // m321_3 = W*in
   wire signed [9:0] m321_3;
   assign m321_3 =10'b0;

   // m321_4 = W*in
   wire signed [9:0] m321_4;
   assign m321_4 ={ {4{in321[5]}} , in321[5:0] };

   // m321_5 = W*in
   wire signed [9:0] m321_5;
   assign m321_5 =10'b0;

   // m321_6 = W*in
   wire signed [9:0] m321_6;
   assign m321_6 =10'b0;

   // m321_7 = W*in
   wire signed [9:0] m321_7;
   assign m321_7 =10'b0;

   // m321_8 = W*in
   wire signed [9:0] m321_8;
   assign m321_8 =10'b0;

   // m321_9 = W*in
   wire signed [9:0] m321_9;
   assign m321_9 =10'b0;

   // m321_10 = W*in
   wire signed [9:0] m321_10;
   assign m321_10 =10'b0;

   // m321_11 = W*in
   wire signed [9:0] m321_11;
   assign m321_11 ={ {4{in321[5]}} , in321[5:0] };

   // m321_12 = W*in
   wire signed [9:0] m321_12;
   assign m321_12 =10'b0;

   // m321_13 = W*in
   wire signed [9:0] m321_13;
   assign m321_13 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_14 = W*in
   wire signed [9:0] m321_14;
   assign m321_14 =10'b0;

   // m321_15 = W*in
   wire signed [9:0] m321_15;
   assign m321_15 ={ {4{in321[5]}} , in321[5:0] };

   // m321_16 = W*in
   wire signed [9:0] m321_16;
   assign m321_16 =10'b0;

   // m321_17 = W*in
   wire signed [9:0] m321_17;
   assign m321_17 ={ {5{in321[5]}} , in321[5:1] };

   // m321_18 = W*in
   wire signed [9:0] m321_18;
   assign m321_18 =10'b0;

   // m321_19 = W*in
   wire signed [9:0] m321_19;
   assign m321_19 =10'b0;

   // m321_20 = W*in
   wire signed [9:0] m321_20;
   assign m321_20 =10'b0;

   // m321_21 = W*in
   wire signed [9:0] m321_21;
   assign m321_21 =10'b0;

   // m321_22 = W*in
   wire signed [9:0] m321_22;
   assign m321_22 =10'b0;

   // m321_23 = W*in
   wire signed [9:0] m321_23;
   assign m321_23 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_24 = W*in
   wire signed [9:0] m321_24;
   assign m321_24 =10'b0;

   // m321_25 = W*in
   wire signed [9:0] m321_25;
   assign m321_25 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_26 = W*in
   wire signed [9:0] m321_26;
   assign m321_26 ={ {5{neg321[5]}} , neg321[5:1] };

   // m321_27 = W*in
   wire signed [9:0] m321_27;
   assign m321_27 =10'b0;

   // m321_28 = W*in
   wire signed [9:0] m321_28;
   assign m321_28 ={ {5{neg321[5]}} , neg321[5:1] };

   // m321_29 = W*in
   wire signed [9:0] m321_29;
   assign m321_29 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_30 = W*in
   wire signed [9:0] m321_30;
   assign m321_30 =10'b0;

   // m321_31 = W*in
   wire signed [9:0] m321_31;
   assign m321_31 =10'b0;

   // m321_32 = W*in
   wire signed [9:0] m321_32;
   assign m321_32 =10'b0;

   // m321_33 = W*in
   wire signed [9:0] m321_33;
   assign m321_33 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_34 = W*in
   wire signed [9:0] m321_34;
   assign m321_34 =10'b0;

   // m321_35 = W*in
   wire signed [9:0] m321_35;
   assign m321_35 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_36 = W*in
   wire signed [9:0] m321_36;
   assign m321_36 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_37 = W*in
   wire signed [9:0] m321_37;
   assign m321_37 ={ {4{in321[5]}} , in321[5:0] };

   // m321_38 = W*in
   wire signed [9:0] m321_38;
   assign m321_38 =10'b0;

   // m321_39 = W*in
   wire signed [9:0] m321_39;
   assign m321_39 =10'b0;

   // m321_40 = W*in
   wire signed [9:0] m321_40;
   assign m321_40 =10'b0;

   // m321_41 = W*in
   wire signed [9:0] m321_41;
   assign m321_41 =10'b0;

   // m321_42 = W*in
   wire signed [9:0] m321_42;
   assign m321_42 =10'b0;

   // m321_43 = W*in
   wire signed [9:0] m321_43;
   assign m321_43 =10'b0;

   // m321_44 = W*in
   wire signed [9:0] m321_44;
   assign m321_44 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_45 = W*in
   wire signed [9:0] m321_45;
   assign m321_45 =10'b0;

   // m321_46 = W*in
   wire signed [9:0] m321_46;
   assign m321_46 =10'b0;

   // m321_47 = W*in
   wire signed [9:0] m321_47;
   assign m321_47 =10'b0;

   // m321_48 = W*in
   wire signed [9:0] m321_48;
   assign m321_48 =10'b0;

   // m321_49 = W*in
   wire signed [9:0] m321_49;
   assign m321_49 =10'b0;

   // m321_50 = W*in
   wire signed [9:0] m321_50;
   assign m321_50 ={ {4{in321[5]}} , in321[5:0] };

   // m321_51 = W*in
   wire signed [9:0] m321_51;
   assign m321_51 =10'b0;

   // m321_52 = W*in
   wire signed [9:0] m321_52;
   assign m321_52 ={ {4{in321[5]}} , in321[5:0] };

   // m321_53 = W*in
   wire signed [9:0] m321_53;
   assign m321_53 =10'b0;

   // m321_54 = W*in
   wire signed [9:0] m321_54;
   assign m321_54 =10'b0;

   // m321_55 = W*in
   wire signed [9:0] m321_55;
   assign m321_55 =10'b0;

   // m321_56 = W*in
   wire signed [9:0] m321_56;
   assign m321_56 =10'b0;

   // m321_57 = W*in
   wire signed [9:0] m321_57;
   assign m321_57 =10'b0;

   // m321_58 = W*in
   wire signed [9:0] m321_58;
   assign m321_58 =10'b0;

   // m321_59 = W*in
   wire signed [9:0] m321_59;
   assign m321_59 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_60 = W*in
   wire signed [9:0] m321_60;
   assign m321_60 =10'b0;

   // m321_61 = W*in
   wire signed [9:0] m321_61;
   assign m321_61 =10'b0;

   // m321_62 = W*in
   wire signed [9:0] m321_62;
   assign m321_62 ={ {4{in321[5]}} , in321[5:0] };

   // m321_63 = W*in
   wire signed [9:0] m321_63;
   assign m321_63 =10'b0;

   // m321_64 = W*in
   wire signed [9:0] m321_64;
   assign m321_64 =10'b0;

   // m321_65 = W*in
   wire signed [9:0] m321_65;
   assign m321_65 =10'b0;

   // m321_66 = W*in
   wire signed [9:0] m321_66;
   assign m321_66 ={ {5{neg321[5]}} , neg321[5:1] };

   // m321_67 = W*in
   wire signed [9:0] m321_67;
   assign m321_67 =10'b0;

   // m321_68 = W*in
   wire signed [9:0] m321_68;
   assign m321_68 =10'b0;

   // m321_69 = W*in
   wire signed [9:0] m321_69;
   assign m321_69 =10'b0;

   // m321_70 = W*in
   wire signed [9:0] m321_70;
   assign m321_70 =10'b0;

   // m321_71 = W*in
   wire signed [9:0] m321_71;
   assign m321_71 =10'b0;

   // m321_72 = W*in
   wire signed [9:0] m321_72;
   assign m321_72 =10'b0;

   // m321_73 = W*in
   wire signed [9:0] m321_73;
   assign m321_73 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_74 = W*in
   wire signed [9:0] m321_74;
   assign m321_74 =10'b0;

   // m321_75 = W*in
   wire signed [9:0] m321_75;
   assign m321_75 =10'b0;

   // m321_76 = W*in
   wire signed [9:0] m321_76;
   assign m321_76 ={ {4{in321[5]}} , in321[5:0] };

   // m321_77 = W*in
   wire signed [9:0] m321_77;
   assign m321_77 ={ {4{in321[5]}} , in321[5:0] };

   // m321_78 = W*in
   wire signed [9:0] m321_78;
   assign m321_78 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_79 = W*in
   wire signed [9:0] m321_79;
   assign m321_79 =10'b0;

   // m321_80 = W*in
   wire signed [9:0] m321_80;
   assign m321_80 =10'b0;

   // m321_81 = W*in
   wire signed [9:0] m321_81;
   assign m321_81 ={ {5{in321[5]}} , in321[5:1] };

   // m321_82 = W*in
   wire signed [9:0] m321_82;
   assign m321_82 =10'b0;

   // m321_83 = W*in
   wire signed [9:0] m321_83;
   assign m321_83 ={ {4{in321[5]}} , in321[5:0] };

   // m321_84 = W*in
   wire signed [9:0] m321_84;
   assign m321_84 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_85 = W*in
   wire signed [9:0] m321_85;
   assign m321_85 =10'b0;

   // m321_86 = W*in
   wire signed [9:0] m321_86;
   assign m321_86 =10'b0;

   // m321_87 = W*in
   wire signed [9:0] m321_87;
   assign m321_87 ={ {4{in321[5]}} , in321[5:0] };

   // m321_88 = W*in
   wire signed [9:0] m321_88;
   assign m321_88 =10'b0;

   // m321_89 = W*in
   wire signed [9:0] m321_89;
   assign m321_89 =10'b0;

   // m321_90 = W*in
   wire signed [9:0] m321_90;
   assign m321_90 =10'b0;

   // m321_91 = W*in
   wire signed [9:0] m321_91;
   assign m321_91 =10'b0;

   // m321_92 = W*in
   wire signed [9:0] m321_92;
   assign m321_92 ={ {4{in321[5]}} , in321[5:0] };

   // m321_93 = W*in
   wire signed [9:0] m321_93;
   assign m321_93 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_94 = W*in
   wire signed [9:0] m321_94;
   assign m321_94 =10'b0;

   // m321_95 = W*in
   wire signed [9:0] m321_95;
   assign m321_95 =10'b0;

   // m321_96 = W*in
   wire signed [9:0] m321_96;
   assign m321_96 =10'b0;

   // m321_97 = W*in
   wire signed [9:0] m321_97;
   assign m321_97 =10'b0;

   // m321_98 = W*in
   wire signed [9:0] m321_98;
   assign m321_98 ={ {4{in321[5]}} , in321[5:0] };

   // m321_99 = W*in
   wire signed [9:0] m321_99;
   assign m321_99 =10'b0;

   // m321_100 = W*in
   wire signed [9:0] m321_100;
   assign m321_100 =10'b0;

   // m321_101 = W*in
   wire signed [9:0] m321_101;
   assign m321_101 =10'b0;

   // m321_102 = W*in
   wire signed [9:0] m321_102;
   assign m321_102 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_103 = W*in
   wire signed [9:0] m321_103;
   assign m321_103 =10'b0;

   // m321_104 = W*in
   wire signed [9:0] m321_104;
   assign m321_104 =10'b0;

   // m321_105 = W*in
   wire signed [9:0] m321_105;
   assign m321_105 =10'b0;

   // m321_106 = W*in
   wire signed [9:0] m321_106;
   assign m321_106 =10'b0;

   // m321_107 = W*in
   wire signed [9:0] m321_107;
   assign m321_107 =10'b0;

   // m321_108 = W*in
   wire signed [9:0] m321_108;
   assign m321_108 ={ {5{neg321[5]}} , neg321[5:1] };

   // m321_109 = W*in
   wire signed [9:0] m321_109;
   assign m321_109 ={ {5{neg321[5]}} , neg321[5:1] };

   // m321_110 = W*in
   wire signed [9:0] m321_110;
   assign m321_110 =10'b0;

   // m321_111 = W*in
   wire signed [9:0] m321_111;
   assign m321_111 ={ {4{neg321[5]}} , neg321[5:0] };

   // m321_112 = W*in
   wire signed [9:0] m321_112;
   assign m321_112 =10'b0;

   // m321_113 = W*in
   wire signed [9:0] m321_113;
   assign m321_113 =10'b0;

   // m321_114 = W*in
   wire signed [9:0] m321_114;
   assign m321_114 =10'b0;

   // m321_115 = W*in
   wire signed [9:0] m321_115;
   assign m321_115 =10'b0;

   // m321_116 = W*in
   wire signed [9:0] m321_116;
   assign m321_116 =10'b0;

   // m321_117 = W*in
   wire signed [9:0] m321_117;
   assign m321_117 ={ {4{neg321[5]}} , neg321[5:0] };

   // m322_1 = W*in
   wire signed [9:0] m322_1;
   assign m322_1 =10'b0;

   // m322_2 = W*in
   wire signed [9:0] m322_2;
   assign m322_2 =10'b0;

   // m322_3 = W*in
   wire signed [9:0] m322_3;
   assign m322_3 ={ {4{in322[5]}} , in322[5:0] };

   // m322_4 = W*in
   wire signed [9:0] m322_4;
   assign m322_4 =10'b0;

   // m322_5 = W*in
   wire signed [9:0] m322_5;
   assign m322_5 =10'b0;

   // m322_6 = W*in
   wire signed [9:0] m322_6;
   assign m322_6 =10'b0;

   // m322_7 = W*in
   wire signed [9:0] m322_7;
   assign m322_7 =10'b0;

   // m322_8 = W*in
   wire signed [9:0] m322_8;
   assign m322_8 =10'b0;

   // m322_9 = W*in
   wire signed [9:0] m322_9;
   assign m322_9 =10'b0;

   // m322_10 = W*in
   wire signed [9:0] m322_10;
   assign m322_10 =10'b0;

   // m322_11 = W*in
   wire signed [9:0] m322_11;
   assign m322_11 =10'b0;

   // m322_12 = W*in
   wire signed [9:0] m322_12;
   assign m322_12 =10'b0;

   // m322_13 = W*in
   wire signed [9:0] m322_13;
   assign m322_13 =10'b0;

   // m322_14 = W*in
   wire signed [9:0] m322_14;
   assign m322_14 =10'b0;

   // m322_15 = W*in
   wire signed [9:0] m322_15;
   assign m322_15 =10'b0;

   // m322_16 = W*in
   wire signed [9:0] m322_16;
   assign m322_16 =10'b0;

   // m322_17 = W*in
   wire signed [9:0] m322_17;
   assign m322_17 ={ {5{in322[5]}} , in322[5:1] };

   // m322_18 = W*in
   wire signed [9:0] m322_18;
   assign m322_18 =10'b0;

   // m322_19 = W*in
   wire signed [9:0] m322_19;
   assign m322_19 =10'b0;

   // m322_20 = W*in
   wire signed [9:0] m322_20;
   assign m322_20 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_21 = W*in
   wire signed [9:0] m322_21;
   assign m322_21 =10'b0;

   // m322_22 = W*in
   wire signed [9:0] m322_22;
   assign m322_22 =10'b0;

   // m322_23 = W*in
   wire signed [9:0] m322_23;
   assign m322_23 =10'b0;

   // m322_24 = W*in
   wire signed [9:0] m322_24;
   assign m322_24 =10'b0;

   // m322_25 = W*in
   wire signed [9:0] m322_25;
   assign m322_25 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_26 = W*in
   wire signed [9:0] m322_26;
   assign m322_26 =10'b0;

   // m322_27 = W*in
   wire signed [9:0] m322_27;
   assign m322_27 ={ {5{in322[5]}} , in322[5:1] };

   // m322_28 = W*in
   wire signed [9:0] m322_28;
   assign m322_28 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_29 = W*in
   wire signed [9:0] m322_29;
   assign m322_29 =10'b0;

   // m322_30 = W*in
   wire signed [9:0] m322_30;
   assign m322_30 =10'b0;

   // m322_31 = W*in
   wire signed [9:0] m322_31;
   assign m322_31 =10'b0;

   // m322_32 = W*in
   wire signed [9:0] m322_32;
   assign m322_32 =10'b0;

   // m322_33 = W*in
   wire signed [9:0] m322_33;
   assign m322_33 =10'b0;

   // m322_34 = W*in
   wire signed [9:0] m322_34;
   assign m322_34 =10'b0;

   // m322_35 = W*in
   wire signed [9:0] m322_35;
   assign m322_35 ={ {5{neg322[5]}} , neg322[5:1] };

   // m322_36 = W*in
   wire signed [9:0] m322_36;
   assign m322_36 =10'b0;

   // m322_37 = W*in
   wire signed [9:0] m322_37;
   assign m322_37 =10'b0;

   // m322_38 = W*in
   wire signed [9:0] m322_38;
   assign m322_38 =10'b0;

   // m322_39 = W*in
   wire signed [9:0] m322_39;
   assign m322_39 =10'b0;

   // m322_40 = W*in
   wire signed [9:0] m322_40;
   assign m322_40 =10'b0;

   // m322_41 = W*in
   wire signed [9:0] m322_41;
   assign m322_41 =10'b0;

   // m322_42 = W*in
   wire signed [9:0] m322_42;
   assign m322_42 =10'b0;

   // m322_43 = W*in
   wire signed [9:0] m322_43;
   assign m322_43 =10'b0;

   // m322_44 = W*in
   wire signed [9:0] m322_44;
   assign m322_44 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_45 = W*in
   wire signed [9:0] m322_45;
   assign m322_45 =10'b0;

   // m322_46 = W*in
   wire signed [9:0] m322_46;
   assign m322_46 =10'b0;

   // m322_47 = W*in
   wire signed [9:0] m322_47;
   assign m322_47 =10'b0;

   // m322_48 = W*in
   wire signed [9:0] m322_48;
   assign m322_48 =10'b0;

   // m322_49 = W*in
   wire signed [9:0] m322_49;
   assign m322_49 =10'b0;

   // m322_50 = W*in
   wire signed [9:0] m322_50;
   assign m322_50 =10'b0;

   // m322_51 = W*in
   wire signed [9:0] m322_51;
   assign m322_51 =10'b0;

   // m322_52 = W*in
   wire signed [9:0] m322_52;
   assign m322_52 ={ {4{in322[5]}} , in322[5:0] };

   // m322_53 = W*in
   wire signed [9:0] m322_53;
   assign m322_53 =10'b0;

   // m322_54 = W*in
   wire signed [9:0] m322_54;
   assign m322_54 =10'b0;

   // m322_55 = W*in
   wire signed [9:0] m322_55;
   assign m322_55 =10'b0;

   // m322_56 = W*in
   wire signed [9:0] m322_56;
   assign m322_56 =10'b0;

   // m322_57 = W*in
   wire signed [9:0] m322_57;
   assign m322_57 =10'b0;

   // m322_58 = W*in
   wire signed [9:0] m322_58;
   assign m322_58 =10'b0;

   // m322_59 = W*in
   wire signed [9:0] m322_59;
   assign m322_59 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_60 = W*in
   wire signed [9:0] m322_60;
   assign m322_60 =10'b0;

   // m322_61 = W*in
   wire signed [9:0] m322_61;
   assign m322_61 =10'b0;

   // m322_62 = W*in
   wire signed [9:0] m322_62;
   assign m322_62 =10'b0;

   // m322_63 = W*in
   wire signed [9:0] m322_63;
   assign m322_63 =10'b0;

   // m322_64 = W*in
   wire signed [9:0] m322_64;
   assign m322_64 ={ {5{neg322[5]}} , neg322[5:1] };

   // m322_65 = W*in
   wire signed [9:0] m322_65;
   assign m322_65 ={ {5{neg322[5]}} , neg322[5:1] };

   // m322_66 = W*in
   wire signed [9:0] m322_66;
   assign m322_66 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_67 = W*in
   wire signed [9:0] m322_67;
   assign m322_67 =10'b0;

   // m322_68 = W*in
   wire signed [9:0] m322_68;
   assign m322_68 =10'b0;

   // m322_69 = W*in
   wire signed [9:0] m322_69;
   assign m322_69 =10'b0;

   // m322_70 = W*in
   wire signed [9:0] m322_70;
   assign m322_70 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_71 = W*in
   wire signed [9:0] m322_71;
   assign m322_71 ={ {4{in322[5]}} , in322[5:0] };

   // m322_72 = W*in
   wire signed [9:0] m322_72;
   assign m322_72 ={ {5{in322[5]}} , in322[5:1] };

   // m322_73 = W*in
   wire signed [9:0] m322_73;
   assign m322_73 ={ {5{neg322[5]}} , neg322[5:1] };

   // m322_74 = W*in
   wire signed [9:0] m322_74;
   assign m322_74 =10'b0;

   // m322_75 = W*in
   wire signed [9:0] m322_75;
   assign m322_75 =10'b0;

   // m322_76 = W*in
   wire signed [9:0] m322_76;
   assign m322_76 =10'b0;

   // m322_77 = W*in
   wire signed [9:0] m322_77;
   assign m322_77 =10'b0;

   // m322_78 = W*in
   wire signed [9:0] m322_78;
   assign m322_78 =10'b0;

   // m322_79 = W*in
   wire signed [9:0] m322_79;
   assign m322_79 =10'b0;

   // m322_80 = W*in
   wire signed [9:0] m322_80;
   assign m322_80 ={ {4{in322[5]}} , in322[5:0] };

   // m322_81 = W*in
   wire signed [9:0] m322_81;
   assign m322_81 =10'b0;

   // m322_82 = W*in
   wire signed [9:0] m322_82;
   assign m322_82 =10'b0;

   // m322_83 = W*in
   wire signed [9:0] m322_83;
   assign m322_83 ={ {5{in322[5]}} , in322[5:1] };

   // m322_84 = W*in
   wire signed [9:0] m322_84;
   assign m322_84 =10'b0;

   // m322_85 = W*in
   wire signed [9:0] m322_85;
   assign m322_85 =10'b0;

   // m322_86 = W*in
   wire signed [9:0] m322_86;
   assign m322_86 =10'b0;

   // m322_87 = W*in
   wire signed [9:0] m322_87;
   assign m322_87 =10'b0;

   // m322_88 = W*in
   wire signed [9:0] m322_88;
   assign m322_88 =10'b0;

   // m322_89 = W*in
   wire signed [9:0] m322_89;
   assign m322_89 =10'b0;

   // m322_90 = W*in
   wire signed [9:0] m322_90;
   assign m322_90 =10'b0;

   // m322_91 = W*in
   wire signed [9:0] m322_91;
   assign m322_91 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_92 = W*in
   wire signed [9:0] m322_92;
   assign m322_92 =10'b0;

   // m322_93 = W*in
   wire signed [9:0] m322_93;
   assign m322_93 =10'b0;

   // m322_94 = W*in
   wire signed [9:0] m322_94;
   assign m322_94 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_95 = W*in
   wire signed [9:0] m322_95;
   assign m322_95 =10'b0;

   // m322_96 = W*in
   wire signed [9:0] m322_96;
   assign m322_96 =10'b0;

   // m322_97 = W*in
   wire signed [9:0] m322_97;
   assign m322_97 =10'b0;

   // m322_98 = W*in
   wire signed [9:0] m322_98;
   assign m322_98 ={ {4{in322[5]}} , in322[5:0] };

   // m322_99 = W*in
   wire signed [9:0] m322_99;
   assign m322_99 =10'b0;

   // m322_100 = W*in
   wire signed [9:0] m322_100;
   assign m322_100 =10'b0;

   // m322_101 = W*in
   wire signed [9:0] m322_101;
   assign m322_101 =10'b0;

   // m322_102 = W*in
   wire signed [9:0] m322_102;
   assign m322_102 =10'b0;

   // m322_103 = W*in
   wire signed [9:0] m322_103;
   assign m322_103 =10'b0;

   // m322_104 = W*in
   wire signed [9:0] m322_104;
   assign m322_104 =10'b0;

   // m322_105 = W*in
   wire signed [9:0] m322_105;
   assign m322_105 ={ {4{in322[5]}} , in322[5:0] };

   // m322_106 = W*in
   wire signed [9:0] m322_106;
   assign m322_106 ={ {4{neg322[5]}} , neg322[5:0] };

   // m322_107 = W*in
   wire signed [9:0] m322_107;
   assign m322_107 ={ {4{in322[5]}} , in322[5:0] };

   // m322_108 = W*in
   wire signed [9:0] m322_108;
   assign m322_108 =10'b0;

   // m322_109 = W*in
   wire signed [9:0] m322_109;
   assign m322_109 =10'b0;

   // m322_110 = W*in
   wire signed [9:0] m322_110;
   assign m322_110 =10'b0;

   // m322_111 = W*in
   wire signed [9:0] m322_111;
   assign m322_111 =10'b0;

   // m322_112 = W*in
   wire signed [9:0] m322_112;
   assign m322_112 =10'b0;

   // m322_113 = W*in
   wire signed [9:0] m322_113;
   assign m322_113 =10'b0;

   // m322_114 = W*in
   wire signed [9:0] m322_114;
   assign m322_114 =10'b0;

   // m322_115 = W*in
   wire signed [9:0] m322_115;
   assign m322_115 =10'b0;

   // m322_116 = W*in
   wire signed [9:0] m322_116;
   assign m322_116 =10'b0;

   // m322_117 = W*in
   wire signed [9:0] m322_117;
   assign m322_117 =10'b0;

   // m323_1 = W*in
   wire signed [9:0] m323_1;
   assign m323_1 =10'b0;

   // m323_2 = W*in
   wire signed [9:0] m323_2;
   assign m323_2 =10'b0;

   // m323_3 = W*in
   wire signed [9:0] m323_3;
   assign m323_3 =10'b0;

   // m323_4 = W*in
   wire signed [9:0] m323_4;
   assign m323_4 =10'b0;

   // m323_5 = W*in
   wire signed [9:0] m323_5;
   assign m323_5 =10'b0;

   // m323_6 = W*in
   wire signed [9:0] m323_6;
   assign m323_6 =10'b0;

   // m323_7 = W*in
   wire signed [9:0] m323_7;
   assign m323_7 ={ {4{in323[5]}} , in323[5:0] };

   // m323_8 = W*in
   wire signed [9:0] m323_8;
   assign m323_8 =10'b0;

   // m323_9 = W*in
   wire signed [9:0] m323_9;
   assign m323_9 =10'b0;

   // m323_10 = W*in
   wire signed [9:0] m323_10;
   assign m323_10 =10'b0;

   // m323_11 = W*in
   wire signed [9:0] m323_11;
   assign m323_11 =10'b0;

   // m323_12 = W*in
   wire signed [9:0] m323_12;
   assign m323_12 =10'b0;

   // m323_13 = W*in
   wire signed [9:0] m323_13;
   assign m323_13 =10'b0;

   // m323_14 = W*in
   wire signed [9:0] m323_14;
   assign m323_14 =10'b0;

   // m323_15 = W*in
   wire signed [9:0] m323_15;
   assign m323_15 =10'b0;

   // m323_16 = W*in
   wire signed [9:0] m323_16;
   assign m323_16 ={ {5{in323[5]}} , in323[5:1] };

   // m323_17 = W*in
   wire signed [9:0] m323_17;
   assign m323_17 ={ {5{in323[5]}} , in323[5:1] };

   // m323_18 = W*in
   wire signed [9:0] m323_18;
   assign m323_18 ={ {5{neg323[5]}} , neg323[5:1] };

   // m323_19 = W*in
   wire signed [9:0] m323_19;
   assign m323_19 =10'b0;

   // m323_20 = W*in
   wire signed [9:0] m323_20;
   assign m323_20 =10'b0;

   // m323_21 = W*in
   wire signed [9:0] m323_21;
   assign m323_21 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_22 = W*in
   wire signed [9:0] m323_22;
   assign m323_22 =10'b0;

   // m323_23 = W*in
   wire signed [9:0] m323_23;
   assign m323_23 =10'b0;

   // m323_24 = W*in
   wire signed [9:0] m323_24;
   assign m323_24 =10'b0;

   // m323_25 = W*in
   wire signed [9:0] m323_25;
   assign m323_25 =10'b0;

   // m323_26 = W*in
   wire signed [9:0] m323_26;
   assign m323_26 =10'b0;

   // m323_27 = W*in
   wire signed [9:0] m323_27;
   assign m323_27 ={ {5{in323[5]}} , in323[5:1] };

   // m323_28 = W*in
   wire signed [9:0] m323_28;
   assign m323_28 =10'b0;

   // m323_29 = W*in
   wire signed [9:0] m323_29;
   assign m323_29 =10'b0;

   // m323_30 = W*in
   wire signed [9:0] m323_30;
   assign m323_30 ={ {5{neg323[5]}} , neg323[5:1] };

   // m323_31 = W*in
   wire signed [9:0] m323_31;
   assign m323_31 =10'b0;

   // m323_32 = W*in
   wire signed [9:0] m323_32;
   assign m323_32 =10'b0;

   // m323_33 = W*in
   wire signed [9:0] m323_33;
   assign m323_33 =10'b0;

   // m323_34 = W*in
   wire signed [9:0] m323_34;
   assign m323_34 =10'b0;

   // m323_35 = W*in
   wire signed [9:0] m323_35;
   assign m323_35 =10'b0;

   // m323_36 = W*in
   wire signed [9:0] m323_36;
   assign m323_36 =10'b0;

   // m323_37 = W*in
   wire signed [9:0] m323_37;
   assign m323_37 =10'b0;

   // m323_38 = W*in
   wire signed [9:0] m323_38;
   assign m323_38 =10'b0;

   // m323_39 = W*in
   wire signed [9:0] m323_39;
   assign m323_39 =10'b0;

   // m323_40 = W*in
   wire signed [9:0] m323_40;
   assign m323_40 =10'b0;

   // m323_41 = W*in
   wire signed [9:0] m323_41;
   assign m323_41 =10'b0;

   // m323_42 = W*in
   wire signed [9:0] m323_42;
   assign m323_42 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_43 = W*in
   wire signed [9:0] m323_43;
   assign m323_43 =10'b0;

   // m323_44 = W*in
   wire signed [9:0] m323_44;
   assign m323_44 =10'b0;

   // m323_45 = W*in
   wire signed [9:0] m323_45;
   assign m323_45 ={ {4{in323[5]}} , in323[5:0] };

   // m323_46 = W*in
   wire signed [9:0] m323_46;
   assign m323_46 =10'b0;

   // m323_47 = W*in
   wire signed [9:0] m323_47;
   assign m323_47 =10'b0;

   // m323_48 = W*in
   wire signed [9:0] m323_48;
   assign m323_48 =10'b0;

   // m323_49 = W*in
   wire signed [9:0] m323_49;
   assign m323_49 =10'b0;

   // m323_50 = W*in
   wire signed [9:0] m323_50;
   assign m323_50 =10'b0;

   // m323_51 = W*in
   wire signed [9:0] m323_51;
   assign m323_51 =10'b0;

   // m323_52 = W*in
   wire signed [9:0] m323_52;
   assign m323_52 =10'b0;

   // m323_53 = W*in
   wire signed [9:0] m323_53;
   assign m323_53 =10'b0;

   // m323_54 = W*in
   wire signed [9:0] m323_54;
   assign m323_54 =10'b0;

   // m323_55 = W*in
   wire signed [9:0] m323_55;
   assign m323_55 =10'b0;

   // m323_56 = W*in
   wire signed [9:0] m323_56;
   assign m323_56 ={ {4{in323[5]}} , in323[5:0] };

   // m323_57 = W*in
   wire signed [9:0] m323_57;
   assign m323_57 =10'b0;

   // m323_58 = W*in
   wire signed [9:0] m323_58;
   assign m323_58 =10'b0;

   // m323_59 = W*in
   wire signed [9:0] m323_59;
   assign m323_59 =10'b0;

   // m323_60 = W*in
   wire signed [9:0] m323_60;
   assign m323_60 =10'b0;

   // m323_61 = W*in
   wire signed [9:0] m323_61;
   assign m323_61 =10'b0;

   // m323_62 = W*in
   wire signed [9:0] m323_62;
   assign m323_62 =10'b0;

   // m323_63 = W*in
   wire signed [9:0] m323_63;
   assign m323_63 =10'b0;

   // m323_64 = W*in
   wire signed [9:0] m323_64;
   assign m323_64 ={ {5{in323[5]}} , in323[5:1] };

   // m323_65 = W*in
   wire signed [9:0] m323_65;
   assign m323_65 ={ {5{in323[5]}} , in323[5:1] };

   // m323_66 = W*in
   wire signed [9:0] m323_66;
   assign m323_66 =10'b0;

   // m323_67 = W*in
   wire signed [9:0] m323_67;
   assign m323_67 =10'b0;

   // m323_68 = W*in
   wire signed [9:0] m323_68;
   assign m323_68 =10'b0;

   // m323_69 = W*in
   wire signed [9:0] m323_69;
   assign m323_69 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_70 = W*in
   wire signed [9:0] m323_70;
   assign m323_70 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_71 = W*in
   wire signed [9:0] m323_71;
   assign m323_71 =10'b0;

   // m323_72 = W*in
   wire signed [9:0] m323_72;
   assign m323_72 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_73 = W*in
   wire signed [9:0] m323_73;
   assign m323_73 =10'b0;

   // m323_74 = W*in
   wire signed [9:0] m323_74;
   assign m323_74 ={ {5{neg323[5]}} , neg323[5:1] };

   // m323_75 = W*in
   wire signed [9:0] m323_75;
   assign m323_75 =10'b0;

   // m323_76 = W*in
   wire signed [9:0] m323_76;
   assign m323_76 =10'b0;

   // m323_77 = W*in
   wire signed [9:0] m323_77;
   assign m323_77 =10'b0;

   // m323_78 = W*in
   wire signed [9:0] m323_78;
   assign m323_78 =10'b0;

   // m323_79 = W*in
   wire signed [9:0] m323_79;
   assign m323_79 =10'b0;

   // m323_80 = W*in
   wire signed [9:0] m323_80;
   assign m323_80 =10'b0;

   // m323_81 = W*in
   wire signed [9:0] m323_81;
   assign m323_81 =10'b0;

   // m323_82 = W*in
   wire signed [9:0] m323_82;
   assign m323_82 =10'b0;

   // m323_83 = W*in
   wire signed [9:0] m323_83;
   assign m323_83 =10'b0;

   // m323_84 = W*in
   wire signed [9:0] m323_84;
   assign m323_84 =10'b0;

   // m323_85 = W*in
   wire signed [9:0] m323_85;
   assign m323_85 =10'b0;

   // m323_86 = W*in
   wire signed [9:0] m323_86;
   assign m323_86 =10'b0;

   // m323_87 = W*in
   wire signed [9:0] m323_87;
   assign m323_87 =10'b0;

   // m323_88 = W*in
   wire signed [9:0] m323_88;
   assign m323_88 =10'b0;

   // m323_89 = W*in
   wire signed [9:0] m323_89;
   assign m323_89 =10'b0;

   // m323_90 = W*in
   wire signed [9:0] m323_90;
   assign m323_90 =10'b0;

   // m323_91 = W*in
   wire signed [9:0] m323_91;
   assign m323_91 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_92 = W*in
   wire signed [9:0] m323_92;
   assign m323_92 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_93 = W*in
   wire signed [9:0] m323_93;
   assign m323_93 =10'b0;

   // m323_94 = W*in
   wire signed [9:0] m323_94;
   assign m323_94 =10'b0;

   // m323_95 = W*in
   wire signed [9:0] m323_95;
   assign m323_95 =10'b0;

   // m323_96 = W*in
   wire signed [9:0] m323_96;
   assign m323_96 =10'b0;

   // m323_97 = W*in
   wire signed [9:0] m323_97;
   assign m323_97 =10'b0;

   // m323_98 = W*in
   wire signed [9:0] m323_98;
   assign m323_98 =10'b0;

   // m323_99 = W*in
   wire signed [9:0] m323_99;
   assign m323_99 ={ {4{neg323[5]}} , neg323[5:0] };

   // m323_100 = W*in
   wire signed [9:0] m323_100;
   assign m323_100 =10'b0;

   // m323_101 = W*in
   wire signed [9:0] m323_101;
   assign m323_101 =10'b0;

   // m323_102 = W*in
   wire signed [9:0] m323_102;
   assign m323_102 =10'b0;

   // m323_103 = W*in
   wire signed [9:0] m323_103;
   assign m323_103 =10'b0;

   // m323_104 = W*in
   wire signed [9:0] m323_104;
   assign m323_104 ={ {4{in323[5]}} , in323[5:0] };

   // m323_105 = W*in
   wire signed [9:0] m323_105;
   assign m323_105 =10'b0;

   // m323_106 = W*in
   wire signed [9:0] m323_106;
   assign m323_106 =10'b0;

   // m323_107 = W*in
   wire signed [9:0] m323_107;
   assign m323_107 =10'b0;

   // m323_108 = W*in
   wire signed [9:0] m323_108;
   assign m323_108 =10'b0;

   // m323_109 = W*in
   wire signed [9:0] m323_109;
   assign m323_109 =10'b0;

   // m323_110 = W*in
   wire signed [9:0] m323_110;
   assign m323_110 =10'b0;

   // m323_111 = W*in
   wire signed [9:0] m323_111;
   assign m323_111 =10'b0;

   // m323_112 = W*in
   wire signed [9:0] m323_112;
   assign m323_112 =10'b0;

   // m323_113 = W*in
   wire signed [9:0] m323_113;
   assign m323_113 =10'b0;

   // m323_114 = W*in
   wire signed [9:0] m323_114;
   assign m323_114 =10'b0;

   // m323_115 = W*in
   wire signed [9:0] m323_115;
   assign m323_115 =10'b0;

   // m323_116 = W*in
   wire signed [9:0] m323_116;
   assign m323_116 =10'b0;

   // m323_117 = W*in
   wire signed [9:0] m323_117;
   assign m323_117 =10'b0;

   // m324_1 = W*in
   wire signed [9:0] m324_1;
   assign m324_1 =10'b0;

   // m324_2 = W*in
   wire signed [9:0] m324_2;
   assign m324_2 =10'b0;

   // m324_3 = W*in
   wire signed [9:0] m324_3;
   assign m324_3 =10'b0;

   // m324_4 = W*in
   wire signed [9:0] m324_4;
   assign m324_4 =10'b0;

   // m324_5 = W*in
   wire signed [9:0] m324_5;
   assign m324_5 =10'b0;

   // m324_6 = W*in
   wire signed [9:0] m324_6;
   assign m324_6 =10'b0;

   // m324_7 = W*in
   wire signed [9:0] m324_7;
   assign m324_7 =10'b0;

   // m324_8 = W*in
   wire signed [9:0] m324_8;
   assign m324_8 =10'b0;

   // m324_9 = W*in
   wire signed [9:0] m324_9;
   assign m324_9 =10'b0;

   // m324_10 = W*in
   wire signed [9:0] m324_10;
   assign m324_10 =10'b0;

   // m324_11 = W*in
   wire signed [9:0] m324_11;
   assign m324_11 =10'b0;

   // m324_12 = W*in
   wire signed [9:0] m324_12;
   assign m324_12 =10'b0;

   // m324_13 = W*in
   wire signed [9:0] m324_13;
   assign m324_13 =10'b0;

   // m324_14 = W*in
   wire signed [9:0] m324_14;
   assign m324_14 =10'b0;

   // m324_15 = W*in
   wire signed [9:0] m324_15;
   assign m324_15 =10'b0;

   // m324_16 = W*in
   wire signed [9:0] m324_16;
   assign m324_16 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_17 = W*in
   wire signed [9:0] m324_17;
   assign m324_17 =10'b0;

   // m324_18 = W*in
   wire signed [9:0] m324_18;
   assign m324_18 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_19 = W*in
   wire signed [9:0] m324_19;
   assign m324_19 =10'b0;

   // m324_20 = W*in
   wire signed [9:0] m324_20;
   assign m324_20 =10'b0;

   // m324_21 = W*in
   wire signed [9:0] m324_21;
   assign m324_21 =10'b0;

   // m324_22 = W*in
   wire signed [9:0] m324_22;
   assign m324_22 =10'b0;

   // m324_23 = W*in
   wire signed [9:0] m324_23;
   assign m324_23 =10'b0;

   // m324_24 = W*in
   wire signed [9:0] m324_24;
   assign m324_24 =10'b0;

   // m324_25 = W*in
   wire signed [9:0] m324_25;
   assign m324_25 ={ {5{in324[5]}} , in324[5:1] };

   // m324_26 = W*in
   wire signed [9:0] m324_26;
   assign m324_26 =10'b0;

   // m324_27 = W*in
   wire signed [9:0] m324_27;
   assign m324_27 =10'b0;

   // m324_28 = W*in
   wire signed [9:0] m324_28;
   assign m324_28 =10'b0;

   // m324_29 = W*in
   wire signed [9:0] m324_29;
   assign m324_29 =10'b0;

   // m324_30 = W*in
   wire signed [9:0] m324_30;
   assign m324_30 =10'b0;

   // m324_31 = W*in
   wire signed [9:0] m324_31;
   assign m324_31 =10'b0;

   // m324_32 = W*in
   wire signed [9:0] m324_32;
   assign m324_32 =10'b0;

   // m324_33 = W*in
   wire signed [9:0] m324_33;
   assign m324_33 =10'b0;

   // m324_34 = W*in
   wire signed [9:0] m324_34;
   assign m324_34 =10'b0;

   // m324_35 = W*in
   wire signed [9:0] m324_35;
   assign m324_35 =10'b0;

   // m324_36 = W*in
   wire signed [9:0] m324_36;
   assign m324_36 =10'b0;

   // m324_37 = W*in
   wire signed [9:0] m324_37;
   assign m324_37 =10'b0;

   // m324_38 = W*in
   wire signed [9:0] m324_38;
   assign m324_38 ={ {4{neg324[5]}} , neg324[5:0] };

   // m324_39 = W*in
   wire signed [9:0] m324_39;
   assign m324_39 =10'b0;

   // m324_40 = W*in
   wire signed [9:0] m324_40;
   assign m324_40 =10'b0;

   // m324_41 = W*in
   wire signed [9:0] m324_41;
   assign m324_41 =10'b0;

   // m324_42 = W*in
   wire signed [9:0] m324_42;
   assign m324_42 =10'b0;

   // m324_43 = W*in
   wire signed [9:0] m324_43;
   assign m324_43 =10'b0;

   // m324_44 = W*in
   wire signed [9:0] m324_44;
   assign m324_44 =10'b0;

   // m324_45 = W*in
   wire signed [9:0] m324_45;
   assign m324_45 =10'b0;

   // m324_46 = W*in
   wire signed [9:0] m324_46;
   assign m324_46 =10'b0;

   // m324_47 = W*in
   wire signed [9:0] m324_47;
   assign m324_47 =10'b0;

   // m324_48 = W*in
   wire signed [9:0] m324_48;
   assign m324_48 =10'b0;

   // m324_49 = W*in
   wire signed [9:0] m324_49;
   assign m324_49 =10'b0;

   // m324_50 = W*in
   wire signed [9:0] m324_50;
   assign m324_50 =10'b0;

   // m324_51 = W*in
   wire signed [9:0] m324_51;
   assign m324_51 =10'b0;

   // m324_52 = W*in
   wire signed [9:0] m324_52;
   assign m324_52 =10'b0;

   // m324_53 = W*in
   wire signed [9:0] m324_53;
   assign m324_53 =10'b0;

   // m324_54 = W*in
   wire signed [9:0] m324_54;
   assign m324_54 =10'b0;

   // m324_55 = W*in
   wire signed [9:0] m324_55;
   assign m324_55 =10'b0;

   // m324_56 = W*in
   wire signed [9:0] m324_56;
   assign m324_56 =10'b0;

   // m324_57 = W*in
   wire signed [9:0] m324_57;
   assign m324_57 =10'b0;

   // m324_58 = W*in
   wire signed [9:0] m324_58;
   assign m324_58 =10'b0;

   // m324_59 = W*in
   wire signed [9:0] m324_59;
   assign m324_59 =10'b0;

   // m324_60 = W*in
   wire signed [9:0] m324_60;
   assign m324_60 =10'b0;

   // m324_61 = W*in
   wire signed [9:0] m324_61;
   assign m324_61 =10'b0;

   // m324_62 = W*in
   wire signed [9:0] m324_62;
   assign m324_62 =10'b0;

   // m324_63 = W*in
   wire signed [9:0] m324_63;
   assign m324_63 =10'b0;

   // m324_64 = W*in
   wire signed [9:0] m324_64;
   assign m324_64 =10'b0;

   // m324_65 = W*in
   wire signed [9:0] m324_65;
   assign m324_65 =10'b0;

   // m324_66 = W*in
   wire signed [9:0] m324_66;
   assign m324_66 =10'b0;

   // m324_67 = W*in
   wire signed [9:0] m324_67;
   assign m324_67 =10'b0;

   // m324_68 = W*in
   wire signed [9:0] m324_68;
   assign m324_68 =10'b0;

   // m324_69 = W*in
   wire signed [9:0] m324_69;
   assign m324_69 ={ {5{in324[5]}} , in324[5:1] };

   // m324_70 = W*in
   wire signed [9:0] m324_70;
   assign m324_70 =10'b0;

   // m324_71 = W*in
   wire signed [9:0] m324_71;
   assign m324_71 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_72 = W*in
   wire signed [9:0] m324_72;
   assign m324_72 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_73 = W*in
   wire signed [9:0] m324_73;
   assign m324_73 ={ {5{in324[5]}} , in324[5:1] };

   // m324_74 = W*in
   wire signed [9:0] m324_74;
   assign m324_74 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_75 = W*in
   wire signed [9:0] m324_75;
   assign m324_75 =10'b0;

   // m324_76 = W*in
   wire signed [9:0] m324_76;
   assign m324_76 =10'b0;

   // m324_77 = W*in
   wire signed [9:0] m324_77;
   assign m324_77 =10'b0;

   // m324_78 = W*in
   wire signed [9:0] m324_78;
   assign m324_78 =10'b0;

   // m324_79 = W*in
   wire signed [9:0] m324_79;
   assign m324_79 =10'b0;

   // m324_80 = W*in
   wire signed [9:0] m324_80;
   assign m324_80 =10'b0;

   // m324_81 = W*in
   wire signed [9:0] m324_81;
   assign m324_81 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_82 = W*in
   wire signed [9:0] m324_82;
   assign m324_82 ={ {4{in324[5]}} , in324[5:0] };

   // m324_83 = W*in
   wire signed [9:0] m324_83;
   assign m324_83 ={ {5{neg324[5]}} , neg324[5:1] };

   // m324_84 = W*in
   wire signed [9:0] m324_84;
   assign m324_84 =10'b0;

   // m324_85 = W*in
   wire signed [9:0] m324_85;
   assign m324_85 =10'b0;

   // m324_86 = W*in
   wire signed [9:0] m324_86;
   assign m324_86 =10'b0;

   // m324_87 = W*in
   wire signed [9:0] m324_87;
   assign m324_87 =10'b0;

   // m324_88 = W*in
   wire signed [9:0] m324_88;
   assign m324_88 =10'b0;

   // m324_89 = W*in
   wire signed [9:0] m324_89;
   assign m324_89 =10'b0;

   // m324_90 = W*in
   wire signed [9:0] m324_90;
   assign m324_90 =10'b0;

   // m324_91 = W*in
   wire signed [9:0] m324_91;
   assign m324_91 =10'b0;

   // m324_92 = W*in
   wire signed [9:0] m324_92;
   assign m324_92 =10'b0;

   // m324_93 = W*in
   wire signed [9:0] m324_93;
   assign m324_93 =10'b0;

   // m324_94 = W*in
   wire signed [9:0] m324_94;
   assign m324_94 =10'b0;

   // m324_95 = W*in
   wire signed [9:0] m324_95;
   assign m324_95 =10'b0;

   // m324_96 = W*in
   wire signed [9:0] m324_96;
   assign m324_96 =10'b0;

   // m324_97 = W*in
   wire signed [9:0] m324_97;
   assign m324_97 =10'b0;

   // m324_98 = W*in
   wire signed [9:0] m324_98;
   assign m324_98 =10'b0;

   // m324_99 = W*in
   wire signed [9:0] m324_99;
   assign m324_99 =10'b0;

   // m324_100 = W*in
   wire signed [9:0] m324_100;
   assign m324_100 =10'b0;

   // m324_101 = W*in
   wire signed [9:0] m324_101;
   assign m324_101 =10'b0;

   // m324_102 = W*in
   wire signed [9:0] m324_102;
   assign m324_102 =10'b0;

   // m324_103 = W*in
   wire signed [9:0] m324_103;
   assign m324_103 =10'b0;

   // m324_104 = W*in
   wire signed [9:0] m324_104;
   assign m324_104 =10'b0;

   // m324_105 = W*in
   wire signed [9:0] m324_105;
   assign m324_105 =10'b0;

   // m324_106 = W*in
   wire signed [9:0] m324_106;
   assign m324_106 =10'b0;

   // m324_107 = W*in
   wire signed [9:0] m324_107;
   assign m324_107 =10'b0;

   // m324_108 = W*in
   wire signed [9:0] m324_108;
   assign m324_108 ={ {5{in324[5]}} , in324[5:1] };

   // m324_109 = W*in
   wire signed [9:0] m324_109;
   assign m324_109 ={ {4{in324[5]}} , in324[5:0] };

   // m324_110 = W*in
   wire signed [9:0] m324_110;
   assign m324_110 =10'b0;

   // m324_111 = W*in
   wire signed [9:0] m324_111;
   assign m324_111 =10'b0;

   // m324_112 = W*in
   wire signed [9:0] m324_112;
   assign m324_112 =10'b0;

   // m324_113 = W*in
   wire signed [9:0] m324_113;
   assign m324_113 =10'b0;

   // m324_114 = W*in
   wire signed [9:0] m324_114;
   assign m324_114 =10'b0;

   // m324_115 = W*in
   wire signed [9:0] m324_115;
   assign m324_115 =10'b0;

   // m324_116 = W*in
   wire signed [9:0] m324_116;
   assign m324_116 =10'b0;

   // m324_117 = W*in
   wire signed [9:0] m324_117;
   assign m324_117 =10'b0;

   // m325_1 = W*in
   wire signed [9:0] m325_1;
   assign m325_1 =10'b0;

   // m325_2 = W*in
   wire signed [9:0] m325_2;
   assign m325_2 =10'b0;

   // m325_3 = W*in
   wire signed [9:0] m325_3;
   assign m325_3 =10'b0;

   // m325_4 = W*in
   wire signed [9:0] m325_4;
   assign m325_4 =10'b0;

   // m325_5 = W*in
   wire signed [9:0] m325_5;
   assign m325_5 =10'b0;

   // m325_6 = W*in
   wire signed [9:0] m325_6;
   assign m325_6 =10'b0;

   // m325_7 = W*in
   wire signed [9:0] m325_7;
   assign m325_7 =10'b0;

   // m325_8 = W*in
   wire signed [9:0] m325_8;
   assign m325_8 ={ {4{in325[5]}} , in325[5:0] };

   // m325_9 = W*in
   wire signed [9:0] m325_9;
   assign m325_9 =10'b0;

   // m325_10 = W*in
   wire signed [9:0] m325_10;
   assign m325_10 =10'b0;

   // m325_11 = W*in
   wire signed [9:0] m325_11;
   assign m325_11 =10'b0;

   // m325_12 = W*in
   wire signed [9:0] m325_12;
   assign m325_12 =10'b0;

   // m325_13 = W*in
   wire signed [9:0] m325_13;
   assign m325_13 =10'b0;

   // m325_14 = W*in
   wire signed [9:0] m325_14;
   assign m325_14 =10'b0;

   // m325_15 = W*in
   wire signed [9:0] m325_15;
   assign m325_15 =10'b0;

   // m325_16 = W*in
   wire signed [9:0] m325_16;
   assign m325_16 =10'b0;

   // m325_17 = W*in
   wire signed [9:0] m325_17;
   assign m325_17 =10'b0;

   // m325_18 = W*in
   wire signed [9:0] m325_18;
   assign m325_18 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_19 = W*in
   wire signed [9:0] m325_19;
   assign m325_19 =10'b0;

   // m325_20 = W*in
   wire signed [9:0] m325_20;
   assign m325_20 =10'b0;

   // m325_21 = W*in
   wire signed [9:0] m325_21;
   assign m325_21 ={ {5{neg325[5]}} , neg325[5:1] };

   // m325_22 = W*in
   wire signed [9:0] m325_22;
   assign m325_22 =10'b0;

   // m325_23 = W*in
   wire signed [9:0] m325_23;
   assign m325_23 =10'b0;

   // m325_24 = W*in
   wire signed [9:0] m325_24;
   assign m325_24 =10'b0;

   // m325_25 = W*in
   wire signed [9:0] m325_25;
   assign m325_25 =10'b0;

   // m325_26 = W*in
   wire signed [9:0] m325_26;
   assign m325_26 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_27 = W*in
   wire signed [9:0] m325_27;
   assign m325_27 ={ {5{in325[5]}} , in325[5:1] };

   // m325_28 = W*in
   wire signed [9:0] m325_28;
   assign m325_28 =10'b0;

   // m325_29 = W*in
   wire signed [9:0] m325_29;
   assign m325_29 =10'b0;

   // m325_30 = W*in
   wire signed [9:0] m325_30;
   assign m325_30 =10'b0;

   // m325_31 = W*in
   wire signed [9:0] m325_31;
   assign m325_31 =10'b0;

   // m325_32 = W*in
   wire signed [9:0] m325_32;
   assign m325_32 =10'b0;

   // m325_33 = W*in
   wire signed [9:0] m325_33;
   assign m325_33 =10'b0;

   // m325_34 = W*in
   wire signed [9:0] m325_34;
   assign m325_34 ={ {4{in325[5]}} , in325[5:0] };

   // m325_35 = W*in
   wire signed [9:0] m325_35;
   assign m325_35 =10'b0;

   // m325_36 = W*in
   wire signed [9:0] m325_36;
   assign m325_36 =10'b0;

   // m325_37 = W*in
   wire signed [9:0] m325_37;
   assign m325_37 =10'b0;

   // m325_38 = W*in
   wire signed [9:0] m325_38;
   assign m325_38 =10'b0;

   // m325_39 = W*in
   wire signed [9:0] m325_39;
   assign m325_39 =10'b0;

   // m325_40 = W*in
   wire signed [9:0] m325_40;
   assign m325_40 =10'b0;

   // m325_41 = W*in
   wire signed [9:0] m325_41;
   assign m325_41 =10'b0;

   // m325_42 = W*in
   wire signed [9:0] m325_42;
   assign m325_42 =10'b0;

   // m325_43 = W*in
   wire signed [9:0] m325_43;
   assign m325_43 =10'b0;

   // m325_44 = W*in
   wire signed [9:0] m325_44;
   assign m325_44 =10'b0;

   // m325_45 = W*in
   wire signed [9:0] m325_45;
   assign m325_45 =10'b0;

   // m325_46 = W*in
   wire signed [9:0] m325_46;
   assign m325_46 =10'b0;

   // m325_47 = W*in
   wire signed [9:0] m325_47;
   assign m325_47 =10'b0;

   // m325_48 = W*in
   wire signed [9:0] m325_48;
   assign m325_48 =10'b0;

   // m325_49 = W*in
   wire signed [9:0] m325_49;
   assign m325_49 =10'b0;

   // m325_50 = W*in
   wire signed [9:0] m325_50;
   assign m325_50 =10'b0;

   // m325_51 = W*in
   wire signed [9:0] m325_51;
   assign m325_51 =10'b0;

   // m325_52 = W*in
   wire signed [9:0] m325_52;
   assign m325_52 =10'b0;

   // m325_53 = W*in
   wire signed [9:0] m325_53;
   assign m325_53 =10'b0;

   // m325_54 = W*in
   wire signed [9:0] m325_54;
   assign m325_54 =10'b0;

   // m325_55 = W*in
   wire signed [9:0] m325_55;
   assign m325_55 =10'b0;

   // m325_56 = W*in
   wire signed [9:0] m325_56;
   assign m325_56 =10'b0;

   // m325_57 = W*in
   wire signed [9:0] m325_57;
   assign m325_57 =10'b0;

   // m325_58 = W*in
   wire signed [9:0] m325_58;
   assign m325_58 =10'b0;

   // m325_59 = W*in
   wire signed [9:0] m325_59;
   assign m325_59 =10'b0;

   // m325_60 = W*in
   wire signed [9:0] m325_60;
   assign m325_60 =10'b0;

   // m325_61 = W*in
   wire signed [9:0] m325_61;
   assign m325_61 =10'b0;

   // m325_62 = W*in
   wire signed [9:0] m325_62;
   assign m325_62 =10'b0;

   // m325_63 = W*in
   wire signed [9:0] m325_63;
   assign m325_63 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_64 = W*in
   wire signed [9:0] m325_64;
   assign m325_64 =10'b0;

   // m325_65 = W*in
   wire signed [9:0] m325_65;
   assign m325_65 ={ {5{neg325[5]}} , neg325[5:1] };

   // m325_66 = W*in
   wire signed [9:0] m325_66;
   assign m325_66 =10'b0;

   // m325_67 = W*in
   wire signed [9:0] m325_67;
   assign m325_67 =10'b0;

   // m325_68 = W*in
   wire signed [9:0] m325_68;
   assign m325_68 =10'b0;

   // m325_69 = W*in
   wire signed [9:0] m325_69;
   assign m325_69 ={ {5{neg325[5]}} , neg325[5:1] };

   // m325_70 = W*in
   wire signed [9:0] m325_70;
   assign m325_70 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_71 = W*in
   wire signed [9:0] m325_71;
   assign m325_71 =10'b0;

   // m325_72 = W*in
   wire signed [9:0] m325_72;
   assign m325_72 =10'b0;

   // m325_73 = W*in
   wire signed [9:0] m325_73;
   assign m325_73 ={ {5{in325[5]}} , in325[5:1] };

   // m325_74 = W*in
   wire signed [9:0] m325_74;
   assign m325_74 =10'b0;

   // m325_75 = W*in
   wire signed [9:0] m325_75;
   assign m325_75 ={ {4{in325[5]}} , in325[5:0] };

   // m325_76 = W*in
   wire signed [9:0] m325_76;
   assign m325_76 =10'b0;

   // m325_77 = W*in
   wire signed [9:0] m325_77;
   assign m325_77 ={ {4{in325[5]}} , in325[5:0] };

   // m325_78 = W*in
   wire signed [9:0] m325_78;
   assign m325_78 =10'b0;

   // m325_79 = W*in
   wire signed [9:0] m325_79;
   assign m325_79 =10'b0;

   // m325_80 = W*in
   wire signed [9:0] m325_80;
   assign m325_80 ={ {5{in325[5]}} , in325[5:1] };

   // m325_81 = W*in
   wire signed [9:0] m325_81;
   assign m325_81 ={ {5{in325[5]}} , in325[5:1] };

   // m325_82 = W*in
   wire signed [9:0] m325_82;
   assign m325_82 =10'b0;

   // m325_83 = W*in
   wire signed [9:0] m325_83;
   assign m325_83 =10'b0;

   // m325_84 = W*in
   wire signed [9:0] m325_84;
   assign m325_84 =10'b0;

   // m325_85 = W*in
   wire signed [9:0] m325_85;
   assign m325_85 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_86 = W*in
   wire signed [9:0] m325_86;
   assign m325_86 =10'b0;

   // m325_87 = W*in
   wire signed [9:0] m325_87;
   assign m325_87 =10'b0;

   // m325_88 = W*in
   wire signed [9:0] m325_88;
   assign m325_88 =10'b0;

   // m325_89 = W*in
   wire signed [9:0] m325_89;
   assign m325_89 =10'b0;

   // m325_90 = W*in
   wire signed [9:0] m325_90;
   assign m325_90 =10'b0;

   // m325_91 = W*in
   wire signed [9:0] m325_91;
   assign m325_91 =10'b0;

   // m325_92 = W*in
   wire signed [9:0] m325_92;
   assign m325_92 =10'b0;

   // m325_93 = W*in
   wire signed [9:0] m325_93;
   assign m325_93 =10'b0;

   // m325_94 = W*in
   wire signed [9:0] m325_94;
   assign m325_94 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_95 = W*in
   wire signed [9:0] m325_95;
   assign m325_95 =10'b0;

   // m325_96 = W*in
   wire signed [9:0] m325_96;
   assign m325_96 =10'b0;

   // m325_97 = W*in
   wire signed [9:0] m325_97;
   assign m325_97 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_98 = W*in
   wire signed [9:0] m325_98;
   assign m325_98 =10'b0;

   // m325_99 = W*in
   wire signed [9:0] m325_99;
   assign m325_99 =10'b0;

   // m325_100 = W*in
   wire signed [9:0] m325_100;
   assign m325_100 =10'b0;

   // m325_101 = W*in
   wire signed [9:0] m325_101;
   assign m325_101 =10'b0;

   // m325_102 = W*in
   wire signed [9:0] m325_102;
   assign m325_102 =10'b0;

   // m325_103 = W*in
   wire signed [9:0] m325_103;
   assign m325_103 =10'b0;

   // m325_104 = W*in
   wire signed [9:0] m325_104;
   assign m325_104 =10'b0;

   // m325_105 = W*in
   wire signed [9:0] m325_105;
   assign m325_105 =10'b0;

   // m325_106 = W*in
   wire signed [9:0] m325_106;
   assign m325_106 =10'b0;

   // m325_107 = W*in
   wire signed [9:0] m325_107;
   assign m325_107 =10'b0;

   // m325_108 = W*in
   wire signed [9:0] m325_108;
   assign m325_108 =10'b0;

   // m325_109 = W*in
   wire signed [9:0] m325_109;
   assign m325_109 =10'b0;

   // m325_110 = W*in
   wire signed [9:0] m325_110;
   assign m325_110 =10'b0;

   // m325_111 = W*in
   wire signed [9:0] m325_111;
   assign m325_111 =10'b0;

   // m325_112 = W*in
   wire signed [9:0] m325_112;
   assign m325_112 =10'b0;

   // m325_113 = W*in
   wire signed [9:0] m325_113;
   assign m325_113 =10'b0;

   // m325_114 = W*in
   wire signed [9:0] m325_114;
   assign m325_114 ={ {5{in325[5]}} , in325[5:1] };

   // m325_115 = W*in
   wire signed [9:0] m325_115;
   assign m325_115 ={ {5{in325[5]}} , in325[5:1] };

   // m325_116 = W*in
   wire signed [9:0] m325_116;
   assign m325_116 ={ {4{neg325[5]}} , neg325[5:0] };

   // m325_117 = W*in
   wire signed [9:0] m325_117;
   assign m325_117 =10'b0;

   // m326_1 = W*in
   wire signed [9:0] m326_1;
   assign m326_1 ={ {4{in326[5]}} , in326[5:0] };

   // m326_2 = W*in
   wire signed [9:0] m326_2;
   assign m326_2 =10'b0;

   // m326_3 = W*in
   wire signed [9:0] m326_3;
   assign m326_3 =10'b0;

   // m326_4 = W*in
   wire signed [9:0] m326_4;
   assign m326_4 ={ {4{in326[5]}} , in326[5:0] };

   // m326_5 = W*in
   wire signed [9:0] m326_5;
   assign m326_5 =10'b0;

   // m326_6 = W*in
   wire signed [9:0] m326_6;
   assign m326_6 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_7 = W*in
   wire signed [9:0] m326_7;
   assign m326_7 =10'b0;

   // m326_8 = W*in
   wire signed [9:0] m326_8;
   assign m326_8 =10'b0;

   // m326_9 = W*in
   wire signed [9:0] m326_9;
   assign m326_9 =10'b0;

   // m326_10 = W*in
   wire signed [9:0] m326_10;
   assign m326_10 =10'b0;

   // m326_11 = W*in
   wire signed [9:0] m326_11;
   assign m326_11 ={ {4{in326[5]}} , in326[5:0] };

   // m326_12 = W*in
   wire signed [9:0] m326_12;
   assign m326_12 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_13 = W*in
   wire signed [9:0] m326_13;
   assign m326_13 =10'b0;

   // m326_14 = W*in
   wire signed [9:0] m326_14;
   assign m326_14 =10'b0;

   // m326_15 = W*in
   wire signed [9:0] m326_15;
   assign m326_15 ={ {4{in326[5]}} , in326[5:0] };

   // m326_16 = W*in
   wire signed [9:0] m326_16;
   assign m326_16 ={ {4{in326[5]}} , in326[5:0] };

   // m326_17 = W*in
   wire signed [9:0] m326_17;
   assign m326_17 =10'b0;

   // m326_18 = W*in
   wire signed [9:0] m326_18;
   assign m326_18 =10'b0;

   // m326_19 = W*in
   wire signed [9:0] m326_19;
   assign m326_19 =10'b0;

   // m326_20 = W*in
   wire signed [9:0] m326_20;
   assign m326_20 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_21 = W*in
   wire signed [9:0] m326_21;
   assign m326_21 ={ {5{neg326[5]}} , neg326[5:1] };

   // m326_22 = W*in
   wire signed [9:0] m326_22;
   assign m326_22 =10'b0;

   // m326_23 = W*in
   wire signed [9:0] m326_23;
   assign m326_23 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_24 = W*in
   wire signed [9:0] m326_24;
   assign m326_24 =10'b0;

   // m326_25 = W*in
   wire signed [9:0] m326_25;
   assign m326_25 =10'b0;

   // m326_26 = W*in
   wire signed [9:0] m326_26;
   assign m326_26 =10'b0;

   // m326_27 = W*in
   wire signed [9:0] m326_27;
   assign m326_27 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_28 = W*in
   wire signed [9:0] m326_28;
   assign m326_28 =10'b0;

   // m326_29 = W*in
   wire signed [9:0] m326_29;
   assign m326_29 =10'b0;

   // m326_30 = W*in
   wire signed [9:0] m326_30;
   assign m326_30 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_31 = W*in
   wire signed [9:0] m326_31;
   assign m326_31 =10'b0;

   // m326_32 = W*in
   wire signed [9:0] m326_32;
   assign m326_32 =10'b0;

   // m326_33 = W*in
   wire signed [9:0] m326_33;
   assign m326_33 =10'b0;

   // m326_34 = W*in
   wire signed [9:0] m326_34;
   assign m326_34 =10'b0;

   // m326_35 = W*in
   wire signed [9:0] m326_35;
   assign m326_35 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_36 = W*in
   wire signed [9:0] m326_36;
   assign m326_36 =10'b0;

   // m326_37 = W*in
   wire signed [9:0] m326_37;
   assign m326_37 ={ {4{in326[5]}} , in326[5:0] };

   // m326_38 = W*in
   wire signed [9:0] m326_38;
   assign m326_38 =10'b0;

   // m326_39 = W*in
   wire signed [9:0] m326_39;
   assign m326_39 =10'b0;

   // m326_40 = W*in
   wire signed [9:0] m326_40;
   assign m326_40 =10'b0;

   // m326_41 = W*in
   wire signed [9:0] m326_41;
   assign m326_41 =10'b0;

   // m326_42 = W*in
   wire signed [9:0] m326_42;
   assign m326_42 =10'b0;

   // m326_43 = W*in
   wire signed [9:0] m326_43;
   assign m326_43 =10'b0;

   // m326_44 = W*in
   wire signed [9:0] m326_44;
   assign m326_44 =10'b0;

   // m326_45 = W*in
   wire signed [9:0] m326_45;
   assign m326_45 ={ {4{in326[5]}} , in326[5:0] };

   // m326_46 = W*in
   wire signed [9:0] m326_46;
   assign m326_46 =10'b0;

   // m326_47 = W*in
   wire signed [9:0] m326_47;
   assign m326_47 =10'b0;

   // m326_48 = W*in
   wire signed [9:0] m326_48;
   assign m326_48 ={ {3{in326[5]}} , in326 , {1{1'b0}} };

   // m326_49 = W*in
   wire signed [9:0] m326_49;
   assign m326_49 =10'b0;

   // m326_50 = W*in
   wire signed [9:0] m326_50;
   assign m326_50 ={ {4{in326[5]}} , in326[5:0] };

   // m326_51 = W*in
   wire signed [9:0] m326_51;
   assign m326_51 ={ {4{in326[5]}} , in326[5:0] };

   // m326_52 = W*in
   wire signed [9:0] m326_52;
   assign m326_52 =10'b0;

   // m326_53 = W*in
   wire signed [9:0] m326_53;
   assign m326_53 =10'b0;

   // m326_54 = W*in
   wire signed [9:0] m326_54;
   assign m326_54 =10'b0;

   // m326_55 = W*in
   wire signed [9:0] m326_55;
   assign m326_55 =10'b0;

   // m326_56 = W*in
   wire signed [9:0] m326_56;
   assign m326_56 =10'b0;

   // m326_57 = W*in
   wire signed [9:0] m326_57;
   assign m326_57 =10'b0;

   // m326_58 = W*in
   wire signed [9:0] m326_58;
   assign m326_58 =10'b0;

   // m326_59 = W*in
   wire signed [9:0] m326_59;
   assign m326_59 =10'b0;

   // m326_60 = W*in
   wire signed [9:0] m326_60;
   assign m326_60 =10'b0;

   // m326_61 = W*in
   wire signed [9:0] m326_61;
   assign m326_61 =10'b0;

   // m326_62 = W*in
   wire signed [9:0] m326_62;
   assign m326_62 ={ {4{in326[5]}} , in326[5:0] };

   // m326_63 = W*in
   wire signed [9:0] m326_63;
   assign m326_63 =10'b0;

   // m326_64 = W*in
   wire signed [9:0] m326_64;
   assign m326_64 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_65 = W*in
   wire signed [9:0] m326_65;
   assign m326_65 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_66 = W*in
   wire signed [9:0] m326_66;
   assign m326_66 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_67 = W*in
   wire signed [9:0] m326_67;
   assign m326_67 =10'b0;

   // m326_68 = W*in
   wire signed [9:0] m326_68;
   assign m326_68 =10'b0;

   // m326_69 = W*in
   wire signed [9:0] m326_69;
   assign m326_69 =10'b0;

   // m326_70 = W*in
   wire signed [9:0] m326_70;
   assign m326_70 =10'b0;

   // m326_71 = W*in
   wire signed [9:0] m326_71;
   assign m326_71 =10'b0;

   // m326_72 = W*in
   wire signed [9:0] m326_72;
   assign m326_72 ={ {3{in326[5]}} , in326 , {1{1'b0}} };

   // m326_73 = W*in
   wire signed [9:0] m326_73;
   assign m326_73 =10'b0;

   // m326_74 = W*in
   wire signed [9:0] m326_74;
   assign m326_74 =10'b0;

   // m326_75 = W*in
   wire signed [9:0] m326_75;
   assign m326_75 =10'b0;

   // m326_76 = W*in
   wire signed [9:0] m326_76;
   assign m326_76 ={ {4{in326[5]}} , in326[5:0] };

   // m326_77 = W*in
   wire signed [9:0] m326_77;
   assign m326_77 ={ {4{in326[5]}} , in326[5:0] };

   // m326_78 = W*in
   wire signed [9:0] m326_78;
   assign m326_78 =10'b0;

   // m326_79 = W*in
   wire signed [9:0] m326_79;
   assign m326_79 =10'b0;

   // m326_80 = W*in
   wire signed [9:0] m326_80;
   assign m326_80 =10'b0;

   // m326_81 = W*in
   wire signed [9:0] m326_81;
   assign m326_81 =10'b0;

   // m326_82 = W*in
   wire signed [9:0] m326_82;
   assign m326_82 =10'b0;

   // m326_83 = W*in
   wire signed [9:0] m326_83;
   assign m326_83 ={ {4{in326[5]}} , in326[5:0] };

   // m326_84 = W*in
   wire signed [9:0] m326_84;
   assign m326_84 ={ {3{in326[5]}} , in326 , {1{1'b0}} };

   // m326_85 = W*in
   wire signed [9:0] m326_85;
   assign m326_85 =10'b0;

   // m326_86 = W*in
   wire signed [9:0] m326_86;
   assign m326_86 =10'b0;

   // m326_87 = W*in
   wire signed [9:0] m326_87;
   assign m326_87 ={ {4{in326[5]}} , in326[5:0] };

   // m326_88 = W*in
   wire signed [9:0] m326_88;
   assign m326_88 ={ {4{in326[5]}} , in326[5:0] };

   // m326_89 = W*in
   wire signed [9:0] m326_89;
   assign m326_89 =10'b0;

   // m326_90 = W*in
   wire signed [9:0] m326_90;
   assign m326_90 ={ {4{in326[5]}} , in326[5:0] };

   // m326_91 = W*in
   wire signed [9:0] m326_91;
   assign m326_91 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_92 = W*in
   wire signed [9:0] m326_92;
   assign m326_92 ={ {4{in326[5]}} , in326[5:0] };

   // m326_93 = W*in
   wire signed [9:0] m326_93;
   assign m326_93 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_94 = W*in
   wire signed [9:0] m326_94;
   assign m326_94 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_95 = W*in
   wire signed [9:0] m326_95;
   assign m326_95 ={ {4{in326[5]}} , in326[5:0] };

   // m326_96 = W*in
   wire signed [9:0] m326_96;
   assign m326_96 =10'b0;

   // m326_97 = W*in
   wire signed [9:0] m326_97;
   assign m326_97 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_98 = W*in
   wire signed [9:0] m326_98;
   assign m326_98 =10'b0;

   // m326_99 = W*in
   wire signed [9:0] m326_99;
   assign m326_99 =10'b0;

   // m326_100 = W*in
   wire signed [9:0] m326_100;
   assign m326_100 =10'b0;

   // m326_101 = W*in
   wire signed [9:0] m326_101;
   assign m326_101 =10'b0;

   // m326_102 = W*in
   wire signed [9:0] m326_102;
   assign m326_102 =10'b0;

   // m326_103 = W*in
   wire signed [9:0] m326_103;
   assign m326_103 =10'b0;

   // m326_104 = W*in
   wire signed [9:0] m326_104;
   assign m326_104 =10'b0;

   // m326_105 = W*in
   wire signed [9:0] m326_105;
   assign m326_105 =10'b0;

   // m326_106 = W*in
   wire signed [9:0] m326_106;
   assign m326_106 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_107 = W*in
   wire signed [9:0] m326_107;
   assign m326_107 ={ {4{in326[5]}} , in326[5:0] };

   // m326_108 = W*in
   wire signed [9:0] m326_108;
   assign m326_108 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_109 = W*in
   wire signed [9:0] m326_109;
   assign m326_109 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_110 = W*in
   wire signed [9:0] m326_110;
   assign m326_110 =10'b0;

   // m326_111 = W*in
   wire signed [9:0] m326_111;
   assign m326_111 ={ {4{in326[5]}} , in326[5:0] };

   // m326_112 = W*in
   wire signed [9:0] m326_112;
   assign m326_112 ={ {4{neg326[5]}} , neg326[5:0] };

   // m326_113 = W*in
   wire signed [9:0] m326_113;
   assign m326_113 ={ {4{in326[5]}} , in326[5:0] };

   // m326_114 = W*in
   wire signed [9:0] m326_114;
   assign m326_114 ={ {5{neg326[5]}} , neg326[5:1] };

   // m326_115 = W*in
   wire signed [9:0] m326_115;
   assign m326_115 =10'b0;

   // m326_116 = W*in
   wire signed [9:0] m326_116;
   assign m326_116 =10'b0;

   // m326_117 = W*in
   wire signed [9:0] m326_117;
   assign m326_117 ={ {4{neg326[5]}} , neg326[5:0] };

   // m327_1 = W*in
   wire signed [9:0] m327_1;
   assign m327_1 =10'b0;

   // m327_2 = W*in
   wire signed [9:0] m327_2;
   assign m327_2 =10'b0;

   // m327_3 = W*in
   wire signed [9:0] m327_3;
   assign m327_3 =10'b0;

   // m327_4 = W*in
   wire signed [9:0] m327_4;
   assign m327_4 =10'b0;

   // m327_5 = W*in
   wire signed [9:0] m327_5;
   assign m327_5 =10'b0;

   // m327_6 = W*in
   wire signed [9:0] m327_6;
   assign m327_6 =10'b0;

   // m327_7 = W*in
   wire signed [9:0] m327_7;
   assign m327_7 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_8 = W*in
   wire signed [9:0] m327_8;
   assign m327_8 =10'b0;

   // m327_9 = W*in
   wire signed [9:0] m327_9;
   assign m327_9 =10'b0;

   // m327_10 = W*in
   wire signed [9:0] m327_10;
   assign m327_10 =10'b0;

   // m327_11 = W*in
   wire signed [9:0] m327_11;
   assign m327_11 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_12 = W*in
   wire signed [9:0] m327_12;
   assign m327_12 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_13 = W*in
   wire signed [9:0] m327_13;
   assign m327_13 =10'b0;

   // m327_14 = W*in
   wire signed [9:0] m327_14;
   assign m327_14 =10'b0;

   // m327_15 = W*in
   wire signed [9:0] m327_15;
   assign m327_15 =10'b0;

   // m327_16 = W*in
   wire signed [9:0] m327_16;
   assign m327_16 ={ {4{in327[5]}} , in327[5:0] };

   // m327_17 = W*in
   wire signed [9:0] m327_17;
   assign m327_17 =10'b0;

   // m327_18 = W*in
   wire signed [9:0] m327_18;
   assign m327_18 =10'b0;

   // m327_19 = W*in
   wire signed [9:0] m327_19;
   assign m327_19 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_20 = W*in
   wire signed [9:0] m327_20;
   assign m327_20 ={ {4{in327[5]}} , in327[5:0] };

   // m327_21 = W*in
   wire signed [9:0] m327_21;
   assign m327_21 ={ {5{in327[5]}} , in327[5:1] };

   // m327_22 = W*in
   wire signed [9:0] m327_22;
   assign m327_22 =10'b0;

   // m327_23 = W*in
   wire signed [9:0] m327_23;
   assign m327_23 =10'b0;

   // m327_24 = W*in
   wire signed [9:0] m327_24;
   assign m327_24 =10'b0;

   // m327_25 = W*in
   wire signed [9:0] m327_25;
   assign m327_25 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_26 = W*in
   wire signed [9:0] m327_26;
   assign m327_26 =10'b0;

   // m327_27 = W*in
   wire signed [9:0] m327_27;
   assign m327_27 =10'b0;

   // m327_28 = W*in
   wire signed [9:0] m327_28;
   assign m327_28 =10'b0;

   // m327_29 = W*in
   wire signed [9:0] m327_29;
   assign m327_29 =10'b0;

   // m327_30 = W*in
   wire signed [9:0] m327_30;
   assign m327_30 =10'b0;

   // m327_31 = W*in
   wire signed [9:0] m327_31;
   assign m327_31 =10'b0;

   // m327_32 = W*in
   wire signed [9:0] m327_32;
   assign m327_32 =10'b0;

   // m327_33 = W*in
   wire signed [9:0] m327_33;
   assign m327_33 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_34 = W*in
   wire signed [9:0] m327_34;
   assign m327_34 ={ {4{in327[5]}} , in327[5:0] };

   // m327_35 = W*in
   wire signed [9:0] m327_35;
   assign m327_35 =10'b0;

   // m327_36 = W*in
   wire signed [9:0] m327_36;
   assign m327_36 =10'b0;

   // m327_37 = W*in
   wire signed [9:0] m327_37;
   assign m327_37 =10'b0;

   // m327_38 = W*in
   wire signed [9:0] m327_38;
   assign m327_38 =10'b0;

   // m327_39 = W*in
   wire signed [9:0] m327_39;
   assign m327_39 =10'b0;

   // m327_40 = W*in
   wire signed [9:0] m327_40;
   assign m327_40 =10'b0;

   // m327_41 = W*in
   wire signed [9:0] m327_41;
   assign m327_41 =10'b0;

   // m327_42 = W*in
   wire signed [9:0] m327_42;
   assign m327_42 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_43 = W*in
   wire signed [9:0] m327_43;
   assign m327_43 =10'b0;

   // m327_44 = W*in
   wire signed [9:0] m327_44;
   assign m327_44 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_45 = W*in
   wire signed [9:0] m327_45;
   assign m327_45 =10'b0;

   // m327_46 = W*in
   wire signed [9:0] m327_46;
   assign m327_46 =10'b0;

   // m327_47 = W*in
   wire signed [9:0] m327_47;
   assign m327_47 =10'b0;

   // m327_48 = W*in
   wire signed [9:0] m327_48;
   assign m327_48 =10'b0;

   // m327_49 = W*in
   wire signed [9:0] m327_49;
   assign m327_49 =10'b0;

   // m327_50 = W*in
   wire signed [9:0] m327_50;
   assign m327_50 =10'b0;

   // m327_51 = W*in
   wire signed [9:0] m327_51;
   assign m327_51 =10'b0;

   // m327_52 = W*in
   wire signed [9:0] m327_52;
   assign m327_52 =10'b0;

   // m327_53 = W*in
   wire signed [9:0] m327_53;
   assign m327_53 =10'b0;

   // m327_54 = W*in
   wire signed [9:0] m327_54;
   assign m327_54 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_55 = W*in
   wire signed [9:0] m327_55;
   assign m327_55 =10'b0;

   // m327_56 = W*in
   wire signed [9:0] m327_56;
   assign m327_56 =10'b0;

   // m327_57 = W*in
   wire signed [9:0] m327_57;
   assign m327_57 =10'b0;

   // m327_58 = W*in
   wire signed [9:0] m327_58;
   assign m327_58 =10'b0;

   // m327_59 = W*in
   wire signed [9:0] m327_59;
   assign m327_59 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_60 = W*in
   wire signed [9:0] m327_60;
   assign m327_60 =10'b0;

   // m327_61 = W*in
   wire signed [9:0] m327_61;
   assign m327_61 =10'b0;

   // m327_62 = W*in
   wire signed [9:0] m327_62;
   assign m327_62 =10'b0;

   // m327_63 = W*in
   wire signed [9:0] m327_63;
   assign m327_63 =10'b0;

   // m327_64 = W*in
   wire signed [9:0] m327_64;
   assign m327_64 =10'b0;

   // m327_65 = W*in
   wire signed [9:0] m327_65;
   assign m327_65 =10'b0;

   // m327_66 = W*in
   wire signed [9:0] m327_66;
   assign m327_66 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_67 = W*in
   wire signed [9:0] m327_67;
   assign m327_67 =10'b0;

   // m327_68 = W*in
   wire signed [9:0] m327_68;
   assign m327_68 =10'b0;

   // m327_69 = W*in
   wire signed [9:0] m327_69;
   assign m327_69 ={ {5{in327[5]}} , in327[5:1] };

   // m327_70 = W*in
   wire signed [9:0] m327_70;
   assign m327_70 ={ {4{in327[5]}} , in327[5:0] };

   // m327_71 = W*in
   wire signed [9:0] m327_71;
   assign m327_71 =10'b0;

   // m327_72 = W*in
   wire signed [9:0] m327_72;
   assign m327_72 ={ {3{in327[5]}} , in327 , {1{1'b0}} };

   // m327_73 = W*in
   wire signed [9:0] m327_73;
   assign m327_73 =10'b0;

   // m327_74 = W*in
   wire signed [9:0] m327_74;
   assign m327_74 ={ {5{in327[5]}} , in327[5:1] };

   // m327_75 = W*in
   wire signed [9:0] m327_75;
   assign m327_75 =10'b0;

   // m327_76 = W*in
   wire signed [9:0] m327_76;
   assign m327_76 ={ {4{in327[5]}} , in327[5:0] };

   // m327_77 = W*in
   wire signed [9:0] m327_77;
   assign m327_77 =10'b0;

   // m327_78 = W*in
   wire signed [9:0] m327_78;
   assign m327_78 =10'b0;

   // m327_79 = W*in
   wire signed [9:0] m327_79;
   assign m327_79 =10'b0;

   // m327_80 = W*in
   wire signed [9:0] m327_80;
   assign m327_80 =10'b0;

   // m327_81 = W*in
   wire signed [9:0] m327_81;
   assign m327_81 =10'b0;

   // m327_82 = W*in
   wire signed [9:0] m327_82;
   assign m327_82 =10'b0;

   // m327_83 = W*in
   wire signed [9:0] m327_83;
   assign m327_83 =10'b0;

   // m327_84 = W*in
   wire signed [9:0] m327_84;
   assign m327_84 ={ {4{in327[5]}} , in327[5:0] };

   // m327_85 = W*in
   wire signed [9:0] m327_85;
   assign m327_85 =10'b0;

   // m327_86 = W*in
   wire signed [9:0] m327_86;
   assign m327_86 =10'b0;

   // m327_87 = W*in
   wire signed [9:0] m327_87;
   assign m327_87 ={ {4{in327[5]}} , in327[5:0] };

   // m327_88 = W*in
   wire signed [9:0] m327_88;
   assign m327_88 ={ {4{in327[5]}} , in327[5:0] };

   // m327_89 = W*in
   wire signed [9:0] m327_89;
   assign m327_89 =10'b0;

   // m327_90 = W*in
   wire signed [9:0] m327_90;
   assign m327_90 ={ {4{in327[5]}} , in327[5:0] };

   // m327_91 = W*in
   wire signed [9:0] m327_91;
   assign m327_91 ={ {3{neg327[5]}} , neg327 , {1{1'b0}} };

   // m327_92 = W*in
   wire signed [9:0] m327_92;
   assign m327_92 ={ {4{in327[5]}} , in327[5:0] };

   // m327_93 = W*in
   wire signed [9:0] m327_93;
   assign m327_93 =10'b0;

   // m327_94 = W*in
   wire signed [9:0] m327_94;
   assign m327_94 =10'b0;

   // m327_95 = W*in
   wire signed [9:0] m327_95;
   assign m327_95 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_96 = W*in
   wire signed [9:0] m327_96;
   assign m327_96 =10'b0;

   // m327_97 = W*in
   wire signed [9:0] m327_97;
   assign m327_97 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_98 = W*in
   wire signed [9:0] m327_98;
   assign m327_98 =10'b0;

   // m327_99 = W*in
   wire signed [9:0] m327_99;
   assign m327_99 ={ {4{in327[5]}} , in327[5:0] };

   // m327_100 = W*in
   wire signed [9:0] m327_100;
   assign m327_100 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_101 = W*in
   wire signed [9:0] m327_101;
   assign m327_101 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_102 = W*in
   wire signed [9:0] m327_102;
   assign m327_102 =10'b0;

   // m327_103 = W*in
   wire signed [9:0] m327_103;
   assign m327_103 =10'b0;

   // m327_104 = W*in
   wire signed [9:0] m327_104;
   assign m327_104 =10'b0;

   // m327_105 = W*in
   wire signed [9:0] m327_105;
   assign m327_105 =10'b0;

   // m327_106 = W*in
   wire signed [9:0] m327_106;
   assign m327_106 =10'b0;

   // m327_107 = W*in
   wire signed [9:0] m327_107;
   assign m327_107 =10'b0;

   // m327_108 = W*in
   wire signed [9:0] m327_108;
   assign m327_108 =10'b0;

   // m327_109 = W*in
   wire signed [9:0] m327_109;
   assign m327_109 =10'b0;

   // m327_110 = W*in
   wire signed [9:0] m327_110;
   assign m327_110 =10'b0;

   // m327_111 = W*in
   wire signed [9:0] m327_111;
   assign m327_111 =10'b0;

   // m327_112 = W*in
   wire signed [9:0] m327_112;
   assign m327_112 ={ {4{neg327[5]}} , neg327[5:0] };

   // m327_113 = W*in
   wire signed [9:0] m327_113;
   assign m327_113 =10'b0;

   // m327_114 = W*in
   wire signed [9:0] m327_114;
   assign m327_114 ={ {5{in327[5]}} , in327[5:1] };

   // m327_115 = W*in
   wire signed [9:0] m327_115;
   assign m327_115 ={ {5{in327[5]}} , in327[5:1] };

   // m327_116 = W*in
   wire signed [9:0] m327_116;
   assign m327_116 =10'b0;

   // m327_117 = W*in
   wire signed [9:0] m327_117;
   assign m327_117 =10'b0;

   // m328_1 = W*in
   wire signed [9:0] m328_1;
   assign m328_1 =10'b0;

   // m328_2 = W*in
   wire signed [9:0] m328_2;
   assign m328_2 =10'b0;

   // m328_3 = W*in
   wire signed [9:0] m328_3;
   assign m328_3 =10'b0;

   // m328_4 = W*in
   wire signed [9:0] m328_4;
   assign m328_4 =10'b0;

   // m328_5 = W*in
   wire signed [9:0] m328_5;
   assign m328_5 =10'b0;

   // m328_6 = W*in
   wire signed [9:0] m328_6;
   assign m328_6 =10'b0;

   // m328_7 = W*in
   wire signed [9:0] m328_7;
   assign m328_7 =10'b0;

   // m328_8 = W*in
   wire signed [9:0] m328_8;
   assign m328_8 =10'b0;

   // m328_9 = W*in
   wire signed [9:0] m328_9;
   assign m328_9 =10'b0;

   // m328_10 = W*in
   wire signed [9:0] m328_10;
   assign m328_10 =10'b0;

   // m328_11 = W*in
   wire signed [9:0] m328_11;
   assign m328_11 =10'b0;

   // m328_12 = W*in
   wire signed [9:0] m328_12;
   assign m328_12 =10'b0;

   // m328_13 = W*in
   wire signed [9:0] m328_13;
   assign m328_13 =10'b0;

   // m328_14 = W*in
   wire signed [9:0] m328_14;
   assign m328_14 =10'b0;

   // m328_15 = W*in
   wire signed [9:0] m328_15;
   assign m328_15 =10'b0;

   // m328_16 = W*in
   wire signed [9:0] m328_16;
   assign m328_16 ={ {5{in328[5]}} , in328[5:1] };

   // m328_17 = W*in
   wire signed [9:0] m328_17;
   assign m328_17 =10'b0;

   // m328_18 = W*in
   wire signed [9:0] m328_18;
   assign m328_18 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_19 = W*in
   wire signed [9:0] m328_19;
   assign m328_19 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_20 = W*in
   wire signed [9:0] m328_20;
   assign m328_20 ={ {5{in328[5]}} , in328[5:1] };

   // m328_21 = W*in
   wire signed [9:0] m328_21;
   assign m328_21 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_22 = W*in
   wire signed [9:0] m328_22;
   assign m328_22 =10'b0;

   // m328_23 = W*in
   wire signed [9:0] m328_23;
   assign m328_23 =10'b0;

   // m328_24 = W*in
   wire signed [9:0] m328_24;
   assign m328_24 =10'b0;

   // m328_25 = W*in
   wire signed [9:0] m328_25;
   assign m328_25 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_26 = W*in
   wire signed [9:0] m328_26;
   assign m328_26 =10'b0;

   // m328_27 = W*in
   wire signed [9:0] m328_27;
   assign m328_27 =10'b0;

   // m328_28 = W*in
   wire signed [9:0] m328_28;
   assign m328_28 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_29 = W*in
   wire signed [9:0] m328_29;
   assign m328_29 =10'b0;

   // m328_30 = W*in
   wire signed [9:0] m328_30;
   assign m328_30 =10'b0;

   // m328_31 = W*in
   wire signed [9:0] m328_31;
   assign m328_31 =10'b0;

   // m328_32 = W*in
   wire signed [9:0] m328_32;
   assign m328_32 =10'b0;

   // m328_33 = W*in
   wire signed [9:0] m328_33;
   assign m328_33 =10'b0;

   // m328_34 = W*in
   wire signed [9:0] m328_34;
   assign m328_34 ={ {5{in328[5]}} , in328[5:1] };

   // m328_35 = W*in
   wire signed [9:0] m328_35;
   assign m328_35 ={ {5{in328[5]}} , in328[5:1] };

   // m328_36 = W*in
   wire signed [9:0] m328_36;
   assign m328_36 ={ {4{in328[5]}} , in328[5:0] };

   // m328_37 = W*in
   wire signed [9:0] m328_37;
   assign m328_37 =10'b0;

   // m328_38 = W*in
   wire signed [9:0] m328_38;
   assign m328_38 =10'b0;

   // m328_39 = W*in
   wire signed [9:0] m328_39;
   assign m328_39 =10'b0;

   // m328_40 = W*in
   wire signed [9:0] m328_40;
   assign m328_40 =10'b0;

   // m328_41 = W*in
   wire signed [9:0] m328_41;
   assign m328_41 =10'b0;

   // m328_42 = W*in
   wire signed [9:0] m328_42;
   assign m328_42 =10'b0;

   // m328_43 = W*in
   wire signed [9:0] m328_43;
   assign m328_43 =10'b0;

   // m328_44 = W*in
   wire signed [9:0] m328_44;
   assign m328_44 ={ {4{neg328[5]}} , neg328[5:0] };

   // m328_45 = W*in
   wire signed [9:0] m328_45;
   assign m328_45 =10'b0;

   // m328_46 = W*in
   wire signed [9:0] m328_46;
   assign m328_46 =10'b0;

   // m328_47 = W*in
   wire signed [9:0] m328_47;
   assign m328_47 =10'b0;

   // m328_48 = W*in
   wire signed [9:0] m328_48;
   assign m328_48 =10'b0;

   // m328_49 = W*in
   wire signed [9:0] m328_49;
   assign m328_49 =10'b0;

   // m328_50 = W*in
   wire signed [9:0] m328_50;
   assign m328_50 =10'b0;

   // m328_51 = W*in
   wire signed [9:0] m328_51;
   assign m328_51 =10'b0;

   // m328_52 = W*in
   wire signed [9:0] m328_52;
   assign m328_52 =10'b0;

   // m328_53 = W*in
   wire signed [9:0] m328_53;
   assign m328_53 =10'b0;

   // m328_54 = W*in
   wire signed [9:0] m328_54;
   assign m328_54 =10'b0;

   // m328_55 = W*in
   wire signed [9:0] m328_55;
   assign m328_55 =10'b0;

   // m328_56 = W*in
   wire signed [9:0] m328_56;
   assign m328_56 =10'b0;

   // m328_57 = W*in
   wire signed [9:0] m328_57;
   assign m328_57 =10'b0;

   // m328_58 = W*in
   wire signed [9:0] m328_58;
   assign m328_58 =10'b0;

   // m328_59 = W*in
   wire signed [9:0] m328_59;
   assign m328_59 =10'b0;

   // m328_60 = W*in
   wire signed [9:0] m328_60;
   assign m328_60 =10'b0;

   // m328_61 = W*in
   wire signed [9:0] m328_61;
   assign m328_61 =10'b0;

   // m328_62 = W*in
   wire signed [9:0] m328_62;
   assign m328_62 =10'b0;

   // m328_63 = W*in
   wire signed [9:0] m328_63;
   assign m328_63 =10'b0;

   // m328_64 = W*in
   wire signed [9:0] m328_64;
   assign m328_64 ={ {5{in328[5]}} , in328[5:1] };

   // m328_65 = W*in
   wire signed [9:0] m328_65;
   assign m328_65 =10'b0;

   // m328_66 = W*in
   wire signed [9:0] m328_66;
   assign m328_66 ={ {4{neg328[5]}} , neg328[5:0] };

   // m328_67 = W*in
   wire signed [9:0] m328_67;
   assign m328_67 =10'b0;

   // m328_68 = W*in
   wire signed [9:0] m328_68;
   assign m328_68 =10'b0;

   // m328_69 = W*in
   wire signed [9:0] m328_69;
   assign m328_69 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_70 = W*in
   wire signed [9:0] m328_70;
   assign m328_70 ={ {4{neg328[5]}} , neg328[5:0] };

   // m328_71 = W*in
   wire signed [9:0] m328_71;
   assign m328_71 =10'b0;

   // m328_72 = W*in
   wire signed [9:0] m328_72;
   assign m328_72 =10'b0;

   // m328_73 = W*in
   wire signed [9:0] m328_73;
   assign m328_73 ={ {5{in328[5]}} , in328[5:1] };

   // m328_74 = W*in
   wire signed [9:0] m328_74;
   assign m328_74 ={ {5{neg328[5]}} , neg328[5:1] };

   // m328_75 = W*in
   wire signed [9:0] m328_75;
   assign m328_75 =10'b0;

   // m328_76 = W*in
   wire signed [9:0] m328_76;
   assign m328_76 =10'b0;

   // m328_77 = W*in
   wire signed [9:0] m328_77;
   assign m328_77 =10'b0;

   // m328_78 = W*in
   wire signed [9:0] m328_78;
   assign m328_78 =10'b0;

   // m328_79 = W*in
   wire signed [9:0] m328_79;
   assign m328_79 =10'b0;

   // m328_80 = W*in
   wire signed [9:0] m328_80;
   assign m328_80 =10'b0;

   // m328_81 = W*in
   wire signed [9:0] m328_81;
   assign m328_81 ={ {5{in328[5]}} , in328[5:1] };

   // m328_82 = W*in
   wire signed [9:0] m328_82;
   assign m328_82 =10'b0;

   // m328_83 = W*in
   wire signed [9:0] m328_83;
   assign m328_83 =10'b0;

   // m328_84 = W*in
   wire signed [9:0] m328_84;
   assign m328_84 =10'b0;

   // m328_85 = W*in
   wire signed [9:0] m328_85;
   assign m328_85 =10'b0;

   // m328_86 = W*in
   wire signed [9:0] m328_86;
   assign m328_86 =10'b0;

   // m328_87 = W*in
   wire signed [9:0] m328_87;
   assign m328_87 =10'b0;

   // m328_88 = W*in
   wire signed [9:0] m328_88;
   assign m328_88 =10'b0;

   // m328_89 = W*in
   wire signed [9:0] m328_89;
   assign m328_89 =10'b0;

   // m328_90 = W*in
   wire signed [9:0] m328_90;
   assign m328_90 =10'b0;

   // m328_91 = W*in
   wire signed [9:0] m328_91;
   assign m328_91 ={ {4{neg328[5]}} , neg328[5:0] };

   // m328_92 = W*in
   wire signed [9:0] m328_92;
   assign m328_92 =10'b0;

   // m328_93 = W*in
   wire signed [9:0] m328_93;
   assign m328_93 =10'b0;

   // m328_94 = W*in
   wire signed [9:0] m328_94;
   assign m328_94 =10'b0;

   // m328_95 = W*in
   wire signed [9:0] m328_95;
   assign m328_95 =10'b0;

   // m328_96 = W*in
   wire signed [9:0] m328_96;
   assign m328_96 =10'b0;

   // m328_97 = W*in
   wire signed [9:0] m328_97;
   assign m328_97 ={ {4{neg328[5]}} , neg328[5:0] };

   // m328_98 = W*in
   wire signed [9:0] m328_98;
   assign m328_98 =10'b0;

   // m328_99 = W*in
   wire signed [9:0] m328_99;
   assign m328_99 =10'b0;

   // m328_100 = W*in
   wire signed [9:0] m328_100;
   assign m328_100 =10'b0;

   // m328_101 = W*in
   wire signed [9:0] m328_101;
   assign m328_101 =10'b0;

   // m328_102 = W*in
   wire signed [9:0] m328_102;
   assign m328_102 =10'b0;

   // m328_103 = W*in
   wire signed [9:0] m328_103;
   assign m328_103 =10'b0;

   // m328_104 = W*in
   wire signed [9:0] m328_104;
   assign m328_104 =10'b0;

   // m328_105 = W*in
   wire signed [9:0] m328_105;
   assign m328_105 =10'b0;

   // m328_106 = W*in
   wire signed [9:0] m328_106;
   assign m328_106 =10'b0;

   // m328_107 = W*in
   wire signed [9:0] m328_107;
   assign m328_107 =10'b0;

   // m328_108 = W*in
   wire signed [9:0] m328_108;
   assign m328_108 =10'b0;

   // m328_109 = W*in
   wire signed [9:0] m328_109;
   assign m328_109 =10'b0;

   // m328_110 = W*in
   wire signed [9:0] m328_110;
   assign m328_110 =10'b0;

   // m328_111 = W*in
   wire signed [9:0] m328_111;
   assign m328_111 =10'b0;

   // m328_112 = W*in
   wire signed [9:0] m328_112;
   assign m328_112 =10'b0;

   // m328_113 = W*in
   wire signed [9:0] m328_113;
   assign m328_113 =10'b0;

   // m328_114 = W*in
   wire signed [9:0] m328_114;
   assign m328_114 ={ {5{in328[5]}} , in328[5:1] };

   // m328_115 = W*in
   wire signed [9:0] m328_115;
   assign m328_115 ={ {5{in328[5]}} , in328[5:1] };

   // m328_116 = W*in
   wire signed [9:0] m328_116;
   assign m328_116 =10'b0;

   // m328_117 = W*in
   wire signed [9:0] m328_117;
   assign m328_117 =10'b0;

   // m329_1 = W*in
   wire signed [9:0] m329_1;
   assign m329_1 =10'b0;

   // m329_2 = W*in
   wire signed [9:0] m329_2;
   assign m329_2 =10'b0;

   // m329_3 = W*in
   wire signed [9:0] m329_3;
   assign m329_3 =10'b0;

   // m329_4 = W*in
   wire signed [9:0] m329_4;
   assign m329_4 =10'b0;

   // m329_5 = W*in
   wire signed [9:0] m329_5;
   assign m329_5 =10'b0;

   // m329_6 = W*in
   wire signed [9:0] m329_6;
   assign m329_6 =10'b0;

   // m329_7 = W*in
   wire signed [9:0] m329_7;
   assign m329_7 =10'b0;

   // m329_8 = W*in
   wire signed [9:0] m329_8;
   assign m329_8 =10'b0;

   // m329_9 = W*in
   wire signed [9:0] m329_9;
   assign m329_9 =10'b0;

   // m329_10 = W*in
   wire signed [9:0] m329_10;
   assign m329_10 =10'b0;

   // m329_11 = W*in
   wire signed [9:0] m329_11;
   assign m329_11 =10'b0;

   // m329_12 = W*in
   wire signed [9:0] m329_12;
   assign m329_12 =10'b0;

   // m329_13 = W*in
   wire signed [9:0] m329_13;
   assign m329_13 =10'b0;

   // m329_14 = W*in
   wire signed [9:0] m329_14;
   assign m329_14 =10'b0;

   // m329_15 = W*in
   wire signed [9:0] m329_15;
   assign m329_15 =10'b0;

   // m329_16 = W*in
   wire signed [9:0] m329_16;
   assign m329_16 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_17 = W*in
   wire signed [9:0] m329_17;
   assign m329_17 =10'b0;

   // m329_18 = W*in
   wire signed [9:0] m329_18;
   assign m329_18 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_19 = W*in
   wire signed [9:0] m329_19;
   assign m329_19 =10'b0;

   // m329_20 = W*in
   wire signed [9:0] m329_20;
   assign m329_20 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_21 = W*in
   wire signed [9:0] m329_21;
   assign m329_21 =10'b0;

   // m329_22 = W*in
   wire signed [9:0] m329_22;
   assign m329_22 =10'b0;

   // m329_23 = W*in
   wire signed [9:0] m329_23;
   assign m329_23 =10'b0;

   // m329_24 = W*in
   wire signed [9:0] m329_24;
   assign m329_24 =10'b0;

   // m329_25 = W*in
   wire signed [9:0] m329_25;
   assign m329_25 ={ {4{in329[5]}} , in329[5:0] };

   // m329_26 = W*in
   wire signed [9:0] m329_26;
   assign m329_26 =10'b0;

   // m329_27 = W*in
   wire signed [9:0] m329_27;
   assign m329_27 =10'b0;

   // m329_28 = W*in
   wire signed [9:0] m329_28;
   assign m329_28 ={ {5{in329[5]}} , in329[5:1] };

   // m329_29 = W*in
   wire signed [9:0] m329_29;
   assign m329_29 =10'b0;

   // m329_30 = W*in
   wire signed [9:0] m329_30;
   assign m329_30 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_31 = W*in
   wire signed [9:0] m329_31;
   assign m329_31 =10'b0;

   // m329_32 = W*in
   wire signed [9:0] m329_32;
   assign m329_32 =10'b0;

   // m329_33 = W*in
   wire signed [9:0] m329_33;
   assign m329_33 =10'b0;

   // m329_34 = W*in
   wire signed [9:0] m329_34;
   assign m329_34 =10'b0;

   // m329_35 = W*in
   wire signed [9:0] m329_35;
   assign m329_35 =10'b0;

   // m329_36 = W*in
   wire signed [9:0] m329_36;
   assign m329_36 =10'b0;

   // m329_37 = W*in
   wire signed [9:0] m329_37;
   assign m329_37 =10'b0;

   // m329_38 = W*in
   wire signed [9:0] m329_38;
   assign m329_38 =10'b0;

   // m329_39 = W*in
   wire signed [9:0] m329_39;
   assign m329_39 =10'b0;

   // m329_40 = W*in
   wire signed [9:0] m329_40;
   assign m329_40 =10'b0;

   // m329_41 = W*in
   wire signed [9:0] m329_41;
   assign m329_41 =10'b0;

   // m329_42 = W*in
   wire signed [9:0] m329_42;
   assign m329_42 ={ {4{neg329[5]}} , neg329[5:0] };

   // m329_43 = W*in
   wire signed [9:0] m329_43;
   assign m329_43 =10'b0;

   // m329_44 = W*in
   wire signed [9:0] m329_44;
   assign m329_44 =10'b0;

   // m329_45 = W*in
   wire signed [9:0] m329_45;
   assign m329_45 =10'b0;

   // m329_46 = W*in
   wire signed [9:0] m329_46;
   assign m329_46 =10'b0;

   // m329_47 = W*in
   wire signed [9:0] m329_47;
   assign m329_47 =10'b0;

   // m329_48 = W*in
   wire signed [9:0] m329_48;
   assign m329_48 =10'b0;

   // m329_49 = W*in
   wire signed [9:0] m329_49;
   assign m329_49 =10'b0;

   // m329_50 = W*in
   wire signed [9:0] m329_50;
   assign m329_50 =10'b0;

   // m329_51 = W*in
   wire signed [9:0] m329_51;
   assign m329_51 =10'b0;

   // m329_52 = W*in
   wire signed [9:0] m329_52;
   assign m329_52 =10'b0;

   // m329_53 = W*in
   wire signed [9:0] m329_53;
   assign m329_53 =10'b0;

   // m329_54 = W*in
   wire signed [9:0] m329_54;
   assign m329_54 =10'b0;

   // m329_55 = W*in
   wire signed [9:0] m329_55;
   assign m329_55 =10'b0;

   // m329_56 = W*in
   wire signed [9:0] m329_56;
   assign m329_56 =10'b0;

   // m329_57 = W*in
   wire signed [9:0] m329_57;
   assign m329_57 =10'b0;

   // m329_58 = W*in
   wire signed [9:0] m329_58;
   assign m329_58 =10'b0;

   // m329_59 = W*in
   wire signed [9:0] m329_59;
   assign m329_59 ={ {4{in329[5]}} , in329[5:0] };

   // m329_60 = W*in
   wire signed [9:0] m329_60;
   assign m329_60 =10'b0;

   // m329_61 = W*in
   wire signed [9:0] m329_61;
   assign m329_61 =10'b0;

   // m329_62 = W*in
   wire signed [9:0] m329_62;
   assign m329_62 =10'b0;

   // m329_63 = W*in
   wire signed [9:0] m329_63;
   assign m329_63 =10'b0;

   // m329_64 = W*in
   wire signed [9:0] m329_64;
   assign m329_64 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_65 = W*in
   wire signed [9:0] m329_65;
   assign m329_65 =10'b0;

   // m329_66 = W*in
   wire signed [9:0] m329_66;
   assign m329_66 =10'b0;

   // m329_67 = W*in
   wire signed [9:0] m329_67;
   assign m329_67 =10'b0;

   // m329_68 = W*in
   wire signed [9:0] m329_68;
   assign m329_68 =10'b0;

   // m329_69 = W*in
   wire signed [9:0] m329_69;
   assign m329_69 =10'b0;

   // m329_70 = W*in
   wire signed [9:0] m329_70;
   assign m329_70 =10'b0;

   // m329_71 = W*in
   wire signed [9:0] m329_71;
   assign m329_71 =10'b0;

   // m329_72 = W*in
   wire signed [9:0] m329_72;
   assign m329_72 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_73 = W*in
   wire signed [9:0] m329_73;
   assign m329_73 =10'b0;

   // m329_74 = W*in
   wire signed [9:0] m329_74;
   assign m329_74 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_75 = W*in
   wire signed [9:0] m329_75;
   assign m329_75 =10'b0;

   // m329_76 = W*in
   wire signed [9:0] m329_76;
   assign m329_76 =10'b0;

   // m329_77 = W*in
   wire signed [9:0] m329_77;
   assign m329_77 =10'b0;

   // m329_78 = W*in
   wire signed [9:0] m329_78;
   assign m329_78 =10'b0;

   // m329_79 = W*in
   wire signed [9:0] m329_79;
   assign m329_79 =10'b0;

   // m329_80 = W*in
   wire signed [9:0] m329_80;
   assign m329_80 =10'b0;

   // m329_81 = W*in
   wire signed [9:0] m329_81;
   assign m329_81 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_82 = W*in
   wire signed [9:0] m329_82;
   assign m329_82 =10'b0;

   // m329_83 = W*in
   wire signed [9:0] m329_83;
   assign m329_83 =10'b0;

   // m329_84 = W*in
   wire signed [9:0] m329_84;
   assign m329_84 =10'b0;

   // m329_85 = W*in
   wire signed [9:0] m329_85;
   assign m329_85 =10'b0;

   // m329_86 = W*in
   wire signed [9:0] m329_86;
   assign m329_86 =10'b0;

   // m329_87 = W*in
   wire signed [9:0] m329_87;
   assign m329_87 =10'b0;

   // m329_88 = W*in
   wire signed [9:0] m329_88;
   assign m329_88 =10'b0;

   // m329_89 = W*in
   wire signed [9:0] m329_89;
   assign m329_89 =10'b0;

   // m329_90 = W*in
   wire signed [9:0] m329_90;
   assign m329_90 =10'b0;

   // m329_91 = W*in
   wire signed [9:0] m329_91;
   assign m329_91 =10'b0;

   // m329_92 = W*in
   wire signed [9:0] m329_92;
   assign m329_92 =10'b0;

   // m329_93 = W*in
   wire signed [9:0] m329_93;
   assign m329_93 =10'b0;

   // m329_94 = W*in
   wire signed [9:0] m329_94;
   assign m329_94 =10'b0;

   // m329_95 = W*in
   wire signed [9:0] m329_95;
   assign m329_95 =10'b0;

   // m329_96 = W*in
   wire signed [9:0] m329_96;
   assign m329_96 =10'b0;

   // m329_97 = W*in
   wire signed [9:0] m329_97;
   assign m329_97 =10'b0;

   // m329_98 = W*in
   wire signed [9:0] m329_98;
   assign m329_98 =10'b0;

   // m329_99 = W*in
   wire signed [9:0] m329_99;
   assign m329_99 =10'b0;

   // m329_100 = W*in
   wire signed [9:0] m329_100;
   assign m329_100 =10'b0;

   // m329_101 = W*in
   wire signed [9:0] m329_101;
   assign m329_101 =10'b0;

   // m329_102 = W*in
   wire signed [9:0] m329_102;
   assign m329_102 =10'b0;

   // m329_103 = W*in
   wire signed [9:0] m329_103;
   assign m329_103 =10'b0;

   // m329_104 = W*in
   wire signed [9:0] m329_104;
   assign m329_104 =10'b0;

   // m329_105 = W*in
   wire signed [9:0] m329_105;
   assign m329_105 =10'b0;

   // m329_106 = W*in
   wire signed [9:0] m329_106;
   assign m329_106 =10'b0;

   // m329_107 = W*in
   wire signed [9:0] m329_107;
   assign m329_107 =10'b0;

   // m329_108 = W*in
   wire signed [9:0] m329_108;
   assign m329_108 =10'b0;

   // m329_109 = W*in
   wire signed [9:0] m329_109;
   assign m329_109 ={ {5{in329[5]}} , in329[5:1] };

   // m329_110 = W*in
   wire signed [9:0] m329_110;
   assign m329_110 =10'b0;

   // m329_111 = W*in
   wire signed [9:0] m329_111;
   assign m329_111 =10'b0;

   // m329_112 = W*in
   wire signed [9:0] m329_112;
   assign m329_112 =10'b0;

   // m329_113 = W*in
   wire signed [9:0] m329_113;
   assign m329_113 =10'b0;

   // m329_114 = W*in
   wire signed [9:0] m329_114;
   assign m329_114 =10'b0;

   // m329_115 = W*in
   wire signed [9:0] m329_115;
   assign m329_115 ={ {5{neg329[5]}} , neg329[5:1] };

   // m329_116 = W*in
   wire signed [9:0] m329_116;
   assign m329_116 =10'b0;

   // m329_117 = W*in
   wire signed [9:0] m329_117;
   assign m329_117 =10'b0;

   // m330_1 = W*in
   wire signed [9:0] m330_1;
   assign m330_1 ={ {4{in330[5]}} , in330[5:0] };

   // m330_2 = W*in
   wire signed [9:0] m330_2;
   assign m330_2 ={ {4{in330[5]}} , in330[5:0] };

   // m330_3 = W*in
   wire signed [9:0] m330_3;
   assign m330_3 =10'b0;

   // m330_4 = W*in
   wire signed [9:0] m330_4;
   assign m330_4 =10'b0;

   // m330_5 = W*in
   wire signed [9:0] m330_5;
   assign m330_5 =10'b0;

   // m330_6 = W*in
   wire signed [9:0] m330_6;
   assign m330_6 =10'b0;

   // m330_7 = W*in
   wire signed [9:0] m330_7;
   assign m330_7 ={ {4{in330[5]}} , in330[5:0] };

   // m330_8 = W*in
   wire signed [9:0] m330_8;
   assign m330_8 =10'b0;

   // m330_9 = W*in
   wire signed [9:0] m330_9;
   assign m330_9 =10'b0;

   // m330_10 = W*in
   wire signed [9:0] m330_10;
   assign m330_10 =10'b0;

   // m330_11 = W*in
   wire signed [9:0] m330_11;
   assign m330_11 ={ {4{in330[5]}} , in330[5:0] };

   // m330_12 = W*in
   wire signed [9:0] m330_12;
   assign m330_12 =10'b0;

   // m330_13 = W*in
   wire signed [9:0] m330_13;
   assign m330_13 =10'b0;

   // m330_14 = W*in
   wire signed [9:0] m330_14;
   assign m330_14 =10'b0;

   // m330_15 = W*in
   wire signed [9:0] m330_15;
   assign m330_15 =10'b0;

   // m330_16 = W*in
   wire signed [9:0] m330_16;
   assign m330_16 ={ {5{in330[5]}} , in330[5:1] };

   // m330_17 = W*in
   wire signed [9:0] m330_17;
   assign m330_17 ={ {5{in330[5]}} , in330[5:1] };

   // m330_18 = W*in
   wire signed [9:0] m330_18;
   assign m330_18 ={ {5{neg330[5]}} , neg330[5:1] };

   // m330_19 = W*in
   wire signed [9:0] m330_19;
   assign m330_19 =10'b0;

   // m330_20 = W*in
   wire signed [9:0] m330_20;
   assign m330_20 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_21 = W*in
   wire signed [9:0] m330_21;
   assign m330_21 =10'b0;

   // m330_22 = W*in
   wire signed [9:0] m330_22;
   assign m330_22 =10'b0;

   // m330_23 = W*in
   wire signed [9:0] m330_23;
   assign m330_23 =10'b0;

   // m330_24 = W*in
   wire signed [9:0] m330_24;
   assign m330_24 =10'b0;

   // m330_25 = W*in
   wire signed [9:0] m330_25;
   assign m330_25 ={ {4{in330[5]}} , in330[5:0] };

   // m330_26 = W*in
   wire signed [9:0] m330_26;
   assign m330_26 =10'b0;

   // m330_27 = W*in
   wire signed [9:0] m330_27;
   assign m330_27 =10'b0;

   // m330_28 = W*in
   wire signed [9:0] m330_28;
   assign m330_28 =10'b0;

   // m330_29 = W*in
   wire signed [9:0] m330_29;
   assign m330_29 =10'b0;

   // m330_30 = W*in
   wire signed [9:0] m330_30;
   assign m330_30 ={ {5{neg330[5]}} , neg330[5:1] };

   // m330_31 = W*in
   wire signed [9:0] m330_31;
   assign m330_31 =10'b0;

   // m330_32 = W*in
   wire signed [9:0] m330_32;
   assign m330_32 =10'b0;

   // m330_33 = W*in
   wire signed [9:0] m330_33;
   assign m330_33 =10'b0;

   // m330_34 = W*in
   wire signed [9:0] m330_34;
   assign m330_34 =10'b0;

   // m330_35 = W*in
   wire signed [9:0] m330_35;
   assign m330_35 ={ {5{neg330[5]}} , neg330[5:1] };

   // m330_36 = W*in
   wire signed [9:0] m330_36;
   assign m330_36 =10'b0;

   // m330_37 = W*in
   wire signed [9:0] m330_37;
   assign m330_37 =10'b0;

   // m330_38 = W*in
   wire signed [9:0] m330_38;
   assign m330_38 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_39 = W*in
   wire signed [9:0] m330_39;
   assign m330_39 =10'b0;

   // m330_40 = W*in
   wire signed [9:0] m330_40;
   assign m330_40 =10'b0;

   // m330_41 = W*in
   wire signed [9:0] m330_41;
   assign m330_41 =10'b0;

   // m330_42 = W*in
   wire signed [9:0] m330_42;
   assign m330_42 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_43 = W*in
   wire signed [9:0] m330_43;
   assign m330_43 =10'b0;

   // m330_44 = W*in
   wire signed [9:0] m330_44;
   assign m330_44 =10'b0;

   // m330_45 = W*in
   wire signed [9:0] m330_45;
   assign m330_45 =10'b0;

   // m330_46 = W*in
   wire signed [9:0] m330_46;
   assign m330_46 =10'b0;

   // m330_47 = W*in
   wire signed [9:0] m330_47;
   assign m330_47 =10'b0;

   // m330_48 = W*in
   wire signed [9:0] m330_48;
   assign m330_48 =10'b0;

   // m330_49 = W*in
   wire signed [9:0] m330_49;
   assign m330_49 =10'b0;

   // m330_50 = W*in
   wire signed [9:0] m330_50;
   assign m330_50 =10'b0;

   // m330_51 = W*in
   wire signed [9:0] m330_51;
   assign m330_51 =10'b0;

   // m330_52 = W*in
   wire signed [9:0] m330_52;
   assign m330_52 =10'b0;

   // m330_53 = W*in
   wire signed [9:0] m330_53;
   assign m330_53 =10'b0;

   // m330_54 = W*in
   wire signed [9:0] m330_54;
   assign m330_54 =10'b0;

   // m330_55 = W*in
   wire signed [9:0] m330_55;
   assign m330_55 =10'b0;

   // m330_56 = W*in
   wire signed [9:0] m330_56;
   assign m330_56 =10'b0;

   // m330_57 = W*in
   wire signed [9:0] m330_57;
   assign m330_57 =10'b0;

   // m330_58 = W*in
   wire signed [9:0] m330_58;
   assign m330_58 =10'b0;

   // m330_59 = W*in
   wire signed [9:0] m330_59;
   assign m330_59 ={ {4{in330[5]}} , in330[5:0] };

   // m330_60 = W*in
   wire signed [9:0] m330_60;
   assign m330_60 =10'b0;

   // m330_61 = W*in
   wire signed [9:0] m330_61;
   assign m330_61 =10'b0;

   // m330_62 = W*in
   wire signed [9:0] m330_62;
   assign m330_62 =10'b0;

   // m330_63 = W*in
   wire signed [9:0] m330_63;
   assign m330_63 =10'b0;

   // m330_64 = W*in
   wire signed [9:0] m330_64;
   assign m330_64 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_65 = W*in
   wire signed [9:0] m330_65;
   assign m330_65 =10'b0;

   // m330_66 = W*in
   wire signed [9:0] m330_66;
   assign m330_66 =10'b0;

   // m330_67 = W*in
   wire signed [9:0] m330_67;
   assign m330_67 =10'b0;

   // m330_68 = W*in
   wire signed [9:0] m330_68;
   assign m330_68 =10'b0;

   // m330_69 = W*in
   wire signed [9:0] m330_69;
   assign m330_69 =10'b0;

   // m330_70 = W*in
   wire signed [9:0] m330_70;
   assign m330_70 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_71 = W*in
   wire signed [9:0] m330_71;
   assign m330_71 =10'b0;

   // m330_72 = W*in
   wire signed [9:0] m330_72;
   assign m330_72 =10'b0;

   // m330_73 = W*in
   wire signed [9:0] m330_73;
   assign m330_73 ={ {4{in330[5]}} , in330[5:0] };

   // m330_74 = W*in
   wire signed [9:0] m330_74;
   assign m330_74 ={ {5{neg330[5]}} , neg330[5:1] };

   // m330_75 = W*in
   wire signed [9:0] m330_75;
   assign m330_75 =10'b0;

   // m330_76 = W*in
   wire signed [9:0] m330_76;
   assign m330_76 =10'b0;

   // m330_77 = W*in
   wire signed [9:0] m330_77;
   assign m330_77 =10'b0;

   // m330_78 = W*in
   wire signed [9:0] m330_78;
   assign m330_78 =10'b0;

   // m330_79 = W*in
   wire signed [9:0] m330_79;
   assign m330_79 =10'b0;

   // m330_80 = W*in
   wire signed [9:0] m330_80;
   assign m330_80 =10'b0;

   // m330_81 = W*in
   wire signed [9:0] m330_81;
   assign m330_81 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_82 = W*in
   wire signed [9:0] m330_82;
   assign m330_82 =10'b0;

   // m330_83 = W*in
   wire signed [9:0] m330_83;
   assign m330_83 ={ {5{in330[5]}} , in330[5:1] };

   // m330_84 = W*in
   wire signed [9:0] m330_84;
   assign m330_84 ={ {5{in330[5]}} , in330[5:1] };

   // m330_85 = W*in
   wire signed [9:0] m330_85;
   assign m330_85 =10'b0;

   // m330_86 = W*in
   wire signed [9:0] m330_86;
   assign m330_86 =10'b0;

   // m330_87 = W*in
   wire signed [9:0] m330_87;
   assign m330_87 =10'b0;

   // m330_88 = W*in
   wire signed [9:0] m330_88;
   assign m330_88 =10'b0;

   // m330_89 = W*in
   wire signed [9:0] m330_89;
   assign m330_89 =10'b0;

   // m330_90 = W*in
   wire signed [9:0] m330_90;
   assign m330_90 =10'b0;

   // m330_91 = W*in
   wire signed [9:0] m330_91;
   assign m330_91 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_92 = W*in
   wire signed [9:0] m330_92;
   assign m330_92 =10'b0;

   // m330_93 = W*in
   wire signed [9:0] m330_93;
   assign m330_93 =10'b0;

   // m330_94 = W*in
   wire signed [9:0] m330_94;
   assign m330_94 =10'b0;

   // m330_95 = W*in
   wire signed [9:0] m330_95;
   assign m330_95 ={ {4{in330[5]}} , in330[5:0] };

   // m330_96 = W*in
   wire signed [9:0] m330_96;
   assign m330_96 =10'b0;

   // m330_97 = W*in
   wire signed [9:0] m330_97;
   assign m330_97 =10'b0;

   // m330_98 = W*in
   wire signed [9:0] m330_98;
   assign m330_98 =10'b0;

   // m330_99 = W*in
   wire signed [9:0] m330_99;
   assign m330_99 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_100 = W*in
   wire signed [9:0] m330_100;
   assign m330_100 ={ {4{neg330[5]}} , neg330[5:0] };

   // m330_101 = W*in
   wire signed [9:0] m330_101;
   assign m330_101 =10'b0;

   // m330_102 = W*in
   wire signed [9:0] m330_102;
   assign m330_102 =10'b0;

   // m330_103 = W*in
   wire signed [9:0] m330_103;
   assign m330_103 =10'b0;

   // m330_104 = W*in
   wire signed [9:0] m330_104;
   assign m330_104 =10'b0;

   // m330_105 = W*in
   wire signed [9:0] m330_105;
   assign m330_105 =10'b0;

   // m330_106 = W*in
   wire signed [9:0] m330_106;
   assign m330_106 =10'b0;

   // m330_107 = W*in
   wire signed [9:0] m330_107;
   assign m330_107 =10'b0;

   // m330_108 = W*in
   wire signed [9:0] m330_108;
   assign m330_108 =10'b0;

   // m330_109 = W*in
   wire signed [9:0] m330_109;
   assign m330_109 =10'b0;

   // m330_110 = W*in
   wire signed [9:0] m330_110;
   assign m330_110 =10'b0;

   // m330_111 = W*in
   wire signed [9:0] m330_111;
   assign m330_111 =10'b0;

   // m330_112 = W*in
   wire signed [9:0] m330_112;
   assign m330_112 =10'b0;

   // m330_113 = W*in
   wire signed [9:0] m330_113;
   assign m330_113 =10'b0;

   // m330_114 = W*in
   wire signed [9:0] m330_114;
   assign m330_114 =10'b0;

   // m330_115 = W*in
   wire signed [9:0] m330_115;
   assign m330_115 =10'b0;

   // m330_116 = W*in
   wire signed [9:0] m330_116;
   assign m330_116 =10'b0;

   // m330_117 = W*in
   wire signed [9:0] m330_117;
   assign m330_117 =10'b0;

   // m331_1 = W*in
   wire signed [9:0] m331_1;
   assign m331_1 ={ {4{in331[5]}} , in331[5:0] };

   // m331_2 = W*in
   wire signed [9:0] m331_2;
   assign m331_2 ={ {4{in331[5]}} , in331[5:0] };

   // m331_3 = W*in
   wire signed [9:0] m331_3;
   assign m331_3 =10'b0;

   // m331_4 = W*in
   wire signed [9:0] m331_4;
   assign m331_4 =10'b0;

   // m331_5 = W*in
   wire signed [9:0] m331_5;
   assign m331_5 =10'b0;

   // m331_6 = W*in
   wire signed [9:0] m331_6;
   assign m331_6 =10'b0;

   // m331_7 = W*in
   wire signed [9:0] m331_7;
   assign m331_7 =10'b0;

   // m331_8 = W*in
   wire signed [9:0] m331_8;
   assign m331_8 ={ {4{in331[5]}} , in331[5:0] };

   // m331_9 = W*in
   wire signed [9:0] m331_9;
   assign m331_9 =10'b0;

   // m331_10 = W*in
   wire signed [9:0] m331_10;
   assign m331_10 =10'b0;

   // m331_11 = W*in
   wire signed [9:0] m331_11;
   assign m331_11 ={ {5{neg331[5]}} , neg331[5:1] };

   // m331_12 = W*in
   wire signed [9:0] m331_12;
   assign m331_12 =10'b0;

   // m331_13 = W*in
   wire signed [9:0] m331_13;
   assign m331_13 =10'b0;

   // m331_14 = W*in
   wire signed [9:0] m331_14;
   assign m331_14 =10'b0;

   // m331_15 = W*in
   wire signed [9:0] m331_15;
   assign m331_15 ={ {4{in331[5]}} , in331[5:0] };

   // m331_16 = W*in
   wire signed [9:0] m331_16;
   assign m331_16 ={ {4{in331[5]}} , in331[5:0] };

   // m331_17 = W*in
   wire signed [9:0] m331_17;
   assign m331_17 ={ {5{in331[5]}} , in331[5:1] };

   // m331_18 = W*in
   wire signed [9:0] m331_18;
   assign m331_18 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_19 = W*in
   wire signed [9:0] m331_19;
   assign m331_19 =10'b0;

   // m331_20 = W*in
   wire signed [9:0] m331_20;
   assign m331_20 ={ {5{in331[5]}} , in331[5:1] };

   // m331_21 = W*in
   wire signed [9:0] m331_21;
   assign m331_21 ={ {5{neg331[5]}} , neg331[5:1] };

   // m331_22 = W*in
   wire signed [9:0] m331_22;
   assign m331_22 ={ {4{in331[5]}} , in331[5:0] };

   // m331_23 = W*in
   wire signed [9:0] m331_23;
   assign m331_23 =10'b0;

   // m331_24 = W*in
   wire signed [9:0] m331_24;
   assign m331_24 =10'b0;

   // m331_25 = W*in
   wire signed [9:0] m331_25;
   assign m331_25 =10'b0;

   // m331_26 = W*in
   wire signed [9:0] m331_26;
   assign m331_26 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_27 = W*in
   wire signed [9:0] m331_27;
   assign m331_27 =10'b0;

   // m331_28 = W*in
   wire signed [9:0] m331_28;
   assign m331_28 ={ {5{in331[5]}} , in331[5:1] };

   // m331_29 = W*in
   wire signed [9:0] m331_29;
   assign m331_29 =10'b0;

   // m331_30 = W*in
   wire signed [9:0] m331_30;
   assign m331_30 =10'b0;

   // m331_31 = W*in
   wire signed [9:0] m331_31;
   assign m331_31 ={ {4{in331[5]}} , in331[5:0] };

   // m331_32 = W*in
   wire signed [9:0] m331_32;
   assign m331_32 =10'b0;

   // m331_33 = W*in
   wire signed [9:0] m331_33;
   assign m331_33 =10'b0;

   // m331_34 = W*in
   wire signed [9:0] m331_34;
   assign m331_34 ={ {4{in331[5]}} , in331[5:0] };

   // m331_35 = W*in
   wire signed [9:0] m331_35;
   assign m331_35 ={ {5{in331[5]}} , in331[5:1] };

   // m331_36 = W*in
   wire signed [9:0] m331_36;
   assign m331_36 =10'b0;

   // m331_37 = W*in
   wire signed [9:0] m331_37;
   assign m331_37 =10'b0;

   // m331_38 = W*in
   wire signed [9:0] m331_38;
   assign m331_38 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_39 = W*in
   wire signed [9:0] m331_39;
   assign m331_39 =10'b0;

   // m331_40 = W*in
   wire signed [9:0] m331_40;
   assign m331_40 =10'b0;

   // m331_41 = W*in
   wire signed [9:0] m331_41;
   assign m331_41 =10'b0;

   // m331_42 = W*in
   wire signed [9:0] m331_42;
   assign m331_42 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_43 = W*in
   wire signed [9:0] m331_43;
   assign m331_43 =10'b0;

   // m331_44 = W*in
   wire signed [9:0] m331_44;
   assign m331_44 =10'b0;

   // m331_45 = W*in
   wire signed [9:0] m331_45;
   assign m331_45 ={ {4{in331[5]}} , in331[5:0] };

   // m331_46 = W*in
   wire signed [9:0] m331_46;
   assign m331_46 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_47 = W*in
   wire signed [9:0] m331_47;
   assign m331_47 =10'b0;

   // m331_48 = W*in
   wire signed [9:0] m331_48;
   assign m331_48 ={ {4{in331[5]}} , in331[5:0] };

   // m331_49 = W*in
   wire signed [9:0] m331_49;
   assign m331_49 =10'b0;

   // m331_50 = W*in
   wire signed [9:0] m331_50;
   assign m331_50 ={ {4{in331[5]}} , in331[5:0] };

   // m331_51 = W*in
   wire signed [9:0] m331_51;
   assign m331_51 ={ {4{in331[5]}} , in331[5:0] };

   // m331_52 = W*in
   wire signed [9:0] m331_52;
   assign m331_52 ={ {4{in331[5]}} , in331[5:0] };

   // m331_53 = W*in
   wire signed [9:0] m331_53;
   assign m331_53 =10'b0;

   // m331_54 = W*in
   wire signed [9:0] m331_54;
   assign m331_54 =10'b0;

   // m331_55 = W*in
   wire signed [9:0] m331_55;
   assign m331_55 =10'b0;

   // m331_56 = W*in
   wire signed [9:0] m331_56;
   assign m331_56 ={ {4{in331[5]}} , in331[5:0] };

   // m331_57 = W*in
   wire signed [9:0] m331_57;
   assign m331_57 =10'b0;

   // m331_58 = W*in
   wire signed [9:0] m331_58;
   assign m331_58 =10'b0;

   // m331_59 = W*in
   wire signed [9:0] m331_59;
   assign m331_59 =10'b0;

   // m331_60 = W*in
   wire signed [9:0] m331_60;
   assign m331_60 =10'b0;

   // m331_61 = W*in
   wire signed [9:0] m331_61;
   assign m331_61 =10'b0;

   // m331_62 = W*in
   wire signed [9:0] m331_62;
   assign m331_62 =10'b0;

   // m331_63 = W*in
   wire signed [9:0] m331_63;
   assign m331_63 =10'b0;

   // m331_64 = W*in
   wire signed [9:0] m331_64;
   assign m331_64 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_65 = W*in
   wire signed [9:0] m331_65;
   assign m331_65 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_66 = W*in
   wire signed [9:0] m331_66;
   assign m331_66 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_67 = W*in
   wire signed [9:0] m331_67;
   assign m331_67 =10'b0;

   // m331_68 = W*in
   wire signed [9:0] m331_68;
   assign m331_68 ={ {4{in331[5]}} , in331[5:0] };

   // m331_69 = W*in
   wire signed [9:0] m331_69;
   assign m331_69 ={ {4{in331[5]}} , in331[5:0] };

   // m331_70 = W*in
   wire signed [9:0] m331_70;
   assign m331_70 =10'b0;

   // m331_71 = W*in
   wire signed [9:0] m331_71;
   assign m331_71 =10'b0;

   // m331_72 = W*in
   wire signed [9:0] m331_72;
   assign m331_72 =10'b0;

   // m331_73 = W*in
   wire signed [9:0] m331_73;
   assign m331_73 ={ {4{in331[5]}} , in331[5:0] };

   // m331_74 = W*in
   wire signed [9:0] m331_74;
   assign m331_74 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_75 = W*in
   wire signed [9:0] m331_75;
   assign m331_75 =10'b0;

   // m331_76 = W*in
   wire signed [9:0] m331_76;
   assign m331_76 ={ {4{in331[5]}} , in331[5:0] };

   // m331_77 = W*in
   wire signed [9:0] m331_77;
   assign m331_77 =10'b0;

   // m331_78 = W*in
   wire signed [9:0] m331_78;
   assign m331_78 =10'b0;

   // m331_79 = W*in
   wire signed [9:0] m331_79;
   assign m331_79 =10'b0;

   // m331_80 = W*in
   wire signed [9:0] m331_80;
   assign m331_80 =10'b0;

   // m331_81 = W*in
   wire signed [9:0] m331_81;
   assign m331_81 =10'b0;

   // m331_82 = W*in
   wire signed [9:0] m331_82;
   assign m331_82 =10'b0;

   // m331_83 = W*in
   wire signed [9:0] m331_83;
   assign m331_83 ={ {4{in331[5]}} , in331[5:0] };

   // m331_84 = W*in
   wire signed [9:0] m331_84;
   assign m331_84 ={ {4{in331[5]}} , in331[5:0] };

   // m331_85 = W*in
   wire signed [9:0] m331_85;
   assign m331_85 =10'b0;

   // m331_86 = W*in
   wire signed [9:0] m331_86;
   assign m331_86 =10'b0;

   // m331_87 = W*in
   wire signed [9:0] m331_87;
   assign m331_87 =10'b0;

   // m331_88 = W*in
   wire signed [9:0] m331_88;
   assign m331_88 =10'b0;

   // m331_89 = W*in
   wire signed [9:0] m331_89;
   assign m331_89 =10'b0;

   // m331_90 = W*in
   wire signed [9:0] m331_90;
   assign m331_90 ={ {3{in331[5]}} , in331 , {1{1'b0}} };

   // m331_91 = W*in
   wire signed [9:0] m331_91;
   assign m331_91 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_92 = W*in
   wire signed [9:0] m331_92;
   assign m331_92 ={ {4{in331[5]}} , in331[5:0] };

   // m331_93 = W*in
   wire signed [9:0] m331_93;
   assign m331_93 =10'b0;

   // m331_94 = W*in
   wire signed [9:0] m331_94;
   assign m331_94 ={ {3{neg331[5]}} , neg331 , {1{1'b0}} };

   // m331_95 = W*in
   wire signed [9:0] m331_95;
   assign m331_95 =10'b0;

   // m331_96 = W*in
   wire signed [9:0] m331_96;
   assign m331_96 =10'b0;

   // m331_97 = W*in
   wire signed [9:0] m331_97;
   assign m331_97 =10'b0;

   // m331_98 = W*in
   wire signed [9:0] m331_98;
   assign m331_98 =10'b0;

   // m331_99 = W*in
   wire signed [9:0] m331_99;
   assign m331_99 =10'b0;

   // m331_100 = W*in
   wire signed [9:0] m331_100;
   assign m331_100 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_101 = W*in
   wire signed [9:0] m331_101;
   assign m331_101 =10'b0;

   // m331_102 = W*in
   wire signed [9:0] m331_102;
   assign m331_102 ={ {4{in331[5]}} , in331[5:0] };

   // m331_103 = W*in
   wire signed [9:0] m331_103;
   assign m331_103 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_104 = W*in
   wire signed [9:0] m331_104;
   assign m331_104 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_105 = W*in
   wire signed [9:0] m331_105;
   assign m331_105 =10'b0;

   // m331_106 = W*in
   wire signed [9:0] m331_106;
   assign m331_106 =10'b0;

   // m331_107 = W*in
   wire signed [9:0] m331_107;
   assign m331_107 ={ {4{in331[5]}} , in331[5:0] };

   // m331_108 = W*in
   wire signed [9:0] m331_108;
   assign m331_108 =10'b0;

   // m331_109 = W*in
   wire signed [9:0] m331_109;
   assign m331_109 ={ {5{neg331[5]}} , neg331[5:1] };

   // m331_110 = W*in
   wire signed [9:0] m331_110;
   assign m331_110 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_111 = W*in
   wire signed [9:0] m331_111;
   assign m331_111 ={ {4{in331[5]}} , in331[5:0] };

   // m331_112 = W*in
   wire signed [9:0] m331_112;
   assign m331_112 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_113 = W*in
   wire signed [9:0] m331_113;
   assign m331_113 ={ {4{in331[5]}} , in331[5:0] };

   // m331_114 = W*in
   wire signed [9:0] m331_114;
   assign m331_114 =10'b0;

   // m331_115 = W*in
   wire signed [9:0] m331_115;
   assign m331_115 =10'b0;

   // m331_116 = W*in
   wire signed [9:0] m331_116;
   assign m331_116 ={ {4{neg331[5]}} , neg331[5:0] };

   // m331_117 = W*in
   wire signed [9:0] m331_117;
   assign m331_117 =10'b0;

   // m332_1 = W*in
   wire signed [9:0] m332_1;
   assign m332_1 =10'b0;

   // m332_2 = W*in
   wire signed [9:0] m332_2;
   assign m332_2 =10'b0;

   // m332_3 = W*in
   wire signed [9:0] m332_3;
   assign m332_3 =10'b0;

   // m332_4 = W*in
   wire signed [9:0] m332_4;
   assign m332_4 =10'b0;

   // m332_5 = W*in
   wire signed [9:0] m332_5;
   assign m332_5 =10'b0;

   // m332_6 = W*in
   wire signed [9:0] m332_6;
   assign m332_6 =10'b0;

   // m332_7 = W*in
   wire signed [9:0] m332_7;
   assign m332_7 =10'b0;

   // m332_8 = W*in
   wire signed [9:0] m332_8;
   assign m332_8 ={ {4{in332[5]}} , in332[5:0] };

   // m332_9 = W*in
   wire signed [9:0] m332_9;
   assign m332_9 =10'b0;

   // m332_10 = W*in
   wire signed [9:0] m332_10;
   assign m332_10 =10'b0;

   // m332_11 = W*in
   wire signed [9:0] m332_11;
   assign m332_11 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_12 = W*in
   wire signed [9:0] m332_12;
   assign m332_12 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_13 = W*in
   wire signed [9:0] m332_13;
   assign m332_13 =10'b0;

   // m332_14 = W*in
   wire signed [9:0] m332_14;
   assign m332_14 =10'b0;

   // m332_15 = W*in
   wire signed [9:0] m332_15;
   assign m332_15 ={ {4{in332[5]}} , in332[5:0] };

   // m332_16 = W*in
   wire signed [9:0] m332_16;
   assign m332_16 =10'b0;

   // m332_17 = W*in
   wire signed [9:0] m332_17;
   assign m332_17 =10'b0;

   // m332_18 = W*in
   wire signed [9:0] m332_18;
   assign m332_18 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_19 = W*in
   wire signed [9:0] m332_19;
   assign m332_19 =10'b0;

   // m332_20 = W*in
   wire signed [9:0] m332_20;
   assign m332_20 ={ {4{in332[5]}} , in332[5:0] };

   // m332_21 = W*in
   wire signed [9:0] m332_21;
   assign m332_21 ={ {5{in332[5]}} , in332[5:1] };

   // m332_22 = W*in
   wire signed [9:0] m332_22;
   assign m332_22 =10'b0;

   // m332_23 = W*in
   wire signed [9:0] m332_23;
   assign m332_23 ={ {4{in332[5]}} , in332[5:0] };

   // m332_24 = W*in
   wire signed [9:0] m332_24;
   assign m332_24 =10'b0;

   // m332_25 = W*in
   wire signed [9:0] m332_25;
   assign m332_25 =10'b0;

   // m332_26 = W*in
   wire signed [9:0] m332_26;
   assign m332_26 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_27 = W*in
   wire signed [9:0] m332_27;
   assign m332_27 ={ {4{in332[5]}} , in332[5:0] };

   // m332_28 = W*in
   wire signed [9:0] m332_28;
   assign m332_28 =10'b0;

   // m332_29 = W*in
   wire signed [9:0] m332_29;
   assign m332_29 =10'b0;

   // m332_30 = W*in
   wire signed [9:0] m332_30;
   assign m332_30 ={ {5{neg332[5]}} , neg332[5:1] };

   // m332_31 = W*in
   wire signed [9:0] m332_31;
   assign m332_31 ={ {4{in332[5]}} , in332[5:0] };

   // m332_32 = W*in
   wire signed [9:0] m332_32;
   assign m332_32 =10'b0;

   // m332_33 = W*in
   wire signed [9:0] m332_33;
   assign m332_33 =10'b0;

   // m332_34 = W*in
   wire signed [9:0] m332_34;
   assign m332_34 ={ {4{in332[5]}} , in332[5:0] };

   // m332_35 = W*in
   wire signed [9:0] m332_35;
   assign m332_35 ={ {5{in332[5]}} , in332[5:1] };

   // m332_36 = W*in
   wire signed [9:0] m332_36;
   assign m332_36 =10'b0;

   // m332_37 = W*in
   wire signed [9:0] m332_37;
   assign m332_37 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_38 = W*in
   wire signed [9:0] m332_38;
   assign m332_38 =10'b0;

   // m332_39 = W*in
   wire signed [9:0] m332_39;
   assign m332_39 =10'b0;

   // m332_40 = W*in
   wire signed [9:0] m332_40;
   assign m332_40 =10'b0;

   // m332_41 = W*in
   wire signed [9:0] m332_41;
   assign m332_41 =10'b0;

   // m332_42 = W*in
   wire signed [9:0] m332_42;
   assign m332_42 =10'b0;

   // m332_43 = W*in
   wire signed [9:0] m332_43;
   assign m332_43 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_44 = W*in
   wire signed [9:0] m332_44;
   assign m332_44 =10'b0;

   // m332_45 = W*in
   wire signed [9:0] m332_45;
   assign m332_45 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_46 = W*in
   wire signed [9:0] m332_46;
   assign m332_46 =10'b0;

   // m332_47 = W*in
   wire signed [9:0] m332_47;
   assign m332_47 =10'b0;

   // m332_48 = W*in
   wire signed [9:0] m332_48;
   assign m332_48 =10'b0;

   // m332_49 = W*in
   wire signed [9:0] m332_49;
   assign m332_49 =10'b0;

   // m332_50 = W*in
   wire signed [9:0] m332_50;
   assign m332_50 =10'b0;

   // m332_51 = W*in
   wire signed [9:0] m332_51;
   assign m332_51 =10'b0;

   // m332_52 = W*in
   wire signed [9:0] m332_52;
   assign m332_52 =10'b0;

   // m332_53 = W*in
   wire signed [9:0] m332_53;
   assign m332_53 =10'b0;

   // m332_54 = W*in
   wire signed [9:0] m332_54;
   assign m332_54 =10'b0;

   // m332_55 = W*in
   wire signed [9:0] m332_55;
   assign m332_55 =10'b0;

   // m332_56 = W*in
   wire signed [9:0] m332_56;
   assign m332_56 =10'b0;

   // m332_57 = W*in
   wire signed [9:0] m332_57;
   assign m332_57 =10'b0;

   // m332_58 = W*in
   wire signed [9:0] m332_58;
   assign m332_58 =10'b0;

   // m332_59 = W*in
   wire signed [9:0] m332_59;
   assign m332_59 =10'b0;

   // m332_60 = W*in
   wire signed [9:0] m332_60;
   assign m332_60 =10'b0;

   // m332_61 = W*in
   wire signed [9:0] m332_61;
   assign m332_61 =10'b0;

   // m332_62 = W*in
   wire signed [9:0] m332_62;
   assign m332_62 =10'b0;

   // m332_63 = W*in
   wire signed [9:0] m332_63;
   assign m332_63 =10'b0;

   // m332_64 = W*in
   wire signed [9:0] m332_64;
   assign m332_64 =10'b0;

   // m332_65 = W*in
   wire signed [9:0] m332_65;
   assign m332_65 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_66 = W*in
   wire signed [9:0] m332_66;
   assign m332_66 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_67 = W*in
   wire signed [9:0] m332_67;
   assign m332_67 =10'b0;

   // m332_68 = W*in
   wire signed [9:0] m332_68;
   assign m332_68 ={ {4{in332[5]}} , in332[5:0] };

   // m332_69 = W*in
   wire signed [9:0] m332_69;
   assign m332_69 =10'b0;

   // m332_70 = W*in
   wire signed [9:0] m332_70;
   assign m332_70 ={ {5{in332[5]}} , in332[5:1] };

   // m332_71 = W*in
   wire signed [9:0] m332_71;
   assign m332_71 =10'b0;

   // m332_72 = W*in
   wire signed [9:0] m332_72;
   assign m332_72 =10'b0;

   // m332_73 = W*in
   wire signed [9:0] m332_73;
   assign m332_73 ={ {4{in332[5]}} , in332[5:0] };

   // m332_74 = W*in
   wire signed [9:0] m332_74;
   assign m332_74 =10'b0;

   // m332_75 = W*in
   wire signed [9:0] m332_75;
   assign m332_75 =10'b0;

   // m332_76 = W*in
   wire signed [9:0] m332_76;
   assign m332_76 =10'b0;

   // m332_77 = W*in
   wire signed [9:0] m332_77;
   assign m332_77 =10'b0;

   // m332_78 = W*in
   wire signed [9:0] m332_78;
   assign m332_78 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_79 = W*in
   wire signed [9:0] m332_79;
   assign m332_79 =10'b0;

   // m332_80 = W*in
   wire signed [9:0] m332_80;
   assign m332_80 ={ {4{in332[5]}} , in332[5:0] };

   // m332_81 = W*in
   wire signed [9:0] m332_81;
   assign m332_81 ={ {5{neg332[5]}} , neg332[5:1] };

   // m332_82 = W*in
   wire signed [9:0] m332_82;
   assign m332_82 =10'b0;

   // m332_83 = W*in
   wire signed [9:0] m332_83;
   assign m332_83 ={ {5{neg332[5]}} , neg332[5:1] };

   // m332_84 = W*in
   wire signed [9:0] m332_84;
   assign m332_84 ={ {5{neg332[5]}} , neg332[5:1] };

   // m332_85 = W*in
   wire signed [9:0] m332_85;
   assign m332_85 =10'b0;

   // m332_86 = W*in
   wire signed [9:0] m332_86;
   assign m332_86 =10'b0;

   // m332_87 = W*in
   wire signed [9:0] m332_87;
   assign m332_87 =10'b0;

   // m332_88 = W*in
   wire signed [9:0] m332_88;
   assign m332_88 ={ {4{in332[5]}} , in332[5:0] };

   // m332_89 = W*in
   wire signed [9:0] m332_89;
   assign m332_89 =10'b0;

   // m332_90 = W*in
   wire signed [9:0] m332_90;
   assign m332_90 ={ {3{in332[5]}} , in332 , {1{1'b0}} };

   // m332_91 = W*in
   wire signed [9:0] m332_91;
   assign m332_91 =10'b0;

   // m332_92 = W*in
   wire signed [9:0] m332_92;
   assign m332_92 =10'b0;

   // m332_93 = W*in
   wire signed [9:0] m332_93;
   assign m332_93 =10'b0;

   // m332_94 = W*in
   wire signed [9:0] m332_94;
   assign m332_94 =10'b0;

   // m332_95 = W*in
   wire signed [9:0] m332_95;
   assign m332_95 =10'b0;

   // m332_96 = W*in
   wire signed [9:0] m332_96;
   assign m332_96 =10'b0;

   // m332_97 = W*in
   wire signed [9:0] m332_97;
   assign m332_97 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_98 = W*in
   wire signed [9:0] m332_98;
   assign m332_98 =10'b0;

   // m332_99 = W*in
   wire signed [9:0] m332_99;
   assign m332_99 =10'b0;

   // m332_100 = W*in
   wire signed [9:0] m332_100;
   assign m332_100 =10'b0;

   // m332_101 = W*in
   wire signed [9:0] m332_101;
   assign m332_101 =10'b0;

   // m332_102 = W*in
   wire signed [9:0] m332_102;
   assign m332_102 =10'b0;

   // m332_103 = W*in
   wire signed [9:0] m332_103;
   assign m332_103 =10'b0;

   // m332_104 = W*in
   wire signed [9:0] m332_104;
   assign m332_104 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_105 = W*in
   wire signed [9:0] m332_105;
   assign m332_105 =10'b0;

   // m332_106 = W*in
   wire signed [9:0] m332_106;
   assign m332_106 =10'b0;

   // m332_107 = W*in
   wire signed [9:0] m332_107;
   assign m332_107 =10'b0;

   // m332_108 = W*in
   wire signed [9:0] m332_108;
   assign m332_108 =10'b0;

   // m332_109 = W*in
   wire signed [9:0] m332_109;
   assign m332_109 =10'b0;

   // m332_110 = W*in
   wire signed [9:0] m332_110;
   assign m332_110 =10'b0;

   // m332_111 = W*in
   wire signed [9:0] m332_111;
   assign m332_111 =10'b0;

   // m332_112 = W*in
   wire signed [9:0] m332_112;
   assign m332_112 ={ {4{neg332[5]}} , neg332[5:0] };

   // m332_113 = W*in
   wire signed [9:0] m332_113;
   assign m332_113 =10'b0;

   // m332_114 = W*in
   wire signed [9:0] m332_114;
   assign m332_114 ={ {5{in332[5]}} , in332[5:1] };

   // m332_115 = W*in
   wire signed [9:0] m332_115;
   assign m332_115 =10'b0;

   // m332_116 = W*in
   wire signed [9:0] m332_116;
   assign m332_116 =10'b0;

   // m332_117 = W*in
   wire signed [9:0] m332_117;
   assign m332_117 =10'b0;

   // m333_1 = W*in
   wire signed [9:0] m333_1;
   assign m333_1 =10'b0;

   // m333_2 = W*in
   wire signed [9:0] m333_2;
   assign m333_2 =10'b0;

   // m333_3 = W*in
   wire signed [9:0] m333_3;
   assign m333_3 =10'b0;

   // m333_4 = W*in
   wire signed [9:0] m333_4;
   assign m333_4 =10'b0;

   // m333_5 = W*in
   wire signed [9:0] m333_5;
   assign m333_5 =10'b0;

   // m333_6 = W*in
   wire signed [9:0] m333_6;
   assign m333_6 =10'b0;

   // m333_7 = W*in
   wire signed [9:0] m333_7;
   assign m333_7 =10'b0;

   // m333_8 = W*in
   wire signed [9:0] m333_8;
   assign m333_8 =10'b0;

   // m333_9 = W*in
   wire signed [9:0] m333_9;
   assign m333_9 =10'b0;

   // m333_10 = W*in
   wire signed [9:0] m333_10;
   assign m333_10 =10'b0;

   // m333_11 = W*in
   wire signed [9:0] m333_11;
   assign m333_11 =10'b0;

   // m333_12 = W*in
   wire signed [9:0] m333_12;
   assign m333_12 =10'b0;

   // m333_13 = W*in
   wire signed [9:0] m333_13;
   assign m333_13 =10'b0;

   // m333_14 = W*in
   wire signed [9:0] m333_14;
   assign m333_14 =10'b0;

   // m333_15 = W*in
   wire signed [9:0] m333_15;
   assign m333_15 =10'b0;

   // m333_16 = W*in
   wire signed [9:0] m333_16;
   assign m333_16 =10'b0;

   // m333_17 = W*in
   wire signed [9:0] m333_17;
   assign m333_17 =10'b0;

   // m333_18 = W*in
   wire signed [9:0] m333_18;
   assign m333_18 =10'b0;

   // m333_19 = W*in
   wire signed [9:0] m333_19;
   assign m333_19 ={ {5{neg333[5]}} , neg333[5:1] };

   // m333_20 = W*in
   wire signed [9:0] m333_20;
   assign m333_20 =10'b0;

   // m333_21 = W*in
   wire signed [9:0] m333_21;
   assign m333_21 =10'b0;

   // m333_22 = W*in
   wire signed [9:0] m333_22;
   assign m333_22 =10'b0;

   // m333_23 = W*in
   wire signed [9:0] m333_23;
   assign m333_23 =10'b0;

   // m333_24 = W*in
   wire signed [9:0] m333_24;
   assign m333_24 =10'b0;

   // m333_25 = W*in
   wire signed [9:0] m333_25;
   assign m333_25 =10'b0;

   // m333_26 = W*in
   wire signed [9:0] m333_26;
   assign m333_26 =10'b0;

   // m333_27 = W*in
   wire signed [9:0] m333_27;
   assign m333_27 =10'b0;

   // m333_28 = W*in
   wire signed [9:0] m333_28;
   assign m333_28 =10'b0;

   // m333_29 = W*in
   wire signed [9:0] m333_29;
   assign m333_29 =10'b0;

   // m333_30 = W*in
   wire signed [9:0] m333_30;
   assign m333_30 ={ {5{neg333[5]}} , neg333[5:1] };

   // m333_31 = W*in
   wire signed [9:0] m333_31;
   assign m333_31 =10'b0;

   // m333_32 = W*in
   wire signed [9:0] m333_32;
   assign m333_32 =10'b0;

   // m333_33 = W*in
   wire signed [9:0] m333_33;
   assign m333_33 =10'b0;

   // m333_34 = W*in
   wire signed [9:0] m333_34;
   assign m333_34 =10'b0;

   // m333_35 = W*in
   wire signed [9:0] m333_35;
   assign m333_35 =10'b0;

   // m333_36 = W*in
   wire signed [9:0] m333_36;
   assign m333_36 =10'b0;

   // m333_37 = W*in
   wire signed [9:0] m333_37;
   assign m333_37 =10'b0;

   // m333_38 = W*in
   wire signed [9:0] m333_38;
   assign m333_38 =10'b0;

   // m333_39 = W*in
   wire signed [9:0] m333_39;
   assign m333_39 =10'b0;

   // m333_40 = W*in
   wire signed [9:0] m333_40;
   assign m333_40 =10'b0;

   // m333_41 = W*in
   wire signed [9:0] m333_41;
   assign m333_41 ={ {4{neg333[5]}} , neg333[5:0] };

   // m333_42 = W*in
   wire signed [9:0] m333_42;
   assign m333_42 =10'b0;

   // m333_43 = W*in
   wire signed [9:0] m333_43;
   assign m333_43 =10'b0;

   // m333_44 = W*in
   wire signed [9:0] m333_44;
   assign m333_44 =10'b0;

   // m333_45 = W*in
   wire signed [9:0] m333_45;
   assign m333_45 =10'b0;

   // m333_46 = W*in
   wire signed [9:0] m333_46;
   assign m333_46 =10'b0;

   // m333_47 = W*in
   wire signed [9:0] m333_47;
   assign m333_47 =10'b0;

   // m333_48 = W*in
   wire signed [9:0] m333_48;
   assign m333_48 =10'b0;

   // m333_49 = W*in
   wire signed [9:0] m333_49;
   assign m333_49 =10'b0;

   // m333_50 = W*in
   wire signed [9:0] m333_50;
   assign m333_50 =10'b0;

   // m333_51 = W*in
   wire signed [9:0] m333_51;
   assign m333_51 =10'b0;

   // m333_52 = W*in
   wire signed [9:0] m333_52;
   assign m333_52 =10'b0;

   // m333_53 = W*in
   wire signed [9:0] m333_53;
   assign m333_53 =10'b0;

   // m333_54 = W*in
   wire signed [9:0] m333_54;
   assign m333_54 =10'b0;

   // m333_55 = W*in
   wire signed [9:0] m333_55;
   assign m333_55 =10'b0;

   // m333_56 = W*in
   wire signed [9:0] m333_56;
   assign m333_56 =10'b0;

   // m333_57 = W*in
   wire signed [9:0] m333_57;
   assign m333_57 =10'b0;

   // m333_58 = W*in
   wire signed [9:0] m333_58;
   assign m333_58 =10'b0;

   // m333_59 = W*in
   wire signed [9:0] m333_59;
   assign m333_59 =10'b0;

   // m333_60 = W*in
   wire signed [9:0] m333_60;
   assign m333_60 =10'b0;

   // m333_61 = W*in
   wire signed [9:0] m333_61;
   assign m333_61 =10'b0;

   // m333_62 = W*in
   wire signed [9:0] m333_62;
   assign m333_62 =10'b0;

   // m333_63 = W*in
   wire signed [9:0] m333_63;
   assign m333_63 =10'b0;

   // m333_64 = W*in
   wire signed [9:0] m333_64;
   assign m333_64 =10'b0;

   // m333_65 = W*in
   wire signed [9:0] m333_65;
   assign m333_65 ={ {5{neg333[5]}} , neg333[5:1] };

   // m333_66 = W*in
   wire signed [9:0] m333_66;
   assign m333_66 ={ {5{neg333[5]}} , neg333[5:1] };

   // m333_67 = W*in
   wire signed [9:0] m333_67;
   assign m333_67 =10'b0;

   // m333_68 = W*in
   wire signed [9:0] m333_68;
   assign m333_68 =10'b0;

   // m333_69 = W*in
   wire signed [9:0] m333_69;
   assign m333_69 =10'b0;

   // m333_70 = W*in
   wire signed [9:0] m333_70;
   assign m333_70 =10'b0;

   // m333_71 = W*in
   wire signed [9:0] m333_71;
   assign m333_71 =10'b0;

   // m333_72 = W*in
   wire signed [9:0] m333_72;
   assign m333_72 =10'b0;

   // m333_73 = W*in
   wire signed [9:0] m333_73;
   assign m333_73 =10'b0;

   // m333_74 = W*in
   wire signed [9:0] m333_74;
   assign m333_74 =10'b0;

   // m333_75 = W*in
   wire signed [9:0] m333_75;
   assign m333_75 =10'b0;

   // m333_76 = W*in
   wire signed [9:0] m333_76;
   assign m333_76 =10'b0;

   // m333_77 = W*in
   wire signed [9:0] m333_77;
   assign m333_77 ={ {5{in333[5]}} , in333[5:1] };

   // m333_78 = W*in
   wire signed [9:0] m333_78;
   assign m333_78 =10'b0;

   // m333_79 = W*in
   wire signed [9:0] m333_79;
   assign m333_79 =10'b0;

   // m333_80 = W*in
   wire signed [9:0] m333_80;
   assign m333_80 ={ {5{in333[5]}} , in333[5:1] };

   // m333_81 = W*in
   wire signed [9:0] m333_81;
   assign m333_81 =10'b0;

   // m333_82 = W*in
   wire signed [9:0] m333_82;
   assign m333_82 =10'b0;

   // m333_83 = W*in
   wire signed [9:0] m333_83;
   assign m333_83 =10'b0;

   // m333_84 = W*in
   wire signed [9:0] m333_84;
   assign m333_84 =10'b0;

   // m333_85 = W*in
   wire signed [9:0] m333_85;
   assign m333_85 =10'b0;

   // m333_86 = W*in
   wire signed [9:0] m333_86;
   assign m333_86 =10'b0;

   // m333_87 = W*in
   wire signed [9:0] m333_87;
   assign m333_87 =10'b0;

   // m333_88 = W*in
   wire signed [9:0] m333_88;
   assign m333_88 =10'b0;

   // m333_89 = W*in
   wire signed [9:0] m333_89;
   assign m333_89 =10'b0;

   // m333_90 = W*in
   wire signed [9:0] m333_90;
   assign m333_90 =10'b0;

   // m333_91 = W*in
   wire signed [9:0] m333_91;
   assign m333_91 =10'b0;

   // m333_92 = W*in
   wire signed [9:0] m333_92;
   assign m333_92 =10'b0;

   // m333_93 = W*in
   wire signed [9:0] m333_93;
   assign m333_93 =10'b0;

   // m333_94 = W*in
   wire signed [9:0] m333_94;
   assign m333_94 ={ {4{neg333[5]}} , neg333[5:0] };

   // m333_95 = W*in
   wire signed [9:0] m333_95;
   assign m333_95 =10'b0;

   // m333_96 = W*in
   wire signed [9:0] m333_96;
   assign m333_96 =10'b0;

   // m333_97 = W*in
   wire signed [9:0] m333_97;
   assign m333_97 =10'b0;

   // m333_98 = W*in
   wire signed [9:0] m333_98;
   assign m333_98 =10'b0;

   // m333_99 = W*in
   wire signed [9:0] m333_99;
   assign m333_99 =10'b0;

   // m333_100 = W*in
   wire signed [9:0] m333_100;
   assign m333_100 =10'b0;

   // m333_101 = W*in
   wire signed [9:0] m333_101;
   assign m333_101 =10'b0;

   // m333_102 = W*in
   wire signed [9:0] m333_102;
   assign m333_102 =10'b0;

   // m333_103 = W*in
   wire signed [9:0] m333_103;
   assign m333_103 =10'b0;

   // m333_104 = W*in
   wire signed [9:0] m333_104;
   assign m333_104 =10'b0;

   // m333_105 = W*in
   wire signed [9:0] m333_105;
   assign m333_105 =10'b0;

   // m333_106 = W*in
   wire signed [9:0] m333_106;
   assign m333_106 =10'b0;

   // m333_107 = W*in
   wire signed [9:0] m333_107;
   assign m333_107 =10'b0;

   // m333_108 = W*in
   wire signed [9:0] m333_108;
   assign m333_108 ={ {5{neg333[5]}} , neg333[5:1] };

   // m333_109 = W*in
   wire signed [9:0] m333_109;
   assign m333_109 =10'b0;

   // m333_110 = W*in
   wire signed [9:0] m333_110;
   assign m333_110 =10'b0;

   // m333_111 = W*in
   wire signed [9:0] m333_111;
   assign m333_111 =10'b0;

   // m333_112 = W*in
   wire signed [9:0] m333_112;
   assign m333_112 =10'b0;

   // m333_113 = W*in
   wire signed [9:0] m333_113;
   assign m333_113 =10'b0;

   // m333_114 = W*in
   wire signed [9:0] m333_114;
   assign m333_114 =10'b0;

   // m333_115 = W*in
   wire signed [9:0] m333_115;
   assign m333_115 =10'b0;

   // m333_116 = W*in
   wire signed [9:0] m333_116;
   assign m333_116 =10'b0;

   // m333_117 = W*in
   wire signed [9:0] m333_117;
   assign m333_117 =10'b0;

   // m334_1 = W*in
   wire signed [9:0] m334_1;
   assign m334_1 =10'b0;

   // m334_2 = W*in
   wire signed [9:0] m334_2;
   assign m334_2 =10'b0;

   // m334_3 = W*in
   wire signed [9:0] m334_3;
   assign m334_3 =10'b0;

   // m334_4 = W*in
   wire signed [9:0] m334_4;
   assign m334_4 =10'b0;

   // m334_5 = W*in
   wire signed [9:0] m334_5;
   assign m334_5 =10'b0;

   // m334_6 = W*in
   wire signed [9:0] m334_6;
   assign m334_6 =10'b0;

   // m334_7 = W*in
   wire signed [9:0] m334_7;
   assign m334_7 =10'b0;

   // m334_8 = W*in
   wire signed [9:0] m334_8;
   assign m334_8 =10'b0;

   // m334_9 = W*in
   wire signed [9:0] m334_9;
   assign m334_9 =10'b0;

   // m334_10 = W*in
   wire signed [9:0] m334_10;
   assign m334_10 =10'b0;

   // m334_11 = W*in
   wire signed [9:0] m334_11;
   assign m334_11 =10'b0;

   // m334_12 = W*in
   wire signed [9:0] m334_12;
   assign m334_12 =10'b0;

   // m334_13 = W*in
   wire signed [9:0] m334_13;
   assign m334_13 =10'b0;

   // m334_14 = W*in
   wire signed [9:0] m334_14;
   assign m334_14 =10'b0;

   // m334_15 = W*in
   wire signed [9:0] m334_15;
   assign m334_15 =10'b0;

   // m334_16 = W*in
   wire signed [9:0] m334_16;
   assign m334_16 =10'b0;

   // m334_17 = W*in
   wire signed [9:0] m334_17;
   assign m334_17 =10'b0;

   // m334_18 = W*in
   wire signed [9:0] m334_18;
   assign m334_18 =10'b0;

   // m334_19 = W*in
   wire signed [9:0] m334_19;
   assign m334_19 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_20 = W*in
   wire signed [9:0] m334_20;
   assign m334_20 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_21 = W*in
   wire signed [9:0] m334_21;
   assign m334_21 ={ {5{in334[5]}} , in334[5:1] };

   // m334_22 = W*in
   wire signed [9:0] m334_22;
   assign m334_22 =10'b0;

   // m334_23 = W*in
   wire signed [9:0] m334_23;
   assign m334_23 =10'b0;

   // m334_24 = W*in
   wire signed [9:0] m334_24;
   assign m334_24 =10'b0;

   // m334_25 = W*in
   wire signed [9:0] m334_25;
   assign m334_25 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_26 = W*in
   wire signed [9:0] m334_26;
   assign m334_26 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_27 = W*in
   wire signed [9:0] m334_27;
   assign m334_27 =10'b0;

   // m334_28 = W*in
   wire signed [9:0] m334_28;
   assign m334_28 =10'b0;

   // m334_29 = W*in
   wire signed [9:0] m334_29;
   assign m334_29 =10'b0;

   // m334_30 = W*in
   wire signed [9:0] m334_30;
   assign m334_30 =10'b0;

   // m334_31 = W*in
   wire signed [9:0] m334_31;
   assign m334_31 =10'b0;

   // m334_32 = W*in
   wire signed [9:0] m334_32;
   assign m334_32 =10'b0;

   // m334_33 = W*in
   wire signed [9:0] m334_33;
   assign m334_33 =10'b0;

   // m334_34 = W*in
   wire signed [9:0] m334_34;
   assign m334_34 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_35 = W*in
   wire signed [9:0] m334_35;
   assign m334_35 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_36 = W*in
   wire signed [9:0] m334_36;
   assign m334_36 =10'b0;

   // m334_37 = W*in
   wire signed [9:0] m334_37;
   assign m334_37 =10'b0;

   // m334_38 = W*in
   wire signed [9:0] m334_38;
   assign m334_38 =10'b0;

   // m334_39 = W*in
   wire signed [9:0] m334_39;
   assign m334_39 =10'b0;

   // m334_40 = W*in
   wire signed [9:0] m334_40;
   assign m334_40 =10'b0;

   // m334_41 = W*in
   wire signed [9:0] m334_41;
   assign m334_41 =10'b0;

   // m334_42 = W*in
   wire signed [9:0] m334_42;
   assign m334_42 =10'b0;

   // m334_43 = W*in
   wire signed [9:0] m334_43;
   assign m334_43 =10'b0;

   // m334_44 = W*in
   wire signed [9:0] m334_44;
   assign m334_44 =10'b0;

   // m334_45 = W*in
   wire signed [9:0] m334_45;
   assign m334_45 =10'b0;

   // m334_46 = W*in
   wire signed [9:0] m334_46;
   assign m334_46 =10'b0;

   // m334_47 = W*in
   wire signed [9:0] m334_47;
   assign m334_47 =10'b0;

   // m334_48 = W*in
   wire signed [9:0] m334_48;
   assign m334_48 =10'b0;

   // m334_49 = W*in
   wire signed [9:0] m334_49;
   assign m334_49 =10'b0;

   // m334_50 = W*in
   wire signed [9:0] m334_50;
   assign m334_50 =10'b0;

   // m334_51 = W*in
   wire signed [9:0] m334_51;
   assign m334_51 =10'b0;

   // m334_52 = W*in
   wire signed [9:0] m334_52;
   assign m334_52 =10'b0;

   // m334_53 = W*in
   wire signed [9:0] m334_53;
   assign m334_53 =10'b0;

   // m334_54 = W*in
   wire signed [9:0] m334_54;
   assign m334_54 =10'b0;

   // m334_55 = W*in
   wire signed [9:0] m334_55;
   assign m334_55 =10'b0;

   // m334_56 = W*in
   wire signed [9:0] m334_56;
   assign m334_56 =10'b0;

   // m334_57 = W*in
   wire signed [9:0] m334_57;
   assign m334_57 =10'b0;

   // m334_58 = W*in
   wire signed [9:0] m334_58;
   assign m334_58 =10'b0;

   // m334_59 = W*in
   wire signed [9:0] m334_59;
   assign m334_59 =10'b0;

   // m334_60 = W*in
   wire signed [9:0] m334_60;
   assign m334_60 =10'b0;

   // m334_61 = W*in
   wire signed [9:0] m334_61;
   assign m334_61 =10'b0;

   // m334_62 = W*in
   wire signed [9:0] m334_62;
   assign m334_62 =10'b0;

   // m334_63 = W*in
   wire signed [9:0] m334_63;
   assign m334_63 =10'b0;

   // m334_64 = W*in
   wire signed [9:0] m334_64;
   assign m334_64 =10'b0;

   // m334_65 = W*in
   wire signed [9:0] m334_65;
   assign m334_65 ={ {5{in334[5]}} , in334[5:1] };

   // m334_66 = W*in
   wire signed [9:0] m334_66;
   assign m334_66 ={ {5{in334[5]}} , in334[5:1] };

   // m334_67 = W*in
   wire signed [9:0] m334_67;
   assign m334_67 =10'b0;

   // m334_68 = W*in
   wire signed [9:0] m334_68;
   assign m334_68 =10'b0;

   // m334_69 = W*in
   wire signed [9:0] m334_69;
   assign m334_69 =10'b0;

   // m334_70 = W*in
   wire signed [9:0] m334_70;
   assign m334_70 =10'b0;

   // m334_71 = W*in
   wire signed [9:0] m334_71;
   assign m334_71 =10'b0;

   // m334_72 = W*in
   wire signed [9:0] m334_72;
   assign m334_72 =10'b0;

   // m334_73 = W*in
   wire signed [9:0] m334_73;
   assign m334_73 =10'b0;

   // m334_74 = W*in
   wire signed [9:0] m334_74;
   assign m334_74 =10'b0;

   // m334_75 = W*in
   wire signed [9:0] m334_75;
   assign m334_75 =10'b0;

   // m334_76 = W*in
   wire signed [9:0] m334_76;
   assign m334_76 =10'b0;

   // m334_77 = W*in
   wire signed [9:0] m334_77;
   assign m334_77 =10'b0;

   // m334_78 = W*in
   wire signed [9:0] m334_78;
   assign m334_78 =10'b0;

   // m334_79 = W*in
   wire signed [9:0] m334_79;
   assign m334_79 =10'b0;

   // m334_80 = W*in
   wire signed [9:0] m334_80;
   assign m334_80 =10'b0;

   // m334_81 = W*in
   wire signed [9:0] m334_81;
   assign m334_81 =10'b0;

   // m334_82 = W*in
   wire signed [9:0] m334_82;
   assign m334_82 =10'b0;

   // m334_83 = W*in
   wire signed [9:0] m334_83;
   assign m334_83 =10'b0;

   // m334_84 = W*in
   wire signed [9:0] m334_84;
   assign m334_84 =10'b0;

   // m334_85 = W*in
   wire signed [9:0] m334_85;
   assign m334_85 ={ {5{in334[5]}} , in334[5:1] };

   // m334_86 = W*in
   wire signed [9:0] m334_86;
   assign m334_86 =10'b0;

   // m334_87 = W*in
   wire signed [9:0] m334_87;
   assign m334_87 =10'b0;

   // m334_88 = W*in
   wire signed [9:0] m334_88;
   assign m334_88 =10'b0;

   // m334_89 = W*in
   wire signed [9:0] m334_89;
   assign m334_89 =10'b0;

   // m334_90 = W*in
   wire signed [9:0] m334_90;
   assign m334_90 =10'b0;

   // m334_91 = W*in
   wire signed [9:0] m334_91;
   assign m334_91 =10'b0;

   // m334_92 = W*in
   wire signed [9:0] m334_92;
   assign m334_92 =10'b0;

   // m334_93 = W*in
   wire signed [9:0] m334_93;
   assign m334_93 =10'b0;

   // m334_94 = W*in
   wire signed [9:0] m334_94;
   assign m334_94 =10'b0;

   // m334_95 = W*in
   wire signed [9:0] m334_95;
   assign m334_95 =10'b0;

   // m334_96 = W*in
   wire signed [9:0] m334_96;
   assign m334_96 =10'b0;

   // m334_97 = W*in
   wire signed [9:0] m334_97;
   assign m334_97 =10'b0;

   // m334_98 = W*in
   wire signed [9:0] m334_98;
   assign m334_98 =10'b0;

   // m334_99 = W*in
   wire signed [9:0] m334_99;
   assign m334_99 =10'b0;

   // m334_100 = W*in
   wire signed [9:0] m334_100;
   assign m334_100 =10'b0;

   // m334_101 = W*in
   wire signed [9:0] m334_101;
   assign m334_101 =10'b0;

   // m334_102 = W*in
   wire signed [9:0] m334_102;
   assign m334_102 =10'b0;

   // m334_103 = W*in
   wire signed [9:0] m334_103;
   assign m334_103 =10'b0;

   // m334_104 = W*in
   wire signed [9:0] m334_104;
   assign m334_104 =10'b0;

   // m334_105 = W*in
   wire signed [9:0] m334_105;
   assign m334_105 =10'b0;

   // m334_106 = W*in
   wire signed [9:0] m334_106;
   assign m334_106 =10'b0;

   // m334_107 = W*in
   wire signed [9:0] m334_107;
   assign m334_107 =10'b0;

   // m334_108 = W*in
   wire signed [9:0] m334_108;
   assign m334_108 ={ {5{in334[5]}} , in334[5:1] };

   // m334_109 = W*in
   wire signed [9:0] m334_109;
   assign m334_109 ={ {5{in334[5]}} , in334[5:1] };

   // m334_110 = W*in
   wire signed [9:0] m334_110;
   assign m334_110 =10'b0;

   // m334_111 = W*in
   wire signed [9:0] m334_111;
   assign m334_111 =10'b0;

   // m334_112 = W*in
   wire signed [9:0] m334_112;
   assign m334_112 =10'b0;

   // m334_113 = W*in
   wire signed [9:0] m334_113;
   assign m334_113 =10'b0;

   // m334_114 = W*in
   wire signed [9:0] m334_114;
   assign m334_114 =10'b0;

   // m334_115 = W*in
   wire signed [9:0] m334_115;
   assign m334_115 ={ {5{neg334[5]}} , neg334[5:1] };

   // m334_116 = W*in
   wire signed [9:0] m334_116;
   assign m334_116 ={ {4{in334[5]}} , in334[5:0] };

   // m334_117 = W*in
   wire signed [9:0] m334_117;
   assign m334_117 =10'b0;

   // m335_1 = W*in
   wire signed [9:0] m335_1;
   assign m335_1 =10'b0;

   // m335_2 = W*in
   wire signed [9:0] m335_2;
   assign m335_2 =10'b0;

   // m335_3 = W*in
   wire signed [9:0] m335_3;
   assign m335_3 =10'b0;

   // m335_4 = W*in
   wire signed [9:0] m335_4;
   assign m335_4 =10'b0;

   // m335_5 = W*in
   wire signed [9:0] m335_5;
   assign m335_5 =10'b0;

   // m335_6 = W*in
   wire signed [9:0] m335_6;
   assign m335_6 =10'b0;

   // m335_7 = W*in
   wire signed [9:0] m335_7;
   assign m335_7 =10'b0;

   // m335_8 = W*in
   wire signed [9:0] m335_8;
   assign m335_8 =10'b0;

   // m335_9 = W*in
   wire signed [9:0] m335_9;
   assign m335_9 =10'b0;

   // m335_10 = W*in
   wire signed [9:0] m335_10;
   assign m335_10 =10'b0;

   // m335_11 = W*in
   wire signed [9:0] m335_11;
   assign m335_11 =10'b0;

   // m335_12 = W*in
   wire signed [9:0] m335_12;
   assign m335_12 =10'b0;

   // m335_13 = W*in
   wire signed [9:0] m335_13;
   assign m335_13 =10'b0;

   // m335_14 = W*in
   wire signed [9:0] m335_14;
   assign m335_14 =10'b0;

   // m335_15 = W*in
   wire signed [9:0] m335_15;
   assign m335_15 =10'b0;

   // m335_16 = W*in
   wire signed [9:0] m335_16;
   assign m335_16 ={ {5{in335[5]}} , in335[5:1] };

   // m335_17 = W*in
   wire signed [9:0] m335_17;
   assign m335_17 =10'b0;

   // m335_18 = W*in
   wire signed [9:0] m335_18;
   assign m335_18 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_19 = W*in
   wire signed [9:0] m335_19;
   assign m335_19 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_20 = W*in
   wire signed [9:0] m335_20;
   assign m335_20 =10'b0;

   // m335_21 = W*in
   wire signed [9:0] m335_21;
   assign m335_21 =10'b0;

   // m335_22 = W*in
   wire signed [9:0] m335_22;
   assign m335_22 =10'b0;

   // m335_23 = W*in
   wire signed [9:0] m335_23;
   assign m335_23 =10'b0;

   // m335_24 = W*in
   wire signed [9:0] m335_24;
   assign m335_24 =10'b0;

   // m335_25 = W*in
   wire signed [9:0] m335_25;
   assign m335_25 =10'b0;

   // m335_26 = W*in
   wire signed [9:0] m335_26;
   assign m335_26 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_27 = W*in
   wire signed [9:0] m335_27;
   assign m335_27 =10'b0;

   // m335_28 = W*in
   wire signed [9:0] m335_28;
   assign m335_28 =10'b0;

   // m335_29 = W*in
   wire signed [9:0] m335_29;
   assign m335_29 =10'b0;

   // m335_30 = W*in
   wire signed [9:0] m335_30;
   assign m335_30 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_31 = W*in
   wire signed [9:0] m335_31;
   assign m335_31 =10'b0;

   // m335_32 = W*in
   wire signed [9:0] m335_32;
   assign m335_32 =10'b0;

   // m335_33 = W*in
   wire signed [9:0] m335_33;
   assign m335_33 =10'b0;

   // m335_34 = W*in
   wire signed [9:0] m335_34;
   assign m335_34 =10'b0;

   // m335_35 = W*in
   wire signed [9:0] m335_35;
   assign m335_35 =10'b0;

   // m335_36 = W*in
   wire signed [9:0] m335_36;
   assign m335_36 =10'b0;

   // m335_37 = W*in
   wire signed [9:0] m335_37;
   assign m335_37 =10'b0;

   // m335_38 = W*in
   wire signed [9:0] m335_38;
   assign m335_38 =10'b0;

   // m335_39 = W*in
   wire signed [9:0] m335_39;
   assign m335_39 =10'b0;

   // m335_40 = W*in
   wire signed [9:0] m335_40;
   assign m335_40 =10'b0;

   // m335_41 = W*in
   wire signed [9:0] m335_41;
   assign m335_41 =10'b0;

   // m335_42 = W*in
   wire signed [9:0] m335_42;
   assign m335_42 =10'b0;

   // m335_43 = W*in
   wire signed [9:0] m335_43;
   assign m335_43 =10'b0;

   // m335_44 = W*in
   wire signed [9:0] m335_44;
   assign m335_44 =10'b0;

   // m335_45 = W*in
   wire signed [9:0] m335_45;
   assign m335_45 =10'b0;

   // m335_46 = W*in
   wire signed [9:0] m335_46;
   assign m335_46 =10'b0;

   // m335_47 = W*in
   wire signed [9:0] m335_47;
   assign m335_47 =10'b0;

   // m335_48 = W*in
   wire signed [9:0] m335_48;
   assign m335_48 =10'b0;

   // m335_49 = W*in
   wire signed [9:0] m335_49;
   assign m335_49 =10'b0;

   // m335_50 = W*in
   wire signed [9:0] m335_50;
   assign m335_50 =10'b0;

   // m335_51 = W*in
   wire signed [9:0] m335_51;
   assign m335_51 =10'b0;

   // m335_52 = W*in
   wire signed [9:0] m335_52;
   assign m335_52 =10'b0;

   // m335_53 = W*in
   wire signed [9:0] m335_53;
   assign m335_53 =10'b0;

   // m335_54 = W*in
   wire signed [9:0] m335_54;
   assign m335_54 =10'b0;

   // m335_55 = W*in
   wire signed [9:0] m335_55;
   assign m335_55 =10'b0;

   // m335_56 = W*in
   wire signed [9:0] m335_56;
   assign m335_56 =10'b0;

   // m335_57 = W*in
   wire signed [9:0] m335_57;
   assign m335_57 =10'b0;

   // m335_58 = W*in
   wire signed [9:0] m335_58;
   assign m335_58 =10'b0;

   // m335_59 = W*in
   wire signed [9:0] m335_59;
   assign m335_59 =10'b0;

   // m335_60 = W*in
   wire signed [9:0] m335_60;
   assign m335_60 =10'b0;

   // m335_61 = W*in
   wire signed [9:0] m335_61;
   assign m335_61 =10'b0;

   // m335_62 = W*in
   wire signed [9:0] m335_62;
   assign m335_62 =10'b0;

   // m335_63 = W*in
   wire signed [9:0] m335_63;
   assign m335_63 =10'b0;

   // m335_64 = W*in
   wire signed [9:0] m335_64;
   assign m335_64 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_65 = W*in
   wire signed [9:0] m335_65;
   assign m335_65 =10'b0;

   // m335_66 = W*in
   wire signed [9:0] m335_66;
   assign m335_66 =10'b0;

   // m335_67 = W*in
   wire signed [9:0] m335_67;
   assign m335_67 =10'b0;

   // m335_68 = W*in
   wire signed [9:0] m335_68;
   assign m335_68 =10'b0;

   // m335_69 = W*in
   wire signed [9:0] m335_69;
   assign m335_69 =10'b0;

   // m335_70 = W*in
   wire signed [9:0] m335_70;
   assign m335_70 ={ {4{in335[5]}} , in335[5:0] };

   // m335_71 = W*in
   wire signed [9:0] m335_71;
   assign m335_71 =10'b0;

   // m335_72 = W*in
   wire signed [9:0] m335_72;
   assign m335_72 =10'b0;

   // m335_73 = W*in
   wire signed [9:0] m335_73;
   assign m335_73 =10'b0;

   // m335_74 = W*in
   wire signed [9:0] m335_74;
   assign m335_74 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_75 = W*in
   wire signed [9:0] m335_75;
   assign m335_75 =10'b0;

   // m335_76 = W*in
   wire signed [9:0] m335_76;
   assign m335_76 =10'b0;

   // m335_77 = W*in
   wire signed [9:0] m335_77;
   assign m335_77 =10'b0;

   // m335_78 = W*in
   wire signed [9:0] m335_78;
   assign m335_78 =10'b0;

   // m335_79 = W*in
   wire signed [9:0] m335_79;
   assign m335_79 =10'b0;

   // m335_80 = W*in
   wire signed [9:0] m335_80;
   assign m335_80 =10'b0;

   // m335_81 = W*in
   wire signed [9:0] m335_81;
   assign m335_81 =10'b0;

   // m335_82 = W*in
   wire signed [9:0] m335_82;
   assign m335_82 =10'b0;

   // m335_83 = W*in
   wire signed [9:0] m335_83;
   assign m335_83 ={ {5{in335[5]}} , in335[5:1] };

   // m335_84 = W*in
   wire signed [9:0] m335_84;
   assign m335_84 =10'b0;

   // m335_85 = W*in
   wire signed [9:0] m335_85;
   assign m335_85 ={ {5{in335[5]}} , in335[5:1] };

   // m335_86 = W*in
   wire signed [9:0] m335_86;
   assign m335_86 =10'b0;

   // m335_87 = W*in
   wire signed [9:0] m335_87;
   assign m335_87 =10'b0;

   // m335_88 = W*in
   wire signed [9:0] m335_88;
   assign m335_88 =10'b0;

   // m335_89 = W*in
   wire signed [9:0] m335_89;
   assign m335_89 =10'b0;

   // m335_90 = W*in
   wire signed [9:0] m335_90;
   assign m335_90 =10'b0;

   // m335_91 = W*in
   wire signed [9:0] m335_91;
   assign m335_91 =10'b0;

   // m335_92 = W*in
   wire signed [9:0] m335_92;
   assign m335_92 =10'b0;

   // m335_93 = W*in
   wire signed [9:0] m335_93;
   assign m335_93 =10'b0;

   // m335_94 = W*in
   wire signed [9:0] m335_94;
   assign m335_94 ={ {4{neg335[5]}} , neg335[5:0] };

   // m335_95 = W*in
   wire signed [9:0] m335_95;
   assign m335_95 =10'b0;

   // m335_96 = W*in
   wire signed [9:0] m335_96;
   assign m335_96 =10'b0;

   // m335_97 = W*in
   wire signed [9:0] m335_97;
   assign m335_97 =10'b0;

   // m335_98 = W*in
   wire signed [9:0] m335_98;
   assign m335_98 =10'b0;

   // m335_99 = W*in
   wire signed [9:0] m335_99;
   assign m335_99 =10'b0;

   // m335_100 = W*in
   wire signed [9:0] m335_100;
   assign m335_100 =10'b0;

   // m335_101 = W*in
   wire signed [9:0] m335_101;
   assign m335_101 =10'b0;

   // m335_102 = W*in
   wire signed [9:0] m335_102;
   assign m335_102 =10'b0;

   // m335_103 = W*in
   wire signed [9:0] m335_103;
   assign m335_103 =10'b0;

   // m335_104 = W*in
   wire signed [9:0] m335_104;
   assign m335_104 =10'b0;

   // m335_105 = W*in
   wire signed [9:0] m335_105;
   assign m335_105 =10'b0;

   // m335_106 = W*in
   wire signed [9:0] m335_106;
   assign m335_106 =10'b0;

   // m335_107 = W*in
   wire signed [9:0] m335_107;
   assign m335_107 =10'b0;

   // m335_108 = W*in
   wire signed [9:0] m335_108;
   assign m335_108 =10'b0;

   // m335_109 = W*in
   wire signed [9:0] m335_109;
   assign m335_109 ={ {5{in335[5]}} , in335[5:1] };

   // m335_110 = W*in
   wire signed [9:0] m335_110;
   assign m335_110 =10'b0;

   // m335_111 = W*in
   wire signed [9:0] m335_111;
   assign m335_111 =10'b0;

   // m335_112 = W*in
   wire signed [9:0] m335_112;
   assign m335_112 =10'b0;

   // m335_113 = W*in
   wire signed [9:0] m335_113;
   assign m335_113 =10'b0;

   // m335_114 = W*in
   wire signed [9:0] m335_114;
   assign m335_114 =10'b0;

   // m335_115 = W*in
   wire signed [9:0] m335_115;
   assign m335_115 ={ {5{neg335[5]}} , neg335[5:1] };

   // m335_116 = W*in
   wire signed [9:0] m335_116;
   assign m335_116 =10'b0;

   // m335_117 = W*in
   wire signed [9:0] m335_117;
   assign m335_117 =10'b0;

   // m336_1 = W*in
   wire signed [9:0] m336_1;
   assign m336_1 =10'b0;

   // m336_2 = W*in
   wire signed [9:0] m336_2;
   assign m336_2 =10'b0;

   // m336_3 = W*in
   wire signed [9:0] m336_3;
   assign m336_3 =10'b0;

   // m336_4 = W*in
   wire signed [9:0] m336_4;
   assign m336_4 =10'b0;

   // m336_5 = W*in
   wire signed [9:0] m336_5;
   assign m336_5 =10'b0;

   // m336_6 = W*in
   wire signed [9:0] m336_6;
   assign m336_6 =10'b0;

   // m336_7 = W*in
   wire signed [9:0] m336_7;
   assign m336_7 =10'b0;

   // m336_8 = W*in
   wire signed [9:0] m336_8;
   assign m336_8 =10'b0;

   // m336_9 = W*in
   wire signed [9:0] m336_9;
   assign m336_9 =10'b0;

   // m336_10 = W*in
   wire signed [9:0] m336_10;
   assign m336_10 =10'b0;

   // m336_11 = W*in
   wire signed [9:0] m336_11;
   assign m336_11 =10'b0;

   // m336_12 = W*in
   wire signed [9:0] m336_12;
   assign m336_12 =10'b0;

   // m336_13 = W*in
   wire signed [9:0] m336_13;
   assign m336_13 =10'b0;

   // m336_14 = W*in
   wire signed [9:0] m336_14;
   assign m336_14 =10'b0;

   // m336_15 = W*in
   wire signed [9:0] m336_15;
   assign m336_15 =10'b0;

   // m336_16 = W*in
   wire signed [9:0] m336_16;
   assign m336_16 =10'b0;

   // m336_17 = W*in
   wire signed [9:0] m336_17;
   assign m336_17 =10'b0;

   // m336_18 = W*in
   wire signed [9:0] m336_18;
   assign m336_18 =10'b0;

   // m336_19 = W*in
   wire signed [9:0] m336_19;
   assign m336_19 =10'b0;

   // m336_20 = W*in
   wire signed [9:0] m336_20;
   assign m336_20 ={ {5{neg336[5]}} , neg336[5:1] };

   // m336_21 = W*in
   wire signed [9:0] m336_21;
   assign m336_21 =10'b0;

   // m336_22 = W*in
   wire signed [9:0] m336_22;
   assign m336_22 =10'b0;

   // m336_23 = W*in
   wire signed [9:0] m336_23;
   assign m336_23 =10'b0;

   // m336_24 = W*in
   wire signed [9:0] m336_24;
   assign m336_24 =10'b0;

   // m336_25 = W*in
   wire signed [9:0] m336_25;
   assign m336_25 =10'b0;

   // m336_26 = W*in
   wire signed [9:0] m336_26;
   assign m336_26 =10'b0;

   // m336_27 = W*in
   wire signed [9:0] m336_27;
   assign m336_27 ={ {5{neg336[5]}} , neg336[5:1] };

   // m336_28 = W*in
   wire signed [9:0] m336_28;
   assign m336_28 =10'b0;

   // m336_29 = W*in
   wire signed [9:0] m336_29;
   assign m336_29 ={ {4{in336[5]}} , in336[5:0] };

   // m336_30 = W*in
   wire signed [9:0] m336_30;
   assign m336_30 ={ {5{neg336[5]}} , neg336[5:1] };

   // m336_31 = W*in
   wire signed [9:0] m336_31;
   assign m336_31 =10'b0;

   // m336_32 = W*in
   wire signed [9:0] m336_32;
   assign m336_32 =10'b0;

   // m336_33 = W*in
   wire signed [9:0] m336_33;
   assign m336_33 =10'b0;

   // m336_34 = W*in
   wire signed [9:0] m336_34;
   assign m336_34 =10'b0;

   // m336_35 = W*in
   wire signed [9:0] m336_35;
   assign m336_35 =10'b0;

   // m336_36 = W*in
   wire signed [9:0] m336_36;
   assign m336_36 =10'b0;

   // m336_37 = W*in
   wire signed [9:0] m336_37;
   assign m336_37 =10'b0;

   // m336_38 = W*in
   wire signed [9:0] m336_38;
   assign m336_38 =10'b0;

   // m336_39 = W*in
   wire signed [9:0] m336_39;
   assign m336_39 =10'b0;

   // m336_40 = W*in
   wire signed [9:0] m336_40;
   assign m336_40 =10'b0;

   // m336_41 = W*in
   wire signed [9:0] m336_41;
   assign m336_41 =10'b0;

   // m336_42 = W*in
   wire signed [9:0] m336_42;
   assign m336_42 =10'b0;

   // m336_43 = W*in
   wire signed [9:0] m336_43;
   assign m336_43 =10'b0;

   // m336_44 = W*in
   wire signed [9:0] m336_44;
   assign m336_44 =10'b0;

   // m336_45 = W*in
   wire signed [9:0] m336_45;
   assign m336_45 =10'b0;

   // m336_46 = W*in
   wire signed [9:0] m336_46;
   assign m336_46 =10'b0;

   // m336_47 = W*in
   wire signed [9:0] m336_47;
   assign m336_47 =10'b0;

   // m336_48 = W*in
   wire signed [9:0] m336_48;
   assign m336_48 =10'b0;

   // m336_49 = W*in
   wire signed [9:0] m336_49;
   assign m336_49 =10'b0;

   // m336_50 = W*in
   wire signed [9:0] m336_50;
   assign m336_50 =10'b0;

   // m336_51 = W*in
   wire signed [9:0] m336_51;
   assign m336_51 =10'b0;

   // m336_52 = W*in
   wire signed [9:0] m336_52;
   assign m336_52 =10'b0;

   // m336_53 = W*in
   wire signed [9:0] m336_53;
   assign m336_53 =10'b0;

   // m336_54 = W*in
   wire signed [9:0] m336_54;
   assign m336_54 =10'b0;

   // m336_55 = W*in
   wire signed [9:0] m336_55;
   assign m336_55 =10'b0;

   // m336_56 = W*in
   wire signed [9:0] m336_56;
   assign m336_56 =10'b0;

   // m336_57 = W*in
   wire signed [9:0] m336_57;
   assign m336_57 =10'b0;

   // m336_58 = W*in
   wire signed [9:0] m336_58;
   assign m336_58 =10'b0;

   // m336_59 = W*in
   wire signed [9:0] m336_59;
   assign m336_59 =10'b0;

   // m336_60 = W*in
   wire signed [9:0] m336_60;
   assign m336_60 =10'b0;

   // m336_61 = W*in
   wire signed [9:0] m336_61;
   assign m336_61 =10'b0;

   // m336_62 = W*in
   wire signed [9:0] m336_62;
   assign m336_62 =10'b0;

   // m336_63 = W*in
   wire signed [9:0] m336_63;
   assign m336_63 =10'b0;

   // m336_64 = W*in
   wire signed [9:0] m336_64;
   assign m336_64 =10'b0;

   // m336_65 = W*in
   wire signed [9:0] m336_65;
   assign m336_65 =10'b0;

   // m336_66 = W*in
   wire signed [9:0] m336_66;
   assign m336_66 =10'b0;

   // m336_67 = W*in
   wire signed [9:0] m336_67;
   assign m336_67 =10'b0;

   // m336_68 = W*in
   wire signed [9:0] m336_68;
   assign m336_68 =10'b0;

   // m336_69 = W*in
   wire signed [9:0] m336_69;
   assign m336_69 =10'b0;

   // m336_70 = W*in
   wire signed [9:0] m336_70;
   assign m336_70 ={ {5{in336[5]}} , in336[5:1] };

   // m336_71 = W*in
   wire signed [9:0] m336_71;
   assign m336_71 ={ {5{neg336[5]}} , neg336[5:1] };

   // m336_72 = W*in
   wire signed [9:0] m336_72;
   assign m336_72 =10'b0;

   // m336_73 = W*in
   wire signed [9:0] m336_73;
   assign m336_73 =10'b0;

   // m336_74 = W*in
   wire signed [9:0] m336_74;
   assign m336_74 =10'b0;

   // m336_75 = W*in
   wire signed [9:0] m336_75;
   assign m336_75 =10'b0;

   // m336_76 = W*in
   wire signed [9:0] m336_76;
   assign m336_76 =10'b0;

   // m336_77 = W*in
   wire signed [9:0] m336_77;
   assign m336_77 =10'b0;

   // m336_78 = W*in
   wire signed [9:0] m336_78;
   assign m336_78 =10'b0;

   // m336_79 = W*in
   wire signed [9:0] m336_79;
   assign m336_79 =10'b0;

   // m336_80 = W*in
   wire signed [9:0] m336_80;
   assign m336_80 =10'b0;

   // m336_81 = W*in
   wire signed [9:0] m336_81;
   assign m336_81 =10'b0;

   // m336_82 = W*in
   wire signed [9:0] m336_82;
   assign m336_82 =10'b0;

   // m336_83 = W*in
   wire signed [9:0] m336_83;
   assign m336_83 =10'b0;

   // m336_84 = W*in
   wire signed [9:0] m336_84;
   assign m336_84 =10'b0;

   // m336_85 = W*in
   wire signed [9:0] m336_85;
   assign m336_85 =10'b0;

   // m336_86 = W*in
   wire signed [9:0] m336_86;
   assign m336_86 =10'b0;

   // m336_87 = W*in
   wire signed [9:0] m336_87;
   assign m336_87 =10'b0;

   // m336_88 = W*in
   wire signed [9:0] m336_88;
   assign m336_88 =10'b0;

   // m336_89 = W*in
   wire signed [9:0] m336_89;
   assign m336_89 =10'b0;

   // m336_90 = W*in
   wire signed [9:0] m336_90;
   assign m336_90 =10'b0;

   // m336_91 = W*in
   wire signed [9:0] m336_91;
   assign m336_91 =10'b0;

   // m336_92 = W*in
   wire signed [9:0] m336_92;
   assign m336_92 =10'b0;

   // m336_93 = W*in
   wire signed [9:0] m336_93;
   assign m336_93 =10'b0;

   // m336_94 = W*in
   wire signed [9:0] m336_94;
   assign m336_94 =10'b0;

   // m336_95 = W*in
   wire signed [9:0] m336_95;
   assign m336_95 =10'b0;

   // m336_96 = W*in
   wire signed [9:0] m336_96;
   assign m336_96 =10'b0;

   // m336_97 = W*in
   wire signed [9:0] m336_97;
   assign m336_97 =10'b0;

   // m336_98 = W*in
   wire signed [9:0] m336_98;
   assign m336_98 =10'b0;

   // m336_99 = W*in
   wire signed [9:0] m336_99;
   assign m336_99 =10'b0;

   // m336_100 = W*in
   wire signed [9:0] m336_100;
   assign m336_100 =10'b0;

   // m336_101 = W*in
   wire signed [9:0] m336_101;
   assign m336_101 =10'b0;

   // m336_102 = W*in
   wire signed [9:0] m336_102;
   assign m336_102 =10'b0;

   // m336_103 = W*in
   wire signed [9:0] m336_103;
   assign m336_103 =10'b0;

   // m336_104 = W*in
   wire signed [9:0] m336_104;
   assign m336_104 =10'b0;

   // m336_105 = W*in
   wire signed [9:0] m336_105;
   assign m336_105 =10'b0;

   // m336_106 = W*in
   wire signed [9:0] m336_106;
   assign m336_106 =10'b0;

   // m336_107 = W*in
   wire signed [9:0] m336_107;
   assign m336_107 =10'b0;

   // m336_108 = W*in
   wire signed [9:0] m336_108;
   assign m336_108 =10'b0;

   // m336_109 = W*in
   wire signed [9:0] m336_109;
   assign m336_109 =10'b0;

   // m336_110 = W*in
   wire signed [9:0] m336_110;
   assign m336_110 =10'b0;

   // m336_111 = W*in
   wire signed [9:0] m336_111;
   assign m336_111 =10'b0;

   // m336_112 = W*in
   wire signed [9:0] m336_112;
   assign m336_112 =10'b0;

   // m336_113 = W*in
   wire signed [9:0] m336_113;
   assign m336_113 =10'b0;

   // m336_114 = W*in
   wire signed [9:0] m336_114;
   assign m336_114 =10'b0;

   // m336_115 = W*in
   wire signed [9:0] m336_115;
   assign m336_115 ={ {5{neg336[5]}} , neg336[5:1] };

   // m336_116 = W*in
   wire signed [9:0] m336_116;
   assign m336_116 =10'b0;

   // m336_117 = W*in
   wire signed [9:0] m336_117;
   assign m336_117 =10'b0;

   // m337_1 = W*in
   wire signed [9:0] m337_1;
   assign m337_1 =10'b0;

   // m337_2 = W*in
   wire signed [9:0] m337_2;
   assign m337_2 =10'b0;

   // m337_3 = W*in
   wire signed [9:0] m337_3;
   assign m337_3 =10'b0;

   // m337_4 = W*in
   wire signed [9:0] m337_4;
   assign m337_4 =10'b0;

   // m337_5 = W*in
   wire signed [9:0] m337_5;
   assign m337_5 =10'b0;

   // m337_6 = W*in
   wire signed [9:0] m337_6;
   assign m337_6 =10'b0;

   // m337_7 = W*in
   wire signed [9:0] m337_7;
   assign m337_7 =10'b0;

   // m337_8 = W*in
   wire signed [9:0] m337_8;
   assign m337_8 =10'b0;

   // m337_9 = W*in
   wire signed [9:0] m337_9;
   assign m337_9 =10'b0;

   // m337_10 = W*in
   wire signed [9:0] m337_10;
   assign m337_10 =10'b0;

   // m337_11 = W*in
   wire signed [9:0] m337_11;
   assign m337_11 =10'b0;

   // m337_12 = W*in
   wire signed [9:0] m337_12;
   assign m337_12 =10'b0;

   // m337_13 = W*in
   wire signed [9:0] m337_13;
   assign m337_13 =10'b0;

   // m337_14 = W*in
   wire signed [9:0] m337_14;
   assign m337_14 =10'b0;

   // m337_15 = W*in
   wire signed [9:0] m337_15;
   assign m337_15 =10'b0;

   // m337_16 = W*in
   wire signed [9:0] m337_16;
   assign m337_16 =10'b0;

   // m337_17 = W*in
   wire signed [9:0] m337_17;
   assign m337_17 =10'b0;

   // m337_18 = W*in
   wire signed [9:0] m337_18;
   assign m337_18 =10'b0;

   // m337_19 = W*in
   wire signed [9:0] m337_19;
   assign m337_19 ={ {4{neg337[5]}} , neg337[5:0] };

   // m337_20 = W*in
   wire signed [9:0] m337_20;
   assign m337_20 =10'b0;

   // m337_21 = W*in
   wire signed [9:0] m337_21;
   assign m337_21 ={ {5{in337[5]}} , in337[5:1] };

   // m337_22 = W*in
   wire signed [9:0] m337_22;
   assign m337_22 =10'b0;

   // m337_23 = W*in
   wire signed [9:0] m337_23;
   assign m337_23 =10'b0;

   // m337_24 = W*in
   wire signed [9:0] m337_24;
   assign m337_24 =10'b0;

   // m337_25 = W*in
   wire signed [9:0] m337_25;
   assign m337_25 ={ {5{neg337[5]}} , neg337[5:1] };

   // m337_26 = W*in
   wire signed [9:0] m337_26;
   assign m337_26 =10'b0;

   // m337_27 = W*in
   wire signed [9:0] m337_27;
   assign m337_27 =10'b0;

   // m337_28 = W*in
   wire signed [9:0] m337_28;
   assign m337_28 ={ {5{neg337[5]}} , neg337[5:1] };

   // m337_29 = W*in
   wire signed [9:0] m337_29;
   assign m337_29 =10'b0;

   // m337_30 = W*in
   wire signed [9:0] m337_30;
   assign m337_30 =10'b0;

   // m337_31 = W*in
   wire signed [9:0] m337_31;
   assign m337_31 =10'b0;

   // m337_32 = W*in
   wire signed [9:0] m337_32;
   assign m337_32 =10'b0;

   // m337_33 = W*in
   wire signed [9:0] m337_33;
   assign m337_33 =10'b0;

   // m337_34 = W*in
   wire signed [9:0] m337_34;
   assign m337_34 =10'b0;

   // m337_35 = W*in
   wire signed [9:0] m337_35;
   assign m337_35 =10'b0;

   // m337_36 = W*in
   wire signed [9:0] m337_36;
   assign m337_36 =10'b0;

   // m337_37 = W*in
   wire signed [9:0] m337_37;
   assign m337_37 =10'b0;

   // m337_38 = W*in
   wire signed [9:0] m337_38;
   assign m337_38 =10'b0;

   // m337_39 = W*in
   wire signed [9:0] m337_39;
   assign m337_39 =10'b0;

   // m337_40 = W*in
   wire signed [9:0] m337_40;
   assign m337_40 =10'b0;

   // m337_41 = W*in
   wire signed [9:0] m337_41;
   assign m337_41 =10'b0;

   // m337_42 = W*in
   wire signed [9:0] m337_42;
   assign m337_42 =10'b0;

   // m337_43 = W*in
   wire signed [9:0] m337_43;
   assign m337_43 =10'b0;

   // m337_44 = W*in
   wire signed [9:0] m337_44;
   assign m337_44 =10'b0;

   // m337_45 = W*in
   wire signed [9:0] m337_45;
   assign m337_45 =10'b0;

   // m337_46 = W*in
   wire signed [9:0] m337_46;
   assign m337_46 =10'b0;

   // m337_47 = W*in
   wire signed [9:0] m337_47;
   assign m337_47 =10'b0;

   // m337_48 = W*in
   wire signed [9:0] m337_48;
   assign m337_48 =10'b0;

   // m337_49 = W*in
   wire signed [9:0] m337_49;
   assign m337_49 ={ {5{neg337[5]}} , neg337[5:1] };

   // m337_50 = W*in
   wire signed [9:0] m337_50;
   assign m337_50 =10'b0;

   // m337_51 = W*in
   wire signed [9:0] m337_51;
   assign m337_51 =10'b0;

   // m337_52 = W*in
   wire signed [9:0] m337_52;
   assign m337_52 =10'b0;

   // m337_53 = W*in
   wire signed [9:0] m337_53;
   assign m337_53 =10'b0;

   // m337_54 = W*in
   wire signed [9:0] m337_54;
   assign m337_54 =10'b0;

   // m337_55 = W*in
   wire signed [9:0] m337_55;
   assign m337_55 =10'b0;

   // m337_56 = W*in
   wire signed [9:0] m337_56;
   assign m337_56 =10'b0;

   // m337_57 = W*in
   wire signed [9:0] m337_57;
   assign m337_57 =10'b0;

   // m337_58 = W*in
   wire signed [9:0] m337_58;
   assign m337_58 =10'b0;

   // m337_59 = W*in
   wire signed [9:0] m337_59;
   assign m337_59 =10'b0;

   // m337_60 = W*in
   wire signed [9:0] m337_60;
   assign m337_60 =10'b0;

   // m337_61 = W*in
   wire signed [9:0] m337_61;
   assign m337_61 =10'b0;

   // m337_62 = W*in
   wire signed [9:0] m337_62;
   assign m337_62 =10'b0;

   // m337_63 = W*in
   wire signed [9:0] m337_63;
   assign m337_63 =10'b0;

   // m337_64 = W*in
   wire signed [9:0] m337_64;
   assign m337_64 ={ {5{in337[5]}} , in337[5:1] };

   // m337_65 = W*in
   wire signed [9:0] m337_65;
   assign m337_65 =10'b0;

   // m337_66 = W*in
   wire signed [9:0] m337_66;
   assign m337_66 =10'b0;

   // m337_67 = W*in
   wire signed [9:0] m337_67;
   assign m337_67 =10'b0;

   // m337_68 = W*in
   wire signed [9:0] m337_68;
   assign m337_68 =10'b0;

   // m337_69 = W*in
   wire signed [9:0] m337_69;
   assign m337_69 ={ {5{in337[5]}} , in337[5:1] };

   // m337_70 = W*in
   wire signed [9:0] m337_70;
   assign m337_70 =10'b0;

   // m337_71 = W*in
   wire signed [9:0] m337_71;
   assign m337_71 =10'b0;

   // m337_72 = W*in
   wire signed [9:0] m337_72;
   assign m337_72 =10'b0;

   // m337_73 = W*in
   wire signed [9:0] m337_73;
   assign m337_73 =10'b0;

   // m337_74 = W*in
   wire signed [9:0] m337_74;
   assign m337_74 =10'b0;

   // m337_75 = W*in
   wire signed [9:0] m337_75;
   assign m337_75 =10'b0;

   // m337_76 = W*in
   wire signed [9:0] m337_76;
   assign m337_76 =10'b0;

   // m337_77 = W*in
   wire signed [9:0] m337_77;
   assign m337_77 =10'b0;

   // m337_78 = W*in
   wire signed [9:0] m337_78;
   assign m337_78 =10'b0;

   // m337_79 = W*in
   wire signed [9:0] m337_79;
   assign m337_79 =10'b0;

   // m337_80 = W*in
   wire signed [9:0] m337_80;
   assign m337_80 =10'b0;

   // m337_81 = W*in
   wire signed [9:0] m337_81;
   assign m337_81 =10'b0;

   // m337_82 = W*in
   wire signed [9:0] m337_82;
   assign m337_82 =10'b0;

   // m337_83 = W*in
   wire signed [9:0] m337_83;
   assign m337_83 =10'b0;

   // m337_84 = W*in
   wire signed [9:0] m337_84;
   assign m337_84 ={ {5{in337[5]}} , in337[5:1] };

   // m337_85 = W*in
   wire signed [9:0] m337_85;
   assign m337_85 =10'b0;

   // m337_86 = W*in
   wire signed [9:0] m337_86;
   assign m337_86 =10'b0;

   // m337_87 = W*in
   wire signed [9:0] m337_87;
   assign m337_87 =10'b0;

   // m337_88 = W*in
   wire signed [9:0] m337_88;
   assign m337_88 =10'b0;

   // m337_89 = W*in
   wire signed [9:0] m337_89;
   assign m337_89 =10'b0;

   // m337_90 = W*in
   wire signed [9:0] m337_90;
   assign m337_90 =10'b0;

   // m337_91 = W*in
   wire signed [9:0] m337_91;
   assign m337_91 =10'b0;

   // m337_92 = W*in
   wire signed [9:0] m337_92;
   assign m337_92 =10'b0;

   // m337_93 = W*in
   wire signed [9:0] m337_93;
   assign m337_93 =10'b0;

   // m337_94 = W*in
   wire signed [9:0] m337_94;
   assign m337_94 =10'b0;

   // m337_95 = W*in
   wire signed [9:0] m337_95;
   assign m337_95 =10'b0;

   // m337_96 = W*in
   wire signed [9:0] m337_96;
   assign m337_96 =10'b0;

   // m337_97 = W*in
   wire signed [9:0] m337_97;
   assign m337_97 =10'b0;

   // m337_98 = W*in
   wire signed [9:0] m337_98;
   assign m337_98 =10'b0;

   // m337_99 = W*in
   wire signed [9:0] m337_99;
   assign m337_99 =10'b0;

   // m337_100 = W*in
   wire signed [9:0] m337_100;
   assign m337_100 =10'b0;

   // m337_101 = W*in
   wire signed [9:0] m337_101;
   assign m337_101 =10'b0;

   // m337_102 = W*in
   wire signed [9:0] m337_102;
   assign m337_102 =10'b0;

   // m337_103 = W*in
   wire signed [9:0] m337_103;
   assign m337_103 =10'b0;

   // m337_104 = W*in
   wire signed [9:0] m337_104;
   assign m337_104 =10'b0;

   // m337_105 = W*in
   wire signed [9:0] m337_105;
   assign m337_105 =10'b0;

   // m337_106 = W*in
   wire signed [9:0] m337_106;
   assign m337_106 =10'b0;

   // m337_107 = W*in
   wire signed [9:0] m337_107;
   assign m337_107 =10'b0;

   // m337_108 = W*in
   wire signed [9:0] m337_108;
   assign m337_108 =10'b0;

   // m337_109 = W*in
   wire signed [9:0] m337_109;
   assign m337_109 ={ {5{in337[5]}} , in337[5:1] };

   // m337_110 = W*in
   wire signed [9:0] m337_110;
   assign m337_110 =10'b0;

   // m337_111 = W*in
   wire signed [9:0] m337_111;
   assign m337_111 =10'b0;

   // m337_112 = W*in
   wire signed [9:0] m337_112;
   assign m337_112 =10'b0;

   // m337_113 = W*in
   wire signed [9:0] m337_113;
   assign m337_113 =10'b0;

   // m337_114 = W*in
   wire signed [9:0] m337_114;
   assign m337_114 =10'b0;

   // m337_115 = W*in
   wire signed [9:0] m337_115;
   assign m337_115 =10'b0;

   // m337_116 = W*in
   wire signed [9:0] m337_116;
   assign m337_116 ={ {4{in337[5]}} , in337[5:0] };

   // m337_117 = W*in
   wire signed [9:0] m337_117;
   assign m337_117 =10'b0;

   // m338_1 = W*in
   wire signed [9:0] m338_1;
   assign m338_1 ={ {4{in338[5]}} , in338[5:0] };

   // m338_2 = W*in
   wire signed [9:0] m338_2;
   assign m338_2 =10'b0;

   // m338_3 = W*in
   wire signed [9:0] m338_3;
   assign m338_3 =10'b0;

   // m338_4 = W*in
   wire signed [9:0] m338_4;
   assign m338_4 =10'b0;

   // m338_5 = W*in
   wire signed [9:0] m338_5;
   assign m338_5 =10'b0;

   // m338_6 = W*in
   wire signed [9:0] m338_6;
   assign m338_6 =10'b0;

   // m338_7 = W*in
   wire signed [9:0] m338_7;
   assign m338_7 =10'b0;

   // m338_8 = W*in
   wire signed [9:0] m338_8;
   assign m338_8 =10'b0;

   // m338_9 = W*in
   wire signed [9:0] m338_9;
   assign m338_9 =10'b0;

   // m338_10 = W*in
   wire signed [9:0] m338_10;
   assign m338_10 ={ {4{in338[5]}} , in338[5:0] };

   // m338_11 = W*in
   wire signed [9:0] m338_11;
   assign m338_11 =10'b0;

   // m338_12 = W*in
   wire signed [9:0] m338_12;
   assign m338_12 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_13 = W*in
   wire signed [9:0] m338_13;
   assign m338_13 =10'b0;

   // m338_14 = W*in
   wire signed [9:0] m338_14;
   assign m338_14 =10'b0;

   // m338_15 = W*in
   wire signed [9:0] m338_15;
   assign m338_15 =10'b0;

   // m338_16 = W*in
   wire signed [9:0] m338_16;
   assign m338_16 ={ {4{in338[5]}} , in338[5:0] };

   // m338_17 = W*in
   wire signed [9:0] m338_17;
   assign m338_17 =10'b0;

   // m338_18 = W*in
   wire signed [9:0] m338_18;
   assign m338_18 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_19 = W*in
   wire signed [9:0] m338_19;
   assign m338_19 ={ {5{neg338[5]}} , neg338[5:1] };

   // m338_20 = W*in
   wire signed [9:0] m338_20;
   assign m338_20 =10'b0;

   // m338_21 = W*in
   wire signed [9:0] m338_21;
   assign m338_21 =10'b0;

   // m338_22 = W*in
   wire signed [9:0] m338_22;
   assign m338_22 =10'b0;

   // m338_23 = W*in
   wire signed [9:0] m338_23;
   assign m338_23 =10'b0;

   // m338_24 = W*in
   wire signed [9:0] m338_24;
   assign m338_24 =10'b0;

   // m338_25 = W*in
   wire signed [9:0] m338_25;
   assign m338_25 ={ {5{in338[5]}} , in338[5:1] };

   // m338_26 = W*in
   wire signed [9:0] m338_26;
   assign m338_26 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_27 = W*in
   wire signed [9:0] m338_27;
   assign m338_27 =10'b0;

   // m338_28 = W*in
   wire signed [9:0] m338_28;
   assign m338_28 =10'b0;

   // m338_29 = W*in
   wire signed [9:0] m338_29;
   assign m338_29 =10'b0;

   // m338_30 = W*in
   wire signed [9:0] m338_30;
   assign m338_30 =10'b0;

   // m338_31 = W*in
   wire signed [9:0] m338_31;
   assign m338_31 =10'b0;

   // m338_32 = W*in
   wire signed [9:0] m338_32;
   assign m338_32 =10'b0;

   // m338_33 = W*in
   wire signed [9:0] m338_33;
   assign m338_33 =10'b0;

   // m338_34 = W*in
   wire signed [9:0] m338_34;
   assign m338_34 ={ {5{neg338[5]}} , neg338[5:1] };

   // m338_35 = W*in
   wire signed [9:0] m338_35;
   assign m338_35 ={ {5{neg338[5]}} , neg338[5:1] };

   // m338_36 = W*in
   wire signed [9:0] m338_36;
   assign m338_36 =10'b0;

   // m338_37 = W*in
   wire signed [9:0] m338_37;
   assign m338_37 ={ {4{in338[5]}} , in338[5:0] };

   // m338_38 = W*in
   wire signed [9:0] m338_38;
   assign m338_38 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_39 = W*in
   wire signed [9:0] m338_39;
   assign m338_39 =10'b0;

   // m338_40 = W*in
   wire signed [9:0] m338_40;
   assign m338_40 =10'b0;

   // m338_41 = W*in
   wire signed [9:0] m338_41;
   assign m338_41 ={ {3{in338[5]}} , in338 , {1{1'b0}} };

   // m338_42 = W*in
   wire signed [9:0] m338_42;
   assign m338_42 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_43 = W*in
   wire signed [9:0] m338_43;
   assign m338_43 =10'b0;

   // m338_44 = W*in
   wire signed [9:0] m338_44;
   assign m338_44 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_45 = W*in
   wire signed [9:0] m338_45;
   assign m338_45 ={ {4{in338[5]}} , in338[5:0] };

   // m338_46 = W*in
   wire signed [9:0] m338_46;
   assign m338_46 =10'b0;

   // m338_47 = W*in
   wire signed [9:0] m338_47;
   assign m338_47 =10'b0;

   // m338_48 = W*in
   wire signed [9:0] m338_48;
   assign m338_48 =10'b0;

   // m338_49 = W*in
   wire signed [9:0] m338_49;
   assign m338_49 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_50 = W*in
   wire signed [9:0] m338_50;
   assign m338_50 =10'b0;

   // m338_51 = W*in
   wire signed [9:0] m338_51;
   assign m338_51 =10'b0;

   // m338_52 = W*in
   wire signed [9:0] m338_52;
   assign m338_52 =10'b0;

   // m338_53 = W*in
   wire signed [9:0] m338_53;
   assign m338_53 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_54 = W*in
   wire signed [9:0] m338_54;
   assign m338_54 =10'b0;

   // m338_55 = W*in
   wire signed [9:0] m338_55;
   assign m338_55 =10'b0;

   // m338_56 = W*in
   wire signed [9:0] m338_56;
   assign m338_56 ={ {4{in338[5]}} , in338[5:0] };

   // m338_57 = W*in
   wire signed [9:0] m338_57;
   assign m338_57 =10'b0;

   // m338_58 = W*in
   wire signed [9:0] m338_58;
   assign m338_58 =10'b0;

   // m338_59 = W*in
   wire signed [9:0] m338_59;
   assign m338_59 =10'b0;

   // m338_60 = W*in
   wire signed [9:0] m338_60;
   assign m338_60 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_61 = W*in
   wire signed [9:0] m338_61;
   assign m338_61 =10'b0;

   // m338_62 = W*in
   wire signed [9:0] m338_62;
   assign m338_62 =10'b0;

   // m338_63 = W*in
   wire signed [9:0] m338_63;
   assign m338_63 =10'b0;

   // m338_64 = W*in
   wire signed [9:0] m338_64;
   assign m338_64 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_65 = W*in
   wire signed [9:0] m338_65;
   assign m338_65 =10'b0;

   // m338_66 = W*in
   wire signed [9:0] m338_66;
   assign m338_66 =10'b0;

   // m338_67 = W*in
   wire signed [9:0] m338_67;
   assign m338_67 =10'b0;

   // m338_68 = W*in
   wire signed [9:0] m338_68;
   assign m338_68 =10'b0;

   // m338_69 = W*in
   wire signed [9:0] m338_69;
   assign m338_69 =10'b0;

   // m338_70 = W*in
   wire signed [9:0] m338_70;
   assign m338_70 =10'b0;

   // m338_71 = W*in
   wire signed [9:0] m338_71;
   assign m338_71 ={ {5{neg338[5]}} , neg338[5:1] };

   // m338_72 = W*in
   wire signed [9:0] m338_72;
   assign m338_72 =10'b0;

   // m338_73 = W*in
   wire signed [9:0] m338_73;
   assign m338_73 =10'b0;

   // m338_74 = W*in
   wire signed [9:0] m338_74;
   assign m338_74 =10'b0;

   // m338_75 = W*in
   wire signed [9:0] m338_75;
   assign m338_75 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_76 = W*in
   wire signed [9:0] m338_76;
   assign m338_76 =10'b0;

   // m338_77 = W*in
   wire signed [9:0] m338_77;
   assign m338_77 =10'b0;

   // m338_78 = W*in
   wire signed [9:0] m338_78;
   assign m338_78 =10'b0;

   // m338_79 = W*in
   wire signed [9:0] m338_79;
   assign m338_79 =10'b0;

   // m338_80 = W*in
   wire signed [9:0] m338_80;
   assign m338_80 =10'b0;

   // m338_81 = W*in
   wire signed [9:0] m338_81;
   assign m338_81 =10'b0;

   // m338_82 = W*in
   wire signed [9:0] m338_82;
   assign m338_82 ={ {4{in338[5]}} , in338[5:0] };

   // m338_83 = W*in
   wire signed [9:0] m338_83;
   assign m338_83 =10'b0;

   // m338_84 = W*in
   wire signed [9:0] m338_84;
   assign m338_84 ={ {5{in338[5]}} , in338[5:1] };

   // m338_85 = W*in
   wire signed [9:0] m338_85;
   assign m338_85 ={ {4{in338[5]}} , in338[5:0] };

   // m338_86 = W*in
   wire signed [9:0] m338_86;
   assign m338_86 =10'b0;

   // m338_87 = W*in
   wire signed [9:0] m338_87;
   assign m338_87 =10'b0;

   // m338_88 = W*in
   wire signed [9:0] m338_88;
   assign m338_88 =10'b0;

   // m338_89 = W*in
   wire signed [9:0] m338_89;
   assign m338_89 ={ {4{in338[5]}} , in338[5:0] };

   // m338_90 = W*in
   wire signed [9:0] m338_90;
   assign m338_90 =10'b0;

   // m338_91 = W*in
   wire signed [9:0] m338_91;
   assign m338_91 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_92 = W*in
   wire signed [9:0] m338_92;
   assign m338_92 =10'b0;

   // m338_93 = W*in
   wire signed [9:0] m338_93;
   assign m338_93 =10'b0;

   // m338_94 = W*in
   wire signed [9:0] m338_94;
   assign m338_94 =10'b0;

   // m338_95 = W*in
   wire signed [9:0] m338_95;
   assign m338_95 =10'b0;

   // m338_96 = W*in
   wire signed [9:0] m338_96;
   assign m338_96 ={ {4{in338[5]}} , in338[5:0] };

   // m338_97 = W*in
   wire signed [9:0] m338_97;
   assign m338_97 ={ {4{neg338[5]}} , neg338[5:0] };

   // m338_98 = W*in
   wire signed [9:0] m338_98;
   assign m338_98 =10'b0;

   // m338_99 = W*in
   wire signed [9:0] m338_99;
   assign m338_99 =10'b0;

   // m338_100 = W*in
   wire signed [9:0] m338_100;
   assign m338_100 =10'b0;

   // m338_101 = W*in
   wire signed [9:0] m338_101;
   assign m338_101 =10'b0;

   // m338_102 = W*in
   wire signed [9:0] m338_102;
   assign m338_102 =10'b0;

   // m338_103 = W*in
   wire signed [9:0] m338_103;
   assign m338_103 =10'b0;

   // m338_104 = W*in
   wire signed [9:0] m338_104;
   assign m338_104 =10'b0;

   // m338_105 = W*in
   wire signed [9:0] m338_105;
   assign m338_105 =10'b0;

   // m338_106 = W*in
   wire signed [9:0] m338_106;
   assign m338_106 =10'b0;

   // m338_107 = W*in
   wire signed [9:0] m338_107;
   assign m338_107 =10'b0;

   // m338_108 = W*in
   wire signed [9:0] m338_108;
   assign m338_108 =10'b0;

   // m338_109 = W*in
   wire signed [9:0] m338_109;
   assign m338_109 ={ {4{in338[5]}} , in338[5:0] };

   // m338_110 = W*in
   wire signed [9:0] m338_110;
   assign m338_110 =10'b0;

   // m338_111 = W*in
   wire signed [9:0] m338_111;
   assign m338_111 ={ {4{in338[5]}} , in338[5:0] };

   // m338_112 = W*in
   wire signed [9:0] m338_112;
   assign m338_112 =10'b0;

   // m338_113 = W*in
   wire signed [9:0] m338_113;
   assign m338_113 =10'b0;

   // m338_114 = W*in
   wire signed [9:0] m338_114;
   assign m338_114 =10'b0;

   // m338_115 = W*in
   wire signed [9:0] m338_115;
   assign m338_115 ={ {5{neg338[5]}} , neg338[5:1] };

   // m338_116 = W*in
   wire signed [9:0] m338_116;
   assign m338_116 ={ {4{in338[5]}} , in338[5:0] };

   // m338_117 = W*in
   wire signed [9:0] m338_117;
   assign m338_117 ={ {4{neg338[5]}} , neg338[5:0] };

   // m339_1 = W*in
   wire signed [9:0] m339_1;
   assign m339_1 =10'b0;

   // m339_2 = W*in
   wire signed [9:0] m339_2;
   assign m339_2 =10'b0;

   // m339_3 = W*in
   wire signed [9:0] m339_3;
   assign m339_3 =10'b0;

   // m339_4 = W*in
   wire signed [9:0] m339_4;
   assign m339_4 =10'b0;

   // m339_5 = W*in
   wire signed [9:0] m339_5;
   assign m339_5 =10'b0;

   // m339_6 = W*in
   wire signed [9:0] m339_6;
   assign m339_6 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_7 = W*in
   wire signed [9:0] m339_7;
   assign m339_7 =10'b0;

   // m339_8 = W*in
   wire signed [9:0] m339_8;
   assign m339_8 =10'b0;

   // m339_9 = W*in
   wire signed [9:0] m339_9;
   assign m339_9 =10'b0;

   // m339_10 = W*in
   wire signed [9:0] m339_10;
   assign m339_10 ={ {4{in339[5]}} , in339[5:0] };

   // m339_11 = W*in
   wire signed [9:0] m339_11;
   assign m339_11 =10'b0;

   // m339_12 = W*in
   wire signed [9:0] m339_12;
   assign m339_12 ={ {4{in339[5]}} , in339[5:0] };

   // m339_13 = W*in
   wire signed [9:0] m339_13;
   assign m339_13 =10'b0;

   // m339_14 = W*in
   wire signed [9:0] m339_14;
   assign m339_14 ={ {4{in339[5]}} , in339[5:0] };

   // m339_15 = W*in
   wire signed [9:0] m339_15;
   assign m339_15 =10'b0;

   // m339_16 = W*in
   wire signed [9:0] m339_16;
   assign m339_16 =10'b0;

   // m339_17 = W*in
   wire signed [9:0] m339_17;
   assign m339_17 ={ {5{neg339[5]}} , neg339[5:1] };

   // m339_18 = W*in
   wire signed [9:0] m339_18;
   assign m339_18 ={ {3{in339[5]}} , in339 , {1{1'b0}} };

   // m339_19 = W*in
   wire signed [9:0] m339_19;
   assign m339_19 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_20 = W*in
   wire signed [9:0] m339_20;
   assign m339_20 ={ {3{neg339[5]}} , neg339 , {1{1'b0}} };

   // m339_21 = W*in
   wire signed [9:0] m339_21;
   assign m339_21 ={ {5{in339[5]}} , in339[5:1] };

   // m339_22 = W*in
   wire signed [9:0] m339_22;
   assign m339_22 =10'b0;

   // m339_23 = W*in
   wire signed [9:0] m339_23;
   assign m339_23 =10'b0;

   // m339_24 = W*in
   wire signed [9:0] m339_24;
   assign m339_24 =10'b0;

   // m339_25 = W*in
   wire signed [9:0] m339_25;
   assign m339_25 ={ {5{in339[5]}} , in339[5:1] };

   // m339_26 = W*in
   wire signed [9:0] m339_26;
   assign m339_26 ={ {3{in339[5]}} , in339 , {1{1'b0}} };

   // m339_27 = W*in
   wire signed [9:0] m339_27;
   assign m339_27 =10'b0;

   // m339_28 = W*in
   wire signed [9:0] m339_28;
   assign m339_28 =10'b0;

   // m339_29 = W*in
   wire signed [9:0] m339_29;
   assign m339_29 =10'b0;

   // m339_30 = W*in
   wire signed [9:0] m339_30;
   assign m339_30 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_31 = W*in
   wire signed [9:0] m339_31;
   assign m339_31 =10'b0;

   // m339_32 = W*in
   wire signed [9:0] m339_32;
   assign m339_32 =10'b0;

   // m339_33 = W*in
   wire signed [9:0] m339_33;
   assign m339_33 =10'b0;

   // m339_34 = W*in
   wire signed [9:0] m339_34;
   assign m339_34 ={ {5{neg339[5]}} , neg339[5:1] };

   // m339_35 = W*in
   wire signed [9:0] m339_35;
   assign m339_35 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_36 = W*in
   wire signed [9:0] m339_36;
   assign m339_36 =10'b0;

   // m339_37 = W*in
   wire signed [9:0] m339_37;
   assign m339_37 =10'b0;

   // m339_38 = W*in
   wire signed [9:0] m339_38;
   assign m339_38 =10'b0;

   // m339_39 = W*in
   wire signed [9:0] m339_39;
   assign m339_39 =10'b0;

   // m339_40 = W*in
   wire signed [9:0] m339_40;
   assign m339_40 =10'b0;

   // m339_41 = W*in
   wire signed [9:0] m339_41;
   assign m339_41 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_42 = W*in
   wire signed [9:0] m339_42;
   assign m339_42 ={ {4{in339[5]}} , in339[5:0] };

   // m339_43 = W*in
   wire signed [9:0] m339_43;
   assign m339_43 =10'b0;

   // m339_44 = W*in
   wire signed [9:0] m339_44;
   assign m339_44 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_45 = W*in
   wire signed [9:0] m339_45;
   assign m339_45 =10'b0;

   // m339_46 = W*in
   wire signed [9:0] m339_46;
   assign m339_46 =10'b0;

   // m339_47 = W*in
   wire signed [9:0] m339_47;
   assign m339_47 =10'b0;

   // m339_48 = W*in
   wire signed [9:0] m339_48;
   assign m339_48 =10'b0;

   // m339_49 = W*in
   wire signed [9:0] m339_49;
   assign m339_49 =10'b0;

   // m339_50 = W*in
   wire signed [9:0] m339_50;
   assign m339_50 =10'b0;

   // m339_51 = W*in
   wire signed [9:0] m339_51;
   assign m339_51 ={ {4{in339[5]}} , in339[5:0] };

   // m339_52 = W*in
   wire signed [9:0] m339_52;
   assign m339_52 =10'b0;

   // m339_53 = W*in
   wire signed [9:0] m339_53;
   assign m339_53 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_54 = W*in
   wire signed [9:0] m339_54;
   assign m339_54 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_55 = W*in
   wire signed [9:0] m339_55;
   assign m339_55 ={ {4{in339[5]}} , in339[5:0] };

   // m339_56 = W*in
   wire signed [9:0] m339_56;
   assign m339_56 =10'b0;

   // m339_57 = W*in
   wire signed [9:0] m339_57;
   assign m339_57 =10'b0;

   // m339_58 = W*in
   wire signed [9:0] m339_58;
   assign m339_58 =10'b0;

   // m339_59 = W*in
   wire signed [9:0] m339_59;
   assign m339_59 =10'b0;

   // m339_60 = W*in
   wire signed [9:0] m339_60;
   assign m339_60 ={ {3{neg339[5]}} , neg339 , {1{1'b0}} };

   // m339_61 = W*in
   wire signed [9:0] m339_61;
   assign m339_61 =10'b0;

   // m339_62 = W*in
   wire signed [9:0] m339_62;
   assign m339_62 =10'b0;

   // m339_63 = W*in
   wire signed [9:0] m339_63;
   assign m339_63 =10'b0;

   // m339_64 = W*in
   wire signed [9:0] m339_64;
   assign m339_64 ={ {5{in339[5]}} , in339[5:1] };

   // m339_65 = W*in
   wire signed [9:0] m339_65;
   assign m339_65 =10'b0;

   // m339_66 = W*in
   wire signed [9:0] m339_66;
   assign m339_66 ={ {5{in339[5]}} , in339[5:1] };

   // m339_67 = W*in
   wire signed [9:0] m339_67;
   assign m339_67 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_68 = W*in
   wire signed [9:0] m339_68;
   assign m339_68 =10'b0;

   // m339_69 = W*in
   wire signed [9:0] m339_69;
   assign m339_69 ={ {5{in339[5]}} , in339[5:1] };

   // m339_70 = W*in
   wire signed [9:0] m339_70;
   assign m339_70 ={ {4{in339[5]}} , in339[5:0] };

   // m339_71 = W*in
   wire signed [9:0] m339_71;
   assign m339_71 =10'b0;

   // m339_72 = W*in
   wire signed [9:0] m339_72;
   assign m339_72 ={ {4{in339[5]}} , in339[5:0] };

   // m339_73 = W*in
   wire signed [9:0] m339_73;
   assign m339_73 =10'b0;

   // m339_74 = W*in
   wire signed [9:0] m339_74;
   assign m339_74 =10'b0;

   // m339_75 = W*in
   wire signed [9:0] m339_75;
   assign m339_75 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_76 = W*in
   wire signed [9:0] m339_76;
   assign m339_76 =10'b0;

   // m339_77 = W*in
   wire signed [9:0] m339_77;
   assign m339_77 ={ {3{in339[5]}} , in339 , {1{1'b0}} };

   // m339_78 = W*in
   wire signed [9:0] m339_78;
   assign m339_78 =10'b0;

   // m339_79 = W*in
   wire signed [9:0] m339_79;
   assign m339_79 =10'b0;

   // m339_80 = W*in
   wire signed [9:0] m339_80;
   assign m339_80 ={ {5{neg339[5]}} , neg339[5:1] };

   // m339_81 = W*in
   wire signed [9:0] m339_81;
   assign m339_81 ={ {5{in339[5]}} , in339[5:1] };

   // m339_82 = W*in
   wire signed [9:0] m339_82;
   assign m339_82 =10'b0;

   // m339_83 = W*in
   wire signed [9:0] m339_83;
   assign m339_83 =10'b0;

   // m339_84 = W*in
   wire signed [9:0] m339_84;
   assign m339_84 ={ {4{in339[5]}} , in339[5:0] };

   // m339_85 = W*in
   wire signed [9:0] m339_85;
   assign m339_85 =10'b0;

   // m339_86 = W*in
   wire signed [9:0] m339_86;
   assign m339_86 ={ {3{in339[5]}} , in339 , {1{1'b0}} };

   // m339_87 = W*in
   wire signed [9:0] m339_87;
   assign m339_87 =10'b0;

   // m339_88 = W*in
   wire signed [9:0] m339_88;
   assign m339_88 =10'b0;

   // m339_89 = W*in
   wire signed [9:0] m339_89;
   assign m339_89 =10'b0;

   // m339_90 = W*in
   wire signed [9:0] m339_90;
   assign m339_90 =10'b0;

   // m339_91 = W*in
   wire signed [9:0] m339_91;
   assign m339_91 =10'b0;

   // m339_92 = W*in
   wire signed [9:0] m339_92;
   assign m339_92 =10'b0;

   // m339_93 = W*in
   wire signed [9:0] m339_93;
   assign m339_93 =10'b0;

   // m339_94 = W*in
   wire signed [9:0] m339_94;
   assign m339_94 =10'b0;

   // m339_95 = W*in
   wire signed [9:0] m339_95;
   assign m339_95 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_96 = W*in
   wire signed [9:0] m339_96;
   assign m339_96 ={ {4{in339[5]}} , in339[5:0] };

   // m339_97 = W*in
   wire signed [9:0] m339_97;
   assign m339_97 =10'b0;

   // m339_98 = W*in
   wire signed [9:0] m339_98;
   assign m339_98 =10'b0;

   // m339_99 = W*in
   wire signed [9:0] m339_99;
   assign m339_99 ={ {4{in339[5]}} , in339[5:0] };

   // m339_100 = W*in
   wire signed [9:0] m339_100;
   assign m339_100 ={ {4{in339[5]}} , in339[5:0] };

   // m339_101 = W*in
   wire signed [9:0] m339_101;
   assign m339_101 =10'b0;

   // m339_102 = W*in
   wire signed [9:0] m339_102;
   assign m339_102 =10'b0;

   // m339_103 = W*in
   wire signed [9:0] m339_103;
   assign m339_103 =10'b0;

   // m339_104 = W*in
   wire signed [9:0] m339_104;
   assign m339_104 =10'b0;

   // m339_105 = W*in
   wire signed [9:0] m339_105;
   assign m339_105 =10'b0;

   // m339_106 = W*in
   wire signed [9:0] m339_106;
   assign m339_106 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_107 = W*in
   wire signed [9:0] m339_107;
   assign m339_107 =10'b0;

   // m339_108 = W*in
   wire signed [9:0] m339_108;
   assign m339_108 =10'b0;

   // m339_109 = W*in
   wire signed [9:0] m339_109;
   assign m339_109 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_110 = W*in
   wire signed [9:0] m339_110;
   assign m339_110 ={ {4{in339[5]}} , in339[5:0] };

   // m339_111 = W*in
   wire signed [9:0] m339_111;
   assign m339_111 ={ {4{in339[5]}} , in339[5:0] };

   // m339_112 = W*in
   wire signed [9:0] m339_112;
   assign m339_112 =10'b0;

   // m339_113 = W*in
   wire signed [9:0] m339_113;
   assign m339_113 =10'b0;

   // m339_114 = W*in
   wire signed [9:0] m339_114;
   assign m339_114 =10'b0;

   // m339_115 = W*in
   wire signed [9:0] m339_115;
   assign m339_115 ={ {4{neg339[5]}} , neg339[5:0] };

   // m339_116 = W*in
   wire signed [9:0] m339_116;
   assign m339_116 =10'b0;

   // m339_117 = W*in
   wire signed [9:0] m339_117;
   assign m339_117 ={ {4{neg339[5]}} , neg339[5:0] };

   // m340_1 = W*in
   wire signed [9:0] m340_1;
   assign m340_1 ={ {4{in340[5]}} , in340[5:0] };

   // m340_2 = W*in
   wire signed [9:0] m340_2;
   assign m340_2 =10'b0;

   // m340_3 = W*in
   wire signed [9:0] m340_3;
   assign m340_3 =10'b0;

   // m340_4 = W*in
   wire signed [9:0] m340_4;
   assign m340_4 =10'b0;

   // m340_5 = W*in
   wire signed [9:0] m340_5;
   assign m340_5 =10'b0;

   // m340_6 = W*in
   wire signed [9:0] m340_6;
   assign m340_6 =10'b0;

   // m340_7 = W*in
   wire signed [9:0] m340_7;
   assign m340_7 =10'b0;

   // m340_8 = W*in
   wire signed [9:0] m340_8;
   assign m340_8 =10'b0;

   // m340_9 = W*in
   wire signed [9:0] m340_9;
   assign m340_9 =10'b0;

   // m340_10 = W*in
   wire signed [9:0] m340_10;
   assign m340_10 =10'b0;

   // m340_11 = W*in
   wire signed [9:0] m340_11;
   assign m340_11 =10'b0;

   // m340_12 = W*in
   wire signed [9:0] m340_12;
   assign m340_12 =10'b0;

   // m340_13 = W*in
   wire signed [9:0] m340_13;
   assign m340_13 ={ {4{in340[5]}} , in340[5:0] };

   // m340_14 = W*in
   wire signed [9:0] m340_14;
   assign m340_14 =10'b0;

   // m340_15 = W*in
   wire signed [9:0] m340_15;
   assign m340_15 =10'b0;

   // m340_16 = W*in
   wire signed [9:0] m340_16;
   assign m340_16 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_17 = W*in
   wire signed [9:0] m340_17;
   assign m340_17 =10'b0;

   // m340_18 = W*in
   wire signed [9:0] m340_18;
   assign m340_18 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_19 = W*in
   wire signed [9:0] m340_19;
   assign m340_19 =10'b0;

   // m340_20 = W*in
   wire signed [9:0] m340_20;
   assign m340_20 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_21 = W*in
   wire signed [9:0] m340_21;
   assign m340_21 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_22 = W*in
   wire signed [9:0] m340_22;
   assign m340_22 =10'b0;

   // m340_23 = W*in
   wire signed [9:0] m340_23;
   assign m340_23 =10'b0;

   // m340_24 = W*in
   wire signed [9:0] m340_24;
   assign m340_24 ={ {4{in340[5]}} , in340[5:0] };

   // m340_25 = W*in
   wire signed [9:0] m340_25;
   assign m340_25 ={ {4{in340[5]}} , in340[5:0] };

   // m340_26 = W*in
   wire signed [9:0] m340_26;
   assign m340_26 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_27 = W*in
   wire signed [9:0] m340_27;
   assign m340_27 ={ {5{in340[5]}} , in340[5:1] };

   // m340_28 = W*in
   wire signed [9:0] m340_28;
   assign m340_28 =10'b0;

   // m340_29 = W*in
   wire signed [9:0] m340_29;
   assign m340_29 =10'b0;

   // m340_30 = W*in
   wire signed [9:0] m340_30;
   assign m340_30 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_31 = W*in
   wire signed [9:0] m340_31;
   assign m340_31 =10'b0;

   // m340_32 = W*in
   wire signed [9:0] m340_32;
   assign m340_32 =10'b0;

   // m340_33 = W*in
   wire signed [9:0] m340_33;
   assign m340_33 ={ {4{in340[5]}} , in340[5:0] };

   // m340_34 = W*in
   wire signed [9:0] m340_34;
   assign m340_34 =10'b0;

   // m340_35 = W*in
   wire signed [9:0] m340_35;
   assign m340_35 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_36 = W*in
   wire signed [9:0] m340_36;
   assign m340_36 =10'b0;

   // m340_37 = W*in
   wire signed [9:0] m340_37;
   assign m340_37 =10'b0;

   // m340_38 = W*in
   wire signed [9:0] m340_38;
   assign m340_38 =10'b0;

   // m340_39 = W*in
   wire signed [9:0] m340_39;
   assign m340_39 ={ {4{in340[5]}} , in340[5:0] };

   // m340_40 = W*in
   wire signed [9:0] m340_40;
   assign m340_40 =10'b0;

   // m340_41 = W*in
   wire signed [9:0] m340_41;
   assign m340_41 =10'b0;

   // m340_42 = W*in
   wire signed [9:0] m340_42;
   assign m340_42 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_43 = W*in
   wire signed [9:0] m340_43;
   assign m340_43 =10'b0;

   // m340_44 = W*in
   wire signed [9:0] m340_44;
   assign m340_44 =10'b0;

   // m340_45 = W*in
   wire signed [9:0] m340_45;
   assign m340_45 =10'b0;

   // m340_46 = W*in
   wire signed [9:0] m340_46;
   assign m340_46 ={ {4{in340[5]}} , in340[5:0] };

   // m340_47 = W*in
   wire signed [9:0] m340_47;
   assign m340_47 =10'b0;

   // m340_48 = W*in
   wire signed [9:0] m340_48;
   assign m340_48 =10'b0;

   // m340_49 = W*in
   wire signed [9:0] m340_49;
   assign m340_49 =10'b0;

   // m340_50 = W*in
   wire signed [9:0] m340_50;
   assign m340_50 =10'b0;

   // m340_51 = W*in
   wire signed [9:0] m340_51;
   assign m340_51 =10'b0;

   // m340_52 = W*in
   wire signed [9:0] m340_52;
   assign m340_52 =10'b0;

   // m340_53 = W*in
   wire signed [9:0] m340_53;
   assign m340_53 =10'b0;

   // m340_54 = W*in
   wire signed [9:0] m340_54;
   assign m340_54 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_55 = W*in
   wire signed [9:0] m340_55;
   assign m340_55 =10'b0;

   // m340_56 = W*in
   wire signed [9:0] m340_56;
   assign m340_56 =10'b0;

   // m340_57 = W*in
   wire signed [9:0] m340_57;
   assign m340_57 =10'b0;

   // m340_58 = W*in
   wire signed [9:0] m340_58;
   assign m340_58 =10'b0;

   // m340_59 = W*in
   wire signed [9:0] m340_59;
   assign m340_59 ={ {4{in340[5]}} , in340[5:0] };

   // m340_60 = W*in
   wire signed [9:0] m340_60;
   assign m340_60 =10'b0;

   // m340_61 = W*in
   wire signed [9:0] m340_61;
   assign m340_61 =10'b0;

   // m340_62 = W*in
   wire signed [9:0] m340_62;
   assign m340_62 =10'b0;

   // m340_63 = W*in
   wire signed [9:0] m340_63;
   assign m340_63 =10'b0;

   // m340_64 = W*in
   wire signed [9:0] m340_64;
   assign m340_64 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_65 = W*in
   wire signed [9:0] m340_65;
   assign m340_65 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_66 = W*in
   wire signed [9:0] m340_66;
   assign m340_66 =10'b0;

   // m340_67 = W*in
   wire signed [9:0] m340_67;
   assign m340_67 =10'b0;

   // m340_68 = W*in
   wire signed [9:0] m340_68;
   assign m340_68 =10'b0;

   // m340_69 = W*in
   wire signed [9:0] m340_69;
   assign m340_69 =10'b0;

   // m340_70 = W*in
   wire signed [9:0] m340_70;
   assign m340_70 =10'b0;

   // m340_71 = W*in
   wire signed [9:0] m340_71;
   assign m340_71 =10'b0;

   // m340_72 = W*in
   wire signed [9:0] m340_72;
   assign m340_72 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_73 = W*in
   wire signed [9:0] m340_73;
   assign m340_73 ={ {4{in340[5]}} , in340[5:0] };

   // m340_74 = W*in
   wire signed [9:0] m340_74;
   assign m340_74 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_75 = W*in
   wire signed [9:0] m340_75;
   assign m340_75 =10'b0;

   // m340_76 = W*in
   wire signed [9:0] m340_76;
   assign m340_76 =10'b0;

   // m340_77 = W*in
   wire signed [9:0] m340_77;
   assign m340_77 =10'b0;

   // m340_78 = W*in
   wire signed [9:0] m340_78;
   assign m340_78 =10'b0;

   // m340_79 = W*in
   wire signed [9:0] m340_79;
   assign m340_79 =10'b0;

   // m340_80 = W*in
   wire signed [9:0] m340_80;
   assign m340_80 ={ {4{in340[5]}} , in340[5:0] };

   // m340_81 = W*in
   wire signed [9:0] m340_81;
   assign m340_81 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_82 = W*in
   wire signed [9:0] m340_82;
   assign m340_82 =10'b0;

   // m340_83 = W*in
   wire signed [9:0] m340_83;
   assign m340_83 ={ {5{neg340[5]}} , neg340[5:1] };

   // m340_84 = W*in
   wire signed [9:0] m340_84;
   assign m340_84 =10'b0;

   // m340_85 = W*in
   wire signed [9:0] m340_85;
   assign m340_85 =10'b0;

   // m340_86 = W*in
   wire signed [9:0] m340_86;
   assign m340_86 =10'b0;

   // m340_87 = W*in
   wire signed [9:0] m340_87;
   assign m340_87 =10'b0;

   // m340_88 = W*in
   wire signed [9:0] m340_88;
   assign m340_88 =10'b0;

   // m340_89 = W*in
   wire signed [9:0] m340_89;
   assign m340_89 =10'b0;

   // m340_90 = W*in
   wire signed [9:0] m340_90;
   assign m340_90 =10'b0;

   // m340_91 = W*in
   wire signed [9:0] m340_91;
   assign m340_91 ={ {4{in340[5]}} , in340[5:0] };

   // m340_92 = W*in
   wire signed [9:0] m340_92;
   assign m340_92 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_93 = W*in
   wire signed [9:0] m340_93;
   assign m340_93 =10'b0;

   // m340_94 = W*in
   wire signed [9:0] m340_94;
   assign m340_94 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_95 = W*in
   wire signed [9:0] m340_95;
   assign m340_95 =10'b0;

   // m340_96 = W*in
   wire signed [9:0] m340_96;
   assign m340_96 =10'b0;

   // m340_97 = W*in
   wire signed [9:0] m340_97;
   assign m340_97 =10'b0;

   // m340_98 = W*in
   wire signed [9:0] m340_98;
   assign m340_98 =10'b0;

   // m340_99 = W*in
   wire signed [9:0] m340_99;
   assign m340_99 =10'b0;

   // m340_100 = W*in
   wire signed [9:0] m340_100;
   assign m340_100 =10'b0;

   // m340_101 = W*in
   wire signed [9:0] m340_101;
   assign m340_101 =10'b0;

   // m340_102 = W*in
   wire signed [9:0] m340_102;
   assign m340_102 =10'b0;

   // m340_103 = W*in
   wire signed [9:0] m340_103;
   assign m340_103 =10'b0;

   // m340_104 = W*in
   wire signed [9:0] m340_104;
   assign m340_104 =10'b0;

   // m340_105 = W*in
   wire signed [9:0] m340_105;
   assign m340_105 =10'b0;

   // m340_106 = W*in
   wire signed [9:0] m340_106;
   assign m340_106 =10'b0;

   // m340_107 = W*in
   wire signed [9:0] m340_107;
   assign m340_107 =10'b0;

   // m340_108 = W*in
   wire signed [9:0] m340_108;
   assign m340_108 =10'b0;

   // m340_109 = W*in
   wire signed [9:0] m340_109;
   assign m340_109 ={ {5{in340[5]}} , in340[5:1] };

   // m340_110 = W*in
   wire signed [9:0] m340_110;
   assign m340_110 =10'b0;

   // m340_111 = W*in
   wire signed [9:0] m340_111;
   assign m340_111 =10'b0;

   // m340_112 = W*in
   wire signed [9:0] m340_112;
   assign m340_112 =10'b0;

   // m340_113 = W*in
   wire signed [9:0] m340_113;
   assign m340_113 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_114 = W*in
   wire signed [9:0] m340_114;
   assign m340_114 =10'b0;

   // m340_115 = W*in
   wire signed [9:0] m340_115;
   assign m340_115 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_116 = W*in
   wire signed [9:0] m340_116;
   assign m340_116 ={ {4{neg340[5]}} , neg340[5:0] };

   // m340_117 = W*in
   wire signed [9:0] m340_117;
   assign m340_117 =10'b0;

   // m341_1 = W*in
   wire signed [9:0] m341_1;
   assign m341_1 =10'b0;

   // m341_2 = W*in
   wire signed [9:0] m341_2;
   assign m341_2 =10'b0;

   // m341_3 = W*in
   wire signed [9:0] m341_3;
   assign m341_3 =10'b0;

   // m341_4 = W*in
   wire signed [9:0] m341_4;
   assign m341_4 =10'b0;

   // m341_5 = W*in
   wire signed [9:0] m341_5;
   assign m341_5 =10'b0;

   // m341_6 = W*in
   wire signed [9:0] m341_6;
   assign m341_6 =10'b0;

   // m341_7 = W*in
   wire signed [9:0] m341_7;
   assign m341_7 =10'b0;

   // m341_8 = W*in
   wire signed [9:0] m341_8;
   assign m341_8 =10'b0;

   // m341_9 = W*in
   wire signed [9:0] m341_9;
   assign m341_9 =10'b0;

   // m341_10 = W*in
   wire signed [9:0] m341_10;
   assign m341_10 =10'b0;

   // m341_11 = W*in
   wire signed [9:0] m341_11;
   assign m341_11 =10'b0;

   // m341_12 = W*in
   wire signed [9:0] m341_12;
   assign m341_12 =10'b0;

   // m341_13 = W*in
   wire signed [9:0] m341_13;
   assign m341_13 =10'b0;

   // m341_14 = W*in
   wire signed [9:0] m341_14;
   assign m341_14 =10'b0;

   // m341_15 = W*in
   wire signed [9:0] m341_15;
   assign m341_15 =10'b0;

   // m341_16 = W*in
   wire signed [9:0] m341_16;
   assign m341_16 =10'b0;

   // m341_17 = W*in
   wire signed [9:0] m341_17;
   assign m341_17 =10'b0;

   // m341_18 = W*in
   wire signed [9:0] m341_18;
   assign m341_18 =10'b0;

   // m341_19 = W*in
   wire signed [9:0] m341_19;
   assign m341_19 =10'b0;

   // m341_20 = W*in
   wire signed [9:0] m341_20;
   assign m341_20 =10'b0;

   // m341_21 = W*in
   wire signed [9:0] m341_21;
   assign m341_21 =10'b0;

   // m341_22 = W*in
   wire signed [9:0] m341_22;
   assign m341_22 =10'b0;

   // m341_23 = W*in
   wire signed [9:0] m341_23;
   assign m341_23 =10'b0;

   // m341_24 = W*in
   wire signed [9:0] m341_24;
   assign m341_24 =10'b0;

   // m341_25 = W*in
   wire signed [9:0] m341_25;
   assign m341_25 =10'b0;

   // m341_26 = W*in
   wire signed [9:0] m341_26;
   assign m341_26 =10'b0;

   // m341_27 = W*in
   wire signed [9:0] m341_27;
   assign m341_27 ={ {5{in341[5]}} , in341[5:1] };

   // m341_28 = W*in
   wire signed [9:0] m341_28;
   assign m341_28 =10'b0;

   // m341_29 = W*in
   wire signed [9:0] m341_29;
   assign m341_29 =10'b0;

   // m341_30 = W*in
   wire signed [9:0] m341_30;
   assign m341_30 ={ {5{neg341[5]}} , neg341[5:1] };

   // m341_31 = W*in
   wire signed [9:0] m341_31;
   assign m341_31 =10'b0;

   // m341_32 = W*in
   wire signed [9:0] m341_32;
   assign m341_32 =10'b0;

   // m341_33 = W*in
   wire signed [9:0] m341_33;
   assign m341_33 =10'b0;

   // m341_34 = W*in
   wire signed [9:0] m341_34;
   assign m341_34 ={ {5{in341[5]}} , in341[5:1] };

   // m341_35 = W*in
   wire signed [9:0] m341_35;
   assign m341_35 =10'b0;

   // m341_36 = W*in
   wire signed [9:0] m341_36;
   assign m341_36 =10'b0;

   // m341_37 = W*in
   wire signed [9:0] m341_37;
   assign m341_37 =10'b0;

   // m341_38 = W*in
   wire signed [9:0] m341_38;
   assign m341_38 =10'b0;

   // m341_39 = W*in
   wire signed [9:0] m341_39;
   assign m341_39 =10'b0;

   // m341_40 = W*in
   wire signed [9:0] m341_40;
   assign m341_40 =10'b0;

   // m341_41 = W*in
   wire signed [9:0] m341_41;
   assign m341_41 =10'b0;

   // m341_42 = W*in
   wire signed [9:0] m341_42;
   assign m341_42 =10'b0;

   // m341_43 = W*in
   wire signed [9:0] m341_43;
   assign m341_43 =10'b0;

   // m341_44 = W*in
   wire signed [9:0] m341_44;
   assign m341_44 =10'b0;

   // m341_45 = W*in
   wire signed [9:0] m341_45;
   assign m341_45 =10'b0;

   // m341_46 = W*in
   wire signed [9:0] m341_46;
   assign m341_46 =10'b0;

   // m341_47 = W*in
   wire signed [9:0] m341_47;
   assign m341_47 =10'b0;

   // m341_48 = W*in
   wire signed [9:0] m341_48;
   assign m341_48 =10'b0;

   // m341_49 = W*in
   wire signed [9:0] m341_49;
   assign m341_49 =10'b0;

   // m341_50 = W*in
   wire signed [9:0] m341_50;
   assign m341_50 =10'b0;

   // m341_51 = W*in
   wire signed [9:0] m341_51;
   assign m341_51 =10'b0;

   // m341_52 = W*in
   wire signed [9:0] m341_52;
   assign m341_52 =10'b0;

   // m341_53 = W*in
   wire signed [9:0] m341_53;
   assign m341_53 =10'b0;

   // m341_54 = W*in
   wire signed [9:0] m341_54;
   assign m341_54 =10'b0;

   // m341_55 = W*in
   wire signed [9:0] m341_55;
   assign m341_55 =10'b0;

   // m341_56 = W*in
   wire signed [9:0] m341_56;
   assign m341_56 =10'b0;

   // m341_57 = W*in
   wire signed [9:0] m341_57;
   assign m341_57 =10'b0;

   // m341_58 = W*in
   wire signed [9:0] m341_58;
   assign m341_58 =10'b0;

   // m341_59 = W*in
   wire signed [9:0] m341_59;
   assign m341_59 =10'b0;

   // m341_60 = W*in
   wire signed [9:0] m341_60;
   assign m341_60 =10'b0;

   // m341_61 = W*in
   wire signed [9:0] m341_61;
   assign m341_61 =10'b0;

   // m341_62 = W*in
   wire signed [9:0] m341_62;
   assign m341_62 =10'b0;

   // m341_63 = W*in
   wire signed [9:0] m341_63;
   assign m341_63 =10'b0;

   // m341_64 = W*in
   wire signed [9:0] m341_64;
   assign m341_64 =10'b0;

   // m341_65 = W*in
   wire signed [9:0] m341_65;
   assign m341_65 =10'b0;

   // m341_66 = W*in
   wire signed [9:0] m341_66;
   assign m341_66 ={ {5{neg341[5]}} , neg341[5:1] };

   // m341_67 = W*in
   wire signed [9:0] m341_67;
   assign m341_67 =10'b0;

   // m341_68 = W*in
   wire signed [9:0] m341_68;
   assign m341_68 =10'b0;

   // m341_69 = W*in
   wire signed [9:0] m341_69;
   assign m341_69 =10'b0;

   // m341_70 = W*in
   wire signed [9:0] m341_70;
   assign m341_70 =10'b0;

   // m341_71 = W*in
   wire signed [9:0] m341_71;
   assign m341_71 =10'b0;

   // m341_72 = W*in
   wire signed [9:0] m341_72;
   assign m341_72 =10'b0;

   // m341_73 = W*in
   wire signed [9:0] m341_73;
   assign m341_73 =10'b0;

   // m341_74 = W*in
   wire signed [9:0] m341_74;
   assign m341_74 =10'b0;

   // m341_75 = W*in
   wire signed [9:0] m341_75;
   assign m341_75 =10'b0;

   // m341_76 = W*in
   wire signed [9:0] m341_76;
   assign m341_76 =10'b0;

   // m341_77 = W*in
   wire signed [9:0] m341_77;
   assign m341_77 =10'b0;

   // m341_78 = W*in
   wire signed [9:0] m341_78;
   assign m341_78 =10'b0;

   // m341_79 = W*in
   wire signed [9:0] m341_79;
   assign m341_79 =10'b0;

   // m341_80 = W*in
   wire signed [9:0] m341_80;
   assign m341_80 =10'b0;

   // m341_81 = W*in
   wire signed [9:0] m341_81;
   assign m341_81 =10'b0;

   // m341_82 = W*in
   wire signed [9:0] m341_82;
   assign m341_82 =10'b0;

   // m341_83 = W*in
   wire signed [9:0] m341_83;
   assign m341_83 =10'b0;

   // m341_84 = W*in
   wire signed [9:0] m341_84;
   assign m341_84 =10'b0;

   // m341_85 = W*in
   wire signed [9:0] m341_85;
   assign m341_85 =10'b0;

   // m341_86 = W*in
   wire signed [9:0] m341_86;
   assign m341_86 =10'b0;

   // m341_87 = W*in
   wire signed [9:0] m341_87;
   assign m341_87 =10'b0;

   // m341_88 = W*in
   wire signed [9:0] m341_88;
   assign m341_88 =10'b0;

   // m341_89 = W*in
   wire signed [9:0] m341_89;
   assign m341_89 =10'b0;

   // m341_90 = W*in
   wire signed [9:0] m341_90;
   assign m341_90 =10'b0;

   // m341_91 = W*in
   wire signed [9:0] m341_91;
   assign m341_91 =10'b0;

   // m341_92 = W*in
   wire signed [9:0] m341_92;
   assign m341_92 =10'b0;

   // m341_93 = W*in
   wire signed [9:0] m341_93;
   assign m341_93 =10'b0;

   // m341_94 = W*in
   wire signed [9:0] m341_94;
   assign m341_94 =10'b0;

   // m341_95 = W*in
   wire signed [9:0] m341_95;
   assign m341_95 =10'b0;

   // m341_96 = W*in
   wire signed [9:0] m341_96;
   assign m341_96 =10'b0;

   // m341_97 = W*in
   wire signed [9:0] m341_97;
   assign m341_97 =10'b0;

   // m341_98 = W*in
   wire signed [9:0] m341_98;
   assign m341_98 =10'b0;

   // m341_99 = W*in
   wire signed [9:0] m341_99;
   assign m341_99 =10'b0;

   // m341_100 = W*in
   wire signed [9:0] m341_100;
   assign m341_100 =10'b0;

   // m341_101 = W*in
   wire signed [9:0] m341_101;
   assign m341_101 =10'b0;

   // m341_102 = W*in
   wire signed [9:0] m341_102;
   assign m341_102 =10'b0;

   // m341_103 = W*in
   wire signed [9:0] m341_103;
   assign m341_103 =10'b0;

   // m341_104 = W*in
   wire signed [9:0] m341_104;
   assign m341_104 =10'b0;

   // m341_105 = W*in
   wire signed [9:0] m341_105;
   assign m341_105 =10'b0;

   // m341_106 = W*in
   wire signed [9:0] m341_106;
   assign m341_106 =10'b0;

   // m341_107 = W*in
   wire signed [9:0] m341_107;
   assign m341_107 =10'b0;

   // m341_108 = W*in
   wire signed [9:0] m341_108;
   assign m341_108 =10'b0;

   // m341_109 = W*in
   wire signed [9:0] m341_109;
   assign m341_109 =10'b0;

   // m341_110 = W*in
   wire signed [9:0] m341_110;
   assign m341_110 =10'b0;

   // m341_111 = W*in
   wire signed [9:0] m341_111;
   assign m341_111 =10'b0;

   // m341_112 = W*in
   wire signed [9:0] m341_112;
   assign m341_112 =10'b0;

   // m341_113 = W*in
   wire signed [9:0] m341_113;
   assign m341_113 =10'b0;

   // m341_114 = W*in
   wire signed [9:0] m341_114;
   assign m341_114 =10'b0;

   // m341_115 = W*in
   wire signed [9:0] m341_115;
   assign m341_115 =10'b0;

   // m341_116 = W*in
   wire signed [9:0] m341_116;
   assign m341_116 =10'b0;

   // m341_117 = W*in
   wire signed [9:0] m341_117;
   assign m341_117 =10'b0;

   // m342_1 = W*in
   wire signed [9:0] m342_1;
   assign m342_1 =10'b0;

   // m342_2 = W*in
   wire signed [9:0] m342_2;
   assign m342_2 =10'b0;

   // m342_3 = W*in
   wire signed [9:0] m342_3;
   assign m342_3 =10'b0;

   // m342_4 = W*in
   wire signed [9:0] m342_4;
   assign m342_4 =10'b0;

   // m342_5 = W*in
   wire signed [9:0] m342_5;
   assign m342_5 =10'b0;

   // m342_6 = W*in
   wire signed [9:0] m342_6;
   assign m342_6 =10'b0;

   // m342_7 = W*in
   wire signed [9:0] m342_7;
   assign m342_7 =10'b0;

   // m342_8 = W*in
   wire signed [9:0] m342_8;
   assign m342_8 =10'b0;

   // m342_9 = W*in
   wire signed [9:0] m342_9;
   assign m342_9 =10'b0;

   // m342_10 = W*in
   wire signed [9:0] m342_10;
   assign m342_10 =10'b0;

   // m342_11 = W*in
   wire signed [9:0] m342_11;
   assign m342_11 =10'b0;

   // m342_12 = W*in
   wire signed [9:0] m342_12;
   assign m342_12 =10'b0;

   // m342_13 = W*in
   wire signed [9:0] m342_13;
   assign m342_13 =10'b0;

   // m342_14 = W*in
   wire signed [9:0] m342_14;
   assign m342_14 =10'b0;

   // m342_15 = W*in
   wire signed [9:0] m342_15;
   assign m342_15 =10'b0;

   // m342_16 = W*in
   wire signed [9:0] m342_16;
   assign m342_16 ={ {5{in342[5]}} , in342[5:1] };

   // m342_17 = W*in
   wire signed [9:0] m342_17;
   assign m342_17 ={ {5{neg342[5]}} , neg342[5:1] };

   // m342_18 = W*in
   wire signed [9:0] m342_18;
   assign m342_18 ={ {5{in342[5]}} , in342[5:1] };

   // m342_19 = W*in
   wire signed [9:0] m342_19;
   assign m342_19 ={ {4{neg342[5]}} , neg342[5:0] };

   // m342_20 = W*in
   wire signed [9:0] m342_20;
   assign m342_20 ={ {4{in342[5]}} , in342[5:0] };

   // m342_21 = W*in
   wire signed [9:0] m342_21;
   assign m342_21 =10'b0;

   // m342_22 = W*in
   wire signed [9:0] m342_22;
   assign m342_22 =10'b0;

   // m342_23 = W*in
   wire signed [9:0] m342_23;
   assign m342_23 =10'b0;

   // m342_24 = W*in
   wire signed [9:0] m342_24;
   assign m342_24 =10'b0;

   // m342_25 = W*in
   wire signed [9:0] m342_25;
   assign m342_25 =10'b0;

   // m342_26 = W*in
   wire signed [9:0] m342_26;
   assign m342_26 ={ {5{in342[5]}} , in342[5:1] };

   // m342_27 = W*in
   wire signed [9:0] m342_27;
   assign m342_27 =10'b0;

   // m342_28 = W*in
   wire signed [9:0] m342_28;
   assign m342_28 ={ {5{neg342[5]}} , neg342[5:1] };

   // m342_29 = W*in
   wire signed [9:0] m342_29;
   assign m342_29 =10'b0;

   // m342_30 = W*in
   wire signed [9:0] m342_30;
   assign m342_30 =10'b0;

   // m342_31 = W*in
   wire signed [9:0] m342_31;
   assign m342_31 =10'b0;

   // m342_32 = W*in
   wire signed [9:0] m342_32;
   assign m342_32 =10'b0;

   // m342_33 = W*in
   wire signed [9:0] m342_33;
   assign m342_33 =10'b0;

   // m342_34 = W*in
   wire signed [9:0] m342_34;
   assign m342_34 ={ {4{in342[5]}} , in342[5:0] };

   // m342_35 = W*in
   wire signed [9:0] m342_35;
   assign m342_35 =10'b0;

   // m342_36 = W*in
   wire signed [9:0] m342_36;
   assign m342_36 =10'b0;

   // m342_37 = W*in
   wire signed [9:0] m342_37;
   assign m342_37 =10'b0;

   // m342_38 = W*in
   wire signed [9:0] m342_38;
   assign m342_38 =10'b0;

   // m342_39 = W*in
   wire signed [9:0] m342_39;
   assign m342_39 =10'b0;

   // m342_40 = W*in
   wire signed [9:0] m342_40;
   assign m342_40 =10'b0;

   // m342_41 = W*in
   wire signed [9:0] m342_41;
   assign m342_41 =10'b0;

   // m342_42 = W*in
   wire signed [9:0] m342_42;
   assign m342_42 =10'b0;

   // m342_43 = W*in
   wire signed [9:0] m342_43;
   assign m342_43 =10'b0;

   // m342_44 = W*in
   wire signed [9:0] m342_44;
   assign m342_44 ={ {4{neg342[5]}} , neg342[5:0] };

   // m342_45 = W*in
   wire signed [9:0] m342_45;
   assign m342_45 =10'b0;

   // m342_46 = W*in
   wire signed [9:0] m342_46;
   assign m342_46 =10'b0;

   // m342_47 = W*in
   wire signed [9:0] m342_47;
   assign m342_47 =10'b0;

   // m342_48 = W*in
   wire signed [9:0] m342_48;
   assign m342_48 =10'b0;

   // m342_49 = W*in
   wire signed [9:0] m342_49;
   assign m342_49 ={ {4{neg342[5]}} , neg342[5:0] };

   // m342_50 = W*in
   wire signed [9:0] m342_50;
   assign m342_50 =10'b0;

   // m342_51 = W*in
   wire signed [9:0] m342_51;
   assign m342_51 =10'b0;

   // m342_52 = W*in
   wire signed [9:0] m342_52;
   assign m342_52 =10'b0;

   // m342_53 = W*in
   wire signed [9:0] m342_53;
   assign m342_53 ={ {4{neg342[5]}} , neg342[5:0] };

   // m342_54 = W*in
   wire signed [9:0] m342_54;
   assign m342_54 =10'b0;

   // m342_55 = W*in
   wire signed [9:0] m342_55;
   assign m342_55 =10'b0;

   // m342_56 = W*in
   wire signed [9:0] m342_56;
   assign m342_56 ={ {4{in342[5]}} , in342[5:0] };

   // m342_57 = W*in
   wire signed [9:0] m342_57;
   assign m342_57 =10'b0;

   // m342_58 = W*in
   wire signed [9:0] m342_58;
   assign m342_58 =10'b0;

   // m342_59 = W*in
   wire signed [9:0] m342_59;
   assign m342_59 =10'b0;

   // m342_60 = W*in
   wire signed [9:0] m342_60;
   assign m342_60 =10'b0;

   // m342_61 = W*in
   wire signed [9:0] m342_61;
   assign m342_61 =10'b0;

   // m342_62 = W*in
   wire signed [9:0] m342_62;
   assign m342_62 =10'b0;

   // m342_63 = W*in
   wire signed [9:0] m342_63;
   assign m342_63 =10'b0;

   // m342_64 = W*in
   wire signed [9:0] m342_64;
   assign m342_64 ={ {5{in342[5]}} , in342[5:1] };

   // m342_65 = W*in
   wire signed [9:0] m342_65;
   assign m342_65 =10'b0;

   // m342_66 = W*in
   wire signed [9:0] m342_66;
   assign m342_66 ={ {5{neg342[5]}} , neg342[5:1] };

   // m342_67 = W*in
   wire signed [9:0] m342_67;
   assign m342_67 ={ {4{neg342[5]}} , neg342[5:0] };

   // m342_68 = W*in
   wire signed [9:0] m342_68;
   assign m342_68 =10'b0;

   // m342_69 = W*in
   wire signed [9:0] m342_69;
   assign m342_69 =10'b0;

   // m342_70 = W*in
   wire signed [9:0] m342_70;
   assign m342_70 ={ {5{in342[5]}} , in342[5:1] };

   // m342_71 = W*in
   wire signed [9:0] m342_71;
   assign m342_71 =10'b0;

   // m342_72 = W*in
   wire signed [9:0] m342_72;
   assign m342_72 ={ {5{in342[5]}} , in342[5:1] };

   // m342_73 = W*in
   wire signed [9:0] m342_73;
   assign m342_73 ={ {5{neg342[5]}} , neg342[5:1] };

   // m342_74 = W*in
   wire signed [9:0] m342_74;
   assign m342_74 ={ {5{in342[5]}} , in342[5:1] };

   // m342_75 = W*in
   wire signed [9:0] m342_75;
   assign m342_75 =10'b0;

   // m342_76 = W*in
   wire signed [9:0] m342_76;
   assign m342_76 =10'b0;

   // m342_77 = W*in
   wire signed [9:0] m342_77;
   assign m342_77 =10'b0;

   // m342_78 = W*in
   wire signed [9:0] m342_78;
   assign m342_78 ={ {4{in342[5]}} , in342[5:0] };

   // m342_79 = W*in
   wire signed [9:0] m342_79;
   assign m342_79 =10'b0;

   // m342_80 = W*in
   wire signed [9:0] m342_80;
   assign m342_80 =10'b0;

   // m342_81 = W*in
   wire signed [9:0] m342_81;
   assign m342_81 =10'b0;

   // m342_82 = W*in
   wire signed [9:0] m342_82;
   assign m342_82 =10'b0;

   // m342_83 = W*in
   wire signed [9:0] m342_83;
   assign m342_83 =10'b0;

   // m342_84 = W*in
   wire signed [9:0] m342_84;
   assign m342_84 ={ {5{in342[5]}} , in342[5:1] };

   // m342_85 = W*in
   wire signed [9:0] m342_85;
   assign m342_85 =10'b0;

   // m342_86 = W*in
   wire signed [9:0] m342_86;
   assign m342_86 =10'b0;

   // m342_87 = W*in
   wire signed [9:0] m342_87;
   assign m342_87 ={ {4{in342[5]}} , in342[5:0] };

   // m342_88 = W*in
   wire signed [9:0] m342_88;
   assign m342_88 ={ {4{in342[5]}} , in342[5:0] };

   // m342_89 = W*in
   wire signed [9:0] m342_89;
   assign m342_89 ={ {4{in342[5]}} , in342[5:0] };

   // m342_90 = W*in
   wire signed [9:0] m342_90;
   assign m342_90 =10'b0;

   // m342_91 = W*in
   wire signed [9:0] m342_91;
   assign m342_91 =10'b0;

   // m342_92 = W*in
   wire signed [9:0] m342_92;
   assign m342_92 =10'b0;

   // m342_93 = W*in
   wire signed [9:0] m342_93;
   assign m342_93 =10'b0;

   // m342_94 = W*in
   wire signed [9:0] m342_94;
   assign m342_94 =10'b0;

   // m342_95 = W*in
   wire signed [9:0] m342_95;
   assign m342_95 =10'b0;

   // m342_96 = W*in
   wire signed [9:0] m342_96;
   assign m342_96 =10'b0;

   // m342_97 = W*in
   wire signed [9:0] m342_97;
   assign m342_97 ={ {4{neg342[5]}} , neg342[5:0] };

   // m342_98 = W*in
   wire signed [9:0] m342_98;
   assign m342_98 =10'b0;

   // m342_99 = W*in
   wire signed [9:0] m342_99;
   assign m342_99 =10'b0;

   // m342_100 = W*in
   wire signed [9:0] m342_100;
   assign m342_100 =10'b0;

   // m342_101 = W*in
   wire signed [9:0] m342_101;
   assign m342_101 =10'b0;

   // m342_102 = W*in
   wire signed [9:0] m342_102;
   assign m342_102 =10'b0;

   // m342_103 = W*in
   wire signed [9:0] m342_103;
   assign m342_103 =10'b0;

   // m342_104 = W*in
   wire signed [9:0] m342_104;
   assign m342_104 =10'b0;

   // m342_105 = W*in
   wire signed [9:0] m342_105;
   assign m342_105 =10'b0;

   // m342_106 = W*in
   wire signed [9:0] m342_106;
   assign m342_106 =10'b0;

   // m342_107 = W*in
   wire signed [9:0] m342_107;
   assign m342_107 =10'b0;

   // m342_108 = W*in
   wire signed [9:0] m342_108;
   assign m342_108 =10'b0;

   // m342_109 = W*in
   wire signed [9:0] m342_109;
   assign m342_109 ={ {4{in342[5]}} , in342[5:0] };

   // m342_110 = W*in
   wire signed [9:0] m342_110;
   assign m342_110 =10'b0;

   // m342_111 = W*in
   wire signed [9:0] m342_111;
   assign m342_111 =10'b0;

   // m342_112 = W*in
   wire signed [9:0] m342_112;
   assign m342_112 =10'b0;

   // m342_113 = W*in
   wire signed [9:0] m342_113;
   assign m342_113 =10'b0;

   // m342_114 = W*in
   wire signed [9:0] m342_114;
   assign m342_114 =10'b0;

   // m342_115 = W*in
   wire signed [9:0] m342_115;
   assign m342_115 ={ {5{in342[5]}} , in342[5:1] };

   // m342_116 = W*in
   wire signed [9:0] m342_116;
   assign m342_116 =10'b0;

   // m342_117 = W*in
   wire signed [9:0] m342_117;
   assign m342_117 =10'b0;

   // m343_1 = W*in
   wire signed [9:0] m343_1;
   assign m343_1 =10'b0;

   // m343_2 = W*in
   wire signed [9:0] m343_2;
   assign m343_2 =10'b0;

   // m343_3 = W*in
   wire signed [9:0] m343_3;
   assign m343_3 =10'b0;

   // m343_4 = W*in
   wire signed [9:0] m343_4;
   assign m343_4 =10'b0;

   // m343_5 = W*in
   wire signed [9:0] m343_5;
   assign m343_5 =10'b0;

   // m343_6 = W*in
   wire signed [9:0] m343_6;
   assign m343_6 =10'b0;

   // m343_7 = W*in
   wire signed [9:0] m343_7;
   assign m343_7 =10'b0;

   // m343_8 = W*in
   wire signed [9:0] m343_8;
   assign m343_8 =10'b0;

   // m343_9 = W*in
   wire signed [9:0] m343_9;
   assign m343_9 =10'b0;

   // m343_10 = W*in
   wire signed [9:0] m343_10;
   assign m343_10 =10'b0;

   // m343_11 = W*in
   wire signed [9:0] m343_11;
   assign m343_11 =10'b0;

   // m343_12 = W*in
   wire signed [9:0] m343_12;
   assign m343_12 =10'b0;

   // m343_13 = W*in
   wire signed [9:0] m343_13;
   assign m343_13 =10'b0;

   // m343_14 = W*in
   wire signed [9:0] m343_14;
   assign m343_14 =10'b0;

   // m343_15 = W*in
   wire signed [9:0] m343_15;
   assign m343_15 =10'b0;

   // m343_16 = W*in
   wire signed [9:0] m343_16;
   assign m343_16 ={ {5{in343[5]}} , in343[5:1] };

   // m343_17 = W*in
   wire signed [9:0] m343_17;
   assign m343_17 ={ {5{neg343[5]}} , neg343[5:1] };

   // m343_18 = W*in
   wire signed [9:0] m343_18;
   assign m343_18 =10'b0;

   // m343_19 = W*in
   wire signed [9:0] m343_19;
   assign m343_19 ={ {5{neg343[5]}} , neg343[5:1] };

   // m343_20 = W*in
   wire signed [9:0] m343_20;
   assign m343_20 =10'b0;

   // m343_21 = W*in
   wire signed [9:0] m343_21;
   assign m343_21 ={ {4{in343[5]}} , in343[5:0] };

   // m343_22 = W*in
   wire signed [9:0] m343_22;
   assign m343_22 =10'b0;

   // m343_23 = W*in
   wire signed [9:0] m343_23;
   assign m343_23 =10'b0;

   // m343_24 = W*in
   wire signed [9:0] m343_24;
   assign m343_24 =10'b0;

   // m343_25 = W*in
   wire signed [9:0] m343_25;
   assign m343_25 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_26 = W*in
   wire signed [9:0] m343_26;
   assign m343_26 ={ {4{in343[5]}} , in343[5:0] };

   // m343_27 = W*in
   wire signed [9:0] m343_27;
   assign m343_27 ={ {5{neg343[5]}} , neg343[5:1] };

   // m343_28 = W*in
   wire signed [9:0] m343_28;
   assign m343_28 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_29 = W*in
   wire signed [9:0] m343_29;
   assign m343_29 =10'b0;

   // m343_30 = W*in
   wire signed [9:0] m343_30;
   assign m343_30 =10'b0;

   // m343_31 = W*in
   wire signed [9:0] m343_31;
   assign m343_31 =10'b0;

   // m343_32 = W*in
   wire signed [9:0] m343_32;
   assign m343_32 =10'b0;

   // m343_33 = W*in
   wire signed [9:0] m343_33;
   assign m343_33 =10'b0;

   // m343_34 = W*in
   wire signed [9:0] m343_34;
   assign m343_34 =10'b0;

   // m343_35 = W*in
   wire signed [9:0] m343_35;
   assign m343_35 =10'b0;

   // m343_36 = W*in
   wire signed [9:0] m343_36;
   assign m343_36 =10'b0;

   // m343_37 = W*in
   wire signed [9:0] m343_37;
   assign m343_37 =10'b0;

   // m343_38 = W*in
   wire signed [9:0] m343_38;
   assign m343_38 =10'b0;

   // m343_39 = W*in
   wire signed [9:0] m343_39;
   assign m343_39 =10'b0;

   // m343_40 = W*in
   wire signed [9:0] m343_40;
   assign m343_40 =10'b0;

   // m343_41 = W*in
   wire signed [9:0] m343_41;
   assign m343_41 =10'b0;

   // m343_42 = W*in
   wire signed [9:0] m343_42;
   assign m343_42 =10'b0;

   // m343_43 = W*in
   wire signed [9:0] m343_43;
   assign m343_43 =10'b0;

   // m343_44 = W*in
   wire signed [9:0] m343_44;
   assign m343_44 =10'b0;

   // m343_45 = W*in
   wire signed [9:0] m343_45;
   assign m343_45 =10'b0;

   // m343_46 = W*in
   wire signed [9:0] m343_46;
   assign m343_46 =10'b0;

   // m343_47 = W*in
   wire signed [9:0] m343_47;
   assign m343_47 =10'b0;

   // m343_48 = W*in
   wire signed [9:0] m343_48;
   assign m343_48 =10'b0;

   // m343_49 = W*in
   wire signed [9:0] m343_49;
   assign m343_49 =10'b0;

   // m343_50 = W*in
   wire signed [9:0] m343_50;
   assign m343_50 =10'b0;

   // m343_51 = W*in
   wire signed [9:0] m343_51;
   assign m343_51 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_52 = W*in
   wire signed [9:0] m343_52;
   assign m343_52 =10'b0;

   // m343_53 = W*in
   wire signed [9:0] m343_53;
   assign m343_53 =10'b0;

   // m343_54 = W*in
   wire signed [9:0] m343_54;
   assign m343_54 =10'b0;

   // m343_55 = W*in
   wire signed [9:0] m343_55;
   assign m343_55 =10'b0;

   // m343_56 = W*in
   wire signed [9:0] m343_56;
   assign m343_56 =10'b0;

   // m343_57 = W*in
   wire signed [9:0] m343_57;
   assign m343_57 =10'b0;

   // m343_58 = W*in
   wire signed [9:0] m343_58;
   assign m343_58 =10'b0;

   // m343_59 = W*in
   wire signed [9:0] m343_59;
   assign m343_59 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_60 = W*in
   wire signed [9:0] m343_60;
   assign m343_60 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_61 = W*in
   wire signed [9:0] m343_61;
   assign m343_61 =10'b0;

   // m343_62 = W*in
   wire signed [9:0] m343_62;
   assign m343_62 =10'b0;

   // m343_63 = W*in
   wire signed [9:0] m343_63;
   assign m343_63 =10'b0;

   // m343_64 = W*in
   wire signed [9:0] m343_64;
   assign m343_64 =10'b0;

   // m343_65 = W*in
   wire signed [9:0] m343_65;
   assign m343_65 ={ {5{in343[5]}} , in343[5:1] };

   // m343_66 = W*in
   wire signed [9:0] m343_66;
   assign m343_66 ={ {5{in343[5]}} , in343[5:1] };

   // m343_67 = W*in
   wire signed [9:0] m343_67;
   assign m343_67 =10'b0;

   // m343_68 = W*in
   wire signed [9:0] m343_68;
   assign m343_68 =10'b0;

   // m343_69 = W*in
   wire signed [9:0] m343_69;
   assign m343_69 ={ {4{in343[5]}} , in343[5:0] };

   // m343_70 = W*in
   wire signed [9:0] m343_70;
   assign m343_70 ={ {4{in343[5]}} , in343[5:0] };

   // m343_71 = W*in
   wire signed [9:0] m343_71;
   assign m343_71 =10'b0;

   // m343_72 = W*in
   wire signed [9:0] m343_72;
   assign m343_72 =10'b0;

   // m343_73 = W*in
   wire signed [9:0] m343_73;
   assign m343_73 =10'b0;

   // m343_74 = W*in
   wire signed [9:0] m343_74;
   assign m343_74 ={ {4{in343[5]}} , in343[5:0] };

   // m343_75 = W*in
   wire signed [9:0] m343_75;
   assign m343_75 =10'b0;

   // m343_76 = W*in
   wire signed [9:0] m343_76;
   assign m343_76 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_77 = W*in
   wire signed [9:0] m343_77;
   assign m343_77 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_78 = W*in
   wire signed [9:0] m343_78;
   assign m343_78 ={ {4{in343[5]}} , in343[5:0] };

   // m343_79 = W*in
   wire signed [9:0] m343_79;
   assign m343_79 =10'b0;

   // m343_80 = W*in
   wire signed [9:0] m343_80;
   assign m343_80 =10'b0;

   // m343_81 = W*in
   wire signed [9:0] m343_81;
   assign m343_81 ={ {5{in343[5]}} , in343[5:1] };

   // m343_82 = W*in
   wire signed [9:0] m343_82;
   assign m343_82 =10'b0;

   // m343_83 = W*in
   wire signed [9:0] m343_83;
   assign m343_83 ={ {5{neg343[5]}} , neg343[5:1] };

   // m343_84 = W*in
   wire signed [9:0] m343_84;
   assign m343_84 =10'b0;

   // m343_85 = W*in
   wire signed [9:0] m343_85;
   assign m343_85 =10'b0;

   // m343_86 = W*in
   wire signed [9:0] m343_86;
   assign m343_86 =10'b0;

   // m343_87 = W*in
   wire signed [9:0] m343_87;
   assign m343_87 =10'b0;

   // m343_88 = W*in
   wire signed [9:0] m343_88;
   assign m343_88 =10'b0;

   // m343_89 = W*in
   wire signed [9:0] m343_89;
   assign m343_89 ={ {4{in343[5]}} , in343[5:0] };

   // m343_90 = W*in
   wire signed [9:0] m343_90;
   assign m343_90 =10'b0;

   // m343_91 = W*in
   wire signed [9:0] m343_91;
   assign m343_91 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_92 = W*in
   wire signed [9:0] m343_92;
   assign m343_92 =10'b0;

   // m343_93 = W*in
   wire signed [9:0] m343_93;
   assign m343_93 =10'b0;

   // m343_94 = W*in
   wire signed [9:0] m343_94;
   assign m343_94 =10'b0;

   // m343_95 = W*in
   wire signed [9:0] m343_95;
   assign m343_95 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_96 = W*in
   wire signed [9:0] m343_96;
   assign m343_96 ={ {4{in343[5]}} , in343[5:0] };

   // m343_97 = W*in
   wire signed [9:0] m343_97;
   assign m343_97 =10'b0;

   // m343_98 = W*in
   wire signed [9:0] m343_98;
   assign m343_98 =10'b0;

   // m343_99 = W*in
   wire signed [9:0] m343_99;
   assign m343_99 =10'b0;

   // m343_100 = W*in
   wire signed [9:0] m343_100;
   assign m343_100 =10'b0;

   // m343_101 = W*in
   wire signed [9:0] m343_101;
   assign m343_101 =10'b0;

   // m343_102 = W*in
   wire signed [9:0] m343_102;
   assign m343_102 =10'b0;

   // m343_103 = W*in
   wire signed [9:0] m343_103;
   assign m343_103 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_104 = W*in
   wire signed [9:0] m343_104;
   assign m343_104 ={ {4{neg343[5]}} , neg343[5:0] };

   // m343_105 = W*in
   wire signed [9:0] m343_105;
   assign m343_105 =10'b0;

   // m343_106 = W*in
   wire signed [9:0] m343_106;
   assign m343_106 =10'b0;

   // m343_107 = W*in
   wire signed [9:0] m343_107;
   assign m343_107 =10'b0;

   // m343_108 = W*in
   wire signed [9:0] m343_108;
   assign m343_108 =10'b0;

   // m343_109 = W*in
   wire signed [9:0] m343_109;
   assign m343_109 =10'b0;

   // m343_110 = W*in
   wire signed [9:0] m343_110;
   assign m343_110 =10'b0;

   // m343_111 = W*in
   wire signed [9:0] m343_111;
   assign m343_111 =10'b0;

   // m343_112 = W*in
   wire signed [9:0] m343_112;
   assign m343_112 =10'b0;

   // m343_113 = W*in
   wire signed [9:0] m343_113;
   assign m343_113 =10'b0;

   // m343_114 = W*in
   wire signed [9:0] m343_114;
   assign m343_114 =10'b0;

   // m343_115 = W*in
   wire signed [9:0] m343_115;
   assign m343_115 =10'b0;

   // m343_116 = W*in
   wire signed [9:0] m343_116;
   assign m343_116 =10'b0;

   // m343_117 = W*in
   wire signed [9:0] m343_117;
   assign m343_117 =10'b0;

   // m344_1 = W*in
   wire signed [9:0] m344_1;
   assign m344_1 =10'b0;

   // m344_2 = W*in
   wire signed [9:0] m344_2;
   assign m344_2 =10'b0;

   // m344_3 = W*in
   wire signed [9:0] m344_3;
   assign m344_3 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_4 = W*in
   wire signed [9:0] m344_4;
   assign m344_4 =10'b0;

   // m344_5 = W*in
   wire signed [9:0] m344_5;
   assign m344_5 =10'b0;

   // m344_6 = W*in
   wire signed [9:0] m344_6;
   assign m344_6 =10'b0;

   // m344_7 = W*in
   wire signed [9:0] m344_7;
   assign m344_7 =10'b0;

   // m344_8 = W*in
   wire signed [9:0] m344_8;
   assign m344_8 =10'b0;

   // m344_9 = W*in
   wire signed [9:0] m344_9;
   assign m344_9 =10'b0;

   // m344_10 = W*in
   wire signed [9:0] m344_10;
   assign m344_10 ={ {4{in344[5]}} , in344[5:0] };

   // m344_11 = W*in
   wire signed [9:0] m344_11;
   assign m344_11 =10'b0;

   // m344_12 = W*in
   wire signed [9:0] m344_12;
   assign m344_12 ={ {4{in344[5]}} , in344[5:0] };

   // m344_13 = W*in
   wire signed [9:0] m344_13;
   assign m344_13 =10'b0;

   // m344_14 = W*in
   wire signed [9:0] m344_14;
   assign m344_14 ={ {4{in344[5]}} , in344[5:0] };

   // m344_15 = W*in
   wire signed [9:0] m344_15;
   assign m344_15 =10'b0;

   // m344_16 = W*in
   wire signed [9:0] m344_16;
   assign m344_16 =10'b0;

   // m344_17 = W*in
   wire signed [9:0] m344_17;
   assign m344_17 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_18 = W*in
   wire signed [9:0] m344_18;
   assign m344_18 ={ {4{in344[5]}} , in344[5:0] };

   // m344_19 = W*in
   wire signed [9:0] m344_19;
   assign m344_19 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_20 = W*in
   wire signed [9:0] m344_20;
   assign m344_20 =10'b0;

   // m344_21 = W*in
   wire signed [9:0] m344_21;
   assign m344_21 =10'b0;

   // m344_22 = W*in
   wire signed [9:0] m344_22;
   assign m344_22 =10'b0;

   // m344_23 = W*in
   wire signed [9:0] m344_23;
   assign m344_23 =10'b0;

   // m344_24 = W*in
   wire signed [9:0] m344_24;
   assign m344_24 =10'b0;

   // m344_25 = W*in
   wire signed [9:0] m344_25;
   assign m344_25 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_26 = W*in
   wire signed [9:0] m344_26;
   assign m344_26 ={ {4{in344[5]}} , in344[5:0] };

   // m344_27 = W*in
   wire signed [9:0] m344_27;
   assign m344_27 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_28 = W*in
   wire signed [9:0] m344_28;
   assign m344_28 =10'b0;

   // m344_29 = W*in
   wire signed [9:0] m344_29;
   assign m344_29 =10'b0;

   // m344_30 = W*in
   wire signed [9:0] m344_30;
   assign m344_30 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_31 = W*in
   wire signed [9:0] m344_31;
   assign m344_31 =10'b0;

   // m344_32 = W*in
   wire signed [9:0] m344_32;
   assign m344_32 =10'b0;

   // m344_33 = W*in
   wire signed [9:0] m344_33;
   assign m344_33 =10'b0;

   // m344_34 = W*in
   wire signed [9:0] m344_34;
   assign m344_34 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_35 = W*in
   wire signed [9:0] m344_35;
   assign m344_35 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_36 = W*in
   wire signed [9:0] m344_36;
   assign m344_36 =10'b0;

   // m344_37 = W*in
   wire signed [9:0] m344_37;
   assign m344_37 =10'b0;

   // m344_38 = W*in
   wire signed [9:0] m344_38;
   assign m344_38 =10'b0;

   // m344_39 = W*in
   wire signed [9:0] m344_39;
   assign m344_39 =10'b0;

   // m344_40 = W*in
   wire signed [9:0] m344_40;
   assign m344_40 =10'b0;

   // m344_41 = W*in
   wire signed [9:0] m344_41;
   assign m344_41 =10'b0;

   // m344_42 = W*in
   wire signed [9:0] m344_42;
   assign m344_42 ={ {4{in344[5]}} , in344[5:0] };

   // m344_43 = W*in
   wire signed [9:0] m344_43;
   assign m344_43 =10'b0;

   // m344_44 = W*in
   wire signed [9:0] m344_44;
   assign m344_44 =10'b0;

   // m344_45 = W*in
   wire signed [9:0] m344_45;
   assign m344_45 =10'b0;

   // m344_46 = W*in
   wire signed [9:0] m344_46;
   assign m344_46 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_47 = W*in
   wire signed [9:0] m344_47;
   assign m344_47 =10'b0;

   // m344_48 = W*in
   wire signed [9:0] m344_48;
   assign m344_48 =10'b0;

   // m344_49 = W*in
   wire signed [9:0] m344_49;
   assign m344_49 =10'b0;

   // m344_50 = W*in
   wire signed [9:0] m344_50;
   assign m344_50 =10'b0;

   // m344_51 = W*in
   wire signed [9:0] m344_51;
   assign m344_51 ={ {4{in344[5]}} , in344[5:0] };

   // m344_52 = W*in
   wire signed [9:0] m344_52;
   assign m344_52 =10'b0;

   // m344_53 = W*in
   wire signed [9:0] m344_53;
   assign m344_53 =10'b0;

   // m344_54 = W*in
   wire signed [9:0] m344_54;
   assign m344_54 =10'b0;

   // m344_55 = W*in
   wire signed [9:0] m344_55;
   assign m344_55 =10'b0;

   // m344_56 = W*in
   wire signed [9:0] m344_56;
   assign m344_56 =10'b0;

   // m344_57 = W*in
   wire signed [9:0] m344_57;
   assign m344_57 =10'b0;

   // m344_58 = W*in
   wire signed [9:0] m344_58;
   assign m344_58 =10'b0;

   // m344_59 = W*in
   wire signed [9:0] m344_59;
   assign m344_59 =10'b0;

   // m344_60 = W*in
   wire signed [9:0] m344_60;
   assign m344_60 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_61 = W*in
   wire signed [9:0] m344_61;
   assign m344_61 =10'b0;

   // m344_62 = W*in
   wire signed [9:0] m344_62;
   assign m344_62 =10'b0;

   // m344_63 = W*in
   wire signed [9:0] m344_63;
   assign m344_63 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_64 = W*in
   wire signed [9:0] m344_64;
   assign m344_64 ={ {4{in344[5]}} , in344[5:0] };

   // m344_65 = W*in
   wire signed [9:0] m344_65;
   assign m344_65 =10'b0;

   // m344_66 = W*in
   wire signed [9:0] m344_66;
   assign m344_66 =10'b0;

   // m344_67 = W*in
   wire signed [9:0] m344_67;
   assign m344_67 =10'b0;

   // m344_68 = W*in
   wire signed [9:0] m344_68;
   assign m344_68 =10'b0;

   // m344_69 = W*in
   wire signed [9:0] m344_69;
   assign m344_69 =10'b0;

   // m344_70 = W*in
   wire signed [9:0] m344_70;
   assign m344_70 ={ {4{in344[5]}} , in344[5:0] };

   // m344_71 = W*in
   wire signed [9:0] m344_71;
   assign m344_71 =10'b0;

   // m344_72 = W*in
   wire signed [9:0] m344_72;
   assign m344_72 =10'b0;

   // m344_73 = W*in
   wire signed [9:0] m344_73;
   assign m344_73 =10'b0;

   // m344_74 = W*in
   wire signed [9:0] m344_74;
   assign m344_74 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_75 = W*in
   wire signed [9:0] m344_75;
   assign m344_75 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_76 = W*in
   wire signed [9:0] m344_76;
   assign m344_76 =10'b0;

   // m344_77 = W*in
   wire signed [9:0] m344_77;
   assign m344_77 ={ {4{in344[5]}} , in344[5:0] };

   // m344_78 = W*in
   wire signed [9:0] m344_78;
   assign m344_78 =10'b0;

   // m344_79 = W*in
   wire signed [9:0] m344_79;
   assign m344_79 =10'b0;

   // m344_80 = W*in
   wire signed [9:0] m344_80;
   assign m344_80 =10'b0;

   // m344_81 = W*in
   wire signed [9:0] m344_81;
   assign m344_81 =10'b0;

   // m344_82 = W*in
   wire signed [9:0] m344_82;
   assign m344_82 =10'b0;

   // m344_83 = W*in
   wire signed [9:0] m344_83;
   assign m344_83 =10'b0;

   // m344_84 = W*in
   wire signed [9:0] m344_84;
   assign m344_84 =10'b0;

   // m344_85 = W*in
   wire signed [9:0] m344_85;
   assign m344_85 ={ {4{in344[5]}} , in344[5:0] };

   // m344_86 = W*in
   wire signed [9:0] m344_86;
   assign m344_86 =10'b0;

   // m344_87 = W*in
   wire signed [9:0] m344_87;
   assign m344_87 =10'b0;

   // m344_88 = W*in
   wire signed [9:0] m344_88;
   assign m344_88 =10'b0;

   // m344_89 = W*in
   wire signed [9:0] m344_89;
   assign m344_89 =10'b0;

   // m344_90 = W*in
   wire signed [9:0] m344_90;
   assign m344_90 =10'b0;

   // m344_91 = W*in
   wire signed [9:0] m344_91;
   assign m344_91 =10'b0;

   // m344_92 = W*in
   wire signed [9:0] m344_92;
   assign m344_92 =10'b0;

   // m344_93 = W*in
   wire signed [9:0] m344_93;
   assign m344_93 =10'b0;

   // m344_94 = W*in
   wire signed [9:0] m344_94;
   assign m344_94 =10'b0;

   // m344_95 = W*in
   wire signed [9:0] m344_95;
   assign m344_95 =10'b0;

   // m344_96 = W*in
   wire signed [9:0] m344_96;
   assign m344_96 =10'b0;

   // m344_97 = W*in
   wire signed [9:0] m344_97;
   assign m344_97 =10'b0;

   // m344_98 = W*in
   wire signed [9:0] m344_98;
   assign m344_98 =10'b0;

   // m344_99 = W*in
   wire signed [9:0] m344_99;
   assign m344_99 =10'b0;

   // m344_100 = W*in
   wire signed [9:0] m344_100;
   assign m344_100 =10'b0;

   // m344_101 = W*in
   wire signed [9:0] m344_101;
   assign m344_101 =10'b0;

   // m344_102 = W*in
   wire signed [9:0] m344_102;
   assign m344_102 =10'b0;

   // m344_103 = W*in
   wire signed [9:0] m344_103;
   assign m344_103 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_104 = W*in
   wire signed [9:0] m344_104;
   assign m344_104 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_105 = W*in
   wire signed [9:0] m344_105;
   assign m344_105 =10'b0;

   // m344_106 = W*in
   wire signed [9:0] m344_106;
   assign m344_106 =10'b0;

   // m344_107 = W*in
   wire signed [9:0] m344_107;
   assign m344_107 =10'b0;

   // m344_108 = W*in
   wire signed [9:0] m344_108;
   assign m344_108 =10'b0;

   // m344_109 = W*in
   wire signed [9:0] m344_109;
   assign m344_109 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_110 = W*in
   wire signed [9:0] m344_110;
   assign m344_110 =10'b0;

   // m344_111 = W*in
   wire signed [9:0] m344_111;
   assign m344_111 =10'b0;

   // m344_112 = W*in
   wire signed [9:0] m344_112;
   assign m344_112 ={ {4{in344[5]}} , in344[5:0] };

   // m344_113 = W*in
   wire signed [9:0] m344_113;
   assign m344_113 =10'b0;

   // m344_114 = W*in
   wire signed [9:0] m344_114;
   assign m344_114 =10'b0;

   // m344_115 = W*in
   wire signed [9:0] m344_115;
   assign m344_115 ={ {5{neg344[5]}} , neg344[5:1] };

   // m344_116 = W*in
   wire signed [9:0] m344_116;
   assign m344_116 ={ {4{neg344[5]}} , neg344[5:0] };

   // m344_117 = W*in
   wire signed [9:0] m344_117;
   assign m344_117 =10'b0;

   // m345_1 = W*in
   wire signed [9:0] m345_1;
   assign m345_1 =10'b0;

   // m345_2 = W*in
   wire signed [9:0] m345_2;
   assign m345_2 =10'b0;

   // m345_3 = W*in
   wire signed [9:0] m345_3;
   assign m345_3 =10'b0;

   // m345_4 = W*in
   wire signed [9:0] m345_4;
   assign m345_4 =10'b0;

   // m345_5 = W*in
   wire signed [9:0] m345_5;
   assign m345_5 =10'b0;

   // m345_6 = W*in
   wire signed [9:0] m345_6;
   assign m345_6 =10'b0;

   // m345_7 = W*in
   wire signed [9:0] m345_7;
   assign m345_7 ={ {4{in345[5]}} , in345[5:0] };

   // m345_8 = W*in
   wire signed [9:0] m345_8;
   assign m345_8 =10'b0;

   // m345_9 = W*in
   wire signed [9:0] m345_9;
   assign m345_9 =10'b0;

   // m345_10 = W*in
   wire signed [9:0] m345_10;
   assign m345_10 =10'b0;

   // m345_11 = W*in
   wire signed [9:0] m345_11;
   assign m345_11 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_12 = W*in
   wire signed [9:0] m345_12;
   assign m345_12 =10'b0;

   // m345_13 = W*in
   wire signed [9:0] m345_13;
   assign m345_13 ={ {4{in345[5]}} , in345[5:0] };

   // m345_14 = W*in
   wire signed [9:0] m345_14;
   assign m345_14 =10'b0;

   // m345_15 = W*in
   wire signed [9:0] m345_15;
   assign m345_15 =10'b0;

   // m345_16 = W*in
   wire signed [9:0] m345_16;
   assign m345_16 =10'b0;

   // m345_17 = W*in
   wire signed [9:0] m345_17;
   assign m345_17 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_18 = W*in
   wire signed [9:0] m345_18;
   assign m345_18 =10'b0;

   // m345_19 = W*in
   wire signed [9:0] m345_19;
   assign m345_19 =10'b0;

   // m345_20 = W*in
   wire signed [9:0] m345_20;
   assign m345_20 =10'b0;

   // m345_21 = W*in
   wire signed [9:0] m345_21;
   assign m345_21 ={ {5{neg345[5]}} , neg345[5:1] };

   // m345_22 = W*in
   wire signed [9:0] m345_22;
   assign m345_22 =10'b0;

   // m345_23 = W*in
   wire signed [9:0] m345_23;
   assign m345_23 ={ {4{in345[5]}} , in345[5:0] };

   // m345_24 = W*in
   wire signed [9:0] m345_24;
   assign m345_24 ={ {4{in345[5]}} , in345[5:0] };

   // m345_25 = W*in
   wire signed [9:0] m345_25;
   assign m345_25 =10'b0;

   // m345_26 = W*in
   wire signed [9:0] m345_26;
   assign m345_26 =10'b0;

   // m345_27 = W*in
   wire signed [9:0] m345_27;
   assign m345_27 =10'b0;

   // m345_28 = W*in
   wire signed [9:0] m345_28;
   assign m345_28 =10'b0;

   // m345_29 = W*in
   wire signed [9:0] m345_29;
   assign m345_29 =10'b0;

   // m345_30 = W*in
   wire signed [9:0] m345_30;
   assign m345_30 ={ {5{neg345[5]}} , neg345[5:1] };

   // m345_31 = W*in
   wire signed [9:0] m345_31;
   assign m345_31 =10'b0;

   // m345_32 = W*in
   wire signed [9:0] m345_32;
   assign m345_32 =10'b0;

   // m345_33 = W*in
   wire signed [9:0] m345_33;
   assign m345_33 ={ {4{in345[5]}} , in345[5:0] };

   // m345_34 = W*in
   wire signed [9:0] m345_34;
   assign m345_34 =10'b0;

   // m345_35 = W*in
   wire signed [9:0] m345_35;
   assign m345_35 =10'b0;

   // m345_36 = W*in
   wire signed [9:0] m345_36;
   assign m345_36 =10'b0;

   // m345_37 = W*in
   wire signed [9:0] m345_37;
   assign m345_37 =10'b0;

   // m345_38 = W*in
   wire signed [9:0] m345_38;
   assign m345_38 =10'b0;

   // m345_39 = W*in
   wire signed [9:0] m345_39;
   assign m345_39 ={ {4{in345[5]}} , in345[5:0] };

   // m345_40 = W*in
   wire signed [9:0] m345_40;
   assign m345_40 =10'b0;

   // m345_41 = W*in
   wire signed [9:0] m345_41;
   assign m345_41 =10'b0;

   // m345_42 = W*in
   wire signed [9:0] m345_42;
   assign m345_42 =10'b0;

   // m345_43 = W*in
   wire signed [9:0] m345_43;
   assign m345_43 =10'b0;

   // m345_44 = W*in
   wire signed [9:0] m345_44;
   assign m345_44 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_45 = W*in
   wire signed [9:0] m345_45;
   assign m345_45 ={ {4{in345[5]}} , in345[5:0] };

   // m345_46 = W*in
   wire signed [9:0] m345_46;
   assign m345_46 =10'b0;

   // m345_47 = W*in
   wire signed [9:0] m345_47;
   assign m345_47 =10'b0;

   // m345_48 = W*in
   wire signed [9:0] m345_48;
   assign m345_48 ={ {4{in345[5]}} , in345[5:0] };

   // m345_49 = W*in
   wire signed [9:0] m345_49;
   assign m345_49 =10'b0;

   // m345_50 = W*in
   wire signed [9:0] m345_50;
   assign m345_50 =10'b0;

   // m345_51 = W*in
   wire signed [9:0] m345_51;
   assign m345_51 ={ {4{in345[5]}} , in345[5:0] };

   // m345_52 = W*in
   wire signed [9:0] m345_52;
   assign m345_52 =10'b0;

   // m345_53 = W*in
   wire signed [9:0] m345_53;
   assign m345_53 =10'b0;

   // m345_54 = W*in
   wire signed [9:0] m345_54;
   assign m345_54 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_55 = W*in
   wire signed [9:0] m345_55;
   assign m345_55 =10'b0;

   // m345_56 = W*in
   wire signed [9:0] m345_56;
   assign m345_56 =10'b0;

   // m345_57 = W*in
   wire signed [9:0] m345_57;
   assign m345_57 =10'b0;

   // m345_58 = W*in
   wire signed [9:0] m345_58;
   assign m345_58 =10'b0;

   // m345_59 = W*in
   wire signed [9:0] m345_59;
   assign m345_59 =10'b0;

   // m345_60 = W*in
   wire signed [9:0] m345_60;
   assign m345_60 =10'b0;

   // m345_61 = W*in
   wire signed [9:0] m345_61;
   assign m345_61 =10'b0;

   // m345_62 = W*in
   wire signed [9:0] m345_62;
   assign m345_62 =10'b0;

   // m345_63 = W*in
   wire signed [9:0] m345_63;
   assign m345_63 ={ {5{neg345[5]}} , neg345[5:1] };

   // m345_64 = W*in
   wire signed [9:0] m345_64;
   assign m345_64 =10'b0;

   // m345_65 = W*in
   wire signed [9:0] m345_65;
   assign m345_65 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_66 = W*in
   wire signed [9:0] m345_66;
   assign m345_66 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_67 = W*in
   wire signed [9:0] m345_67;
   assign m345_67 =10'b0;

   // m345_68 = W*in
   wire signed [9:0] m345_68;
   assign m345_68 =10'b0;

   // m345_69 = W*in
   wire signed [9:0] m345_69;
   assign m345_69 =10'b0;

   // m345_70 = W*in
   wire signed [9:0] m345_70;
   assign m345_70 =10'b0;

   // m345_71 = W*in
   wire signed [9:0] m345_71;
   assign m345_71 =10'b0;

   // m345_72 = W*in
   wire signed [9:0] m345_72;
   assign m345_72 ={ {4{in345[5]}} , in345[5:0] };

   // m345_73 = W*in
   wire signed [9:0] m345_73;
   assign m345_73 ={ {4{in345[5]}} , in345[5:0] };

   // m345_74 = W*in
   wire signed [9:0] m345_74;
   assign m345_74 ={ {5{neg345[5]}} , neg345[5:1] };

   // m345_75 = W*in
   wire signed [9:0] m345_75;
   assign m345_75 =10'b0;

   // m345_76 = W*in
   wire signed [9:0] m345_76;
   assign m345_76 =10'b0;

   // m345_77 = W*in
   wire signed [9:0] m345_77;
   assign m345_77 =10'b0;

   // m345_78 = W*in
   wire signed [9:0] m345_78;
   assign m345_78 =10'b0;

   // m345_79 = W*in
   wire signed [9:0] m345_79;
   assign m345_79 =10'b0;

   // m345_80 = W*in
   wire signed [9:0] m345_80;
   assign m345_80 =10'b0;

   // m345_81 = W*in
   wire signed [9:0] m345_81;
   assign m345_81 =10'b0;

   // m345_82 = W*in
   wire signed [9:0] m345_82;
   assign m345_82 =10'b0;

   // m345_83 = W*in
   wire signed [9:0] m345_83;
   assign m345_83 =10'b0;

   // m345_84 = W*in
   wire signed [9:0] m345_84;
   assign m345_84 ={ {4{in345[5]}} , in345[5:0] };

   // m345_85 = W*in
   wire signed [9:0] m345_85;
   assign m345_85 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_86 = W*in
   wire signed [9:0] m345_86;
   assign m345_86 =10'b0;

   // m345_87 = W*in
   wire signed [9:0] m345_87;
   assign m345_87 =10'b0;

   // m345_88 = W*in
   wire signed [9:0] m345_88;
   assign m345_88 =10'b0;

   // m345_89 = W*in
   wire signed [9:0] m345_89;
   assign m345_89 ={ {4{in345[5]}} , in345[5:0] };

   // m345_90 = W*in
   wire signed [9:0] m345_90;
   assign m345_90 =10'b0;

   // m345_91 = W*in
   wire signed [9:0] m345_91;
   assign m345_91 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_92 = W*in
   wire signed [9:0] m345_92;
   assign m345_92 =10'b0;

   // m345_93 = W*in
   wire signed [9:0] m345_93;
   assign m345_93 =10'b0;

   // m345_94 = W*in
   wire signed [9:0] m345_94;
   assign m345_94 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_95 = W*in
   wire signed [9:0] m345_95;
   assign m345_95 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_96 = W*in
   wire signed [9:0] m345_96;
   assign m345_96 =10'b0;

   // m345_97 = W*in
   wire signed [9:0] m345_97;
   assign m345_97 =10'b0;

   // m345_98 = W*in
   wire signed [9:0] m345_98;
   assign m345_98 =10'b0;

   // m345_99 = W*in
   wire signed [9:0] m345_99;
   assign m345_99 =10'b0;

   // m345_100 = W*in
   wire signed [9:0] m345_100;
   assign m345_100 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_101 = W*in
   wire signed [9:0] m345_101;
   assign m345_101 =10'b0;

   // m345_102 = W*in
   wire signed [9:0] m345_102;
   assign m345_102 =10'b0;

   // m345_103 = W*in
   wire signed [9:0] m345_103;
   assign m345_103 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_104 = W*in
   wire signed [9:0] m345_104;
   assign m345_104 =10'b0;

   // m345_105 = W*in
   wire signed [9:0] m345_105;
   assign m345_105 =10'b0;

   // m345_106 = W*in
   wire signed [9:0] m345_106;
   assign m345_106 =10'b0;

   // m345_107 = W*in
   wire signed [9:0] m345_107;
   assign m345_107 =10'b0;

   // m345_108 = W*in
   wire signed [9:0] m345_108;
   assign m345_108 =10'b0;

   // m345_109 = W*in
   wire signed [9:0] m345_109;
   assign m345_109 =10'b0;

   // m345_110 = W*in
   wire signed [9:0] m345_110;
   assign m345_110 =10'b0;

   // m345_111 = W*in
   wire signed [9:0] m345_111;
   assign m345_111 =10'b0;

   // m345_112 = W*in
   wire signed [9:0] m345_112;
   assign m345_112 ={ {4{neg345[5]}} , neg345[5:0] };

   // m345_113 = W*in
   wire signed [9:0] m345_113;
   assign m345_113 =10'b0;

   // m345_114 = W*in
   wire signed [9:0] m345_114;
   assign m345_114 =10'b0;

   // m345_115 = W*in
   wire signed [9:0] m345_115;
   assign m345_115 =10'b0;

   // m345_116 = W*in
   wire signed [9:0] m345_116;
   assign m345_116 =10'b0;

   // m345_117 = W*in
   wire signed [9:0] m345_117;
   assign m345_117 =10'b0;

   // m346_1 = W*in
   wire signed [9:0] m346_1;
   assign m346_1 =10'b0;

   // m346_2 = W*in
   wire signed [9:0] m346_2;
   assign m346_2 =10'b0;

   // m346_3 = W*in
   wire signed [9:0] m346_3;
   assign m346_3 =10'b0;

   // m346_4 = W*in
   wire signed [9:0] m346_4;
   assign m346_4 =10'b0;

   // m346_5 = W*in
   wire signed [9:0] m346_5;
   assign m346_5 =10'b0;

   // m346_6 = W*in
   wire signed [9:0] m346_6;
   assign m346_6 =10'b0;

   // m346_7 = W*in
   wire signed [9:0] m346_7;
   assign m346_7 =10'b0;

   // m346_8 = W*in
   wire signed [9:0] m346_8;
   assign m346_8 =10'b0;

   // m346_9 = W*in
   wire signed [9:0] m346_9;
   assign m346_9 =10'b0;

   // m346_10 = W*in
   wire signed [9:0] m346_10;
   assign m346_10 =10'b0;

   // m346_11 = W*in
   wire signed [9:0] m346_11;
   assign m346_11 =10'b0;

   // m346_12 = W*in
   wire signed [9:0] m346_12;
   assign m346_12 =10'b0;

   // m346_13 = W*in
   wire signed [9:0] m346_13;
   assign m346_13 =10'b0;

   // m346_14 = W*in
   wire signed [9:0] m346_14;
   assign m346_14 =10'b0;

   // m346_15 = W*in
   wire signed [9:0] m346_15;
   assign m346_15 =10'b0;

   // m346_16 = W*in
   wire signed [9:0] m346_16;
   assign m346_16 =10'b0;

   // m346_17 = W*in
   wire signed [9:0] m346_17;
   assign m346_17 =10'b0;

   // m346_18 = W*in
   wire signed [9:0] m346_18;
   assign m346_18 =10'b0;

   // m346_19 = W*in
   wire signed [9:0] m346_19;
   assign m346_19 =10'b0;

   // m346_20 = W*in
   wire signed [9:0] m346_20;
   assign m346_20 ={ {5{in346[5]}} , in346[5:1] };

   // m346_21 = W*in
   wire signed [9:0] m346_21;
   assign m346_21 ={ {5{neg346[5]}} , neg346[5:1] };

   // m346_22 = W*in
   wire signed [9:0] m346_22;
   assign m346_22 ={ {4{in346[5]}} , in346[5:0] };

   // m346_23 = W*in
   wire signed [9:0] m346_23;
   assign m346_23 =10'b0;

   // m346_24 = W*in
   wire signed [9:0] m346_24;
   assign m346_24 =10'b0;

   // m346_25 = W*in
   wire signed [9:0] m346_25;
   assign m346_25 =10'b0;

   // m346_26 = W*in
   wire signed [9:0] m346_26;
   assign m346_26 =10'b0;

   // m346_27 = W*in
   wire signed [9:0] m346_27;
   assign m346_27 ={ {5{in346[5]}} , in346[5:1] };

   // m346_28 = W*in
   wire signed [9:0] m346_28;
   assign m346_28 ={ {5{in346[5]}} , in346[5:1] };

   // m346_29 = W*in
   wire signed [9:0] m346_29;
   assign m346_29 =10'b0;

   // m346_30 = W*in
   wire signed [9:0] m346_30;
   assign m346_30 ={ {5{neg346[5]}} , neg346[5:1] };

   // m346_31 = W*in
   wire signed [9:0] m346_31;
   assign m346_31 =10'b0;

   // m346_32 = W*in
   wire signed [9:0] m346_32;
   assign m346_32 =10'b0;

   // m346_33 = W*in
   wire signed [9:0] m346_33;
   assign m346_33 =10'b0;

   // m346_34 = W*in
   wire signed [9:0] m346_34;
   assign m346_34 ={ {5{in346[5]}} , in346[5:1] };

   // m346_35 = W*in
   wire signed [9:0] m346_35;
   assign m346_35 =10'b0;

   // m346_36 = W*in
   wire signed [9:0] m346_36;
   assign m346_36 =10'b0;

   // m346_37 = W*in
   wire signed [9:0] m346_37;
   assign m346_37 =10'b0;

   // m346_38 = W*in
   wire signed [9:0] m346_38;
   assign m346_38 =10'b0;

   // m346_39 = W*in
   wire signed [9:0] m346_39;
   assign m346_39 =10'b0;

   // m346_40 = W*in
   wire signed [9:0] m346_40;
   assign m346_40 =10'b0;

   // m346_41 = W*in
   wire signed [9:0] m346_41;
   assign m346_41 =10'b0;

   // m346_42 = W*in
   wire signed [9:0] m346_42;
   assign m346_42 ={ {4{neg346[5]}} , neg346[5:0] };

   // m346_43 = W*in
   wire signed [9:0] m346_43;
   assign m346_43 =10'b0;

   // m346_44 = W*in
   wire signed [9:0] m346_44;
   assign m346_44 =10'b0;

   // m346_45 = W*in
   wire signed [9:0] m346_45;
   assign m346_45 =10'b0;

   // m346_46 = W*in
   wire signed [9:0] m346_46;
   assign m346_46 =10'b0;

   // m346_47 = W*in
   wire signed [9:0] m346_47;
   assign m346_47 ={ {4{in346[5]}} , in346[5:0] };

   // m346_48 = W*in
   wire signed [9:0] m346_48;
   assign m346_48 =10'b0;

   // m346_49 = W*in
   wire signed [9:0] m346_49;
   assign m346_49 =10'b0;

   // m346_50 = W*in
   wire signed [9:0] m346_50;
   assign m346_50 =10'b0;

   // m346_51 = W*in
   wire signed [9:0] m346_51;
   assign m346_51 =10'b0;

   // m346_52 = W*in
   wire signed [9:0] m346_52;
   assign m346_52 =10'b0;

   // m346_53 = W*in
   wire signed [9:0] m346_53;
   assign m346_53 =10'b0;

   // m346_54 = W*in
   wire signed [9:0] m346_54;
   assign m346_54 =10'b0;

   // m346_55 = W*in
   wire signed [9:0] m346_55;
   assign m346_55 =10'b0;

   // m346_56 = W*in
   wire signed [9:0] m346_56;
   assign m346_56 =10'b0;

   // m346_57 = W*in
   wire signed [9:0] m346_57;
   assign m346_57 =10'b0;

   // m346_58 = W*in
   wire signed [9:0] m346_58;
   assign m346_58 =10'b0;

   // m346_59 = W*in
   wire signed [9:0] m346_59;
   assign m346_59 =10'b0;

   // m346_60 = W*in
   wire signed [9:0] m346_60;
   assign m346_60 =10'b0;

   // m346_61 = W*in
   wire signed [9:0] m346_61;
   assign m346_61 =10'b0;

   // m346_62 = W*in
   wire signed [9:0] m346_62;
   assign m346_62 =10'b0;

   // m346_63 = W*in
   wire signed [9:0] m346_63;
   assign m346_63 =10'b0;

   // m346_64 = W*in
   wire signed [9:0] m346_64;
   assign m346_64 =10'b0;

   // m346_65 = W*in
   wire signed [9:0] m346_65;
   assign m346_65 ={ {4{neg346[5]}} , neg346[5:0] };

   // m346_66 = W*in
   wire signed [9:0] m346_66;
   assign m346_66 ={ {4{neg346[5]}} , neg346[5:0] };

   // m346_67 = W*in
   wire signed [9:0] m346_67;
   assign m346_67 =10'b0;

   // m346_68 = W*in
   wire signed [9:0] m346_68;
   assign m346_68 =10'b0;

   // m346_69 = W*in
   wire signed [9:0] m346_69;
   assign m346_69 ={ {5{neg346[5]}} , neg346[5:1] };

   // m346_70 = W*in
   wire signed [9:0] m346_70;
   assign m346_70 ={ {5{neg346[5]}} , neg346[5:1] };

   // m346_71 = W*in
   wire signed [9:0] m346_71;
   assign m346_71 =10'b0;

   // m346_72 = W*in
   wire signed [9:0] m346_72;
   assign m346_72 ={ {5{in346[5]}} , in346[5:1] };

   // m346_73 = W*in
   wire signed [9:0] m346_73;
   assign m346_73 =10'b0;

   // m346_74 = W*in
   wire signed [9:0] m346_74;
   assign m346_74 =10'b0;

   // m346_75 = W*in
   wire signed [9:0] m346_75;
   assign m346_75 =10'b0;

   // m346_76 = W*in
   wire signed [9:0] m346_76;
   assign m346_76 =10'b0;

   // m346_77 = W*in
   wire signed [9:0] m346_77;
   assign m346_77 =10'b0;

   // m346_78 = W*in
   wire signed [9:0] m346_78;
   assign m346_78 =10'b0;

   // m346_79 = W*in
   wire signed [9:0] m346_79;
   assign m346_79 =10'b0;

   // m346_80 = W*in
   wire signed [9:0] m346_80;
   assign m346_80 =10'b0;

   // m346_81 = W*in
   wire signed [9:0] m346_81;
   assign m346_81 =10'b0;

   // m346_82 = W*in
   wire signed [9:0] m346_82;
   assign m346_82 =10'b0;

   // m346_83 = W*in
   wire signed [9:0] m346_83;
   assign m346_83 =10'b0;

   // m346_84 = W*in
   wire signed [9:0] m346_84;
   assign m346_84 =10'b0;

   // m346_85 = W*in
   wire signed [9:0] m346_85;
   assign m346_85 =10'b0;

   // m346_86 = W*in
   wire signed [9:0] m346_86;
   assign m346_86 =10'b0;

   // m346_87 = W*in
   wire signed [9:0] m346_87;
   assign m346_87 =10'b0;

   // m346_88 = W*in
   wire signed [9:0] m346_88;
   assign m346_88 =10'b0;

   // m346_89 = W*in
   wire signed [9:0] m346_89;
   assign m346_89 =10'b0;

   // m346_90 = W*in
   wire signed [9:0] m346_90;
   assign m346_90 =10'b0;

   // m346_91 = W*in
   wire signed [9:0] m346_91;
   assign m346_91 =10'b0;

   // m346_92 = W*in
   wire signed [9:0] m346_92;
   assign m346_92 =10'b0;

   // m346_93 = W*in
   wire signed [9:0] m346_93;
   assign m346_93 =10'b0;

   // m346_94 = W*in
   wire signed [9:0] m346_94;
   assign m346_94 ={ {4{neg346[5]}} , neg346[5:0] };

   // m346_95 = W*in
   wire signed [9:0] m346_95;
   assign m346_95 =10'b0;

   // m346_96 = W*in
   wire signed [9:0] m346_96;
   assign m346_96 =10'b0;

   // m346_97 = W*in
   wire signed [9:0] m346_97;
   assign m346_97 =10'b0;

   // m346_98 = W*in
   wire signed [9:0] m346_98;
   assign m346_98 =10'b0;

   // m346_99 = W*in
   wire signed [9:0] m346_99;
   assign m346_99 =10'b0;

   // m346_100 = W*in
   wire signed [9:0] m346_100;
   assign m346_100 ={ {4{neg346[5]}} , neg346[5:0] };

   // m346_101 = W*in
   wire signed [9:0] m346_101;
   assign m346_101 =10'b0;

   // m346_102 = W*in
   wire signed [9:0] m346_102;
   assign m346_102 =10'b0;

   // m346_103 = W*in
   wire signed [9:0] m346_103;
   assign m346_103 =10'b0;

   // m346_104 = W*in
   wire signed [9:0] m346_104;
   assign m346_104 =10'b0;

   // m346_105 = W*in
   wire signed [9:0] m346_105;
   assign m346_105 =10'b0;

   // m346_106 = W*in
   wire signed [9:0] m346_106;
   assign m346_106 =10'b0;

   // m346_107 = W*in
   wire signed [9:0] m346_107;
   assign m346_107 =10'b0;

   // m346_108 = W*in
   wire signed [9:0] m346_108;
   assign m346_108 =10'b0;

   // m346_109 = W*in
   wire signed [9:0] m346_109;
   assign m346_109 =10'b0;

   // m346_110 = W*in
   wire signed [9:0] m346_110;
   assign m346_110 =10'b0;

   // m346_111 = W*in
   wire signed [9:0] m346_111;
   assign m346_111 =10'b0;

   // m346_112 = W*in
   wire signed [9:0] m346_112;
   assign m346_112 =10'b0;

   // m346_113 = W*in
   wire signed [9:0] m346_113;
   assign m346_113 =10'b0;

   // m346_114 = W*in
   wire signed [9:0] m346_114;
   assign m346_114 ={ {4{in346[5]}} , in346[5:0] };

   // m346_115 = W*in
   wire signed [9:0] m346_115;
   assign m346_115 ={ {5{in346[5]}} , in346[5:1] };

   // m346_116 = W*in
   wire signed [9:0] m346_116;
   assign m346_116 =10'b0;

   // m346_117 = W*in
   wire signed [9:0] m346_117;
   assign m346_117 =10'b0;

   // m347_1 = W*in
   wire signed [9:0] m347_1;
   assign m347_1 =10'b0;

   // m347_2 = W*in
   wire signed [9:0] m347_2;
   assign m347_2 =10'b0;

   // m347_3 = W*in
   wire signed [9:0] m347_3;
   assign m347_3 =10'b0;

   // m347_4 = W*in
   wire signed [9:0] m347_4;
   assign m347_4 =10'b0;

   // m347_5 = W*in
   wire signed [9:0] m347_5;
   assign m347_5 =10'b0;

   // m347_6 = W*in
   wire signed [9:0] m347_6;
   assign m347_6 =10'b0;

   // m347_7 = W*in
   wire signed [9:0] m347_7;
   assign m347_7 =10'b0;

   // m347_8 = W*in
   wire signed [9:0] m347_8;
   assign m347_8 =10'b0;

   // m347_9 = W*in
   wire signed [9:0] m347_9;
   assign m347_9 =10'b0;

   // m347_10 = W*in
   wire signed [9:0] m347_10;
   assign m347_10 =10'b0;

   // m347_11 = W*in
   wire signed [9:0] m347_11;
   assign m347_11 =10'b0;

   // m347_12 = W*in
   wire signed [9:0] m347_12;
   assign m347_12 =10'b0;

   // m347_13 = W*in
   wire signed [9:0] m347_13;
   assign m347_13 =10'b0;

   // m347_14 = W*in
   wire signed [9:0] m347_14;
   assign m347_14 =10'b0;

   // m347_15 = W*in
   wire signed [9:0] m347_15;
   assign m347_15 =10'b0;

   // m347_16 = W*in
   wire signed [9:0] m347_16;
   assign m347_16 =10'b0;

   // m347_17 = W*in
   wire signed [9:0] m347_17;
   assign m347_17 =10'b0;

   // m347_18 = W*in
   wire signed [9:0] m347_18;
   assign m347_18 =10'b0;

   // m347_19 = W*in
   wire signed [9:0] m347_19;
   assign m347_19 =10'b0;

   // m347_20 = W*in
   wire signed [9:0] m347_20;
   assign m347_20 ={ {4{in347[5]}} , in347[5:0] };

   // m347_21 = W*in
   wire signed [9:0] m347_21;
   assign m347_21 ={ {4{neg347[5]}} , neg347[5:0] };

   // m347_22 = W*in
   wire signed [9:0] m347_22;
   assign m347_22 ={ {4{in347[5]}} , in347[5:0] };

   // m347_23 = W*in
   wire signed [9:0] m347_23;
   assign m347_23 ={ {4{in347[5]}} , in347[5:0] };

   // m347_24 = W*in
   wire signed [9:0] m347_24;
   assign m347_24 ={ {4{in347[5]}} , in347[5:0] };

   // m347_25 = W*in
   wire signed [9:0] m347_25;
   assign m347_25 ={ {5{in347[5]}} , in347[5:1] };

   // m347_26 = W*in
   wire signed [9:0] m347_26;
   assign m347_26 =10'b0;

   // m347_27 = W*in
   wire signed [9:0] m347_27;
   assign m347_27 ={ {4{in347[5]}} , in347[5:0] };

   // m347_28 = W*in
   wire signed [9:0] m347_28;
   assign m347_28 ={ {5{in347[5]}} , in347[5:1] };

   // m347_29 = W*in
   wire signed [9:0] m347_29;
   assign m347_29 =10'b0;

   // m347_30 = W*in
   wire signed [9:0] m347_30;
   assign m347_30 ={ {5{in347[5]}} , in347[5:1] };

   // m347_31 = W*in
   wire signed [9:0] m347_31;
   assign m347_31 =10'b0;

   // m347_32 = W*in
   wire signed [9:0] m347_32;
   assign m347_32 =10'b0;

   // m347_33 = W*in
   wire signed [9:0] m347_33;
   assign m347_33 =10'b0;

   // m347_34 = W*in
   wire signed [9:0] m347_34;
   assign m347_34 ={ {5{in347[5]}} , in347[5:1] };

   // m347_35 = W*in
   wire signed [9:0] m347_35;
   assign m347_35 =10'b0;

   // m347_36 = W*in
   wire signed [9:0] m347_36;
   assign m347_36 =10'b0;

   // m347_37 = W*in
   wire signed [9:0] m347_37;
   assign m347_37 =10'b0;

   // m347_38 = W*in
   wire signed [9:0] m347_38;
   assign m347_38 =10'b0;

   // m347_39 = W*in
   wire signed [9:0] m347_39;
   assign m347_39 =10'b0;

   // m347_40 = W*in
   wire signed [9:0] m347_40;
   assign m347_40 =10'b0;

   // m347_41 = W*in
   wire signed [9:0] m347_41;
   assign m347_41 =10'b0;

   // m347_42 = W*in
   wire signed [9:0] m347_42;
   assign m347_42 =10'b0;

   // m347_43 = W*in
   wire signed [9:0] m347_43;
   assign m347_43 =10'b0;

   // m347_44 = W*in
   wire signed [9:0] m347_44;
   assign m347_44 =10'b0;

   // m347_45 = W*in
   wire signed [9:0] m347_45;
   assign m347_45 =10'b0;

   // m347_46 = W*in
   wire signed [9:0] m347_46;
   assign m347_46 =10'b0;

   // m347_47 = W*in
   wire signed [9:0] m347_47;
   assign m347_47 =10'b0;

   // m347_48 = W*in
   wire signed [9:0] m347_48;
   assign m347_48 =10'b0;

   // m347_49 = W*in
   wire signed [9:0] m347_49;
   assign m347_49 =10'b0;

   // m347_50 = W*in
   wire signed [9:0] m347_50;
   assign m347_50 =10'b0;

   // m347_51 = W*in
   wire signed [9:0] m347_51;
   assign m347_51 =10'b0;

   // m347_52 = W*in
   wire signed [9:0] m347_52;
   assign m347_52 =10'b0;

   // m347_53 = W*in
   wire signed [9:0] m347_53;
   assign m347_53 =10'b0;

   // m347_54 = W*in
   wire signed [9:0] m347_54;
   assign m347_54 =10'b0;

   // m347_55 = W*in
   wire signed [9:0] m347_55;
   assign m347_55 =10'b0;

   // m347_56 = W*in
   wire signed [9:0] m347_56;
   assign m347_56 =10'b0;

   // m347_57 = W*in
   wire signed [9:0] m347_57;
   assign m347_57 =10'b0;

   // m347_58 = W*in
   wire signed [9:0] m347_58;
   assign m347_58 =10'b0;

   // m347_59 = W*in
   wire signed [9:0] m347_59;
   assign m347_59 =10'b0;

   // m347_60 = W*in
   wire signed [9:0] m347_60;
   assign m347_60 =10'b0;

   // m347_61 = W*in
   wire signed [9:0] m347_61;
   assign m347_61 =10'b0;

   // m347_62 = W*in
   wire signed [9:0] m347_62;
   assign m347_62 =10'b0;

   // m347_63 = W*in
   wire signed [9:0] m347_63;
   assign m347_63 =10'b0;

   // m347_64 = W*in
   wire signed [9:0] m347_64;
   assign m347_64 ={ {5{in347[5]}} , in347[5:1] };

   // m347_65 = W*in
   wire signed [9:0] m347_65;
   assign m347_65 ={ {5{neg347[5]}} , neg347[5:1] };

   // m347_66 = W*in
   wire signed [9:0] m347_66;
   assign m347_66 ={ {5{neg347[5]}} , neg347[5:1] };

   // m347_67 = W*in
   wire signed [9:0] m347_67;
   assign m347_67 ={ {4{neg347[5]}} , neg347[5:0] };

   // m347_68 = W*in
   wire signed [9:0] m347_68;
   assign m347_68 =10'b0;

   // m347_69 = W*in
   wire signed [9:0] m347_69;
   assign m347_69 ={ {4{neg347[5]}} , neg347[5:0] };

   // m347_70 = W*in
   wire signed [9:0] m347_70;
   assign m347_70 ={ {5{neg347[5]}} , neg347[5:1] };

   // m347_71 = W*in
   wire signed [9:0] m347_71;
   assign m347_71 =10'b0;

   // m347_72 = W*in
   wire signed [9:0] m347_72;
   assign m347_72 =10'b0;

   // m347_73 = W*in
   wire signed [9:0] m347_73;
   assign m347_73 =10'b0;

   // m347_74 = W*in
   wire signed [9:0] m347_74;
   assign m347_74 =10'b0;

   // m347_75 = W*in
   wire signed [9:0] m347_75;
   assign m347_75 =10'b0;

   // m347_76 = W*in
   wire signed [9:0] m347_76;
   assign m347_76 =10'b0;

   // m347_77 = W*in
   wire signed [9:0] m347_77;
   assign m347_77 =10'b0;

   // m347_78 = W*in
   wire signed [9:0] m347_78;
   assign m347_78 =10'b0;

   // m347_79 = W*in
   wire signed [9:0] m347_79;
   assign m347_79 =10'b0;

   // m347_80 = W*in
   wire signed [9:0] m347_80;
   assign m347_80 =10'b0;

   // m347_81 = W*in
   wire signed [9:0] m347_81;
   assign m347_81 =10'b0;

   // m347_82 = W*in
   wire signed [9:0] m347_82;
   assign m347_82 =10'b0;

   // m347_83 = W*in
   wire signed [9:0] m347_83;
   assign m347_83 =10'b0;

   // m347_84 = W*in
   wire signed [9:0] m347_84;
   assign m347_84 =10'b0;

   // m347_85 = W*in
   wire signed [9:0] m347_85;
   assign m347_85 =10'b0;

   // m347_86 = W*in
   wire signed [9:0] m347_86;
   assign m347_86 =10'b0;

   // m347_87 = W*in
   wire signed [9:0] m347_87;
   assign m347_87 =10'b0;

   // m347_88 = W*in
   wire signed [9:0] m347_88;
   assign m347_88 =10'b0;

   // m347_89 = W*in
   wire signed [9:0] m347_89;
   assign m347_89 =10'b0;

   // m347_90 = W*in
   wire signed [9:0] m347_90;
   assign m347_90 =10'b0;

   // m347_91 = W*in
   wire signed [9:0] m347_91;
   assign m347_91 =10'b0;

   // m347_92 = W*in
   wire signed [9:0] m347_92;
   assign m347_92 =10'b0;

   // m347_93 = W*in
   wire signed [9:0] m347_93;
   assign m347_93 =10'b0;

   // m347_94 = W*in
   wire signed [9:0] m347_94;
   assign m347_94 =10'b0;

   // m347_95 = W*in
   wire signed [9:0] m347_95;
   assign m347_95 =10'b0;

   // m347_96 = W*in
   wire signed [9:0] m347_96;
   assign m347_96 =10'b0;

   // m347_97 = W*in
   wire signed [9:0] m347_97;
   assign m347_97 =10'b0;

   // m347_98 = W*in
   wire signed [9:0] m347_98;
   assign m347_98 =10'b0;

   // m347_99 = W*in
   wire signed [9:0] m347_99;
   assign m347_99 =10'b0;

   // m347_100 = W*in
   wire signed [9:0] m347_100;
   assign m347_100 =10'b0;

   // m347_101 = W*in
   wire signed [9:0] m347_101;
   assign m347_101 =10'b0;

   // m347_102 = W*in
   wire signed [9:0] m347_102;
   assign m347_102 =10'b0;

   // m347_103 = W*in
   wire signed [9:0] m347_103;
   assign m347_103 =10'b0;

   // m347_104 = W*in
   wire signed [9:0] m347_104;
   assign m347_104 =10'b0;

   // m347_105 = W*in
   wire signed [9:0] m347_105;
   assign m347_105 =10'b0;

   // m347_106 = W*in
   wire signed [9:0] m347_106;
   assign m347_106 =10'b0;

   // m347_107 = W*in
   wire signed [9:0] m347_107;
   assign m347_107 =10'b0;

   // m347_108 = W*in
   wire signed [9:0] m347_108;
   assign m347_108 =10'b0;

   // m347_109 = W*in
   wire signed [9:0] m347_109;
   assign m347_109 =10'b0;

   // m347_110 = W*in
   wire signed [9:0] m347_110;
   assign m347_110 =10'b0;

   // m347_111 = W*in
   wire signed [9:0] m347_111;
   assign m347_111 =10'b0;

   // m347_112 = W*in
   wire signed [9:0] m347_112;
   assign m347_112 =10'b0;

   // m347_113 = W*in
   wire signed [9:0] m347_113;
   assign m347_113 =10'b0;

   // m347_114 = W*in
   wire signed [9:0] m347_114;
   assign m347_114 =10'b0;

   // m347_115 = W*in
   wire signed [9:0] m347_115;
   assign m347_115 ={ {5{in347[5]}} , in347[5:1] };

   // m347_116 = W*in
   wire signed [9:0] m347_116;
   assign m347_116 ={ {4{neg347[5]}} , neg347[5:0] };

   // m347_117 = W*in
   wire signed [9:0] m347_117;
   assign m347_117 ={ {4{in347[5]}} , in347[5:0] };

   // m348_1 = W*in
   wire signed [9:0] m348_1;
   assign m348_1 =10'b0;

   // m348_2 = W*in
   wire signed [9:0] m348_2;
   assign m348_2 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_3 = W*in
   wire signed [9:0] m348_3;
   assign m348_3 =10'b0;

   // m348_4 = W*in
   wire signed [9:0] m348_4;
   assign m348_4 =10'b0;

   // m348_5 = W*in
   wire signed [9:0] m348_5;
   assign m348_5 =10'b0;

   // m348_6 = W*in
   wire signed [9:0] m348_6;
   assign m348_6 ={ {4{in348[5]}} , in348[5:0] };

   // m348_7 = W*in
   wire signed [9:0] m348_7;
   assign m348_7 =10'b0;

   // m348_8 = W*in
   wire signed [9:0] m348_8;
   assign m348_8 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_9 = W*in
   wire signed [9:0] m348_9;
   assign m348_9 =10'b0;

   // m348_10 = W*in
   wire signed [9:0] m348_10;
   assign m348_10 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_11 = W*in
   wire signed [9:0] m348_11;
   assign m348_11 =10'b0;

   // m348_12 = W*in
   wire signed [9:0] m348_12;
   assign m348_12 =10'b0;

   // m348_13 = W*in
   wire signed [9:0] m348_13;
   assign m348_13 =10'b0;

   // m348_14 = W*in
   wire signed [9:0] m348_14;
   assign m348_14 =10'b0;

   // m348_15 = W*in
   wire signed [9:0] m348_15;
   assign m348_15 =10'b0;

   // m348_16 = W*in
   wire signed [9:0] m348_16;
   assign m348_16 ={ {5{neg348[5]}} , neg348[5:1] };

   // m348_17 = W*in
   wire signed [9:0] m348_17;
   assign m348_17 =10'b0;

   // m348_18 = W*in
   wire signed [9:0] m348_18;
   assign m348_18 =10'b0;

   // m348_19 = W*in
   wire signed [9:0] m348_19;
   assign m348_19 =10'b0;

   // m348_20 = W*in
   wire signed [9:0] m348_20;
   assign m348_20 ={ {5{in348[5]}} , in348[5:1] };

   // m348_21 = W*in
   wire signed [9:0] m348_21;
   assign m348_21 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_22 = W*in
   wire signed [9:0] m348_22;
   assign m348_22 ={ {4{in348[5]}} , in348[5:0] };

   // m348_23 = W*in
   wire signed [9:0] m348_23;
   assign m348_23 =10'b0;

   // m348_24 = W*in
   wire signed [9:0] m348_24;
   assign m348_24 =10'b0;

   // m348_25 = W*in
   wire signed [9:0] m348_25;
   assign m348_25 =10'b0;

   // m348_26 = W*in
   wire signed [9:0] m348_26;
   assign m348_26 =10'b0;

   // m348_27 = W*in
   wire signed [9:0] m348_27;
   assign m348_27 =10'b0;

   // m348_28 = W*in
   wire signed [9:0] m348_28;
   assign m348_28 =10'b0;

   // m348_29 = W*in
   wire signed [9:0] m348_29;
   assign m348_29 =10'b0;

   // m348_30 = W*in
   wire signed [9:0] m348_30;
   assign m348_30 =10'b0;

   // m348_31 = W*in
   wire signed [9:0] m348_31;
   assign m348_31 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_32 = W*in
   wire signed [9:0] m348_32;
   assign m348_32 =10'b0;

   // m348_33 = W*in
   wire signed [9:0] m348_33;
   assign m348_33 =10'b0;

   // m348_34 = W*in
   wire signed [9:0] m348_34;
   assign m348_34 =10'b0;

   // m348_35 = W*in
   wire signed [9:0] m348_35;
   assign m348_35 =10'b0;

   // m348_36 = W*in
   wire signed [9:0] m348_36;
   assign m348_36 =10'b0;

   // m348_37 = W*in
   wire signed [9:0] m348_37;
   assign m348_37 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_38 = W*in
   wire signed [9:0] m348_38;
   assign m348_38 =10'b0;

   // m348_39 = W*in
   wire signed [9:0] m348_39;
   assign m348_39 =10'b0;

   // m348_40 = W*in
   wire signed [9:0] m348_40;
   assign m348_40 =10'b0;

   // m348_41 = W*in
   wire signed [9:0] m348_41;
   assign m348_41 =10'b0;

   // m348_42 = W*in
   wire signed [9:0] m348_42;
   assign m348_42 =10'b0;

   // m348_43 = W*in
   wire signed [9:0] m348_43;
   assign m348_43 =10'b0;

   // m348_44 = W*in
   wire signed [9:0] m348_44;
   assign m348_44 =10'b0;

   // m348_45 = W*in
   wire signed [9:0] m348_45;
   assign m348_45 =10'b0;

   // m348_46 = W*in
   wire signed [9:0] m348_46;
   assign m348_46 =10'b0;

   // m348_47 = W*in
   wire signed [9:0] m348_47;
   assign m348_47 =10'b0;

   // m348_48 = W*in
   wire signed [9:0] m348_48;
   assign m348_48 =10'b0;

   // m348_49 = W*in
   wire signed [9:0] m348_49;
   assign m348_49 ={ {4{in348[5]}} , in348[5:0] };

   // m348_50 = W*in
   wire signed [9:0] m348_50;
   assign m348_50 =10'b0;

   // m348_51 = W*in
   wire signed [9:0] m348_51;
   assign m348_51 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_52 = W*in
   wire signed [9:0] m348_52;
   assign m348_52 =10'b0;

   // m348_53 = W*in
   wire signed [9:0] m348_53;
   assign m348_53 =10'b0;

   // m348_54 = W*in
   wire signed [9:0] m348_54;
   assign m348_54 =10'b0;

   // m348_55 = W*in
   wire signed [9:0] m348_55;
   assign m348_55 =10'b0;

   // m348_56 = W*in
   wire signed [9:0] m348_56;
   assign m348_56 =10'b0;

   // m348_57 = W*in
   wire signed [9:0] m348_57;
   assign m348_57 =10'b0;

   // m348_58 = W*in
   wire signed [9:0] m348_58;
   assign m348_58 =10'b0;

   // m348_59 = W*in
   wire signed [9:0] m348_59;
   assign m348_59 =10'b0;

   // m348_60 = W*in
   wire signed [9:0] m348_60;
   assign m348_60 ={ {4{in348[5]}} , in348[5:0] };

   // m348_61 = W*in
   wire signed [9:0] m348_61;
   assign m348_61 =10'b0;

   // m348_62 = W*in
   wire signed [9:0] m348_62;
   assign m348_62 =10'b0;

   // m348_63 = W*in
   wire signed [9:0] m348_63;
   assign m348_63 =10'b0;

   // m348_64 = W*in
   wire signed [9:0] m348_64;
   assign m348_64 =10'b0;

   // m348_65 = W*in
   wire signed [9:0] m348_65;
   assign m348_65 =10'b0;

   // m348_66 = W*in
   wire signed [9:0] m348_66;
   assign m348_66 =10'b0;

   // m348_67 = W*in
   wire signed [9:0] m348_67;
   assign m348_67 =10'b0;

   // m348_68 = W*in
   wire signed [9:0] m348_68;
   assign m348_68 =10'b0;

   // m348_69 = W*in
   wire signed [9:0] m348_69;
   assign m348_69 =10'b0;

   // m348_70 = W*in
   wire signed [9:0] m348_70;
   assign m348_70 ={ {5{neg348[5]}} , neg348[5:1] };

   // m348_71 = W*in
   wire signed [9:0] m348_71;
   assign m348_71 =10'b0;

   // m348_72 = W*in
   wire signed [9:0] m348_72;
   assign m348_72 =10'b0;

   // m348_73 = W*in
   wire signed [9:0] m348_73;
   assign m348_73 =10'b0;

   // m348_74 = W*in
   wire signed [9:0] m348_74;
   assign m348_74 ={ {5{in348[5]}} , in348[5:1] };

   // m348_75 = W*in
   wire signed [9:0] m348_75;
   assign m348_75 =10'b0;

   // m348_76 = W*in
   wire signed [9:0] m348_76;
   assign m348_76 =10'b0;

   // m348_77 = W*in
   wire signed [9:0] m348_77;
   assign m348_77 =10'b0;

   // m348_78 = W*in
   wire signed [9:0] m348_78;
   assign m348_78 =10'b0;

   // m348_79 = W*in
   wire signed [9:0] m348_79;
   assign m348_79 =10'b0;

   // m348_80 = W*in
   wire signed [9:0] m348_80;
   assign m348_80 ={ {5{neg348[5]}} , neg348[5:1] };

   // m348_81 = W*in
   wire signed [9:0] m348_81;
   assign m348_81 ={ {5{in348[5]}} , in348[5:1] };

   // m348_82 = W*in
   wire signed [9:0] m348_82;
   assign m348_82 =10'b0;

   // m348_83 = W*in
   wire signed [9:0] m348_83;
   assign m348_83 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_84 = W*in
   wire signed [9:0] m348_84;
   assign m348_84 =10'b0;

   // m348_85 = W*in
   wire signed [9:0] m348_85;
   assign m348_85 =10'b0;

   // m348_86 = W*in
   wire signed [9:0] m348_86;
   assign m348_86 =10'b0;

   // m348_87 = W*in
   wire signed [9:0] m348_87;
   assign m348_87 =10'b0;

   // m348_88 = W*in
   wire signed [9:0] m348_88;
   assign m348_88 =10'b0;

   // m348_89 = W*in
   wire signed [9:0] m348_89;
   assign m348_89 =10'b0;

   // m348_90 = W*in
   wire signed [9:0] m348_90;
   assign m348_90 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_91 = W*in
   wire signed [9:0] m348_91;
   assign m348_91 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_92 = W*in
   wire signed [9:0] m348_92;
   assign m348_92 =10'b0;

   // m348_93 = W*in
   wire signed [9:0] m348_93;
   assign m348_93 =10'b0;

   // m348_94 = W*in
   wire signed [9:0] m348_94;
   assign m348_94 =10'b0;

   // m348_95 = W*in
   wire signed [9:0] m348_95;
   assign m348_95 =10'b0;

   // m348_96 = W*in
   wire signed [9:0] m348_96;
   assign m348_96 =10'b0;

   // m348_97 = W*in
   wire signed [9:0] m348_97;
   assign m348_97 =10'b0;

   // m348_98 = W*in
   wire signed [9:0] m348_98;
   assign m348_98 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_99 = W*in
   wire signed [9:0] m348_99;
   assign m348_99 =10'b0;

   // m348_100 = W*in
   wire signed [9:0] m348_100;
   assign m348_100 =10'b0;

   // m348_101 = W*in
   wire signed [9:0] m348_101;
   assign m348_101 =10'b0;

   // m348_102 = W*in
   wire signed [9:0] m348_102;
   assign m348_102 =10'b0;

   // m348_103 = W*in
   wire signed [9:0] m348_103;
   assign m348_103 =10'b0;

   // m348_104 = W*in
   wire signed [9:0] m348_104;
   assign m348_104 =10'b0;

   // m348_105 = W*in
   wire signed [9:0] m348_105;
   assign m348_105 ={ {4{neg348[5]}} , neg348[5:0] };

   // m348_106 = W*in
   wire signed [9:0] m348_106;
   assign m348_106 =10'b0;

   // m348_107 = W*in
   wire signed [9:0] m348_107;
   assign m348_107 =10'b0;

   // m348_108 = W*in
   wire signed [9:0] m348_108;
   assign m348_108 =10'b0;

   // m348_109 = W*in
   wire signed [9:0] m348_109;
   assign m348_109 =10'b0;

   // m348_110 = W*in
   wire signed [9:0] m348_110;
   assign m348_110 =10'b0;

   // m348_111 = W*in
   wire signed [9:0] m348_111;
   assign m348_111 =10'b0;

   // m348_112 = W*in
   wire signed [9:0] m348_112;
   assign m348_112 =10'b0;

   // m348_113 = W*in
   wire signed [9:0] m348_113;
   assign m348_113 =10'b0;

   // m348_114 = W*in
   wire signed [9:0] m348_114;
   assign m348_114 =10'b0;

   // m348_115 = W*in
   wire signed [9:0] m348_115;
   assign m348_115 =10'b0;

   // m348_116 = W*in
   wire signed [9:0] m348_116;
   assign m348_116 =10'b0;

   // m348_117 = W*in
   wire signed [9:0] m348_117;
   assign m348_117 ={ {4{in348[5]}} , in348[5:0] };

   // m349_1 = W*in
   wire signed [9:0] m349_1;
   assign m349_1 =10'b0;

   // m349_2 = W*in
   wire signed [9:0] m349_2;
   assign m349_2 =10'b0;

   // m349_3 = W*in
   wire signed [9:0] m349_3;
   assign m349_3 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_4 = W*in
   wire signed [9:0] m349_4;
   assign m349_4 =10'b0;

   // m349_5 = W*in
   wire signed [9:0] m349_5;
   assign m349_5 =10'b0;

   // m349_6 = W*in
   wire signed [9:0] m349_6;
   assign m349_6 =10'b0;

   // m349_7 = W*in
   wire signed [9:0] m349_7;
   assign m349_7 =10'b0;

   // m349_8 = W*in
   wire signed [9:0] m349_8;
   assign m349_8 =10'b0;

   // m349_9 = W*in
   wire signed [9:0] m349_9;
   assign m349_9 =10'b0;

   // m349_10 = W*in
   wire signed [9:0] m349_10;
   assign m349_10 =10'b0;

   // m349_11 = W*in
   wire signed [9:0] m349_11;
   assign m349_11 =10'b0;

   // m349_12 = W*in
   wire signed [9:0] m349_12;
   assign m349_12 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_13 = W*in
   wire signed [9:0] m349_13;
   assign m349_13 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_14 = W*in
   wire signed [9:0] m349_14;
   assign m349_14 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_15 = W*in
   wire signed [9:0] m349_15;
   assign m349_15 =10'b0;

   // m349_16 = W*in
   wire signed [9:0] m349_16;
   assign m349_16 ={ {5{in349[5]}} , in349[5:1] };

   // m349_17 = W*in
   wire signed [9:0] m349_17;
   assign m349_17 =10'b0;

   // m349_18 = W*in
   wire signed [9:0] m349_18;
   assign m349_18 =10'b0;

   // m349_19 = W*in
   wire signed [9:0] m349_19;
   assign m349_19 =10'b0;

   // m349_20 = W*in
   wire signed [9:0] m349_20;
   assign m349_20 ={ {5{in349[5]}} , in349[5:1] };

   // m349_21 = W*in
   wire signed [9:0] m349_21;
   assign m349_21 ={ {5{neg349[5]}} , neg349[5:1] };

   // m349_22 = W*in
   wire signed [9:0] m349_22;
   assign m349_22 =10'b0;

   // m349_23 = W*in
   wire signed [9:0] m349_23;
   assign m349_23 =10'b0;

   // m349_24 = W*in
   wire signed [9:0] m349_24;
   assign m349_24 =10'b0;

   // m349_25 = W*in
   wire signed [9:0] m349_25;
   assign m349_25 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_26 = W*in
   wire signed [9:0] m349_26;
   assign m349_26 =10'b0;

   // m349_27 = W*in
   wire signed [9:0] m349_27;
   assign m349_27 ={ {5{neg349[5]}} , neg349[5:1] };

   // m349_28 = W*in
   wire signed [9:0] m349_28;
   assign m349_28 =10'b0;

   // m349_29 = W*in
   wire signed [9:0] m349_29;
   assign m349_29 =10'b0;

   // m349_30 = W*in
   wire signed [9:0] m349_30;
   assign m349_30 =10'b0;

   // m349_31 = W*in
   wire signed [9:0] m349_31;
   assign m349_31 =10'b0;

   // m349_32 = W*in
   wire signed [9:0] m349_32;
   assign m349_32 ={ {5{in349[5]}} , in349[5:1] };

   // m349_33 = W*in
   wire signed [9:0] m349_33;
   assign m349_33 =10'b0;

   // m349_34 = W*in
   wire signed [9:0] m349_34;
   assign m349_34 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_35 = W*in
   wire signed [9:0] m349_35;
   assign m349_35 =10'b0;

   // m349_36 = W*in
   wire signed [9:0] m349_36;
   assign m349_36 =10'b0;

   // m349_37 = W*in
   wire signed [9:0] m349_37;
   assign m349_37 =10'b0;

   // m349_38 = W*in
   wire signed [9:0] m349_38;
   assign m349_38 =10'b0;

   // m349_39 = W*in
   wire signed [9:0] m349_39;
   assign m349_39 =10'b0;

   // m349_40 = W*in
   wire signed [9:0] m349_40;
   assign m349_40 =10'b0;

   // m349_41 = W*in
   wire signed [9:0] m349_41;
   assign m349_41 =10'b0;

   // m349_42 = W*in
   wire signed [9:0] m349_42;
   assign m349_42 ={ {4{in349[5]}} , in349[5:0] };

   // m349_43 = W*in
   wire signed [9:0] m349_43;
   assign m349_43 =10'b0;

   // m349_44 = W*in
   wire signed [9:0] m349_44;
   assign m349_44 =10'b0;

   // m349_45 = W*in
   wire signed [9:0] m349_45;
   assign m349_45 =10'b0;

   // m349_46 = W*in
   wire signed [9:0] m349_46;
   assign m349_46 =10'b0;

   // m349_47 = W*in
   wire signed [9:0] m349_47;
   assign m349_47 =10'b0;

   // m349_48 = W*in
   wire signed [9:0] m349_48;
   assign m349_48 =10'b0;

   // m349_49 = W*in
   wire signed [9:0] m349_49;
   assign m349_49 =10'b0;

   // m349_50 = W*in
   wire signed [9:0] m349_50;
   assign m349_50 =10'b0;

   // m349_51 = W*in
   wire signed [9:0] m349_51;
   assign m349_51 ={ {4{in349[5]}} , in349[5:0] };

   // m349_52 = W*in
   wire signed [9:0] m349_52;
   assign m349_52 =10'b0;

   // m349_53 = W*in
   wire signed [9:0] m349_53;
   assign m349_53 =10'b0;

   // m349_54 = W*in
   wire signed [9:0] m349_54;
   assign m349_54 =10'b0;

   // m349_55 = W*in
   wire signed [9:0] m349_55;
   assign m349_55 =10'b0;

   // m349_56 = W*in
   wire signed [9:0] m349_56;
   assign m349_56 =10'b0;

   // m349_57 = W*in
   wire signed [9:0] m349_57;
   assign m349_57 =10'b0;

   // m349_58 = W*in
   wire signed [9:0] m349_58;
   assign m349_58 =10'b0;

   // m349_59 = W*in
   wire signed [9:0] m349_59;
   assign m349_59 =10'b0;

   // m349_60 = W*in
   wire signed [9:0] m349_60;
   assign m349_60 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_61 = W*in
   wire signed [9:0] m349_61;
   assign m349_61 ={ {4{in349[5]}} , in349[5:0] };

   // m349_62 = W*in
   wire signed [9:0] m349_62;
   assign m349_62 =10'b0;

   // m349_63 = W*in
   wire signed [9:0] m349_63;
   assign m349_63 =10'b0;

   // m349_64 = W*in
   wire signed [9:0] m349_64;
   assign m349_64 ={ {4{in349[5]}} , in349[5:0] };

   // m349_65 = W*in
   wire signed [9:0] m349_65;
   assign m349_65 ={ {5{in349[5]}} , in349[5:1] };

   // m349_66 = W*in
   wire signed [9:0] m349_66;
   assign m349_66 =10'b0;

   // m349_67 = W*in
   wire signed [9:0] m349_67;
   assign m349_67 =10'b0;

   // m349_68 = W*in
   wire signed [9:0] m349_68;
   assign m349_68 =10'b0;

   // m349_69 = W*in
   wire signed [9:0] m349_69;
   assign m349_69 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_70 = W*in
   wire signed [9:0] m349_70;
   assign m349_70 =10'b0;

   // m349_71 = W*in
   wire signed [9:0] m349_71;
   assign m349_71 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_72 = W*in
   wire signed [9:0] m349_72;
   assign m349_72 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_73 = W*in
   wire signed [9:0] m349_73;
   assign m349_73 ={ {5{neg349[5]}} , neg349[5:1] };

   // m349_74 = W*in
   wire signed [9:0] m349_74;
   assign m349_74 =10'b0;

   // m349_75 = W*in
   wire signed [9:0] m349_75;
   assign m349_75 ={ {4{in349[5]}} , in349[5:0] };

   // m349_76 = W*in
   wire signed [9:0] m349_76;
   assign m349_76 =10'b0;

   // m349_77 = W*in
   wire signed [9:0] m349_77;
   assign m349_77 =10'b0;

   // m349_78 = W*in
   wire signed [9:0] m349_78;
   assign m349_78 =10'b0;

   // m349_79 = W*in
   wire signed [9:0] m349_79;
   assign m349_79 =10'b0;

   // m349_80 = W*in
   wire signed [9:0] m349_80;
   assign m349_80 =10'b0;

   // m349_81 = W*in
   wire signed [9:0] m349_81;
   assign m349_81 ={ {4{in349[5]}} , in349[5:0] };

   // m349_82 = W*in
   wire signed [9:0] m349_82;
   assign m349_82 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_83 = W*in
   wire signed [9:0] m349_83;
   assign m349_83 ={ {4{in349[5]}} , in349[5:0] };

   // m349_84 = W*in
   wire signed [9:0] m349_84;
   assign m349_84 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_85 = W*in
   wire signed [9:0] m349_85;
   assign m349_85 =10'b0;

   // m349_86 = W*in
   wire signed [9:0] m349_86;
   assign m349_86 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_87 = W*in
   wire signed [9:0] m349_87;
   assign m349_87 =10'b0;

   // m349_88 = W*in
   wire signed [9:0] m349_88;
   assign m349_88 =10'b0;

   // m349_89 = W*in
   wire signed [9:0] m349_89;
   assign m349_89 =10'b0;

   // m349_90 = W*in
   wire signed [9:0] m349_90;
   assign m349_90 =10'b0;

   // m349_91 = W*in
   wire signed [9:0] m349_91;
   assign m349_91 ={ {5{neg349[5]}} , neg349[5:1] };

   // m349_92 = W*in
   wire signed [9:0] m349_92;
   assign m349_92 =10'b0;

   // m349_93 = W*in
   wire signed [9:0] m349_93;
   assign m349_93 =10'b0;

   // m349_94 = W*in
   wire signed [9:0] m349_94;
   assign m349_94 ={ {4{in349[5]}} , in349[5:0] };

   // m349_95 = W*in
   wire signed [9:0] m349_95;
   assign m349_95 =10'b0;

   // m349_96 = W*in
   wire signed [9:0] m349_96;
   assign m349_96 =10'b0;

   // m349_97 = W*in
   wire signed [9:0] m349_97;
   assign m349_97 =10'b0;

   // m349_98 = W*in
   wire signed [9:0] m349_98;
   assign m349_98 =10'b0;

   // m349_99 = W*in
   wire signed [9:0] m349_99;
   assign m349_99 =10'b0;

   // m349_100 = W*in
   wire signed [9:0] m349_100;
   assign m349_100 =10'b0;

   // m349_101 = W*in
   wire signed [9:0] m349_101;
   assign m349_101 =10'b0;

   // m349_102 = W*in
   wire signed [9:0] m349_102;
   assign m349_102 =10'b0;

   // m349_103 = W*in
   wire signed [9:0] m349_103;
   assign m349_103 ={ {5{neg349[5]}} , neg349[5:1] };

   // m349_104 = W*in
   wire signed [9:0] m349_104;
   assign m349_104 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_105 = W*in
   wire signed [9:0] m349_105;
   assign m349_105 =10'b0;

   // m349_106 = W*in
   wire signed [9:0] m349_106;
   assign m349_106 =10'b0;

   // m349_107 = W*in
   wire signed [9:0] m349_107;
   assign m349_107 =10'b0;

   // m349_108 = W*in
   wire signed [9:0] m349_108;
   assign m349_108 =10'b0;

   // m349_109 = W*in
   wire signed [9:0] m349_109;
   assign m349_109 =10'b0;

   // m349_110 = W*in
   wire signed [9:0] m349_110;
   assign m349_110 =10'b0;

   // m349_111 = W*in
   wire signed [9:0] m349_111;
   assign m349_111 ={ {4{neg349[5]}} , neg349[5:0] };

   // m349_112 = W*in
   wire signed [9:0] m349_112;
   assign m349_112 =10'b0;

   // m349_113 = W*in
   wire signed [9:0] m349_113;
   assign m349_113 =10'b0;

   // m349_114 = W*in
   wire signed [9:0] m349_114;
   assign m349_114 =10'b0;

   // m349_115 = W*in
   wire signed [9:0] m349_115;
   assign m349_115 ={ {4{in349[5]}} , in349[5:0] };

   // m349_116 = W*in
   wire signed [9:0] m349_116;
   assign m349_116 =10'b0;

   // m349_117 = W*in
   wire signed [9:0] m349_117;
   assign m349_117 =10'b0;

   // m350_1 = W*in
   wire signed [9:0] m350_1;
   assign m350_1 =10'b0;

   // m350_2 = W*in
   wire signed [9:0] m350_2;
   assign m350_2 =10'b0;

   // m350_3 = W*in
   wire signed [9:0] m350_3;
   assign m350_3 =10'b0;

   // m350_4 = W*in
   wire signed [9:0] m350_4;
   assign m350_4 =10'b0;

   // m350_5 = W*in
   wire signed [9:0] m350_5;
   assign m350_5 =10'b0;

   // m350_6 = W*in
   wire signed [9:0] m350_6;
   assign m350_6 =10'b0;

   // m350_7 = W*in
   wire signed [9:0] m350_7;
   assign m350_7 =10'b0;

   // m350_8 = W*in
   wire signed [9:0] m350_8;
   assign m350_8 =10'b0;

   // m350_9 = W*in
   wire signed [9:0] m350_9;
   assign m350_9 =10'b0;

   // m350_10 = W*in
   wire signed [9:0] m350_10;
   assign m350_10 ={ {4{in350[5]}} , in350[5:0] };

   // m350_11 = W*in
   wire signed [9:0] m350_11;
   assign m350_11 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_12 = W*in
   wire signed [9:0] m350_12;
   assign m350_12 =10'b0;

   // m350_13 = W*in
   wire signed [9:0] m350_13;
   assign m350_13 =10'b0;

   // m350_14 = W*in
   wire signed [9:0] m350_14;
   assign m350_14 =10'b0;

   // m350_15 = W*in
   wire signed [9:0] m350_15;
   assign m350_15 =10'b0;

   // m350_16 = W*in
   wire signed [9:0] m350_16;
   assign m350_16 =10'b0;

   // m350_17 = W*in
   wire signed [9:0] m350_17;
   assign m350_17 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_18 = W*in
   wire signed [9:0] m350_18;
   assign m350_18 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_19 = W*in
   wire signed [9:0] m350_19;
   assign m350_19 =10'b0;

   // m350_20 = W*in
   wire signed [9:0] m350_20;
   assign m350_20 =10'b0;

   // m350_21 = W*in
   wire signed [9:0] m350_21;
   assign m350_21 =10'b0;

   // m350_22 = W*in
   wire signed [9:0] m350_22;
   assign m350_22 =10'b0;

   // m350_23 = W*in
   wire signed [9:0] m350_23;
   assign m350_23 =10'b0;

   // m350_24 = W*in
   wire signed [9:0] m350_24;
   assign m350_24 =10'b0;

   // m350_25 = W*in
   wire signed [9:0] m350_25;
   assign m350_25 ={ {4{in350[5]}} , in350[5:0] };

   // m350_26 = W*in
   wire signed [9:0] m350_26;
   assign m350_26 =10'b0;

   // m350_27 = W*in
   wire signed [9:0] m350_27;
   assign m350_27 =10'b0;

   // m350_28 = W*in
   wire signed [9:0] m350_28;
   assign m350_28 =10'b0;

   // m350_29 = W*in
   wire signed [9:0] m350_29;
   assign m350_29 =10'b0;

   // m350_30 = W*in
   wire signed [9:0] m350_30;
   assign m350_30 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_31 = W*in
   wire signed [9:0] m350_31;
   assign m350_31 =10'b0;

   // m350_32 = W*in
   wire signed [9:0] m350_32;
   assign m350_32 ={ {4{in350[5]}} , in350[5:0] };

   // m350_33 = W*in
   wire signed [9:0] m350_33;
   assign m350_33 ={ {4{in350[5]}} , in350[5:0] };

   // m350_34 = W*in
   wire signed [9:0] m350_34;
   assign m350_34 ={ {5{neg350[5]}} , neg350[5:1] };

   // m350_35 = W*in
   wire signed [9:0] m350_35;
   assign m350_35 ={ {5{neg350[5]}} , neg350[5:1] };

   // m350_36 = W*in
   wire signed [9:0] m350_36;
   assign m350_36 =10'b0;

   // m350_37 = W*in
   wire signed [9:0] m350_37;
   assign m350_37 ={ {4{in350[5]}} , in350[5:0] };

   // m350_38 = W*in
   wire signed [9:0] m350_38;
   assign m350_38 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_39 = W*in
   wire signed [9:0] m350_39;
   assign m350_39 =10'b0;

   // m350_40 = W*in
   wire signed [9:0] m350_40;
   assign m350_40 =10'b0;

   // m350_41 = W*in
   wire signed [9:0] m350_41;
   assign m350_41 =10'b0;

   // m350_42 = W*in
   wire signed [9:0] m350_42;
   assign m350_42 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_43 = W*in
   wire signed [9:0] m350_43;
   assign m350_43 =10'b0;

   // m350_44 = W*in
   wire signed [9:0] m350_44;
   assign m350_44 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_45 = W*in
   wire signed [9:0] m350_45;
   assign m350_45 ={ {4{in350[5]}} , in350[5:0] };

   // m350_46 = W*in
   wire signed [9:0] m350_46;
   assign m350_46 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_47 = W*in
   wire signed [9:0] m350_47;
   assign m350_47 =10'b0;

   // m350_48 = W*in
   wire signed [9:0] m350_48;
   assign m350_48 ={ {4{in350[5]}} , in350[5:0] };

   // m350_49 = W*in
   wire signed [9:0] m350_49;
   assign m350_49 =10'b0;

   // m350_50 = W*in
   wire signed [9:0] m350_50;
   assign m350_50 =10'b0;

   // m350_51 = W*in
   wire signed [9:0] m350_51;
   assign m350_51 ={ {4{in350[5]}} , in350[5:0] };

   // m350_52 = W*in
   wire signed [9:0] m350_52;
   assign m350_52 =10'b0;

   // m350_53 = W*in
   wire signed [9:0] m350_53;
   assign m350_53 =10'b0;

   // m350_54 = W*in
   wire signed [9:0] m350_54;
   assign m350_54 =10'b0;

   // m350_55 = W*in
   wire signed [9:0] m350_55;
   assign m350_55 =10'b0;

   // m350_56 = W*in
   wire signed [9:0] m350_56;
   assign m350_56 =10'b0;

   // m350_57 = W*in
   wire signed [9:0] m350_57;
   assign m350_57 =10'b0;

   // m350_58 = W*in
   wire signed [9:0] m350_58;
   assign m350_58 =10'b0;

   // m350_59 = W*in
   wire signed [9:0] m350_59;
   assign m350_59 =10'b0;

   // m350_60 = W*in
   wire signed [9:0] m350_60;
   assign m350_60 =10'b0;

   // m350_61 = W*in
   wire signed [9:0] m350_61;
   assign m350_61 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_62 = W*in
   wire signed [9:0] m350_62;
   assign m350_62 =10'b0;

   // m350_63 = W*in
   wire signed [9:0] m350_63;
   assign m350_63 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_64 = W*in
   wire signed [9:0] m350_64;
   assign m350_64 ={ {5{neg350[5]}} , neg350[5:1] };

   // m350_65 = W*in
   wire signed [9:0] m350_65;
   assign m350_65 ={ {5{neg350[5]}} , neg350[5:1] };

   // m350_66 = W*in
   wire signed [9:0] m350_66;
   assign m350_66 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_67 = W*in
   wire signed [9:0] m350_67;
   assign m350_67 =10'b0;

   // m350_68 = W*in
   wire signed [9:0] m350_68;
   assign m350_68 =10'b0;

   // m350_69 = W*in
   wire signed [9:0] m350_69;
   assign m350_69 =10'b0;

   // m350_70 = W*in
   wire signed [9:0] m350_70;
   assign m350_70 =10'b0;

   // m350_71 = W*in
   wire signed [9:0] m350_71;
   assign m350_71 ={ {5{neg350[5]}} , neg350[5:1] };

   // m350_72 = W*in
   wire signed [9:0] m350_72;
   assign m350_72 =10'b0;

   // m350_73 = W*in
   wire signed [9:0] m350_73;
   assign m350_73 =10'b0;

   // m350_74 = W*in
   wire signed [9:0] m350_74;
   assign m350_74 =10'b0;

   // m350_75 = W*in
   wire signed [9:0] m350_75;
   assign m350_75 =10'b0;

   // m350_76 = W*in
   wire signed [9:0] m350_76;
   assign m350_76 =10'b0;

   // m350_77 = W*in
   wire signed [9:0] m350_77;
   assign m350_77 =10'b0;

   // m350_78 = W*in
   wire signed [9:0] m350_78;
   assign m350_78 =10'b0;

   // m350_79 = W*in
   wire signed [9:0] m350_79;
   assign m350_79 =10'b0;

   // m350_80 = W*in
   wire signed [9:0] m350_80;
   assign m350_80 =10'b0;

   // m350_81 = W*in
   wire signed [9:0] m350_81;
   assign m350_81 =10'b0;

   // m350_82 = W*in
   wire signed [9:0] m350_82;
   assign m350_82 =10'b0;

   // m350_83 = W*in
   wire signed [9:0] m350_83;
   assign m350_83 ={ {4{in350[5]}} , in350[5:0] };

   // m350_84 = W*in
   wire signed [9:0] m350_84;
   assign m350_84 ={ {5{in350[5]}} , in350[5:1] };

   // m350_85 = W*in
   wire signed [9:0] m350_85;
   assign m350_85 =10'b0;

   // m350_86 = W*in
   wire signed [9:0] m350_86;
   assign m350_86 =10'b0;

   // m350_87 = W*in
   wire signed [9:0] m350_87;
   assign m350_87 =10'b0;

   // m350_88 = W*in
   wire signed [9:0] m350_88;
   assign m350_88 =10'b0;

   // m350_89 = W*in
   wire signed [9:0] m350_89;
   assign m350_89 =10'b0;

   // m350_90 = W*in
   wire signed [9:0] m350_90;
   assign m350_90 =10'b0;

   // m350_91 = W*in
   wire signed [9:0] m350_91;
   assign m350_91 ={ {3{neg350[5]}} , neg350 , {1{1'b0}} };

   // m350_92 = W*in
   wire signed [9:0] m350_92;
   assign m350_92 =10'b0;

   // m350_93 = W*in
   wire signed [9:0] m350_93;
   assign m350_93 =10'b0;

   // m350_94 = W*in
   wire signed [9:0] m350_94;
   assign m350_94 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_95 = W*in
   wire signed [9:0] m350_95;
   assign m350_95 =10'b0;

   // m350_96 = W*in
   wire signed [9:0] m350_96;
   assign m350_96 =10'b0;

   // m350_97 = W*in
   wire signed [9:0] m350_97;
   assign m350_97 =10'b0;

   // m350_98 = W*in
   wire signed [9:0] m350_98;
   assign m350_98 =10'b0;

   // m350_99 = W*in
   wire signed [9:0] m350_99;
   assign m350_99 =10'b0;

   // m350_100 = W*in
   wire signed [9:0] m350_100;
   assign m350_100 =10'b0;

   // m350_101 = W*in
   wire signed [9:0] m350_101;
   assign m350_101 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_102 = W*in
   wire signed [9:0] m350_102;
   assign m350_102 =10'b0;

   // m350_103 = W*in
   wire signed [9:0] m350_103;
   assign m350_103 =10'b0;

   // m350_104 = W*in
   wire signed [9:0] m350_104;
   assign m350_104 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_105 = W*in
   wire signed [9:0] m350_105;
   assign m350_105 =10'b0;

   // m350_106 = W*in
   wire signed [9:0] m350_106;
   assign m350_106 =10'b0;

   // m350_107 = W*in
   wire signed [9:0] m350_107;
   assign m350_107 =10'b0;

   // m350_108 = W*in
   wire signed [9:0] m350_108;
   assign m350_108 =10'b0;

   // m350_109 = W*in
   wire signed [9:0] m350_109;
   assign m350_109 =10'b0;

   // m350_110 = W*in
   wire signed [9:0] m350_110;
   assign m350_110 ={ {4{neg350[5]}} , neg350[5:0] };

   // m350_111 = W*in
   wire signed [9:0] m350_111;
   assign m350_111 =10'b0;

   // m350_112 = W*in
   wire signed [9:0] m350_112;
   assign m350_112 =10'b0;

   // m350_113 = W*in
   wire signed [9:0] m350_113;
   assign m350_113 =10'b0;

   // m350_114 = W*in
   wire signed [9:0] m350_114;
   assign m350_114 =10'b0;

   // m350_115 = W*in
   wire signed [9:0] m350_115;
   assign m350_115 =10'b0;

   // m350_116 = W*in
   wire signed [9:0] m350_116;
   assign m350_116 =10'b0;

   // m350_117 = W*in
   wire signed [9:0] m350_117;
   assign m350_117 ={ {4{neg350[5]}} , neg350[5:0] };

   // m351_1 = W*in
   wire signed [9:0] m351_1;
   assign m351_1 =10'b0;

   // m351_2 = W*in
   wire signed [9:0] m351_2;
   assign m351_2 =10'b0;

   // m351_3 = W*in
   wire signed [9:0] m351_3;
   assign m351_3 =10'b0;

   // m351_4 = W*in
   wire signed [9:0] m351_4;
   assign m351_4 =10'b0;

   // m351_5 = W*in
   wire signed [9:0] m351_5;
   assign m351_5 =10'b0;

   // m351_6 = W*in
   wire signed [9:0] m351_6;
   assign m351_6 =10'b0;

   // m351_7 = W*in
   wire signed [9:0] m351_7;
   assign m351_7 =10'b0;

   // m351_8 = W*in
   wire signed [9:0] m351_8;
   assign m351_8 =10'b0;

   // m351_9 = W*in
   wire signed [9:0] m351_9;
   assign m351_9 =10'b0;

   // m351_10 = W*in
   wire signed [9:0] m351_10;
   assign m351_10 =10'b0;

   // m351_11 = W*in
   wire signed [9:0] m351_11;
   assign m351_11 =10'b0;

   // m351_12 = W*in
   wire signed [9:0] m351_12;
   assign m351_12 =10'b0;

   // m351_13 = W*in
   wire signed [9:0] m351_13;
   assign m351_13 =10'b0;

   // m351_14 = W*in
   wire signed [9:0] m351_14;
   assign m351_14 =10'b0;

   // m351_15 = W*in
   wire signed [9:0] m351_15;
   assign m351_15 =10'b0;

   // m351_16 = W*in
   wire signed [9:0] m351_16;
   assign m351_16 =10'b0;

   // m351_17 = W*in
   wire signed [9:0] m351_17;
   assign m351_17 =10'b0;

   // m351_18 = W*in
   wire signed [9:0] m351_18;
   assign m351_18 =10'b0;

   // m351_19 = W*in
   wire signed [9:0] m351_19;
   assign m351_19 =10'b0;

   // m351_20 = W*in
   wire signed [9:0] m351_20;
   assign m351_20 =10'b0;

   // m351_21 = W*in
   wire signed [9:0] m351_21;
   assign m351_21 =10'b0;

   // m351_22 = W*in
   wire signed [9:0] m351_22;
   assign m351_22 =10'b0;

   // m351_23 = W*in
   wire signed [9:0] m351_23;
   assign m351_23 =10'b0;

   // m351_24 = W*in
   wire signed [9:0] m351_24;
   assign m351_24 =10'b0;

   // m351_25 = W*in
   wire signed [9:0] m351_25;
   assign m351_25 ={ {5{in351[5]}} , in351[5:1] };

   // m351_26 = W*in
   wire signed [9:0] m351_26;
   assign m351_26 ={ {5{in351[5]}} , in351[5:1] };

   // m351_27 = W*in
   wire signed [9:0] m351_27;
   assign m351_27 =10'b0;

   // m351_28 = W*in
   wire signed [9:0] m351_28;
   assign m351_28 ={ {5{in351[5]}} , in351[5:1] };

   // m351_29 = W*in
   wire signed [9:0] m351_29;
   assign m351_29 =10'b0;

   // m351_30 = W*in
   wire signed [9:0] m351_30;
   assign m351_30 =10'b0;

   // m351_31 = W*in
   wire signed [9:0] m351_31;
   assign m351_31 =10'b0;

   // m351_32 = W*in
   wire signed [9:0] m351_32;
   assign m351_32 =10'b0;

   // m351_33 = W*in
   wire signed [9:0] m351_33;
   assign m351_33 =10'b0;

   // m351_34 = W*in
   wire signed [9:0] m351_34;
   assign m351_34 =10'b0;

   // m351_35 = W*in
   wire signed [9:0] m351_35;
   assign m351_35 ={ {5{neg351[5]}} , neg351[5:1] };

   // m351_36 = W*in
   wire signed [9:0] m351_36;
   assign m351_36 =10'b0;

   // m351_37 = W*in
   wire signed [9:0] m351_37;
   assign m351_37 =10'b0;

   // m351_38 = W*in
   wire signed [9:0] m351_38;
   assign m351_38 =10'b0;

   // m351_39 = W*in
   wire signed [9:0] m351_39;
   assign m351_39 =10'b0;

   // m351_40 = W*in
   wire signed [9:0] m351_40;
   assign m351_40 =10'b0;

   // m351_41 = W*in
   wire signed [9:0] m351_41;
   assign m351_41 =10'b0;

   // m351_42 = W*in
   wire signed [9:0] m351_42;
   assign m351_42 =10'b0;

   // m351_43 = W*in
   wire signed [9:0] m351_43;
   assign m351_43 =10'b0;

   // m351_44 = W*in
   wire signed [9:0] m351_44;
   assign m351_44 =10'b0;

   // m351_45 = W*in
   wire signed [9:0] m351_45;
   assign m351_45 =10'b0;

   // m351_46 = W*in
   wire signed [9:0] m351_46;
   assign m351_46 =10'b0;

   // m351_47 = W*in
   wire signed [9:0] m351_47;
   assign m351_47 =10'b0;

   // m351_48 = W*in
   wire signed [9:0] m351_48;
   assign m351_48 =10'b0;

   // m351_49 = W*in
   wire signed [9:0] m351_49;
   assign m351_49 =10'b0;

   // m351_50 = W*in
   wire signed [9:0] m351_50;
   assign m351_50 =10'b0;

   // m351_51 = W*in
   wire signed [9:0] m351_51;
   assign m351_51 =10'b0;

   // m351_52 = W*in
   wire signed [9:0] m351_52;
   assign m351_52 =10'b0;

   // m351_53 = W*in
   wire signed [9:0] m351_53;
   assign m351_53 =10'b0;

   // m351_54 = W*in
   wire signed [9:0] m351_54;
   assign m351_54 =10'b0;

   // m351_55 = W*in
   wire signed [9:0] m351_55;
   assign m351_55 =10'b0;

   // m351_56 = W*in
   wire signed [9:0] m351_56;
   assign m351_56 =10'b0;

   // m351_57 = W*in
   wire signed [9:0] m351_57;
   assign m351_57 =10'b0;

   // m351_58 = W*in
   wire signed [9:0] m351_58;
   assign m351_58 =10'b0;

   // m351_59 = W*in
   wire signed [9:0] m351_59;
   assign m351_59 =10'b0;

   // m351_60 = W*in
   wire signed [9:0] m351_60;
   assign m351_60 =10'b0;

   // m351_61 = W*in
   wire signed [9:0] m351_61;
   assign m351_61 =10'b0;

   // m351_62 = W*in
   wire signed [9:0] m351_62;
   assign m351_62 =10'b0;

   // m351_63 = W*in
   wire signed [9:0] m351_63;
   assign m351_63 =10'b0;

   // m351_64 = W*in
   wire signed [9:0] m351_64;
   assign m351_64 =10'b0;

   // m351_65 = W*in
   wire signed [9:0] m351_65;
   assign m351_65 ={ {5{neg351[5]}} , neg351[5:1] };

   // m351_66 = W*in
   wire signed [9:0] m351_66;
   assign m351_66 ={ {5{neg351[5]}} , neg351[5:1] };

   // m351_67 = W*in
   wire signed [9:0] m351_67;
   assign m351_67 =10'b0;

   // m351_68 = W*in
   wire signed [9:0] m351_68;
   assign m351_68 =10'b0;

   // m351_69 = W*in
   wire signed [9:0] m351_69;
   assign m351_69 ={ {5{neg351[5]}} , neg351[5:1] };

   // m351_70 = W*in
   wire signed [9:0] m351_70;
   assign m351_70 =10'b0;

   // m351_71 = W*in
   wire signed [9:0] m351_71;
   assign m351_71 =10'b0;

   // m351_72 = W*in
   wire signed [9:0] m351_72;
   assign m351_72 =10'b0;

   // m351_73 = W*in
   wire signed [9:0] m351_73;
   assign m351_73 =10'b0;

   // m351_74 = W*in
   wire signed [9:0] m351_74;
   assign m351_74 =10'b0;

   // m351_75 = W*in
   wire signed [9:0] m351_75;
   assign m351_75 =10'b0;

   // m351_76 = W*in
   wire signed [9:0] m351_76;
   assign m351_76 =10'b0;

   // m351_77 = W*in
   wire signed [9:0] m351_77;
   assign m351_77 =10'b0;

   // m351_78 = W*in
   wire signed [9:0] m351_78;
   assign m351_78 =10'b0;

   // m351_79 = W*in
   wire signed [9:0] m351_79;
   assign m351_79 =10'b0;

   // m351_80 = W*in
   wire signed [9:0] m351_80;
   assign m351_80 =10'b0;

   // m351_81 = W*in
   wire signed [9:0] m351_81;
   assign m351_81 =10'b0;

   // m351_82 = W*in
   wire signed [9:0] m351_82;
   assign m351_82 =10'b0;

   // m351_83 = W*in
   wire signed [9:0] m351_83;
   assign m351_83 =10'b0;

   // m351_84 = W*in
   wire signed [9:0] m351_84;
   assign m351_84 ={ {5{in351[5]}} , in351[5:1] };

   // m351_85 = W*in
   wire signed [9:0] m351_85;
   assign m351_85 =10'b0;

   // m351_86 = W*in
   wire signed [9:0] m351_86;
   assign m351_86 =10'b0;

   // m351_87 = W*in
   wire signed [9:0] m351_87;
   assign m351_87 =10'b0;

   // m351_88 = W*in
   wire signed [9:0] m351_88;
   assign m351_88 =10'b0;

   // m351_89 = W*in
   wire signed [9:0] m351_89;
   assign m351_89 =10'b0;

   // m351_90 = W*in
   wire signed [9:0] m351_90;
   assign m351_90 =10'b0;

   // m351_91 = W*in
   wire signed [9:0] m351_91;
   assign m351_91 =10'b0;

   // m351_92 = W*in
   wire signed [9:0] m351_92;
   assign m351_92 =10'b0;

   // m351_93 = W*in
   wire signed [9:0] m351_93;
   assign m351_93 =10'b0;

   // m351_94 = W*in
   wire signed [9:0] m351_94;
   assign m351_94 =10'b0;

   // m351_95 = W*in
   wire signed [9:0] m351_95;
   assign m351_95 =10'b0;

   // m351_96 = W*in
   wire signed [9:0] m351_96;
   assign m351_96 =10'b0;

   // m351_97 = W*in
   wire signed [9:0] m351_97;
   assign m351_97 =10'b0;

   // m351_98 = W*in
   wire signed [9:0] m351_98;
   assign m351_98 =10'b0;

   // m351_99 = W*in
   wire signed [9:0] m351_99;
   assign m351_99 =10'b0;

   // m351_100 = W*in
   wire signed [9:0] m351_100;
   assign m351_100 =10'b0;

   // m351_101 = W*in
   wire signed [9:0] m351_101;
   assign m351_101 =10'b0;

   // m351_102 = W*in
   wire signed [9:0] m351_102;
   assign m351_102 =10'b0;

   // m351_103 = W*in
   wire signed [9:0] m351_103;
   assign m351_103 =10'b0;

   // m351_104 = W*in
   wire signed [9:0] m351_104;
   assign m351_104 =10'b0;

   // m351_105 = W*in
   wire signed [9:0] m351_105;
   assign m351_105 =10'b0;

   // m351_106 = W*in
   wire signed [9:0] m351_106;
   assign m351_106 =10'b0;

   // m351_107 = W*in
   wire signed [9:0] m351_107;
   assign m351_107 =10'b0;

   // m351_108 = W*in
   wire signed [9:0] m351_108;
   assign m351_108 =10'b0;

   // m351_109 = W*in
   wire signed [9:0] m351_109;
   assign m351_109 =10'b0;

   // m351_110 = W*in
   wire signed [9:0] m351_110;
   assign m351_110 =10'b0;

   // m351_111 = W*in
   wire signed [9:0] m351_111;
   assign m351_111 =10'b0;

   // m351_112 = W*in
   wire signed [9:0] m351_112;
   assign m351_112 =10'b0;

   // m351_113 = W*in
   wire signed [9:0] m351_113;
   assign m351_113 =10'b0;

   // m351_114 = W*in
   wire signed [9:0] m351_114;
   assign m351_114 =10'b0;

   // m351_115 = W*in
   wire signed [9:0] m351_115;
   assign m351_115 =10'b0;

   // m351_116 = W*in
   wire signed [9:0] m351_116;
   assign m351_116 =10'b0;

   // m351_117 = W*in
   wire signed [9:0] m351_117;
   assign m351_117 =10'b0;

   // m352_1 = W*in
   wire signed [9:0] m352_1;
   assign m352_1 =10'b0;

   // m352_2 = W*in
   wire signed [9:0] m352_2;
   assign m352_2 =10'b0;

   // m352_3 = W*in
   wire signed [9:0] m352_3;
   assign m352_3 =10'b0;

   // m352_4 = W*in
   wire signed [9:0] m352_4;
   assign m352_4 =10'b0;

   // m352_5 = W*in
   wire signed [9:0] m352_5;
   assign m352_5 =10'b0;

   // m352_6 = W*in
   wire signed [9:0] m352_6;
   assign m352_6 =10'b0;

   // m352_7 = W*in
   wire signed [9:0] m352_7;
   assign m352_7 =10'b0;

   // m352_8 = W*in
   wire signed [9:0] m352_8;
   assign m352_8 =10'b0;

   // m352_9 = W*in
   wire signed [9:0] m352_9;
   assign m352_9 =10'b0;

   // m352_10 = W*in
   wire signed [9:0] m352_10;
   assign m352_10 =10'b0;

   // m352_11 = W*in
   wire signed [9:0] m352_11;
   assign m352_11 =10'b0;

   // m352_12 = W*in
   wire signed [9:0] m352_12;
   assign m352_12 =10'b0;

   // m352_13 = W*in
   wire signed [9:0] m352_13;
   assign m352_13 =10'b0;

   // m352_14 = W*in
   wire signed [9:0] m352_14;
   assign m352_14 =10'b0;

   // m352_15 = W*in
   wire signed [9:0] m352_15;
   assign m352_15 =10'b0;

   // m352_16 = W*in
   wire signed [9:0] m352_16;
   assign m352_16 =10'b0;

   // m352_17 = W*in
   wire signed [9:0] m352_17;
   assign m352_17 =10'b0;

   // m352_18 = W*in
   wire signed [9:0] m352_18;
   assign m352_18 =10'b0;

   // m352_19 = W*in
   wire signed [9:0] m352_19;
   assign m352_19 =10'b0;

   // m352_20 = W*in
   wire signed [9:0] m352_20;
   assign m352_20 ={ {5{in352[5]}} , in352[5:1] };

   // m352_21 = W*in
   wire signed [9:0] m352_21;
   assign m352_21 ={ {5{neg352[5]}} , neg352[5:1] };

   // m352_22 = W*in
   wire signed [9:0] m352_22;
   assign m352_22 =10'b0;

   // m352_23 = W*in
   wire signed [9:0] m352_23;
   assign m352_23 =10'b0;

   // m352_24 = W*in
   wire signed [9:0] m352_24;
   assign m352_24 =10'b0;

   // m352_25 = W*in
   wire signed [9:0] m352_25;
   assign m352_25 =10'b0;

   // m352_26 = W*in
   wire signed [9:0] m352_26;
   assign m352_26 =10'b0;

   // m352_27 = W*in
   wire signed [9:0] m352_27;
   assign m352_27 ={ {5{in352[5]}} , in352[5:1] };

   // m352_28 = W*in
   wire signed [9:0] m352_28;
   assign m352_28 =10'b0;

   // m352_29 = W*in
   wire signed [9:0] m352_29;
   assign m352_29 =10'b0;

   // m352_30 = W*in
   wire signed [9:0] m352_30;
   assign m352_30 =10'b0;

   // m352_31 = W*in
   wire signed [9:0] m352_31;
   assign m352_31 =10'b0;

   // m352_32 = W*in
   wire signed [9:0] m352_32;
   assign m352_32 =10'b0;

   // m352_33 = W*in
   wire signed [9:0] m352_33;
   assign m352_33 =10'b0;

   // m352_34 = W*in
   wire signed [9:0] m352_34;
   assign m352_34 ={ {5{in352[5]}} , in352[5:1] };

   // m352_35 = W*in
   wire signed [9:0] m352_35;
   assign m352_35 ={ {5{in352[5]}} , in352[5:1] };

   // m352_36 = W*in
   wire signed [9:0] m352_36;
   assign m352_36 =10'b0;

   // m352_37 = W*in
   wire signed [9:0] m352_37;
   assign m352_37 =10'b0;

   // m352_38 = W*in
   wire signed [9:0] m352_38;
   assign m352_38 =10'b0;

   // m352_39 = W*in
   wire signed [9:0] m352_39;
   assign m352_39 =10'b0;

   // m352_40 = W*in
   wire signed [9:0] m352_40;
   assign m352_40 =10'b0;

   // m352_41 = W*in
   wire signed [9:0] m352_41;
   assign m352_41 =10'b0;

   // m352_42 = W*in
   wire signed [9:0] m352_42;
   assign m352_42 =10'b0;

   // m352_43 = W*in
   wire signed [9:0] m352_43;
   assign m352_43 =10'b0;

   // m352_44 = W*in
   wire signed [9:0] m352_44;
   assign m352_44 =10'b0;

   // m352_45 = W*in
   wire signed [9:0] m352_45;
   assign m352_45 =10'b0;

   // m352_46 = W*in
   wire signed [9:0] m352_46;
   assign m352_46 =10'b0;

   // m352_47 = W*in
   wire signed [9:0] m352_47;
   assign m352_47 =10'b0;

   // m352_48 = W*in
   wire signed [9:0] m352_48;
   assign m352_48 =10'b0;

   // m352_49 = W*in
   wire signed [9:0] m352_49;
   assign m352_49 =10'b0;

   // m352_50 = W*in
   wire signed [9:0] m352_50;
   assign m352_50 =10'b0;

   // m352_51 = W*in
   wire signed [9:0] m352_51;
   assign m352_51 =10'b0;

   // m352_52 = W*in
   wire signed [9:0] m352_52;
   assign m352_52 =10'b0;

   // m352_53 = W*in
   wire signed [9:0] m352_53;
   assign m352_53 =10'b0;

   // m352_54 = W*in
   wire signed [9:0] m352_54;
   assign m352_54 =10'b0;

   // m352_55 = W*in
   wire signed [9:0] m352_55;
   assign m352_55 =10'b0;

   // m352_56 = W*in
   wire signed [9:0] m352_56;
   assign m352_56 =10'b0;

   // m352_57 = W*in
   wire signed [9:0] m352_57;
   assign m352_57 =10'b0;

   // m352_58 = W*in
   wire signed [9:0] m352_58;
   assign m352_58 =10'b0;

   // m352_59 = W*in
   wire signed [9:0] m352_59;
   assign m352_59 =10'b0;

   // m352_60 = W*in
   wire signed [9:0] m352_60;
   assign m352_60 =10'b0;

   // m352_61 = W*in
   wire signed [9:0] m352_61;
   assign m352_61 =10'b0;

   // m352_62 = W*in
   wire signed [9:0] m352_62;
   assign m352_62 =10'b0;

   // m352_63 = W*in
   wire signed [9:0] m352_63;
   assign m352_63 =10'b0;

   // m352_64 = W*in
   wire signed [9:0] m352_64;
   assign m352_64 ={ {5{in352[5]}} , in352[5:1] };

   // m352_65 = W*in
   wire signed [9:0] m352_65;
   assign m352_65 =10'b0;

   // m352_66 = W*in
   wire signed [9:0] m352_66;
   assign m352_66 =10'b0;

   // m352_67 = W*in
   wire signed [9:0] m352_67;
   assign m352_67 =10'b0;

   // m352_68 = W*in
   wire signed [9:0] m352_68;
   assign m352_68 =10'b0;

   // m352_69 = W*in
   wire signed [9:0] m352_69;
   assign m352_69 =10'b0;

   // m352_70 = W*in
   wire signed [9:0] m352_70;
   assign m352_70 =10'b0;

   // m352_71 = W*in
   wire signed [9:0] m352_71;
   assign m352_71 =10'b0;

   // m352_72 = W*in
   wire signed [9:0] m352_72;
   assign m352_72 =10'b0;

   // m352_73 = W*in
   wire signed [9:0] m352_73;
   assign m352_73 =10'b0;

   // m352_74 = W*in
   wire signed [9:0] m352_74;
   assign m352_74 =10'b0;

   // m352_75 = W*in
   wire signed [9:0] m352_75;
   assign m352_75 =10'b0;

   // m352_76 = W*in
   wire signed [9:0] m352_76;
   assign m352_76 =10'b0;

   // m352_77 = W*in
   wire signed [9:0] m352_77;
   assign m352_77 =10'b0;

   // m352_78 = W*in
   wire signed [9:0] m352_78;
   assign m352_78 =10'b0;

   // m352_79 = W*in
   wire signed [9:0] m352_79;
   assign m352_79 =10'b0;

   // m352_80 = W*in
   wire signed [9:0] m352_80;
   assign m352_80 =10'b0;

   // m352_81 = W*in
   wire signed [9:0] m352_81;
   assign m352_81 ={ {5{in352[5]}} , in352[5:1] };

   // m352_82 = W*in
   wire signed [9:0] m352_82;
   assign m352_82 =10'b0;

   // m352_83 = W*in
   wire signed [9:0] m352_83;
   assign m352_83 =10'b0;

   // m352_84 = W*in
   wire signed [9:0] m352_84;
   assign m352_84 =10'b0;

   // m352_85 = W*in
   wire signed [9:0] m352_85;
   assign m352_85 =10'b0;

   // m352_86 = W*in
   wire signed [9:0] m352_86;
   assign m352_86 =10'b0;

   // m352_87 = W*in
   wire signed [9:0] m352_87;
   assign m352_87 =10'b0;

   // m352_88 = W*in
   wire signed [9:0] m352_88;
   assign m352_88 =10'b0;

   // m352_89 = W*in
   wire signed [9:0] m352_89;
   assign m352_89 =10'b0;

   // m352_90 = W*in
   wire signed [9:0] m352_90;
   assign m352_90 =10'b0;

   // m352_91 = W*in
   wire signed [9:0] m352_91;
   assign m352_91 =10'b0;

   // m352_92 = W*in
   wire signed [9:0] m352_92;
   assign m352_92 =10'b0;

   // m352_93 = W*in
   wire signed [9:0] m352_93;
   assign m352_93 =10'b0;

   // m352_94 = W*in
   wire signed [9:0] m352_94;
   assign m352_94 =10'b0;

   // m352_95 = W*in
   wire signed [9:0] m352_95;
   assign m352_95 =10'b0;

   // m352_96 = W*in
   wire signed [9:0] m352_96;
   assign m352_96 =10'b0;

   // m352_97 = W*in
   wire signed [9:0] m352_97;
   assign m352_97 =10'b0;

   // m352_98 = W*in
   wire signed [9:0] m352_98;
   assign m352_98 =10'b0;

   // m352_99 = W*in
   wire signed [9:0] m352_99;
   assign m352_99 =10'b0;

   // m352_100 = W*in
   wire signed [9:0] m352_100;
   assign m352_100 =10'b0;

   // m352_101 = W*in
   wire signed [9:0] m352_101;
   assign m352_101 =10'b0;

   // m352_102 = W*in
   wire signed [9:0] m352_102;
   assign m352_102 =10'b0;

   // m352_103 = W*in
   wire signed [9:0] m352_103;
   assign m352_103 =10'b0;

   // m352_104 = W*in
   wire signed [9:0] m352_104;
   assign m352_104 =10'b0;

   // m352_105 = W*in
   wire signed [9:0] m352_105;
   assign m352_105 =10'b0;

   // m352_106 = W*in
   wire signed [9:0] m352_106;
   assign m352_106 =10'b0;

   // m352_107 = W*in
   wire signed [9:0] m352_107;
   assign m352_107 =10'b0;

   // m352_108 = W*in
   wire signed [9:0] m352_108;
   assign m352_108 =10'b0;

   // m352_109 = W*in
   wire signed [9:0] m352_109;
   assign m352_109 =10'b0;

   // m352_110 = W*in
   wire signed [9:0] m352_110;
   assign m352_110 =10'b0;

   // m352_111 = W*in
   wire signed [9:0] m352_111;
   assign m352_111 =10'b0;

   // m352_112 = W*in
   wire signed [9:0] m352_112;
   assign m352_112 =10'b0;

   // m352_113 = W*in
   wire signed [9:0] m352_113;
   assign m352_113 =10'b0;

   // m352_114 = W*in
   wire signed [9:0] m352_114;
   assign m352_114 =10'b0;

   // m352_115 = W*in
   wire signed [9:0] m352_115;
   assign m352_115 =10'b0;

   // m352_116 = W*in
   wire signed [9:0] m352_116;
   assign m352_116 =10'b0;

   // m352_117 = W*in
   wire signed [9:0] m352_117;
   assign m352_117 =10'b0;

   // m353_1 = W*in
   wire signed [9:0] m353_1;
   assign m353_1 =10'b0;

   // m353_2 = W*in
   wire signed [9:0] m353_2;
   assign m353_2 =10'b0;

   // m353_3 = W*in
   wire signed [9:0] m353_3;
   assign m353_3 =10'b0;

   // m353_4 = W*in
   wire signed [9:0] m353_4;
   assign m353_4 =10'b0;

   // m353_5 = W*in
   wire signed [9:0] m353_5;
   assign m353_5 =10'b0;

   // m353_6 = W*in
   wire signed [9:0] m353_6;
   assign m353_6 =10'b0;

   // m353_7 = W*in
   wire signed [9:0] m353_7;
   assign m353_7 =10'b0;

   // m353_8 = W*in
   wire signed [9:0] m353_8;
   assign m353_8 =10'b0;

   // m353_9 = W*in
   wire signed [9:0] m353_9;
   assign m353_9 =10'b0;

   // m353_10 = W*in
   wire signed [9:0] m353_10;
   assign m353_10 =10'b0;

   // m353_11 = W*in
   wire signed [9:0] m353_11;
   assign m353_11 =10'b0;

   // m353_12 = W*in
   wire signed [9:0] m353_12;
   assign m353_12 =10'b0;

   // m353_13 = W*in
   wire signed [9:0] m353_13;
   assign m353_13 =10'b0;

   // m353_14 = W*in
   wire signed [9:0] m353_14;
   assign m353_14 =10'b0;

   // m353_15 = W*in
   wire signed [9:0] m353_15;
   assign m353_15 ={ {4{neg353[5]}} , neg353[5:0] };

   // m353_16 = W*in
   wire signed [9:0] m353_16;
   assign m353_16 ={ {5{in353[5]}} , in353[5:1] };

   // m353_17 = W*in
   wire signed [9:0] m353_17;
   assign m353_17 ={ {5{in353[5]}} , in353[5:1] };

   // m353_18 = W*in
   wire signed [9:0] m353_18;
   assign m353_18 ={ {5{in353[5]}} , in353[5:1] };

   // m353_19 = W*in
   wire signed [9:0] m353_19;
   assign m353_19 =10'b0;

   // m353_20 = W*in
   wire signed [9:0] m353_20;
   assign m353_20 =10'b0;

   // m353_21 = W*in
   wire signed [9:0] m353_21;
   assign m353_21 =10'b0;

   // m353_22 = W*in
   wire signed [9:0] m353_22;
   assign m353_22 =10'b0;

   // m353_23 = W*in
   wire signed [9:0] m353_23;
   assign m353_23 =10'b0;

   // m353_24 = W*in
   wire signed [9:0] m353_24;
   assign m353_24 =10'b0;

   // m353_25 = W*in
   wire signed [9:0] m353_25;
   assign m353_25 =10'b0;

   // m353_26 = W*in
   wire signed [9:0] m353_26;
   assign m353_26 =10'b0;

   // m353_27 = W*in
   wire signed [9:0] m353_27;
   assign m353_27 =10'b0;

   // m353_28 = W*in
   wire signed [9:0] m353_28;
   assign m353_28 ={ {5{in353[5]}} , in353[5:1] };

   // m353_29 = W*in
   wire signed [9:0] m353_29;
   assign m353_29 =10'b0;

   // m353_30 = W*in
   wire signed [9:0] m353_30;
   assign m353_30 =10'b0;

   // m353_31 = W*in
   wire signed [9:0] m353_31;
   assign m353_31 =10'b0;

   // m353_32 = W*in
   wire signed [9:0] m353_32;
   assign m353_32 =10'b0;

   // m353_33 = W*in
   wire signed [9:0] m353_33;
   assign m353_33 =10'b0;

   // m353_34 = W*in
   wire signed [9:0] m353_34;
   assign m353_34 =10'b0;

   // m353_35 = W*in
   wire signed [9:0] m353_35;
   assign m353_35 =10'b0;

   // m353_36 = W*in
   wire signed [9:0] m353_36;
   assign m353_36 =10'b0;

   // m353_37 = W*in
   wire signed [9:0] m353_37;
   assign m353_37 =10'b0;

   // m353_38 = W*in
   wire signed [9:0] m353_38;
   assign m353_38 =10'b0;

   // m353_39 = W*in
   wire signed [9:0] m353_39;
   assign m353_39 =10'b0;

   // m353_40 = W*in
   wire signed [9:0] m353_40;
   assign m353_40 =10'b0;

   // m353_41 = W*in
   wire signed [9:0] m353_41;
   assign m353_41 =10'b0;

   // m353_42 = W*in
   wire signed [9:0] m353_42;
   assign m353_42 =10'b0;

   // m353_43 = W*in
   wire signed [9:0] m353_43;
   assign m353_43 =10'b0;

   // m353_44 = W*in
   wire signed [9:0] m353_44;
   assign m353_44 =10'b0;

   // m353_45 = W*in
   wire signed [9:0] m353_45;
   assign m353_45 =10'b0;

   // m353_46 = W*in
   wire signed [9:0] m353_46;
   assign m353_46 =10'b0;

   // m353_47 = W*in
   wire signed [9:0] m353_47;
   assign m353_47 =10'b0;

   // m353_48 = W*in
   wire signed [9:0] m353_48;
   assign m353_48 =10'b0;

   // m353_49 = W*in
   wire signed [9:0] m353_49;
   assign m353_49 =10'b0;

   // m353_50 = W*in
   wire signed [9:0] m353_50;
   assign m353_50 =10'b0;

   // m353_51 = W*in
   wire signed [9:0] m353_51;
   assign m353_51 =10'b0;

   // m353_52 = W*in
   wire signed [9:0] m353_52;
   assign m353_52 =10'b0;

   // m353_53 = W*in
   wire signed [9:0] m353_53;
   assign m353_53 =10'b0;

   // m353_54 = W*in
   wire signed [9:0] m353_54;
   assign m353_54 =10'b0;

   // m353_55 = W*in
   wire signed [9:0] m353_55;
   assign m353_55 =10'b0;

   // m353_56 = W*in
   wire signed [9:0] m353_56;
   assign m353_56 =10'b0;

   // m353_57 = W*in
   wire signed [9:0] m353_57;
   assign m353_57 =10'b0;

   // m353_58 = W*in
   wire signed [9:0] m353_58;
   assign m353_58 =10'b0;

   // m353_59 = W*in
   wire signed [9:0] m353_59;
   assign m353_59 =10'b0;

   // m353_60 = W*in
   wire signed [9:0] m353_60;
   assign m353_60 =10'b0;

   // m353_61 = W*in
   wire signed [9:0] m353_61;
   assign m353_61 =10'b0;

   // m353_62 = W*in
   wire signed [9:0] m353_62;
   assign m353_62 =10'b0;

   // m353_63 = W*in
   wire signed [9:0] m353_63;
   assign m353_63 ={ {4{neg353[5]}} , neg353[5:0] };

   // m353_64 = W*in
   wire signed [9:0] m353_64;
   assign m353_64 =10'b0;

   // m353_65 = W*in
   wire signed [9:0] m353_65;
   assign m353_65 =10'b0;

   // m353_66 = W*in
   wire signed [9:0] m353_66;
   assign m353_66 =10'b0;

   // m353_67 = W*in
   wire signed [9:0] m353_67;
   assign m353_67 =10'b0;

   // m353_68 = W*in
   wire signed [9:0] m353_68;
   assign m353_68 =10'b0;

   // m353_69 = W*in
   wire signed [9:0] m353_69;
   assign m353_69 ={ {4{neg353[5]}} , neg353[5:0] };

   // m353_70 = W*in
   wire signed [9:0] m353_70;
   assign m353_70 ={ {4{neg353[5]}} , neg353[5:0] };

   // m353_71 = W*in
   wire signed [9:0] m353_71;
   assign m353_71 ={ {5{in353[5]}} , in353[5:1] };

   // m353_72 = W*in
   wire signed [9:0] m353_72;
   assign m353_72 =10'b0;

   // m353_73 = W*in
   wire signed [9:0] m353_73;
   assign m353_73 =10'b0;

   // m353_74 = W*in
   wire signed [9:0] m353_74;
   assign m353_74 =10'b0;

   // m353_75 = W*in
   wire signed [9:0] m353_75;
   assign m353_75 =10'b0;

   // m353_76 = W*in
   wire signed [9:0] m353_76;
   assign m353_76 =10'b0;

   // m353_77 = W*in
   wire signed [9:0] m353_77;
   assign m353_77 =10'b0;

   // m353_78 = W*in
   wire signed [9:0] m353_78;
   assign m353_78 =10'b0;

   // m353_79 = W*in
   wire signed [9:0] m353_79;
   assign m353_79 =10'b0;

   // m353_80 = W*in
   wire signed [9:0] m353_80;
   assign m353_80 =10'b0;

   // m353_81 = W*in
   wire signed [9:0] m353_81;
   assign m353_81 =10'b0;

   // m353_82 = W*in
   wire signed [9:0] m353_82;
   assign m353_82 ={ {4{neg353[5]}} , neg353[5:0] };

   // m353_83 = W*in
   wire signed [9:0] m353_83;
   assign m353_83 ={ {5{neg353[5]}} , neg353[5:1] };

   // m353_84 = W*in
   wire signed [9:0] m353_84;
   assign m353_84 =10'b0;

   // m353_85 = W*in
   wire signed [9:0] m353_85;
   assign m353_85 =10'b0;

   // m353_86 = W*in
   wire signed [9:0] m353_86;
   assign m353_86 =10'b0;

   // m353_87 = W*in
   wire signed [9:0] m353_87;
   assign m353_87 =10'b0;

   // m353_88 = W*in
   wire signed [9:0] m353_88;
   assign m353_88 =10'b0;

   // m353_89 = W*in
   wire signed [9:0] m353_89;
   assign m353_89 ={ {4{neg353[5]}} , neg353[5:0] };

   // m353_90 = W*in
   wire signed [9:0] m353_90;
   assign m353_90 =10'b0;

   // m353_91 = W*in
   wire signed [9:0] m353_91;
   assign m353_91 =10'b0;

   // m353_92 = W*in
   wire signed [9:0] m353_92;
   assign m353_92 =10'b0;

   // m353_93 = W*in
   wire signed [9:0] m353_93;
   assign m353_93 =10'b0;

   // m353_94 = W*in
   wire signed [9:0] m353_94;
   assign m353_94 =10'b0;

   // m353_95 = W*in
   wire signed [9:0] m353_95;
   assign m353_95 =10'b0;

   // m353_96 = W*in
   wire signed [9:0] m353_96;
   assign m353_96 =10'b0;

   // m353_97 = W*in
   wire signed [9:0] m353_97;
   assign m353_97 ={ {5{in353[5]}} , in353[5:1] };

   // m353_98 = W*in
   wire signed [9:0] m353_98;
   assign m353_98 =10'b0;

   // m353_99 = W*in
   wire signed [9:0] m353_99;
   assign m353_99 =10'b0;

   // m353_100 = W*in
   wire signed [9:0] m353_100;
   assign m353_100 =10'b0;

   // m353_101 = W*in
   wire signed [9:0] m353_101;
   assign m353_101 =10'b0;

   // m353_102 = W*in
   wire signed [9:0] m353_102;
   assign m353_102 =10'b0;

   // m353_103 = W*in
   wire signed [9:0] m353_103;
   assign m353_103 =10'b0;

   // m353_104 = W*in
   wire signed [9:0] m353_104;
   assign m353_104 =10'b0;

   // m353_105 = W*in
   wire signed [9:0] m353_105;
   assign m353_105 =10'b0;

   // m353_106 = W*in
   wire signed [9:0] m353_106;
   assign m353_106 =10'b0;

   // m353_107 = W*in
   wire signed [9:0] m353_107;
   assign m353_107 =10'b0;

   // m353_108 = W*in
   wire signed [9:0] m353_108;
   assign m353_108 =10'b0;

   // m353_109 = W*in
   wire signed [9:0] m353_109;
   assign m353_109 =10'b0;

   // m353_110 = W*in
   wire signed [9:0] m353_110;
   assign m353_110 =10'b0;

   // m353_111 = W*in
   wire signed [9:0] m353_111;
   assign m353_111 =10'b0;

   // m353_112 = W*in
   wire signed [9:0] m353_112;
   assign m353_112 =10'b0;

   // m353_113 = W*in
   wire signed [9:0] m353_113;
   assign m353_113 =10'b0;

   // m353_114 = W*in
   wire signed [9:0] m353_114;
   assign m353_114 =10'b0;

   // m353_115 = W*in
   wire signed [9:0] m353_115;
   assign m353_115 =10'b0;

   // m353_116 = W*in
   wire signed [9:0] m353_116;
   assign m353_116 =10'b0;

   // m353_117 = W*in
   wire signed [9:0] m353_117;
   assign m353_117 =10'b0;

   // m354_1 = W*in
   wire signed [9:0] m354_1;
   assign m354_1 =10'b0;

   // m354_2 = W*in
   wire signed [9:0] m354_2;
   assign m354_2 =10'b0;

   // m354_3 = W*in
   wire signed [9:0] m354_3;
   assign m354_3 =10'b0;

   // m354_4 = W*in
   wire signed [9:0] m354_4;
   assign m354_4 =10'b0;

   // m354_5 = W*in
   wire signed [9:0] m354_5;
   assign m354_5 =10'b0;

   // m354_6 = W*in
   wire signed [9:0] m354_6;
   assign m354_6 =10'b0;

   // m354_7 = W*in
   wire signed [9:0] m354_7;
   assign m354_7 =10'b0;

   // m354_8 = W*in
   wire signed [9:0] m354_8;
   assign m354_8 ={ {4{in354[5]}} , in354[5:0] };

   // m354_9 = W*in
   wire signed [9:0] m354_9;
   assign m354_9 =10'b0;

   // m354_10 = W*in
   wire signed [9:0] m354_10;
   assign m354_10 =10'b0;

   // m354_11 = W*in
   wire signed [9:0] m354_11;
   assign m354_11 =10'b0;

   // m354_12 = W*in
   wire signed [9:0] m354_12;
   assign m354_12 =10'b0;

   // m354_13 = W*in
   wire signed [9:0] m354_13;
   assign m354_13 =10'b0;

   // m354_14 = W*in
   wire signed [9:0] m354_14;
   assign m354_14 =10'b0;

   // m354_15 = W*in
   wire signed [9:0] m354_15;
   assign m354_15 =10'b0;

   // m354_16 = W*in
   wire signed [9:0] m354_16;
   assign m354_16 ={ {5{neg354[5]}} , neg354[5:1] };

   // m354_17 = W*in
   wire signed [9:0] m354_17;
   assign m354_17 =10'b0;

   // m354_18 = W*in
   wire signed [9:0] m354_18;
   assign m354_18 ={ {4{in354[5]}} , in354[5:0] };

   // m354_19 = W*in
   wire signed [9:0] m354_19;
   assign m354_19 =10'b0;

   // m354_20 = W*in
   wire signed [9:0] m354_20;
   assign m354_20 =10'b0;

   // m354_21 = W*in
   wire signed [9:0] m354_21;
   assign m354_21 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_22 = W*in
   wire signed [9:0] m354_22;
   assign m354_22 ={ {4{in354[5]}} , in354[5:0] };

   // m354_23 = W*in
   wire signed [9:0] m354_23;
   assign m354_23 =10'b0;

   // m354_24 = W*in
   wire signed [9:0] m354_24;
   assign m354_24 =10'b0;

   // m354_25 = W*in
   wire signed [9:0] m354_25;
   assign m354_25 =10'b0;

   // m354_26 = W*in
   wire signed [9:0] m354_26;
   assign m354_26 ={ {5{in354[5]}} , in354[5:1] };

   // m354_27 = W*in
   wire signed [9:0] m354_27;
   assign m354_27 ={ {5{neg354[5]}} , neg354[5:1] };

   // m354_28 = W*in
   wire signed [9:0] m354_28;
   assign m354_28 ={ {5{neg354[5]}} , neg354[5:1] };

   // m354_29 = W*in
   wire signed [9:0] m354_29;
   assign m354_29 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_30 = W*in
   wire signed [9:0] m354_30;
   assign m354_30 =10'b0;

   // m354_31 = W*in
   wire signed [9:0] m354_31;
   assign m354_31 =10'b0;

   // m354_32 = W*in
   wire signed [9:0] m354_32;
   assign m354_32 =10'b0;

   // m354_33 = W*in
   wire signed [9:0] m354_33;
   assign m354_33 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_34 = W*in
   wire signed [9:0] m354_34;
   assign m354_34 =10'b0;

   // m354_35 = W*in
   wire signed [9:0] m354_35;
   assign m354_35 =10'b0;

   // m354_36 = W*in
   wire signed [9:0] m354_36;
   assign m354_36 =10'b0;

   // m354_37 = W*in
   wire signed [9:0] m354_37;
   assign m354_37 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_38 = W*in
   wire signed [9:0] m354_38;
   assign m354_38 =10'b0;

   // m354_39 = W*in
   wire signed [9:0] m354_39;
   assign m354_39 =10'b0;

   // m354_40 = W*in
   wire signed [9:0] m354_40;
   assign m354_40 =10'b0;

   // m354_41 = W*in
   wire signed [9:0] m354_41;
   assign m354_41 =10'b0;

   // m354_42 = W*in
   wire signed [9:0] m354_42;
   assign m354_42 =10'b0;

   // m354_43 = W*in
   wire signed [9:0] m354_43;
   assign m354_43 =10'b0;

   // m354_44 = W*in
   wire signed [9:0] m354_44;
   assign m354_44 =10'b0;

   // m354_45 = W*in
   wire signed [9:0] m354_45;
   assign m354_45 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_46 = W*in
   wire signed [9:0] m354_46;
   assign m354_46 =10'b0;

   // m354_47 = W*in
   wire signed [9:0] m354_47;
   assign m354_47 =10'b0;

   // m354_48 = W*in
   wire signed [9:0] m354_48;
   assign m354_48 =10'b0;

   // m354_49 = W*in
   wire signed [9:0] m354_49;
   assign m354_49 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_50 = W*in
   wire signed [9:0] m354_50;
   assign m354_50 =10'b0;

   // m354_51 = W*in
   wire signed [9:0] m354_51;
   assign m354_51 ={ {4{in354[5]}} , in354[5:0] };

   // m354_52 = W*in
   wire signed [9:0] m354_52;
   assign m354_52 =10'b0;

   // m354_53 = W*in
   wire signed [9:0] m354_53;
   assign m354_53 ={ {4{in354[5]}} , in354[5:0] };

   // m354_54 = W*in
   wire signed [9:0] m354_54;
   assign m354_54 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_55 = W*in
   wire signed [9:0] m354_55;
   assign m354_55 =10'b0;

   // m354_56 = W*in
   wire signed [9:0] m354_56;
   assign m354_56 =10'b0;

   // m354_57 = W*in
   wire signed [9:0] m354_57;
   assign m354_57 =10'b0;

   // m354_58 = W*in
   wire signed [9:0] m354_58;
   assign m354_58 =10'b0;

   // m354_59 = W*in
   wire signed [9:0] m354_59;
   assign m354_59 =10'b0;

   // m354_60 = W*in
   wire signed [9:0] m354_60;
   assign m354_60 =10'b0;

   // m354_61 = W*in
   wire signed [9:0] m354_61;
   assign m354_61 =10'b0;

   // m354_62 = W*in
   wire signed [9:0] m354_62;
   assign m354_62 =10'b0;

   // m354_63 = W*in
   wire signed [9:0] m354_63;
   assign m354_63 ={ {5{neg354[5]}} , neg354[5:1] };

   // m354_64 = W*in
   wire signed [9:0] m354_64;
   assign m354_64 ={ {4{in354[5]}} , in354[5:0] };

   // m354_65 = W*in
   wire signed [9:0] m354_65;
   assign m354_65 =10'b0;

   // m354_66 = W*in
   wire signed [9:0] m354_66;
   assign m354_66 =10'b0;

   // m354_67 = W*in
   wire signed [9:0] m354_67;
   assign m354_67 =10'b0;

   // m354_68 = W*in
   wire signed [9:0] m354_68;
   assign m354_68 ={ {4{in354[5]}} , in354[5:0] };

   // m354_69 = W*in
   wire signed [9:0] m354_69;
   assign m354_69 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_70 = W*in
   wire signed [9:0] m354_70;
   assign m354_70 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_71 = W*in
   wire signed [9:0] m354_71;
   assign m354_71 =10'b0;

   // m354_72 = W*in
   wire signed [9:0] m354_72;
   assign m354_72 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_73 = W*in
   wire signed [9:0] m354_73;
   assign m354_73 ={ {4{in354[5]}} , in354[5:0] };

   // m354_74 = W*in
   wire signed [9:0] m354_74;
   assign m354_74 ={ {4{in354[5]}} , in354[5:0] };

   // m354_75 = W*in
   wire signed [9:0] m354_75;
   assign m354_75 =10'b0;

   // m354_76 = W*in
   wire signed [9:0] m354_76;
   assign m354_76 =10'b0;

   // m354_77 = W*in
   wire signed [9:0] m354_77;
   assign m354_77 =10'b0;

   // m354_78 = W*in
   wire signed [9:0] m354_78;
   assign m354_78 =10'b0;

   // m354_79 = W*in
   wire signed [9:0] m354_79;
   assign m354_79 =10'b0;

   // m354_80 = W*in
   wire signed [9:0] m354_80;
   assign m354_80 =10'b0;

   // m354_81 = W*in
   wire signed [9:0] m354_81;
   assign m354_81 ={ {4{in354[5]}} , in354[5:0] };

   // m354_82 = W*in
   wire signed [9:0] m354_82;
   assign m354_82 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_83 = W*in
   wire signed [9:0] m354_83;
   assign m354_83 =10'b0;

   // m354_84 = W*in
   wire signed [9:0] m354_84;
   assign m354_84 ={ {5{neg354[5]}} , neg354[5:1] };

   // m354_85 = W*in
   wire signed [9:0] m354_85;
   assign m354_85 ={ {5{neg354[5]}} , neg354[5:1] };

   // m354_86 = W*in
   wire signed [9:0] m354_86;
   assign m354_86 =10'b0;

   // m354_87 = W*in
   wire signed [9:0] m354_87;
   assign m354_87 =10'b0;

   // m354_88 = W*in
   wire signed [9:0] m354_88;
   assign m354_88 =10'b0;

   // m354_89 = W*in
   wire signed [9:0] m354_89;
   assign m354_89 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_90 = W*in
   wire signed [9:0] m354_90;
   assign m354_90 =10'b0;

   // m354_91 = W*in
   wire signed [9:0] m354_91;
   assign m354_91 =10'b0;

   // m354_92 = W*in
   wire signed [9:0] m354_92;
   assign m354_92 =10'b0;

   // m354_93 = W*in
   wire signed [9:0] m354_93;
   assign m354_93 ={ {4{neg354[5]}} , neg354[5:0] };

   // m354_94 = W*in
   wire signed [9:0] m354_94;
   assign m354_94 =10'b0;

   // m354_95 = W*in
   wire signed [9:0] m354_95;
   assign m354_95 =10'b0;

   // m354_96 = W*in
   wire signed [9:0] m354_96;
   assign m354_96 =10'b0;

   // m354_97 = W*in
   wire signed [9:0] m354_97;
   assign m354_97 =10'b0;

   // m354_98 = W*in
   wire signed [9:0] m354_98;
   assign m354_98 =10'b0;

   // m354_99 = W*in
   wire signed [9:0] m354_99;
   assign m354_99 =10'b0;

   // m354_100 = W*in
   wire signed [9:0] m354_100;
   assign m354_100 =10'b0;

   // m354_101 = W*in
   wire signed [9:0] m354_101;
   assign m354_101 =10'b0;

   // m354_102 = W*in
   wire signed [9:0] m354_102;
   assign m354_102 =10'b0;

   // m354_103 = W*in
   wire signed [9:0] m354_103;
   assign m354_103 =10'b0;

   // m354_104 = W*in
   wire signed [9:0] m354_104;
   assign m354_104 =10'b0;

   // m354_105 = W*in
   wire signed [9:0] m354_105;
   assign m354_105 =10'b0;

   // m354_106 = W*in
   wire signed [9:0] m354_106;
   assign m354_106 =10'b0;

   // m354_107 = W*in
   wire signed [9:0] m354_107;
   assign m354_107 =10'b0;

   // m354_108 = W*in
   wire signed [9:0] m354_108;
   assign m354_108 =10'b0;

   // m354_109 = W*in
   wire signed [9:0] m354_109;
   assign m354_109 =10'b0;

   // m354_110 = W*in
   wire signed [9:0] m354_110;
   assign m354_110 =10'b0;

   // m354_111 = W*in
   wire signed [9:0] m354_111;
   assign m354_111 =10'b0;

   // m354_112 = W*in
   wire signed [9:0] m354_112;
   assign m354_112 =10'b0;

   // m354_113 = W*in
   wire signed [9:0] m354_113;
   assign m354_113 ={ {4{in354[5]}} , in354[5:0] };

   // m354_114 = W*in
   wire signed [9:0] m354_114;
   assign m354_114 =10'b0;

   // m354_115 = W*in
   wire signed [9:0] m354_115;
   assign m354_115 ={ {5{in354[5]}} , in354[5:1] };

   // m354_116 = W*in
   wire signed [9:0] m354_116;
   assign m354_116 =10'b0;

   // m354_117 = W*in
   wire signed [9:0] m354_117;
   assign m354_117 =10'b0;

   // m355_1 = W*in
   wire signed [9:0] m355_1;
   assign m355_1 =10'b0;

   // m355_2 = W*in
   wire signed [9:0] m355_2;
   assign m355_2 =10'b0;

   // m355_3 = W*in
   wire signed [9:0] m355_3;
   assign m355_3 =10'b0;

   // m355_4 = W*in
   wire signed [9:0] m355_4;
   assign m355_4 =10'b0;

   // m355_5 = W*in
   wire signed [9:0] m355_5;
   assign m355_5 =10'b0;

   // m355_6 = W*in
   wire signed [9:0] m355_6;
   assign m355_6 =10'b0;

   // m355_7 = W*in
   wire signed [9:0] m355_7;
   assign m355_7 =10'b0;

   // m355_8 = W*in
   wire signed [9:0] m355_8;
   assign m355_8 =10'b0;

   // m355_9 = W*in
   wire signed [9:0] m355_9;
   assign m355_9 =10'b0;

   // m355_10 = W*in
   wire signed [9:0] m355_10;
   assign m355_10 =10'b0;

   // m355_11 = W*in
   wire signed [9:0] m355_11;
   assign m355_11 =10'b0;

   // m355_12 = W*in
   wire signed [9:0] m355_12;
   assign m355_12 =10'b0;

   // m355_13 = W*in
   wire signed [9:0] m355_13;
   assign m355_13 =10'b0;

   // m355_14 = W*in
   wire signed [9:0] m355_14;
   assign m355_14 =10'b0;

   // m355_15 = W*in
   wire signed [9:0] m355_15;
   assign m355_15 =10'b0;

   // m355_16 = W*in
   wire signed [9:0] m355_16;
   assign m355_16 =10'b0;

   // m355_17 = W*in
   wire signed [9:0] m355_17;
   assign m355_17 ={ {5{neg355[5]}} , neg355[5:1] };

   // m355_18 = W*in
   wire signed [9:0] m355_18;
   assign m355_18 =10'b0;

   // m355_19 = W*in
   wire signed [9:0] m355_19;
   assign m355_19 ={ {5{neg355[5]}} , neg355[5:1] };

   // m355_20 = W*in
   wire signed [9:0] m355_20;
   assign m355_20 =10'b0;

   // m355_21 = W*in
   wire signed [9:0] m355_21;
   assign m355_21 =10'b0;

   // m355_22 = W*in
   wire signed [9:0] m355_22;
   assign m355_22 =10'b0;

   // m355_23 = W*in
   wire signed [9:0] m355_23;
   assign m355_23 =10'b0;

   // m355_24 = W*in
   wire signed [9:0] m355_24;
   assign m355_24 =10'b0;

   // m355_25 = W*in
   wire signed [9:0] m355_25;
   assign m355_25 =10'b0;

   // m355_26 = W*in
   wire signed [9:0] m355_26;
   assign m355_26 =10'b0;

   // m355_27 = W*in
   wire signed [9:0] m355_27;
   assign m355_27 ={ {5{neg355[5]}} , neg355[5:1] };

   // m355_28 = W*in
   wire signed [9:0] m355_28;
   assign m355_28 ={ {4{neg355[5]}} , neg355[5:0] };

   // m355_29 = W*in
   wire signed [9:0] m355_29;
   assign m355_29 ={ {4{neg355[5]}} , neg355[5:0] };

   // m355_30 = W*in
   wire signed [9:0] m355_30;
   assign m355_30 =10'b0;

   // m355_31 = W*in
   wire signed [9:0] m355_31;
   assign m355_31 =10'b0;

   // m355_32 = W*in
   wire signed [9:0] m355_32;
   assign m355_32 =10'b0;

   // m355_33 = W*in
   wire signed [9:0] m355_33;
   assign m355_33 =10'b0;

   // m355_34 = W*in
   wire signed [9:0] m355_34;
   assign m355_34 =10'b0;

   // m355_35 = W*in
   wire signed [9:0] m355_35;
   assign m355_35 ={ {5{neg355[5]}} , neg355[5:1] };

   // m355_36 = W*in
   wire signed [9:0] m355_36;
   assign m355_36 =10'b0;

   // m355_37 = W*in
   wire signed [9:0] m355_37;
   assign m355_37 =10'b0;

   // m355_38 = W*in
   wire signed [9:0] m355_38;
   assign m355_38 =10'b0;

   // m355_39 = W*in
   wire signed [9:0] m355_39;
   assign m355_39 =10'b0;

   // m355_40 = W*in
   wire signed [9:0] m355_40;
   assign m355_40 =10'b0;

   // m355_41 = W*in
   wire signed [9:0] m355_41;
   assign m355_41 =10'b0;

   // m355_42 = W*in
   wire signed [9:0] m355_42;
   assign m355_42 =10'b0;

   // m355_43 = W*in
   wire signed [9:0] m355_43;
   assign m355_43 =10'b0;

   // m355_44 = W*in
   wire signed [9:0] m355_44;
   assign m355_44 =10'b0;

   // m355_45 = W*in
   wire signed [9:0] m355_45;
   assign m355_45 =10'b0;

   // m355_46 = W*in
   wire signed [9:0] m355_46;
   assign m355_46 =10'b0;

   // m355_47 = W*in
   wire signed [9:0] m355_47;
   assign m355_47 =10'b0;

   // m355_48 = W*in
   wire signed [9:0] m355_48;
   assign m355_48 =10'b0;

   // m355_49 = W*in
   wire signed [9:0] m355_49;
   assign m355_49 =10'b0;

   // m355_50 = W*in
   wire signed [9:0] m355_50;
   assign m355_50 =10'b0;

   // m355_51 = W*in
   wire signed [9:0] m355_51;
   assign m355_51 =10'b0;

   // m355_52 = W*in
   wire signed [9:0] m355_52;
   assign m355_52 =10'b0;

   // m355_53 = W*in
   wire signed [9:0] m355_53;
   assign m355_53 =10'b0;

   // m355_54 = W*in
   wire signed [9:0] m355_54;
   assign m355_54 =10'b0;

   // m355_55 = W*in
   wire signed [9:0] m355_55;
   assign m355_55 =10'b0;

   // m355_56 = W*in
   wire signed [9:0] m355_56;
   assign m355_56 =10'b0;

   // m355_57 = W*in
   wire signed [9:0] m355_57;
   assign m355_57 =10'b0;

   // m355_58 = W*in
   wire signed [9:0] m355_58;
   assign m355_58 =10'b0;

   // m355_59 = W*in
   wire signed [9:0] m355_59;
   assign m355_59 =10'b0;

   // m355_60 = W*in
   wire signed [9:0] m355_60;
   assign m355_60 =10'b0;

   // m355_61 = W*in
   wire signed [9:0] m355_61;
   assign m355_61 =10'b0;

   // m355_62 = W*in
   wire signed [9:0] m355_62;
   assign m355_62 =10'b0;

   // m355_63 = W*in
   wire signed [9:0] m355_63;
   assign m355_63 =10'b0;

   // m355_64 = W*in
   wire signed [9:0] m355_64;
   assign m355_64 =10'b0;

   // m355_65 = W*in
   wire signed [9:0] m355_65;
   assign m355_65 =10'b0;

   // m355_66 = W*in
   wire signed [9:0] m355_66;
   assign m355_66 =10'b0;

   // m355_67 = W*in
   wire signed [9:0] m355_67;
   assign m355_67 =10'b0;

   // m355_68 = W*in
   wire signed [9:0] m355_68;
   assign m355_68 =10'b0;

   // m355_69 = W*in
   wire signed [9:0] m355_69;
   assign m355_69 =10'b0;

   // m355_70 = W*in
   wire signed [9:0] m355_70;
   assign m355_70 =10'b0;

   // m355_71 = W*in
   wire signed [9:0] m355_71;
   assign m355_71 =10'b0;

   // m355_72 = W*in
   wire signed [9:0] m355_72;
   assign m355_72 =10'b0;

   // m355_73 = W*in
   wire signed [9:0] m355_73;
   assign m355_73 =10'b0;

   // m355_74 = W*in
   wire signed [9:0] m355_74;
   assign m355_74 =10'b0;

   // m355_75 = W*in
   wire signed [9:0] m355_75;
   assign m355_75 =10'b0;

   // m355_76 = W*in
   wire signed [9:0] m355_76;
   assign m355_76 =10'b0;

   // m355_77 = W*in
   wire signed [9:0] m355_77;
   assign m355_77 =10'b0;

   // m355_78 = W*in
   wire signed [9:0] m355_78;
   assign m355_78 =10'b0;

   // m355_79 = W*in
   wire signed [9:0] m355_79;
   assign m355_79 =10'b0;

   // m355_80 = W*in
   wire signed [9:0] m355_80;
   assign m355_80 =10'b0;

   // m355_81 = W*in
   wire signed [9:0] m355_81;
   assign m355_81 =10'b0;

   // m355_82 = W*in
   wire signed [9:0] m355_82;
   assign m355_82 =10'b0;

   // m355_83 = W*in
   wire signed [9:0] m355_83;
   assign m355_83 =10'b0;

   // m355_84 = W*in
   wire signed [9:0] m355_84;
   assign m355_84 =10'b0;

   // m355_85 = W*in
   wire signed [9:0] m355_85;
   assign m355_85 ={ {4{neg355[5]}} , neg355[5:0] };

   // m355_86 = W*in
   wire signed [9:0] m355_86;
   assign m355_86 =10'b0;

   // m355_87 = W*in
   wire signed [9:0] m355_87;
   assign m355_87 =10'b0;

   // m355_88 = W*in
   wire signed [9:0] m355_88;
   assign m355_88 ={ {4{in355[5]}} , in355[5:0] };

   // m355_89 = W*in
   wire signed [9:0] m355_89;
   assign m355_89 =10'b0;

   // m355_90 = W*in
   wire signed [9:0] m355_90;
   assign m355_90 =10'b0;

   // m355_91 = W*in
   wire signed [9:0] m355_91;
   assign m355_91 =10'b0;

   // m355_92 = W*in
   wire signed [9:0] m355_92;
   assign m355_92 ={ {4{in355[5]}} , in355[5:0] };

   // m355_93 = W*in
   wire signed [9:0] m355_93;
   assign m355_93 =10'b0;

   // m355_94 = W*in
   wire signed [9:0] m355_94;
   assign m355_94 =10'b0;

   // m355_95 = W*in
   wire signed [9:0] m355_95;
   assign m355_95 =10'b0;

   // m355_96 = W*in
   wire signed [9:0] m355_96;
   assign m355_96 =10'b0;

   // m355_97 = W*in
   wire signed [9:0] m355_97;
   assign m355_97 =10'b0;

   // m355_98 = W*in
   wire signed [9:0] m355_98;
   assign m355_98 =10'b0;

   // m355_99 = W*in
   wire signed [9:0] m355_99;
   assign m355_99 =10'b0;

   // m355_100 = W*in
   wire signed [9:0] m355_100;
   assign m355_100 =10'b0;

   // m355_101 = W*in
   wire signed [9:0] m355_101;
   assign m355_101 =10'b0;

   // m355_102 = W*in
   wire signed [9:0] m355_102;
   assign m355_102 ={ {5{neg355[5]}} , neg355[5:1] };

   // m355_103 = W*in
   wire signed [9:0] m355_103;
   assign m355_103 =10'b0;

   // m355_104 = W*in
   wire signed [9:0] m355_104;
   assign m355_104 =10'b0;

   // m355_105 = W*in
   wire signed [9:0] m355_105;
   assign m355_105 =10'b0;

   // m355_106 = W*in
   wire signed [9:0] m355_106;
   assign m355_106 =10'b0;

   // m355_107 = W*in
   wire signed [9:0] m355_107;
   assign m355_107 =10'b0;

   // m355_108 = W*in
   wire signed [9:0] m355_108;
   assign m355_108 =10'b0;

   // m355_109 = W*in
   wire signed [9:0] m355_109;
   assign m355_109 =10'b0;

   // m355_110 = W*in
   wire signed [9:0] m355_110;
   assign m355_110 =10'b0;

   // m355_111 = W*in
   wire signed [9:0] m355_111;
   assign m355_111 =10'b0;

   // m355_112 = W*in
   wire signed [9:0] m355_112;
   assign m355_112 =10'b0;

   // m355_113 = W*in
   wire signed [9:0] m355_113;
   assign m355_113 =10'b0;

   // m355_114 = W*in
   wire signed [9:0] m355_114;
   assign m355_114 =10'b0;

   // m355_115 = W*in
   wire signed [9:0] m355_115;
   assign m355_115 =10'b0;

   // m355_116 = W*in
   wire signed [9:0] m355_116;
   assign m355_116 =10'b0;

   // m355_117 = W*in
   wire signed [9:0] m355_117;
   assign m355_117 =10'b0;

   // m356_1 = W*in
   wire signed [9:0] m356_1;
   assign m356_1 =10'b0;

   // m356_2 = W*in
   wire signed [9:0] m356_2;
   assign m356_2 =10'b0;

   // m356_3 = W*in
   wire signed [9:0] m356_3;
   assign m356_3 =10'b0;

   // m356_4 = W*in
   wire signed [9:0] m356_4;
   assign m356_4 =10'b0;

   // m356_5 = W*in
   wire signed [9:0] m356_5;
   assign m356_5 =10'b0;

   // m356_6 = W*in
   wire signed [9:0] m356_6;
   assign m356_6 =10'b0;

   // m356_7 = W*in
   wire signed [9:0] m356_7;
   assign m356_7 =10'b0;

   // m356_8 = W*in
   wire signed [9:0] m356_8;
   assign m356_8 =10'b0;

   // m356_9 = W*in
   wire signed [9:0] m356_9;
   assign m356_9 =10'b0;

   // m356_10 = W*in
   wire signed [9:0] m356_10;
   assign m356_10 =10'b0;

   // m356_11 = W*in
   wire signed [9:0] m356_11;
   assign m356_11 =10'b0;

   // m356_12 = W*in
   wire signed [9:0] m356_12;
   assign m356_12 =10'b0;

   // m356_13 = W*in
   wire signed [9:0] m356_13;
   assign m356_13 =10'b0;

   // m356_14 = W*in
   wire signed [9:0] m356_14;
   assign m356_14 =10'b0;

   // m356_15 = W*in
   wire signed [9:0] m356_15;
   assign m356_15 =10'b0;

   // m356_16 = W*in
   wire signed [9:0] m356_16;
   assign m356_16 =10'b0;

   // m356_17 = W*in
   wire signed [9:0] m356_17;
   assign m356_17 =10'b0;

   // m356_18 = W*in
   wire signed [9:0] m356_18;
   assign m356_18 =10'b0;

   // m356_19 = W*in
   wire signed [9:0] m356_19;
   assign m356_19 =10'b0;

   // m356_20 = W*in
   wire signed [9:0] m356_20;
   assign m356_20 =10'b0;

   // m356_21 = W*in
   wire signed [9:0] m356_21;
   assign m356_21 =10'b0;

   // m356_22 = W*in
   wire signed [9:0] m356_22;
   assign m356_22 =10'b0;

   // m356_23 = W*in
   wire signed [9:0] m356_23;
   assign m356_23 =10'b0;

   // m356_24 = W*in
   wire signed [9:0] m356_24;
   assign m356_24 =10'b0;

   // m356_25 = W*in
   wire signed [9:0] m356_25;
   assign m356_25 =10'b0;

   // m356_26 = W*in
   wire signed [9:0] m356_26;
   assign m356_26 =10'b0;

   // m356_27 = W*in
   wire signed [9:0] m356_27;
   assign m356_27 =10'b0;

   // m356_28 = W*in
   wire signed [9:0] m356_28;
   assign m356_28 =10'b0;

   // m356_29 = W*in
   wire signed [9:0] m356_29;
   assign m356_29 =10'b0;

   // m356_30 = W*in
   wire signed [9:0] m356_30;
   assign m356_30 ={ {5{neg356[5]}} , neg356[5:1] };

   // m356_31 = W*in
   wire signed [9:0] m356_31;
   assign m356_31 =10'b0;

   // m356_32 = W*in
   wire signed [9:0] m356_32;
   assign m356_32 =10'b0;

   // m356_33 = W*in
   wire signed [9:0] m356_33;
   assign m356_33 =10'b0;

   // m356_34 = W*in
   wire signed [9:0] m356_34;
   assign m356_34 =10'b0;

   // m356_35 = W*in
   wire signed [9:0] m356_35;
   assign m356_35 =10'b0;

   // m356_36 = W*in
   wire signed [9:0] m356_36;
   assign m356_36 =10'b0;

   // m356_37 = W*in
   wire signed [9:0] m356_37;
   assign m356_37 =10'b0;

   // m356_38 = W*in
   wire signed [9:0] m356_38;
   assign m356_38 =10'b0;

   // m356_39 = W*in
   wire signed [9:0] m356_39;
   assign m356_39 =10'b0;

   // m356_40 = W*in
   wire signed [9:0] m356_40;
   assign m356_40 =10'b0;

   // m356_41 = W*in
   wire signed [9:0] m356_41;
   assign m356_41 =10'b0;

   // m356_42 = W*in
   wire signed [9:0] m356_42;
   assign m356_42 =10'b0;

   // m356_43 = W*in
   wire signed [9:0] m356_43;
   assign m356_43 =10'b0;

   // m356_44 = W*in
   wire signed [9:0] m356_44;
   assign m356_44 =10'b0;

   // m356_45 = W*in
   wire signed [9:0] m356_45;
   assign m356_45 =10'b0;

   // m356_46 = W*in
   wire signed [9:0] m356_46;
   assign m356_46 =10'b0;

   // m356_47 = W*in
   wire signed [9:0] m356_47;
   assign m356_47 =10'b0;

   // m356_48 = W*in
   wire signed [9:0] m356_48;
   assign m356_48 ={ {4{in356[5]}} , in356[5:0] };

   // m356_49 = W*in
   wire signed [9:0] m356_49;
   assign m356_49 =10'b0;

   // m356_50 = W*in
   wire signed [9:0] m356_50;
   assign m356_50 =10'b0;

   // m356_51 = W*in
   wire signed [9:0] m356_51;
   assign m356_51 =10'b0;

   // m356_52 = W*in
   wire signed [9:0] m356_52;
   assign m356_52 =10'b0;

   // m356_53 = W*in
   wire signed [9:0] m356_53;
   assign m356_53 =10'b0;

   // m356_54 = W*in
   wire signed [9:0] m356_54;
   assign m356_54 =10'b0;

   // m356_55 = W*in
   wire signed [9:0] m356_55;
   assign m356_55 =10'b0;

   // m356_56 = W*in
   wire signed [9:0] m356_56;
   assign m356_56 =10'b0;

   // m356_57 = W*in
   wire signed [9:0] m356_57;
   assign m356_57 =10'b0;

   // m356_58 = W*in
   wire signed [9:0] m356_58;
   assign m356_58 =10'b0;

   // m356_59 = W*in
   wire signed [9:0] m356_59;
   assign m356_59 =10'b0;

   // m356_60 = W*in
   wire signed [9:0] m356_60;
   assign m356_60 =10'b0;

   // m356_61 = W*in
   wire signed [9:0] m356_61;
   assign m356_61 =10'b0;

   // m356_62 = W*in
   wire signed [9:0] m356_62;
   assign m356_62 =10'b0;

   // m356_63 = W*in
   wire signed [9:0] m356_63;
   assign m356_63 =10'b0;

   // m356_64 = W*in
   wire signed [9:0] m356_64;
   assign m356_64 =10'b0;

   // m356_65 = W*in
   wire signed [9:0] m356_65;
   assign m356_65 =10'b0;

   // m356_66 = W*in
   wire signed [9:0] m356_66;
   assign m356_66 ={ {5{neg356[5]}} , neg356[5:1] };

   // m356_67 = W*in
   wire signed [9:0] m356_67;
   assign m356_67 =10'b0;

   // m356_68 = W*in
   wire signed [9:0] m356_68;
   assign m356_68 =10'b0;

   // m356_69 = W*in
   wire signed [9:0] m356_69;
   assign m356_69 =10'b0;

   // m356_70 = W*in
   wire signed [9:0] m356_70;
   assign m356_70 =10'b0;

   // m356_71 = W*in
   wire signed [9:0] m356_71;
   assign m356_71 =10'b0;

   // m356_72 = W*in
   wire signed [9:0] m356_72;
   assign m356_72 ={ {4{in356[5]}} , in356[5:0] };

   // m356_73 = W*in
   wire signed [9:0] m356_73;
   assign m356_73 =10'b0;

   // m356_74 = W*in
   wire signed [9:0] m356_74;
   assign m356_74 =10'b0;

   // m356_75 = W*in
   wire signed [9:0] m356_75;
   assign m356_75 =10'b0;

   // m356_76 = W*in
   wire signed [9:0] m356_76;
   assign m356_76 =10'b0;

   // m356_77 = W*in
   wire signed [9:0] m356_77;
   assign m356_77 =10'b0;

   // m356_78 = W*in
   wire signed [9:0] m356_78;
   assign m356_78 =10'b0;

   // m356_79 = W*in
   wire signed [9:0] m356_79;
   assign m356_79 =10'b0;

   // m356_80 = W*in
   wire signed [9:0] m356_80;
   assign m356_80 =10'b0;

   // m356_81 = W*in
   wire signed [9:0] m356_81;
   assign m356_81 =10'b0;

   // m356_82 = W*in
   wire signed [9:0] m356_82;
   assign m356_82 =10'b0;

   // m356_83 = W*in
   wire signed [9:0] m356_83;
   assign m356_83 =10'b0;

   // m356_84 = W*in
   wire signed [9:0] m356_84;
   assign m356_84 =10'b0;

   // m356_85 = W*in
   wire signed [9:0] m356_85;
   assign m356_85 =10'b0;

   // m356_86 = W*in
   wire signed [9:0] m356_86;
   assign m356_86 =10'b0;

   // m356_87 = W*in
   wire signed [9:0] m356_87;
   assign m356_87 =10'b0;

   // m356_88 = W*in
   wire signed [9:0] m356_88;
   assign m356_88 =10'b0;

   // m356_89 = W*in
   wire signed [9:0] m356_89;
   assign m356_89 =10'b0;

   // m356_90 = W*in
   wire signed [9:0] m356_90;
   assign m356_90 =10'b0;

   // m356_91 = W*in
   wire signed [9:0] m356_91;
   assign m356_91 =10'b0;

   // m356_92 = W*in
   wire signed [9:0] m356_92;
   assign m356_92 =10'b0;

   // m356_93 = W*in
   wire signed [9:0] m356_93;
   assign m356_93 =10'b0;

   // m356_94 = W*in
   wire signed [9:0] m356_94;
   assign m356_94 =10'b0;

   // m356_95 = W*in
   wire signed [9:0] m356_95;
   assign m356_95 =10'b0;

   // m356_96 = W*in
   wire signed [9:0] m356_96;
   assign m356_96 =10'b0;

   // m356_97 = W*in
   wire signed [9:0] m356_97;
   assign m356_97 =10'b0;

   // m356_98 = W*in
   wire signed [9:0] m356_98;
   assign m356_98 =10'b0;

   // m356_99 = W*in
   wire signed [9:0] m356_99;
   assign m356_99 =10'b0;

   // m356_100 = W*in
   wire signed [9:0] m356_100;
   assign m356_100 =10'b0;

   // m356_101 = W*in
   wire signed [9:0] m356_101;
   assign m356_101 =10'b0;

   // m356_102 = W*in
   wire signed [9:0] m356_102;
   assign m356_102 =10'b0;

   // m356_103 = W*in
   wire signed [9:0] m356_103;
   assign m356_103 =10'b0;

   // m356_104 = W*in
   wire signed [9:0] m356_104;
   assign m356_104 =10'b0;

   // m356_105 = W*in
   wire signed [9:0] m356_105;
   assign m356_105 =10'b0;

   // m356_106 = W*in
   wire signed [9:0] m356_106;
   assign m356_106 =10'b0;

   // m356_107 = W*in
   wire signed [9:0] m356_107;
   assign m356_107 =10'b0;

   // m356_108 = W*in
   wire signed [9:0] m356_108;
   assign m356_108 =10'b0;

   // m356_109 = W*in
   wire signed [9:0] m356_109;
   assign m356_109 =10'b0;

   // m356_110 = W*in
   wire signed [9:0] m356_110;
   assign m356_110 =10'b0;

   // m356_111 = W*in
   wire signed [9:0] m356_111;
   assign m356_111 =10'b0;

   // m356_112 = W*in
   wire signed [9:0] m356_112;
   assign m356_112 =10'b0;

   // m356_113 = W*in
   wire signed [9:0] m356_113;
   assign m356_113 =10'b0;

   // m356_114 = W*in
   wire signed [9:0] m356_114;
   assign m356_114 =10'b0;

   // m356_115 = W*in
   wire signed [9:0] m356_115;
   assign m356_115 =10'b0;

   // m356_116 = W*in
   wire signed [9:0] m356_116;
   assign m356_116 =10'b0;

   // m356_117 = W*in
   wire signed [9:0] m356_117;
   assign m356_117 =10'b0;

   // m357_1 = W*in
   wire signed [9:0] m357_1;
   assign m357_1 =10'b0;

   // m357_2 = W*in
   wire signed [9:0] m357_2;
   assign m357_2 ={ {4{in357[5]}} , in357[5:0] };

   // m357_3 = W*in
   wire signed [9:0] m357_3;
   assign m357_3 =10'b0;

   // m357_4 = W*in
   wire signed [9:0] m357_4;
   assign m357_4 =10'b0;

   // m357_5 = W*in
   wire signed [9:0] m357_5;
   assign m357_5 =10'b0;

   // m357_6 = W*in
   wire signed [9:0] m357_6;
   assign m357_6 =10'b0;

   // m357_7 = W*in
   wire signed [9:0] m357_7;
   assign m357_7 =10'b0;

   // m357_8 = W*in
   wire signed [9:0] m357_8;
   assign m357_8 =10'b0;

   // m357_9 = W*in
   wire signed [9:0] m357_9;
   assign m357_9 =10'b0;

   // m357_10 = W*in
   wire signed [9:0] m357_10;
   assign m357_10 =10'b0;

   // m357_11 = W*in
   wire signed [9:0] m357_11;
   assign m357_11 =10'b0;

   // m357_12 = W*in
   wire signed [9:0] m357_12;
   assign m357_12 =10'b0;

   // m357_13 = W*in
   wire signed [9:0] m357_13;
   assign m357_13 =10'b0;

   // m357_14 = W*in
   wire signed [9:0] m357_14;
   assign m357_14 =10'b0;

   // m357_15 = W*in
   wire signed [9:0] m357_15;
   assign m357_15 =10'b0;

   // m357_16 = W*in
   wire signed [9:0] m357_16;
   assign m357_16 =10'b0;

   // m357_17 = W*in
   wire signed [9:0] m357_17;
   assign m357_17 =10'b0;

   // m357_18 = W*in
   wire signed [9:0] m357_18;
   assign m357_18 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_19 = W*in
   wire signed [9:0] m357_19;
   assign m357_19 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_20 = W*in
   wire signed [9:0] m357_20;
   assign m357_20 =10'b0;

   // m357_21 = W*in
   wire signed [9:0] m357_21;
   assign m357_21 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_22 = W*in
   wire signed [9:0] m357_22;
   assign m357_22 =10'b0;

   // m357_23 = W*in
   wire signed [9:0] m357_23;
   assign m357_23 ={ {5{in357[5]}} , in357[5:1] };

   // m357_24 = W*in
   wire signed [9:0] m357_24;
   assign m357_24 =10'b0;

   // m357_25 = W*in
   wire signed [9:0] m357_25;
   assign m357_25 =10'b0;

   // m357_26 = W*in
   wire signed [9:0] m357_26;
   assign m357_26 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_27 = W*in
   wire signed [9:0] m357_27;
   assign m357_27 =10'b0;

   // m357_28 = W*in
   wire signed [9:0] m357_28;
   assign m357_28 =10'b0;

   // m357_29 = W*in
   wire signed [9:0] m357_29;
   assign m357_29 =10'b0;

   // m357_30 = W*in
   wire signed [9:0] m357_30;
   assign m357_30 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_31 = W*in
   wire signed [9:0] m357_31;
   assign m357_31 =10'b0;

   // m357_32 = W*in
   wire signed [9:0] m357_32;
   assign m357_32 =10'b0;

   // m357_33 = W*in
   wire signed [9:0] m357_33;
   assign m357_33 =10'b0;

   // m357_34 = W*in
   wire signed [9:0] m357_34;
   assign m357_34 ={ {5{in357[5]}} , in357[5:1] };

   // m357_35 = W*in
   wire signed [9:0] m357_35;
   assign m357_35 =10'b0;

   // m357_36 = W*in
   wire signed [9:0] m357_36;
   assign m357_36 =10'b0;

   // m357_37 = W*in
   wire signed [9:0] m357_37;
   assign m357_37 =10'b0;

   // m357_38 = W*in
   wire signed [9:0] m357_38;
   assign m357_38 ={ {4{neg357[5]}} , neg357[5:0] };

   // m357_39 = W*in
   wire signed [9:0] m357_39;
   assign m357_39 =10'b0;

   // m357_40 = W*in
   wire signed [9:0] m357_40;
   assign m357_40 =10'b0;

   // m357_41 = W*in
   wire signed [9:0] m357_41;
   assign m357_41 =10'b0;

   // m357_42 = W*in
   wire signed [9:0] m357_42;
   assign m357_42 =10'b0;

   // m357_43 = W*in
   wire signed [9:0] m357_43;
   assign m357_43 =10'b0;

   // m357_44 = W*in
   wire signed [9:0] m357_44;
   assign m357_44 =10'b0;

   // m357_45 = W*in
   wire signed [9:0] m357_45;
   assign m357_45 =10'b0;

   // m357_46 = W*in
   wire signed [9:0] m357_46;
   assign m357_46 =10'b0;

   // m357_47 = W*in
   wire signed [9:0] m357_47;
   assign m357_47 =10'b0;

   // m357_48 = W*in
   wire signed [9:0] m357_48;
   assign m357_48 =10'b0;

   // m357_49 = W*in
   wire signed [9:0] m357_49;
   assign m357_49 =10'b0;

   // m357_50 = W*in
   wire signed [9:0] m357_50;
   assign m357_50 =10'b0;

   // m357_51 = W*in
   wire signed [9:0] m357_51;
   assign m357_51 ={ {4{in357[5]}} , in357[5:0] };

   // m357_52 = W*in
   wire signed [9:0] m357_52;
   assign m357_52 ={ {4{in357[5]}} , in357[5:0] };

   // m357_53 = W*in
   wire signed [9:0] m357_53;
   assign m357_53 =10'b0;

   // m357_54 = W*in
   wire signed [9:0] m357_54;
   assign m357_54 =10'b0;

   // m357_55 = W*in
   wire signed [9:0] m357_55;
   assign m357_55 =10'b0;

   // m357_56 = W*in
   wire signed [9:0] m357_56;
   assign m357_56 =10'b0;

   // m357_57 = W*in
   wire signed [9:0] m357_57;
   assign m357_57 =10'b0;

   // m357_58 = W*in
   wire signed [9:0] m357_58;
   assign m357_58 =10'b0;

   // m357_59 = W*in
   wire signed [9:0] m357_59;
   assign m357_59 =10'b0;

   // m357_60 = W*in
   wire signed [9:0] m357_60;
   assign m357_60 =10'b0;

   // m357_61 = W*in
   wire signed [9:0] m357_61;
   assign m357_61 =10'b0;

   // m357_62 = W*in
   wire signed [9:0] m357_62;
   assign m357_62 =10'b0;

   // m357_63 = W*in
   wire signed [9:0] m357_63;
   assign m357_63 ={ {4{neg357[5]}} , neg357[5:0] };

   // m357_64 = W*in
   wire signed [9:0] m357_64;
   assign m357_64 =10'b0;

   // m357_65 = W*in
   wire signed [9:0] m357_65;
   assign m357_65 =10'b0;

   // m357_66 = W*in
   wire signed [9:0] m357_66;
   assign m357_66 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_67 = W*in
   wire signed [9:0] m357_67;
   assign m357_67 =10'b0;

   // m357_68 = W*in
   wire signed [9:0] m357_68;
   assign m357_68 =10'b0;

   // m357_69 = W*in
   wire signed [9:0] m357_69;
   assign m357_69 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_70 = W*in
   wire signed [9:0] m357_70;
   assign m357_70 ={ {4{neg357[5]}} , neg357[5:0] };

   // m357_71 = W*in
   wire signed [9:0] m357_71;
   assign m357_71 =10'b0;

   // m357_72 = W*in
   wire signed [9:0] m357_72;
   assign m357_72 ={ {5{neg357[5]}} , neg357[5:1] };

   // m357_73 = W*in
   wire signed [9:0] m357_73;
   assign m357_73 ={ {5{in357[5]}} , in357[5:1] };

   // m357_74 = W*in
   wire signed [9:0] m357_74;
   assign m357_74 ={ {4{neg357[5]}} , neg357[5:0] };

   // m357_75 = W*in
   wire signed [9:0] m357_75;
   assign m357_75 =10'b0;

   // m357_76 = W*in
   wire signed [9:0] m357_76;
   assign m357_76 =10'b0;

   // m357_77 = W*in
   wire signed [9:0] m357_77;
   assign m357_77 =10'b0;

   // m357_78 = W*in
   wire signed [9:0] m357_78;
   assign m357_78 =10'b0;

   // m357_79 = W*in
   wire signed [9:0] m357_79;
   assign m357_79 =10'b0;

   // m357_80 = W*in
   wire signed [9:0] m357_80;
   assign m357_80 ={ {4{in357[5]}} , in357[5:0] };

   // m357_81 = W*in
   wire signed [9:0] m357_81;
   assign m357_81 =10'b0;

   // m357_82 = W*in
   wire signed [9:0] m357_82;
   assign m357_82 =10'b0;

   // m357_83 = W*in
   wire signed [9:0] m357_83;
   assign m357_83 =10'b0;

   // m357_84 = W*in
   wire signed [9:0] m357_84;
   assign m357_84 =10'b0;

   // m357_85 = W*in
   wire signed [9:0] m357_85;
   assign m357_85 =10'b0;

   // m357_86 = W*in
   wire signed [9:0] m357_86;
   assign m357_86 =10'b0;

   // m357_87 = W*in
   wire signed [9:0] m357_87;
   assign m357_87 =10'b0;

   // m357_88 = W*in
   wire signed [9:0] m357_88;
   assign m357_88 =10'b0;

   // m357_89 = W*in
   wire signed [9:0] m357_89;
   assign m357_89 =10'b0;

   // m357_90 = W*in
   wire signed [9:0] m357_90;
   assign m357_90 =10'b0;

   // m357_91 = W*in
   wire signed [9:0] m357_91;
   assign m357_91 ={ {4{neg357[5]}} , neg357[5:0] };

   // m357_92 = W*in
   wire signed [9:0] m357_92;
   assign m357_92 =10'b0;

   // m357_93 = W*in
   wire signed [9:0] m357_93;
   assign m357_93 =10'b0;

   // m357_94 = W*in
   wire signed [9:0] m357_94;
   assign m357_94 =10'b0;

   // m357_95 = W*in
   wire signed [9:0] m357_95;
   assign m357_95 =10'b0;

   // m357_96 = W*in
   wire signed [9:0] m357_96;
   assign m357_96 =10'b0;

   // m357_97 = W*in
   wire signed [9:0] m357_97;
   assign m357_97 =10'b0;

   // m357_98 = W*in
   wire signed [9:0] m357_98;
   assign m357_98 =10'b0;

   // m357_99 = W*in
   wire signed [9:0] m357_99;
   assign m357_99 =10'b0;

   // m357_100 = W*in
   wire signed [9:0] m357_100;
   assign m357_100 =10'b0;

   // m357_101 = W*in
   wire signed [9:0] m357_101;
   assign m357_101 =10'b0;

   // m357_102 = W*in
   wire signed [9:0] m357_102;
   assign m357_102 =10'b0;

   // m357_103 = W*in
   wire signed [9:0] m357_103;
   assign m357_103 =10'b0;

   // m357_104 = W*in
   wire signed [9:0] m357_104;
   assign m357_104 =10'b0;

   // m357_105 = W*in
   wire signed [9:0] m357_105;
   assign m357_105 =10'b0;

   // m357_106 = W*in
   wire signed [9:0] m357_106;
   assign m357_106 =10'b0;

   // m357_107 = W*in
   wire signed [9:0] m357_107;
   assign m357_107 =10'b0;

   // m357_108 = W*in
   wire signed [9:0] m357_108;
   assign m357_108 =10'b0;

   // m357_109 = W*in
   wire signed [9:0] m357_109;
   assign m357_109 =10'b0;

   // m357_110 = W*in
   wire signed [9:0] m357_110;
   assign m357_110 =10'b0;

   // m357_111 = W*in
   wire signed [9:0] m357_111;
   assign m357_111 =10'b0;

   // m357_112 = W*in
   wire signed [9:0] m357_112;
   assign m357_112 =10'b0;

   // m357_113 = W*in
   wire signed [9:0] m357_113;
   assign m357_113 =10'b0;

   // m357_114 = W*in
   wire signed [9:0] m357_114;
   assign m357_114 =10'b0;

   // m357_115 = W*in
   wire signed [9:0] m357_115;
   assign m357_115 =10'b0;

   // m357_116 = W*in
   wire signed [9:0] m357_116;
   assign m357_116 =10'b0;

   // m357_117 = W*in
   wire signed [9:0] m357_117;
   assign m357_117 =10'b0;

   // m358_1 = W*in
   wire signed [9:0] m358_1;
   assign m358_1 =10'b0;

   // m358_2 = W*in
   wire signed [9:0] m358_2;
   assign m358_2 =10'b0;

   // m358_3 = W*in
   wire signed [9:0] m358_3;
   assign m358_3 ={ {4{in358[5]}} , in358[5:0] };

   // m358_4 = W*in
   wire signed [9:0] m358_4;
   assign m358_4 =10'b0;

   // m358_5 = W*in
   wire signed [9:0] m358_5;
   assign m358_5 =10'b0;

   // m358_6 = W*in
   wire signed [9:0] m358_6;
   assign m358_6 =10'b0;

   // m358_7 = W*in
   wire signed [9:0] m358_7;
   assign m358_7 =10'b0;

   // m358_8 = W*in
   wire signed [9:0] m358_8;
   assign m358_8 =10'b0;

   // m358_9 = W*in
   wire signed [9:0] m358_9;
   assign m358_9 =10'b0;

   // m358_10 = W*in
   wire signed [9:0] m358_10;
   assign m358_10 =10'b0;

   // m358_11 = W*in
   wire signed [9:0] m358_11;
   assign m358_11 =10'b0;

   // m358_12 = W*in
   wire signed [9:0] m358_12;
   assign m358_12 ={ {4{in358[5]}} , in358[5:0] };

   // m358_13 = W*in
   wire signed [9:0] m358_13;
   assign m358_13 ={ {4{in358[5]}} , in358[5:0] };

   // m358_14 = W*in
   wire signed [9:0] m358_14;
   assign m358_14 =10'b0;

   // m358_15 = W*in
   wire signed [9:0] m358_15;
   assign m358_15 =10'b0;

   // m358_16 = W*in
   wire signed [9:0] m358_16;
   assign m358_16 ={ {5{neg358[5]}} , neg358[5:1] };

   // m358_17 = W*in
   wire signed [9:0] m358_17;
   assign m358_17 =10'b0;

   // m358_18 = W*in
   wire signed [9:0] m358_18;
   assign m358_18 ={ {5{neg358[5]}} , neg358[5:1] };

   // m358_19 = W*in
   wire signed [9:0] m358_19;
   assign m358_19 =10'b0;

   // m358_20 = W*in
   wire signed [9:0] m358_20;
   assign m358_20 ={ {5{neg358[5]}} , neg358[5:1] };

   // m358_21 = W*in
   wire signed [9:0] m358_21;
   assign m358_21 =10'b0;

   // m358_22 = W*in
   wire signed [9:0] m358_22;
   assign m358_22 =10'b0;

   // m358_23 = W*in
   wire signed [9:0] m358_23;
   assign m358_23 ={ {4{in358[5]}} , in358[5:0] };

   // m358_24 = W*in
   wire signed [9:0] m358_24;
   assign m358_24 ={ {4{in358[5]}} , in358[5:0] };

   // m358_25 = W*in
   wire signed [9:0] m358_25;
   assign m358_25 =10'b0;

   // m358_26 = W*in
   wire signed [9:0] m358_26;
   assign m358_26 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_27 = W*in
   wire signed [9:0] m358_27;
   assign m358_27 ={ {5{in358[5]}} , in358[5:1] };

   // m358_28 = W*in
   wire signed [9:0] m358_28;
   assign m358_28 =10'b0;

   // m358_29 = W*in
   wire signed [9:0] m358_29;
   assign m358_29 =10'b0;

   // m358_30 = W*in
   wire signed [9:0] m358_30;
   assign m358_30 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_31 = W*in
   wire signed [9:0] m358_31;
   assign m358_31 ={ {4{in358[5]}} , in358[5:0] };

   // m358_32 = W*in
   wire signed [9:0] m358_32;
   assign m358_32 =10'b0;

   // m358_33 = W*in
   wire signed [9:0] m358_33;
   assign m358_33 =10'b0;

   // m358_34 = W*in
   wire signed [9:0] m358_34;
   assign m358_34 ={ {5{in358[5]}} , in358[5:1] };

   // m358_35 = W*in
   wire signed [9:0] m358_35;
   assign m358_35 =10'b0;

   // m358_36 = W*in
   wire signed [9:0] m358_36;
   assign m358_36 =10'b0;

   // m358_37 = W*in
   wire signed [9:0] m358_37;
   assign m358_37 =10'b0;

   // m358_38 = W*in
   wire signed [9:0] m358_38;
   assign m358_38 =10'b0;

   // m358_39 = W*in
   wire signed [9:0] m358_39;
   assign m358_39 =10'b0;

   // m358_40 = W*in
   wire signed [9:0] m358_40;
   assign m358_40 =10'b0;

   // m358_41 = W*in
   wire signed [9:0] m358_41;
   assign m358_41 =10'b0;

   // m358_42 = W*in
   wire signed [9:0] m358_42;
   assign m358_42 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_43 = W*in
   wire signed [9:0] m358_43;
   assign m358_43 =10'b0;

   // m358_44 = W*in
   wire signed [9:0] m358_44;
   assign m358_44 =10'b0;

   // m358_45 = W*in
   wire signed [9:0] m358_45;
   assign m358_45 =10'b0;

   // m358_46 = W*in
   wire signed [9:0] m358_46;
   assign m358_46 =10'b0;

   // m358_47 = W*in
   wire signed [9:0] m358_47;
   assign m358_47 =10'b0;

   // m358_48 = W*in
   wire signed [9:0] m358_48;
   assign m358_48 =10'b0;

   // m358_49 = W*in
   wire signed [9:0] m358_49;
   assign m358_49 =10'b0;

   // m358_50 = W*in
   wire signed [9:0] m358_50;
   assign m358_50 =10'b0;

   // m358_51 = W*in
   wire signed [9:0] m358_51;
   assign m358_51 =10'b0;

   // m358_52 = W*in
   wire signed [9:0] m358_52;
   assign m358_52 =10'b0;

   // m358_53 = W*in
   wire signed [9:0] m358_53;
   assign m358_53 =10'b0;

   // m358_54 = W*in
   wire signed [9:0] m358_54;
   assign m358_54 =10'b0;

   // m358_55 = W*in
   wire signed [9:0] m358_55;
   assign m358_55 =10'b0;

   // m358_56 = W*in
   wire signed [9:0] m358_56;
   assign m358_56 =10'b0;

   // m358_57 = W*in
   wire signed [9:0] m358_57;
   assign m358_57 =10'b0;

   // m358_58 = W*in
   wire signed [9:0] m358_58;
   assign m358_58 =10'b0;

   // m358_59 = W*in
   wire signed [9:0] m358_59;
   assign m358_59 =10'b0;

   // m358_60 = W*in
   wire signed [9:0] m358_60;
   assign m358_60 =10'b0;

   // m358_61 = W*in
   wire signed [9:0] m358_61;
   assign m358_61 =10'b0;

   // m358_62 = W*in
   wire signed [9:0] m358_62;
   assign m358_62 =10'b0;

   // m358_63 = W*in
   wire signed [9:0] m358_63;
   assign m358_63 =10'b0;

   // m358_64 = W*in
   wire signed [9:0] m358_64;
   assign m358_64 =10'b0;

   // m358_65 = W*in
   wire signed [9:0] m358_65;
   assign m358_65 =10'b0;

   // m358_66 = W*in
   wire signed [9:0] m358_66;
   assign m358_66 =10'b0;

   // m358_67 = W*in
   wire signed [9:0] m358_67;
   assign m358_67 =10'b0;

   // m358_68 = W*in
   wire signed [9:0] m358_68;
   assign m358_68 ={ {4{in358[5]}} , in358[5:0] };

   // m358_69 = W*in
   wire signed [9:0] m358_69;
   assign m358_69 =10'b0;

   // m358_70 = W*in
   wire signed [9:0] m358_70;
   assign m358_70 =10'b0;

   // m358_71 = W*in
   wire signed [9:0] m358_71;
   assign m358_71 =10'b0;

   // m358_72 = W*in
   wire signed [9:0] m358_72;
   assign m358_72 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_73 = W*in
   wire signed [9:0] m358_73;
   assign m358_73 ={ {4{in358[5]}} , in358[5:0] };

   // m358_74 = W*in
   wire signed [9:0] m358_74;
   assign m358_74 =10'b0;

   // m358_75 = W*in
   wire signed [9:0] m358_75;
   assign m358_75 =10'b0;

   // m358_76 = W*in
   wire signed [9:0] m358_76;
   assign m358_76 =10'b0;

   // m358_77 = W*in
   wire signed [9:0] m358_77;
   assign m358_77 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_78 = W*in
   wire signed [9:0] m358_78;
   assign m358_78 =10'b0;

   // m358_79 = W*in
   wire signed [9:0] m358_79;
   assign m358_79 =10'b0;

   // m358_80 = W*in
   wire signed [9:0] m358_80;
   assign m358_80 ={ {4{in358[5]}} , in358[5:0] };

   // m358_81 = W*in
   wire signed [9:0] m358_81;
   assign m358_81 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_82 = W*in
   wire signed [9:0] m358_82;
   assign m358_82 =10'b0;

   // m358_83 = W*in
   wire signed [9:0] m358_83;
   assign m358_83 ={ {5{neg358[5]}} , neg358[5:1] };

   // m358_84 = W*in
   wire signed [9:0] m358_84;
   assign m358_84 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_85 = W*in
   wire signed [9:0] m358_85;
   assign m358_85 =10'b0;

   // m358_86 = W*in
   wire signed [9:0] m358_86;
   assign m358_86 =10'b0;

   // m358_87 = W*in
   wire signed [9:0] m358_87;
   assign m358_87 =10'b0;

   // m358_88 = W*in
   wire signed [9:0] m358_88;
   assign m358_88 =10'b0;

   // m358_89 = W*in
   wire signed [9:0] m358_89;
   assign m358_89 ={ {4{in358[5]}} , in358[5:0] };

   // m358_90 = W*in
   wire signed [9:0] m358_90;
   assign m358_90 =10'b0;

   // m358_91 = W*in
   wire signed [9:0] m358_91;
   assign m358_91 =10'b0;

   // m358_92 = W*in
   wire signed [9:0] m358_92;
   assign m358_92 =10'b0;

   // m358_93 = W*in
   wire signed [9:0] m358_93;
   assign m358_93 =10'b0;

   // m358_94 = W*in
   wire signed [9:0] m358_94;
   assign m358_94 =10'b0;

   // m358_95 = W*in
   wire signed [9:0] m358_95;
   assign m358_95 =10'b0;

   // m358_96 = W*in
   wire signed [9:0] m358_96;
   assign m358_96 =10'b0;

   // m358_97 = W*in
   wire signed [9:0] m358_97;
   assign m358_97 =10'b0;

   // m358_98 = W*in
   wire signed [9:0] m358_98;
   assign m358_98 =10'b0;

   // m358_99 = W*in
   wire signed [9:0] m358_99;
   assign m358_99 =10'b0;

   // m358_100 = W*in
   wire signed [9:0] m358_100;
   assign m358_100 =10'b0;

   // m358_101 = W*in
   wire signed [9:0] m358_101;
   assign m358_101 =10'b0;

   // m358_102 = W*in
   wire signed [9:0] m358_102;
   assign m358_102 =10'b0;

   // m358_103 = W*in
   wire signed [9:0] m358_103;
   assign m358_103 =10'b0;

   // m358_104 = W*in
   wire signed [9:0] m358_104;
   assign m358_104 =10'b0;

   // m358_105 = W*in
   wire signed [9:0] m358_105;
   assign m358_105 =10'b0;

   // m358_106 = W*in
   wire signed [9:0] m358_106;
   assign m358_106 =10'b0;

   // m358_107 = W*in
   wire signed [9:0] m358_107;
   assign m358_107 ={ {4{in358[5]}} , in358[5:0] };

   // m358_108 = W*in
   wire signed [9:0] m358_108;
   assign m358_108 =10'b0;

   // m358_109 = W*in
   wire signed [9:0] m358_109;
   assign m358_109 ={ {4{in358[5]}} , in358[5:0] };

   // m358_110 = W*in
   wire signed [9:0] m358_110;
   assign m358_110 =10'b0;

   // m358_111 = W*in
   wire signed [9:0] m358_111;
   assign m358_111 =10'b0;

   // m358_112 = W*in
   wire signed [9:0] m358_112;
   assign m358_112 =10'b0;

   // m358_113 = W*in
   wire signed [9:0] m358_113;
   assign m358_113 ={ {4{neg358[5]}} , neg358[5:0] };

   // m358_114 = W*in
   wire signed [9:0] m358_114;
   assign m358_114 =10'b0;

   // m358_115 = W*in
   wire signed [9:0] m358_115;
   assign m358_115 ={ {5{neg358[5]}} , neg358[5:1] };

   // m358_116 = W*in
   wire signed [9:0] m358_116;
   assign m358_116 =10'b0;

   // m358_117 = W*in
   wire signed [9:0] m358_117;
   assign m358_117 =10'b0;

   // m359_1 = W*in
   wire signed [9:0] m359_1;
   assign m359_1 =10'b0;

   // m359_2 = W*in
   wire signed [9:0] m359_2;
   assign m359_2 =10'b0;

   // m359_3 = W*in
   wire signed [9:0] m359_3;
   assign m359_3 =10'b0;

   // m359_4 = W*in
   wire signed [9:0] m359_4;
   assign m359_4 =10'b0;

   // m359_5 = W*in
   wire signed [9:0] m359_5;
   assign m359_5 =10'b0;

   // m359_6 = W*in
   wire signed [9:0] m359_6;
   assign m359_6 =10'b0;

   // m359_7 = W*in
   wire signed [9:0] m359_7;
   assign m359_7 =10'b0;

   // m359_8 = W*in
   wire signed [9:0] m359_8;
   assign m359_8 =10'b0;

   // m359_9 = W*in
   wire signed [9:0] m359_9;
   assign m359_9 =10'b0;

   // m359_10 = W*in
   wire signed [9:0] m359_10;
   assign m359_10 =10'b0;

   // m359_11 = W*in
   wire signed [9:0] m359_11;
   assign m359_11 =10'b0;

   // m359_12 = W*in
   wire signed [9:0] m359_12;
   assign m359_12 =10'b0;

   // m359_13 = W*in
   wire signed [9:0] m359_13;
   assign m359_13 =10'b0;

   // m359_14 = W*in
   wire signed [9:0] m359_14;
   assign m359_14 =10'b0;

   // m359_15 = W*in
   wire signed [9:0] m359_15;
   assign m359_15 =10'b0;

   // m359_16 = W*in
   wire signed [9:0] m359_16;
   assign m359_16 =10'b0;

   // m359_17 = W*in
   wire signed [9:0] m359_17;
   assign m359_17 =10'b0;

   // m359_18 = W*in
   wire signed [9:0] m359_18;
   assign m359_18 =10'b0;

   // m359_19 = W*in
   wire signed [9:0] m359_19;
   assign m359_19 =10'b0;

   // m359_20 = W*in
   wire signed [9:0] m359_20;
   assign m359_20 =10'b0;

   // m359_21 = W*in
   wire signed [9:0] m359_21;
   assign m359_21 =10'b0;

   // m359_22 = W*in
   wire signed [9:0] m359_22;
   assign m359_22 =10'b0;

   // m359_23 = W*in
   wire signed [9:0] m359_23;
   assign m359_23 ={ {4{in359[5]}} , in359[5:0] };

   // m359_24 = W*in
   wire signed [9:0] m359_24;
   assign m359_24 ={ {4{in359[5]}} , in359[5:0] };

   // m359_25 = W*in
   wire signed [9:0] m359_25;
   assign m359_25 =10'b0;

   // m359_26 = W*in
   wire signed [9:0] m359_26;
   assign m359_26 =10'b0;

   // m359_27 = W*in
   wire signed [9:0] m359_27;
   assign m359_27 ={ {5{in359[5]}} , in359[5:1] };

   // m359_28 = W*in
   wire signed [9:0] m359_28;
   assign m359_28 =10'b0;

   // m359_29 = W*in
   wire signed [9:0] m359_29;
   assign m359_29 =10'b0;

   // m359_30 = W*in
   wire signed [9:0] m359_30;
   assign m359_30 ={ {5{neg359[5]}} , neg359[5:1] };

   // m359_31 = W*in
   wire signed [9:0] m359_31;
   assign m359_31 =10'b0;

   // m359_32 = W*in
   wire signed [9:0] m359_32;
   assign m359_32 =10'b0;

   // m359_33 = W*in
   wire signed [9:0] m359_33;
   assign m359_33 =10'b0;

   // m359_34 = W*in
   wire signed [9:0] m359_34;
   assign m359_34 ={ {5{in359[5]}} , in359[5:1] };

   // m359_35 = W*in
   wire signed [9:0] m359_35;
   assign m359_35 ={ {5{neg359[5]}} , neg359[5:1] };

   // m359_36 = W*in
   wire signed [9:0] m359_36;
   assign m359_36 =10'b0;

   // m359_37 = W*in
   wire signed [9:0] m359_37;
   assign m359_37 =10'b0;

   // m359_38 = W*in
   wire signed [9:0] m359_38;
   assign m359_38 =10'b0;

   // m359_39 = W*in
   wire signed [9:0] m359_39;
   assign m359_39 =10'b0;

   // m359_40 = W*in
   wire signed [9:0] m359_40;
   assign m359_40 =10'b0;

   // m359_41 = W*in
   wire signed [9:0] m359_41;
   assign m359_41 =10'b0;

   // m359_42 = W*in
   wire signed [9:0] m359_42;
   assign m359_42 =10'b0;

   // m359_43 = W*in
   wire signed [9:0] m359_43;
   assign m359_43 =10'b0;

   // m359_44 = W*in
   wire signed [9:0] m359_44;
   assign m359_44 =10'b0;

   // m359_45 = W*in
   wire signed [9:0] m359_45;
   assign m359_45 =10'b0;

   // m359_46 = W*in
   wire signed [9:0] m359_46;
   assign m359_46 =10'b0;

   // m359_47 = W*in
   wire signed [9:0] m359_47;
   assign m359_47 =10'b0;

   // m359_48 = W*in
   wire signed [9:0] m359_48;
   assign m359_48 =10'b0;

   // m359_49 = W*in
   wire signed [9:0] m359_49;
   assign m359_49 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_50 = W*in
   wire signed [9:0] m359_50;
   assign m359_50 =10'b0;

   // m359_51 = W*in
   wire signed [9:0] m359_51;
   assign m359_51 =10'b0;

   // m359_52 = W*in
   wire signed [9:0] m359_52;
   assign m359_52 =10'b0;

   // m359_53 = W*in
   wire signed [9:0] m359_53;
   assign m359_53 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_54 = W*in
   wire signed [9:0] m359_54;
   assign m359_54 =10'b0;

   // m359_55 = W*in
   wire signed [9:0] m359_55;
   assign m359_55 =10'b0;

   // m359_56 = W*in
   wire signed [9:0] m359_56;
   assign m359_56 =10'b0;

   // m359_57 = W*in
   wire signed [9:0] m359_57;
   assign m359_57 =10'b0;

   // m359_58 = W*in
   wire signed [9:0] m359_58;
   assign m359_58 =10'b0;

   // m359_59 = W*in
   wire signed [9:0] m359_59;
   assign m359_59 =10'b0;

   // m359_60 = W*in
   wire signed [9:0] m359_60;
   assign m359_60 =10'b0;

   // m359_61 = W*in
   wire signed [9:0] m359_61;
   assign m359_61 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_62 = W*in
   wire signed [9:0] m359_62;
   assign m359_62 =10'b0;

   // m359_63 = W*in
   wire signed [9:0] m359_63;
   assign m359_63 ={ {4{in359[5]}} , in359[5:0] };

   // m359_64 = W*in
   wire signed [9:0] m359_64;
   assign m359_64 =10'b0;

   // m359_65 = W*in
   wire signed [9:0] m359_65;
   assign m359_65 ={ {4{in359[5]}} , in359[5:0] };

   // m359_66 = W*in
   wire signed [9:0] m359_66;
   assign m359_66 =10'b0;

   // m359_67 = W*in
   wire signed [9:0] m359_67;
   assign m359_67 ={ {5{neg359[5]}} , neg359[5:1] };

   // m359_68 = W*in
   wire signed [9:0] m359_68;
   assign m359_68 =10'b0;

   // m359_69 = W*in
   wire signed [9:0] m359_69;
   assign m359_69 =10'b0;

   // m359_70 = W*in
   wire signed [9:0] m359_70;
   assign m359_70 =10'b0;

   // m359_71 = W*in
   wire signed [9:0] m359_71;
   assign m359_71 ={ {5{in359[5]}} , in359[5:1] };

   // m359_72 = W*in
   wire signed [9:0] m359_72;
   assign m359_72 =10'b0;

   // m359_73 = W*in
   wire signed [9:0] m359_73;
   assign m359_73 =10'b0;

   // m359_74 = W*in
   wire signed [9:0] m359_74;
   assign m359_74 =10'b0;

   // m359_75 = W*in
   wire signed [9:0] m359_75;
   assign m359_75 =10'b0;

   // m359_76 = W*in
   wire signed [9:0] m359_76;
   assign m359_76 =10'b0;

   // m359_77 = W*in
   wire signed [9:0] m359_77;
   assign m359_77 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_78 = W*in
   wire signed [9:0] m359_78;
   assign m359_78 =10'b0;

   // m359_79 = W*in
   wire signed [9:0] m359_79;
   assign m359_79 =10'b0;

   // m359_80 = W*in
   wire signed [9:0] m359_80;
   assign m359_80 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_81 = W*in
   wire signed [9:0] m359_81;
   assign m359_81 =10'b0;

   // m359_82 = W*in
   wire signed [9:0] m359_82;
   assign m359_82 =10'b0;

   // m359_83 = W*in
   wire signed [9:0] m359_83;
   assign m359_83 =10'b0;

   // m359_84 = W*in
   wire signed [9:0] m359_84;
   assign m359_84 =10'b0;

   // m359_85 = W*in
   wire signed [9:0] m359_85;
   assign m359_85 =10'b0;

   // m359_86 = W*in
   wire signed [9:0] m359_86;
   assign m359_86 =10'b0;

   // m359_87 = W*in
   wire signed [9:0] m359_87;
   assign m359_87 =10'b0;

   // m359_88 = W*in
   wire signed [9:0] m359_88;
   assign m359_88 =10'b0;

   // m359_89 = W*in
   wire signed [9:0] m359_89;
   assign m359_89 =10'b0;

   // m359_90 = W*in
   wire signed [9:0] m359_90;
   assign m359_90 =10'b0;

   // m359_91 = W*in
   wire signed [9:0] m359_91;
   assign m359_91 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_92 = W*in
   wire signed [9:0] m359_92;
   assign m359_92 =10'b0;

   // m359_93 = W*in
   wire signed [9:0] m359_93;
   assign m359_93 =10'b0;

   // m359_94 = W*in
   wire signed [9:0] m359_94;
   assign m359_94 =10'b0;

   // m359_95 = W*in
   wire signed [9:0] m359_95;
   assign m359_95 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_96 = W*in
   wire signed [9:0] m359_96;
   assign m359_96 =10'b0;

   // m359_97 = W*in
   wire signed [9:0] m359_97;
   assign m359_97 ={ {4{neg359[5]}} , neg359[5:0] };

   // m359_98 = W*in
   wire signed [9:0] m359_98;
   assign m359_98 =10'b0;

   // m359_99 = W*in
   wire signed [9:0] m359_99;
   assign m359_99 =10'b0;

   // m359_100 = W*in
   wire signed [9:0] m359_100;
   assign m359_100 =10'b0;

   // m359_101 = W*in
   wire signed [9:0] m359_101;
   assign m359_101 =10'b0;

   // m359_102 = W*in
   wire signed [9:0] m359_102;
   assign m359_102 =10'b0;

   // m359_103 = W*in
   wire signed [9:0] m359_103;
   assign m359_103 =10'b0;

   // m359_104 = W*in
   wire signed [9:0] m359_104;
   assign m359_104 ={ {5{neg359[5]}} , neg359[5:1] };

   // m359_105 = W*in
   wire signed [9:0] m359_105;
   assign m359_105 =10'b0;

   // m359_106 = W*in
   wire signed [9:0] m359_106;
   assign m359_106 =10'b0;

   // m359_107 = W*in
   wire signed [9:0] m359_107;
   assign m359_107 =10'b0;

   // m359_108 = W*in
   wire signed [9:0] m359_108;
   assign m359_108 =10'b0;

   // m359_109 = W*in
   wire signed [9:0] m359_109;
   assign m359_109 ={ {4{in359[5]}} , in359[5:0] };

   // m359_110 = W*in
   wire signed [9:0] m359_110;
   assign m359_110 =10'b0;

   // m359_111 = W*in
   wire signed [9:0] m359_111;
   assign m359_111 =10'b0;

   // m359_112 = W*in
   wire signed [9:0] m359_112;
   assign m359_112 =10'b0;

   // m359_113 = W*in
   wire signed [9:0] m359_113;
   assign m359_113 =10'b0;

   // m359_114 = W*in
   wire signed [9:0] m359_114;
   assign m359_114 =10'b0;

   // m359_115 = W*in
   wire signed [9:0] m359_115;
   assign m359_115 =10'b0;

   // m359_116 = W*in
   wire signed [9:0] m359_116;
   assign m359_116 =10'b0;

   // m359_117 = W*in
   wire signed [9:0] m359_117;
   assign m359_117 =10'b0;

   // m360_1 = W*in
   wire signed [9:0] m360_1;
   assign m360_1 =10'b0;

   // m360_2 = W*in
   wire signed [9:0] m360_2;
   assign m360_2 =10'b0;

   // m360_3 = W*in
   wire signed [9:0] m360_3;
   assign m360_3 =10'b0;

   // m360_4 = W*in
   wire signed [9:0] m360_4;
   assign m360_4 =10'b0;

   // m360_5 = W*in
   wire signed [9:0] m360_5;
   assign m360_5 =10'b0;

   // m360_6 = W*in
   wire signed [9:0] m360_6;
   assign m360_6 =10'b0;

   // m360_7 = W*in
   wire signed [9:0] m360_7;
   assign m360_7 =10'b0;

   // m360_8 = W*in
   wire signed [9:0] m360_8;
   assign m360_8 =10'b0;

   // m360_9 = W*in
   wire signed [9:0] m360_9;
   assign m360_9 =10'b0;

   // m360_10 = W*in
   wire signed [9:0] m360_10;
   assign m360_10 =10'b0;

   // m360_11 = W*in
   wire signed [9:0] m360_11;
   assign m360_11 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_12 = W*in
   wire signed [9:0] m360_12;
   assign m360_12 =10'b0;

   // m360_13 = W*in
   wire signed [9:0] m360_13;
   assign m360_13 =10'b0;

   // m360_14 = W*in
   wire signed [9:0] m360_14;
   assign m360_14 =10'b0;

   // m360_15 = W*in
   wire signed [9:0] m360_15;
   assign m360_15 =10'b0;

   // m360_16 = W*in
   wire signed [9:0] m360_16;
   assign m360_16 ={ {4{in360[5]}} , in360[5:0] };

   // m360_17 = W*in
   wire signed [9:0] m360_17;
   assign m360_17 =10'b0;

   // m360_18 = W*in
   wire signed [9:0] m360_18;
   assign m360_18 =10'b0;

   // m360_19 = W*in
   wire signed [9:0] m360_19;
   assign m360_19 =10'b0;

   // m360_20 = W*in
   wire signed [9:0] m360_20;
   assign m360_20 =10'b0;

   // m360_21 = W*in
   wire signed [9:0] m360_21;
   assign m360_21 ={ {5{in360[5]}} , in360[5:1] };

   // m360_22 = W*in
   wire signed [9:0] m360_22;
   assign m360_22 =10'b0;

   // m360_23 = W*in
   wire signed [9:0] m360_23;
   assign m360_23 =10'b0;

   // m360_24 = W*in
   wire signed [9:0] m360_24;
   assign m360_24 =10'b0;

   // m360_25 = W*in
   wire signed [9:0] m360_25;
   assign m360_25 =10'b0;

   // m360_26 = W*in
   wire signed [9:0] m360_26;
   assign m360_26 =10'b0;

   // m360_27 = W*in
   wire signed [9:0] m360_27;
   assign m360_27 =10'b0;

   // m360_28 = W*in
   wire signed [9:0] m360_28;
   assign m360_28 =10'b0;

   // m360_29 = W*in
   wire signed [9:0] m360_29;
   assign m360_29 =10'b0;

   // m360_30 = W*in
   wire signed [9:0] m360_30;
   assign m360_30 =10'b0;

   // m360_31 = W*in
   wire signed [9:0] m360_31;
   assign m360_31 =10'b0;

   // m360_32 = W*in
   wire signed [9:0] m360_32;
   assign m360_32 =10'b0;

   // m360_33 = W*in
   wire signed [9:0] m360_33;
   assign m360_33 =10'b0;

   // m360_34 = W*in
   wire signed [9:0] m360_34;
   assign m360_34 =10'b0;

   // m360_35 = W*in
   wire signed [9:0] m360_35;
   assign m360_35 =10'b0;

   // m360_36 = W*in
   wire signed [9:0] m360_36;
   assign m360_36 =10'b0;

   // m360_37 = W*in
   wire signed [9:0] m360_37;
   assign m360_37 =10'b0;

   // m360_38 = W*in
   wire signed [9:0] m360_38;
   assign m360_38 =10'b0;

   // m360_39 = W*in
   wire signed [9:0] m360_39;
   assign m360_39 =10'b0;

   // m360_40 = W*in
   wire signed [9:0] m360_40;
   assign m360_40 =10'b0;

   // m360_41 = W*in
   wire signed [9:0] m360_41;
   assign m360_41 ={ {4{in360[5]}} , in360[5:0] };

   // m360_42 = W*in
   wire signed [9:0] m360_42;
   assign m360_42 =10'b0;

   // m360_43 = W*in
   wire signed [9:0] m360_43;
   assign m360_43 =10'b0;

   // m360_44 = W*in
   wire signed [9:0] m360_44;
   assign m360_44 =10'b0;

   // m360_45 = W*in
   wire signed [9:0] m360_45;
   assign m360_45 =10'b0;

   // m360_46 = W*in
   wire signed [9:0] m360_46;
   assign m360_46 =10'b0;

   // m360_47 = W*in
   wire signed [9:0] m360_47;
   assign m360_47 =10'b0;

   // m360_48 = W*in
   wire signed [9:0] m360_48;
   assign m360_48 =10'b0;

   // m360_49 = W*in
   wire signed [9:0] m360_49;
   assign m360_49 =10'b0;

   // m360_50 = W*in
   wire signed [9:0] m360_50;
   assign m360_50 =10'b0;

   // m360_51 = W*in
   wire signed [9:0] m360_51;
   assign m360_51 =10'b0;

   // m360_52 = W*in
   wire signed [9:0] m360_52;
   assign m360_52 =10'b0;

   // m360_53 = W*in
   wire signed [9:0] m360_53;
   assign m360_53 =10'b0;

   // m360_54 = W*in
   wire signed [9:0] m360_54;
   assign m360_54 =10'b0;

   // m360_55 = W*in
   wire signed [9:0] m360_55;
   assign m360_55 =10'b0;

   // m360_56 = W*in
   wire signed [9:0] m360_56;
   assign m360_56 =10'b0;

   // m360_57 = W*in
   wire signed [9:0] m360_57;
   assign m360_57 =10'b0;

   // m360_58 = W*in
   wire signed [9:0] m360_58;
   assign m360_58 =10'b0;

   // m360_59 = W*in
   wire signed [9:0] m360_59;
   assign m360_59 =10'b0;

   // m360_60 = W*in
   wire signed [9:0] m360_60;
   assign m360_60 =10'b0;

   // m360_61 = W*in
   wire signed [9:0] m360_61;
   assign m360_61 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_62 = W*in
   wire signed [9:0] m360_62;
   assign m360_62 =10'b0;

   // m360_63 = W*in
   wire signed [9:0] m360_63;
   assign m360_63 =10'b0;

   // m360_64 = W*in
   wire signed [9:0] m360_64;
   assign m360_64 =10'b0;

   // m360_65 = W*in
   wire signed [9:0] m360_65;
   assign m360_65 =10'b0;

   // m360_66 = W*in
   wire signed [9:0] m360_66;
   assign m360_66 =10'b0;

   // m360_67 = W*in
   wire signed [9:0] m360_67;
   assign m360_67 =10'b0;

   // m360_68 = W*in
   wire signed [9:0] m360_68;
   assign m360_68 =10'b0;

   // m360_69 = W*in
   wire signed [9:0] m360_69;
   assign m360_69 =10'b0;

   // m360_70 = W*in
   wire signed [9:0] m360_70;
   assign m360_70 =10'b0;

   // m360_71 = W*in
   wire signed [9:0] m360_71;
   assign m360_71 ={ {5{neg360[5]}} , neg360[5:1] };

   // m360_72 = W*in
   wire signed [9:0] m360_72;
   assign m360_72 ={ {5{in360[5]}} , in360[5:1] };

   // m360_73 = W*in
   wire signed [9:0] m360_73;
   assign m360_73 ={ {5{neg360[5]}} , neg360[5:1] };

   // m360_74 = W*in
   wire signed [9:0] m360_74;
   assign m360_74 =10'b0;

   // m360_75 = W*in
   wire signed [9:0] m360_75;
   assign m360_75 =10'b0;

   // m360_76 = W*in
   wire signed [9:0] m360_76;
   assign m360_76 =10'b0;

   // m360_77 = W*in
   wire signed [9:0] m360_77;
   assign m360_77 =10'b0;

   // m360_78 = W*in
   wire signed [9:0] m360_78;
   assign m360_78 =10'b0;

   // m360_79 = W*in
   wire signed [9:0] m360_79;
   assign m360_79 =10'b0;

   // m360_80 = W*in
   wire signed [9:0] m360_80;
   assign m360_80 =10'b0;

   // m360_81 = W*in
   wire signed [9:0] m360_81;
   assign m360_81 =10'b0;

   // m360_82 = W*in
   wire signed [9:0] m360_82;
   assign m360_82 =10'b0;

   // m360_83 = W*in
   wire signed [9:0] m360_83;
   assign m360_83 =10'b0;

   // m360_84 = W*in
   wire signed [9:0] m360_84;
   assign m360_84 =10'b0;

   // m360_85 = W*in
   wire signed [9:0] m360_85;
   assign m360_85 =10'b0;

   // m360_86 = W*in
   wire signed [9:0] m360_86;
   assign m360_86 =10'b0;

   // m360_87 = W*in
   wire signed [9:0] m360_87;
   assign m360_87 =10'b0;

   // m360_88 = W*in
   wire signed [9:0] m360_88;
   assign m360_88 =10'b0;

   // m360_89 = W*in
   wire signed [9:0] m360_89;
   assign m360_89 =10'b0;

   // m360_90 = W*in
   wire signed [9:0] m360_90;
   assign m360_90 =10'b0;

   // m360_91 = W*in
   wire signed [9:0] m360_91;
   assign m360_91 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_92 = W*in
   wire signed [9:0] m360_92;
   assign m360_92 =10'b0;

   // m360_93 = W*in
   wire signed [9:0] m360_93;
   assign m360_93 =10'b0;

   // m360_94 = W*in
   wire signed [9:0] m360_94;
   assign m360_94 =10'b0;

   // m360_95 = W*in
   wire signed [9:0] m360_95;
   assign m360_95 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_96 = W*in
   wire signed [9:0] m360_96;
   assign m360_96 =10'b0;

   // m360_97 = W*in
   wire signed [9:0] m360_97;
   assign m360_97 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_98 = W*in
   wire signed [9:0] m360_98;
   assign m360_98 =10'b0;

   // m360_99 = W*in
   wire signed [9:0] m360_99;
   assign m360_99 =10'b0;

   // m360_100 = W*in
   wire signed [9:0] m360_100;
   assign m360_100 =10'b0;

   // m360_101 = W*in
   wire signed [9:0] m360_101;
   assign m360_101 =10'b0;

   // m360_102 = W*in
   wire signed [9:0] m360_102;
   assign m360_102 =10'b0;

   // m360_103 = W*in
   wire signed [9:0] m360_103;
   assign m360_103 =10'b0;

   // m360_104 = W*in
   wire signed [9:0] m360_104;
   assign m360_104 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_105 = W*in
   wire signed [9:0] m360_105;
   assign m360_105 =10'b0;

   // m360_106 = W*in
   wire signed [9:0] m360_106;
   assign m360_106 ={ {4{in360[5]}} , in360[5:0] };

   // m360_107 = W*in
   wire signed [9:0] m360_107;
   assign m360_107 =10'b0;

   // m360_108 = W*in
   wire signed [9:0] m360_108;
   assign m360_108 ={ {4{in360[5]}} , in360[5:0] };

   // m360_109 = W*in
   wire signed [9:0] m360_109;
   assign m360_109 =10'b0;

   // m360_110 = W*in
   wire signed [9:0] m360_110;
   assign m360_110 ={ {4{neg360[5]}} , neg360[5:0] };

   // m360_111 = W*in
   wire signed [9:0] m360_111;
   assign m360_111 =10'b0;

   // m360_112 = W*in
   wire signed [9:0] m360_112;
   assign m360_112 =10'b0;

   // m360_113 = W*in
   wire signed [9:0] m360_113;
   assign m360_113 =10'b0;

   // m360_114 = W*in
   wire signed [9:0] m360_114;
   assign m360_114 =10'b0;

   // m360_115 = W*in
   wire signed [9:0] m360_115;
   assign m360_115 =10'b0;

   // m360_116 = W*in
   wire signed [9:0] m360_116;
   assign m360_116 ={ {5{in360[5]}} , in360[5:1] };

   // m360_117 = W*in
   wire signed [9:0] m360_117;
   assign m360_117 =10'b0;

   // m361_1 = W*in
   wire signed [9:0] m361_1;
   assign m361_1 =10'b0;

   // m361_2 = W*in
   wire signed [9:0] m361_2;
   assign m361_2 =10'b0;

   // m361_3 = W*in
   wire signed [9:0] m361_3;
   assign m361_3 =10'b0;

   // m361_4 = W*in
   wire signed [9:0] m361_4;
   assign m361_4 =10'b0;

   // m361_5 = W*in
   wire signed [9:0] m361_5;
   assign m361_5 =10'b0;

   // m361_6 = W*in
   wire signed [9:0] m361_6;
   assign m361_6 =10'b0;

   // m361_7 = W*in
   wire signed [9:0] m361_7;
   assign m361_7 =10'b0;

   // m361_8 = W*in
   wire signed [9:0] m361_8;
   assign m361_8 =10'b0;

   // m361_9 = W*in
   wire signed [9:0] m361_9;
   assign m361_9 =10'b0;

   // m361_10 = W*in
   wire signed [9:0] m361_10;
   assign m361_10 =10'b0;

   // m361_11 = W*in
   wire signed [9:0] m361_11;
   assign m361_11 =10'b0;

   // m361_12 = W*in
   wire signed [9:0] m361_12;
   assign m361_12 =10'b0;

   // m361_13 = W*in
   wire signed [9:0] m361_13;
   assign m361_13 =10'b0;

   // m361_14 = W*in
   wire signed [9:0] m361_14;
   assign m361_14 =10'b0;

   // m361_15 = W*in
   wire signed [9:0] m361_15;
   assign m361_15 =10'b0;

   // m361_16 = W*in
   wire signed [9:0] m361_16;
   assign m361_16 =10'b0;

   // m361_17 = W*in
   wire signed [9:0] m361_17;
   assign m361_17 =10'b0;

   // m361_18 = W*in
   wire signed [9:0] m361_18;
   assign m361_18 =10'b0;

   // m361_19 = W*in
   wire signed [9:0] m361_19;
   assign m361_19 =10'b0;

   // m361_20 = W*in
   wire signed [9:0] m361_20;
   assign m361_20 =10'b0;

   // m361_21 = W*in
   wire signed [9:0] m361_21;
   assign m361_21 ={ {5{in361[5]}} , in361[5:1] };

   // m361_22 = W*in
   wire signed [9:0] m361_22;
   assign m361_22 =10'b0;

   // m361_23 = W*in
   wire signed [9:0] m361_23;
   assign m361_23 =10'b0;

   // m361_24 = W*in
   wire signed [9:0] m361_24;
   assign m361_24 =10'b0;

   // m361_25 = W*in
   wire signed [9:0] m361_25;
   assign m361_25 ={ {5{neg361[5]}} , neg361[5:1] };

   // m361_26 = W*in
   wire signed [9:0] m361_26;
   assign m361_26 ={ {5{neg361[5]}} , neg361[5:1] };

   // m361_27 = W*in
   wire signed [9:0] m361_27;
   assign m361_27 ={ {5{neg361[5]}} , neg361[5:1] };

   // m361_28 = W*in
   wire signed [9:0] m361_28;
   assign m361_28 =10'b0;

   // m361_29 = W*in
   wire signed [9:0] m361_29;
   assign m361_29 =10'b0;

   // m361_30 = W*in
   wire signed [9:0] m361_30;
   assign m361_30 =10'b0;

   // m361_31 = W*in
   wire signed [9:0] m361_31;
   assign m361_31 =10'b0;

   // m361_32 = W*in
   wire signed [9:0] m361_32;
   assign m361_32 =10'b0;

   // m361_33 = W*in
   wire signed [9:0] m361_33;
   assign m361_33 =10'b0;

   // m361_34 = W*in
   wire signed [9:0] m361_34;
   assign m361_34 =10'b0;

   // m361_35 = W*in
   wire signed [9:0] m361_35;
   assign m361_35 =10'b0;

   // m361_36 = W*in
   wire signed [9:0] m361_36;
   assign m361_36 =10'b0;

   // m361_37 = W*in
   wire signed [9:0] m361_37;
   assign m361_37 =10'b0;

   // m361_38 = W*in
   wire signed [9:0] m361_38;
   assign m361_38 =10'b0;

   // m361_39 = W*in
   wire signed [9:0] m361_39;
   assign m361_39 =10'b0;

   // m361_40 = W*in
   wire signed [9:0] m361_40;
   assign m361_40 =10'b0;

   // m361_41 = W*in
   wire signed [9:0] m361_41;
   assign m361_41 =10'b0;

   // m361_42 = W*in
   wire signed [9:0] m361_42;
   assign m361_42 =10'b0;

   // m361_43 = W*in
   wire signed [9:0] m361_43;
   assign m361_43 =10'b0;

   // m361_44 = W*in
   wire signed [9:0] m361_44;
   assign m361_44 =10'b0;

   // m361_45 = W*in
   wire signed [9:0] m361_45;
   assign m361_45 =10'b0;

   // m361_46 = W*in
   wire signed [9:0] m361_46;
   assign m361_46 =10'b0;

   // m361_47 = W*in
   wire signed [9:0] m361_47;
   assign m361_47 =10'b0;

   // m361_48 = W*in
   wire signed [9:0] m361_48;
   assign m361_48 ={ {4{neg361[5]}} , neg361[5:0] };

   // m361_49 = W*in
   wire signed [9:0] m361_49;
   assign m361_49 =10'b0;

   // m361_50 = W*in
   wire signed [9:0] m361_50;
   assign m361_50 =10'b0;

   // m361_51 = W*in
   wire signed [9:0] m361_51;
   assign m361_51 =10'b0;

   // m361_52 = W*in
   wire signed [9:0] m361_52;
   assign m361_52 =10'b0;

   // m361_53 = W*in
   wire signed [9:0] m361_53;
   assign m361_53 =10'b0;

   // m361_54 = W*in
   wire signed [9:0] m361_54;
   assign m361_54 ={ {4{neg361[5]}} , neg361[5:0] };

   // m361_55 = W*in
   wire signed [9:0] m361_55;
   assign m361_55 =10'b0;

   // m361_56 = W*in
   wire signed [9:0] m361_56;
   assign m361_56 =10'b0;

   // m361_57 = W*in
   wire signed [9:0] m361_57;
   assign m361_57 =10'b0;

   // m361_58 = W*in
   wire signed [9:0] m361_58;
   assign m361_58 =10'b0;

   // m361_59 = W*in
   wire signed [9:0] m361_59;
   assign m361_59 =10'b0;

   // m361_60 = W*in
   wire signed [9:0] m361_60;
   assign m361_60 =10'b0;

   // m361_61 = W*in
   wire signed [9:0] m361_61;
   assign m361_61 =10'b0;

   // m361_62 = W*in
   wire signed [9:0] m361_62;
   assign m361_62 =10'b0;

   // m361_63 = W*in
   wire signed [9:0] m361_63;
   assign m361_63 ={ {5{neg361[5]}} , neg361[5:1] };

   // m361_64 = W*in
   wire signed [9:0] m361_64;
   assign m361_64 =10'b0;

   // m361_65 = W*in
   wire signed [9:0] m361_65;
   assign m361_65 ={ {5{in361[5]}} , in361[5:1] };

   // m361_66 = W*in
   wire signed [9:0] m361_66;
   assign m361_66 =10'b0;

   // m361_67 = W*in
   wire signed [9:0] m361_67;
   assign m361_67 =10'b0;

   // m361_68 = W*in
   wire signed [9:0] m361_68;
   assign m361_68 =10'b0;

   // m361_69 = W*in
   wire signed [9:0] m361_69;
   assign m361_69 =10'b0;

   // m361_70 = W*in
   wire signed [9:0] m361_70;
   assign m361_70 ={ {5{in361[5]}} , in361[5:1] };

   // m361_71 = W*in
   wire signed [9:0] m361_71;
   assign m361_71 ={ {5{neg361[5]}} , neg361[5:1] };

   // m361_72 = W*in
   wire signed [9:0] m361_72;
   assign m361_72 =10'b0;

   // m361_73 = W*in
   wire signed [9:0] m361_73;
   assign m361_73 ={ {5{neg361[5]}} , neg361[5:1] };

   // m361_74 = W*in
   wire signed [9:0] m361_74;
   assign m361_74 =10'b0;

   // m361_75 = W*in
   wire signed [9:0] m361_75;
   assign m361_75 =10'b0;

   // m361_76 = W*in
   wire signed [9:0] m361_76;
   assign m361_76 =10'b0;

   // m361_77 = W*in
   wire signed [9:0] m361_77;
   assign m361_77 =10'b0;

   // m361_78 = W*in
   wire signed [9:0] m361_78;
   assign m361_78 =10'b0;

   // m361_79 = W*in
   wire signed [9:0] m361_79;
   assign m361_79 =10'b0;

   // m361_80 = W*in
   wire signed [9:0] m361_80;
   assign m361_80 =10'b0;

   // m361_81 = W*in
   wire signed [9:0] m361_81;
   assign m361_81 =10'b0;

   // m361_82 = W*in
   wire signed [9:0] m361_82;
   assign m361_82 =10'b0;

   // m361_83 = W*in
   wire signed [9:0] m361_83;
   assign m361_83 =10'b0;

   // m361_84 = W*in
   wire signed [9:0] m361_84;
   assign m361_84 =10'b0;

   // m361_85 = W*in
   wire signed [9:0] m361_85;
   assign m361_85 =10'b0;

   // m361_86 = W*in
   wire signed [9:0] m361_86;
   assign m361_86 =10'b0;

   // m361_87 = W*in
   wire signed [9:0] m361_87;
   assign m361_87 =10'b0;

   // m361_88 = W*in
   wire signed [9:0] m361_88;
   assign m361_88 =10'b0;

   // m361_89 = W*in
   wire signed [9:0] m361_89;
   assign m361_89 =10'b0;

   // m361_90 = W*in
   wire signed [9:0] m361_90;
   assign m361_90 =10'b0;

   // m361_91 = W*in
   wire signed [9:0] m361_91;
   assign m361_91 =10'b0;

   // m361_92 = W*in
   wire signed [9:0] m361_92;
   assign m361_92 =10'b0;

   // m361_93 = W*in
   wire signed [9:0] m361_93;
   assign m361_93 =10'b0;

   // m361_94 = W*in
   wire signed [9:0] m361_94;
   assign m361_94 =10'b0;

   // m361_95 = W*in
   wire signed [9:0] m361_95;
   assign m361_95 =10'b0;

   // m361_96 = W*in
   wire signed [9:0] m361_96;
   assign m361_96 ={ {5{in361[5]}} , in361[5:1] };

   // m361_97 = W*in
   wire signed [9:0] m361_97;
   assign m361_97 =10'b0;

   // m361_98 = W*in
   wire signed [9:0] m361_98;
   assign m361_98 =10'b0;

   // m361_99 = W*in
   wire signed [9:0] m361_99;
   assign m361_99 =10'b0;

   // m361_100 = W*in
   wire signed [9:0] m361_100;
   assign m361_100 =10'b0;

   // m361_101 = W*in
   wire signed [9:0] m361_101;
   assign m361_101 =10'b0;

   // m361_102 = W*in
   wire signed [9:0] m361_102;
   assign m361_102 =10'b0;

   // m361_103 = W*in
   wire signed [9:0] m361_103;
   assign m361_103 =10'b0;

   // m361_104 = W*in
   wire signed [9:0] m361_104;
   assign m361_104 =10'b0;

   // m361_105 = W*in
   wire signed [9:0] m361_105;
   assign m361_105 =10'b0;

   // m361_106 = W*in
   wire signed [9:0] m361_106;
   assign m361_106 =10'b0;

   // m361_107 = W*in
   wire signed [9:0] m361_107;
   assign m361_107 =10'b0;

   // m361_108 = W*in
   wire signed [9:0] m361_108;
   assign m361_108 ={ {4{in361[5]}} , in361[5:0] };

   // m361_109 = W*in
   wire signed [9:0] m361_109;
   assign m361_109 ={ {4{in361[5]}} , in361[5:0] };

   // m361_110 = W*in
   wire signed [9:0] m361_110;
   assign m361_110 =10'b0;

   // m361_111 = W*in
   wire signed [9:0] m361_111;
   assign m361_111 =10'b0;

   // m361_112 = W*in
   wire signed [9:0] m361_112;
   assign m361_112 =10'b0;

   // m361_113 = W*in
   wire signed [9:0] m361_113;
   assign m361_113 =10'b0;

   // m361_114 = W*in
   wire signed [9:0] m361_114;
   assign m361_114 =10'b0;

   // m361_115 = W*in
   wire signed [9:0] m361_115;
   assign m361_115 =10'b0;

   // m361_116 = W*in
   wire signed [9:0] m361_116;
   assign m361_116 ={ {4{in361[5]}} , in361[5:0] };

   // m361_117 = W*in
   wire signed [9:0] m361_117;
   assign m361_117 =10'b0;

   // m362_1 = W*in
   wire signed [9:0] m362_1;
   assign m362_1 =10'b0;

   // m362_2 = W*in
   wire signed [9:0] m362_2;
   assign m362_2 =10'b0;

   // m362_3 = W*in
   wire signed [9:0] m362_3;
   assign m362_3 =10'b0;

   // m362_4 = W*in
   wire signed [9:0] m362_4;
   assign m362_4 =10'b0;

   // m362_5 = W*in
   wire signed [9:0] m362_5;
   assign m362_5 =10'b0;

   // m362_6 = W*in
   wire signed [9:0] m362_6;
   assign m362_6 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_7 = W*in
   wire signed [9:0] m362_7;
   assign m362_7 =10'b0;

   // m362_8 = W*in
   wire signed [9:0] m362_8;
   assign m362_8 =10'b0;

   // m362_9 = W*in
   wire signed [9:0] m362_9;
   assign m362_9 =10'b0;

   // m362_10 = W*in
   wire signed [9:0] m362_10;
   assign m362_10 =10'b0;

   // m362_11 = W*in
   wire signed [9:0] m362_11;
   assign m362_11 =10'b0;

   // m362_12 = W*in
   wire signed [9:0] m362_12;
   assign m362_12 =10'b0;

   // m362_13 = W*in
   wire signed [9:0] m362_13;
   assign m362_13 =10'b0;

   // m362_14 = W*in
   wire signed [9:0] m362_14;
   assign m362_14 =10'b0;

   // m362_15 = W*in
   wire signed [9:0] m362_15;
   assign m362_15 =10'b0;

   // m362_16 = W*in
   wire signed [9:0] m362_16;
   assign m362_16 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_17 = W*in
   wire signed [9:0] m362_17;
   assign m362_17 ={ {5{in362[5]}} , in362[5:1] };

   // m362_18 = W*in
   wire signed [9:0] m362_18;
   assign m362_18 ={ {5{neg362[5]}} , neg362[5:1] };

   // m362_19 = W*in
   wire signed [9:0] m362_19;
   assign m362_19 ={ {5{in362[5]}} , in362[5:1] };

   // m362_20 = W*in
   wire signed [9:0] m362_20;
   assign m362_20 ={ {5{neg362[5]}} , neg362[5:1] };

   // m362_21 = W*in
   wire signed [9:0] m362_21;
   assign m362_21 =10'b0;

   // m362_22 = W*in
   wire signed [9:0] m362_22;
   assign m362_22 =10'b0;

   // m362_23 = W*in
   wire signed [9:0] m362_23;
   assign m362_23 =10'b0;

   // m362_24 = W*in
   wire signed [9:0] m362_24;
   assign m362_24 =10'b0;

   // m362_25 = W*in
   wire signed [9:0] m362_25;
   assign m362_25 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_26 = W*in
   wire signed [9:0] m362_26;
   assign m362_26 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_27 = W*in
   wire signed [9:0] m362_27;
   assign m362_27 ={ {5{in362[5]}} , in362[5:1] };

   // m362_28 = W*in
   wire signed [9:0] m362_28;
   assign m362_28 =10'b0;

   // m362_29 = W*in
   wire signed [9:0] m362_29;
   assign m362_29 =10'b0;

   // m362_30 = W*in
   wire signed [9:0] m362_30;
   assign m362_30 =10'b0;

   // m362_31 = W*in
   wire signed [9:0] m362_31;
   assign m362_31 =10'b0;

   // m362_32 = W*in
   wire signed [9:0] m362_32;
   assign m362_32 =10'b0;

   // m362_33 = W*in
   wire signed [9:0] m362_33;
   assign m362_33 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_34 = W*in
   wire signed [9:0] m362_34;
   assign m362_34 =10'b0;

   // m362_35 = W*in
   wire signed [9:0] m362_35;
   assign m362_35 =10'b0;

   // m362_36 = W*in
   wire signed [9:0] m362_36;
   assign m362_36 =10'b0;

   // m362_37 = W*in
   wire signed [9:0] m362_37;
   assign m362_37 =10'b0;

   // m362_38 = W*in
   wire signed [9:0] m362_38;
   assign m362_38 =10'b0;

   // m362_39 = W*in
   wire signed [9:0] m362_39;
   assign m362_39 =10'b0;

   // m362_40 = W*in
   wire signed [9:0] m362_40;
   assign m362_40 =10'b0;

   // m362_41 = W*in
   wire signed [9:0] m362_41;
   assign m362_41 =10'b0;

   // m362_42 = W*in
   wire signed [9:0] m362_42;
   assign m362_42 =10'b0;

   // m362_43 = W*in
   wire signed [9:0] m362_43;
   assign m362_43 =10'b0;

   // m362_44 = W*in
   wire signed [9:0] m362_44;
   assign m362_44 ={ {4{in362[5]}} , in362[5:0] };

   // m362_45 = W*in
   wire signed [9:0] m362_45;
   assign m362_45 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_46 = W*in
   wire signed [9:0] m362_46;
   assign m362_46 =10'b0;

   // m362_47 = W*in
   wire signed [9:0] m362_47;
   assign m362_47 =10'b0;

   // m362_48 = W*in
   wire signed [9:0] m362_48;
   assign m362_48 =10'b0;

   // m362_49 = W*in
   wire signed [9:0] m362_49;
   assign m362_49 =10'b0;

   // m362_50 = W*in
   wire signed [9:0] m362_50;
   assign m362_50 =10'b0;

   // m362_51 = W*in
   wire signed [9:0] m362_51;
   assign m362_51 =10'b0;

   // m362_52 = W*in
   wire signed [9:0] m362_52;
   assign m362_52 =10'b0;

   // m362_53 = W*in
   wire signed [9:0] m362_53;
   assign m362_53 =10'b0;

   // m362_54 = W*in
   wire signed [9:0] m362_54;
   assign m362_54 =10'b0;

   // m362_55 = W*in
   wire signed [9:0] m362_55;
   assign m362_55 =10'b0;

   // m362_56 = W*in
   wire signed [9:0] m362_56;
   assign m362_56 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_57 = W*in
   wire signed [9:0] m362_57;
   assign m362_57 =10'b0;

   // m362_58 = W*in
   wire signed [9:0] m362_58;
   assign m362_58 =10'b0;

   // m362_59 = W*in
   wire signed [9:0] m362_59;
   assign m362_59 =10'b0;

   // m362_60 = W*in
   wire signed [9:0] m362_60;
   assign m362_60 =10'b0;

   // m362_61 = W*in
   wire signed [9:0] m362_61;
   assign m362_61 =10'b0;

   // m362_62 = W*in
   wire signed [9:0] m362_62;
   assign m362_62 =10'b0;

   // m362_63 = W*in
   wire signed [9:0] m362_63;
   assign m362_63 =10'b0;

   // m362_64 = W*in
   wire signed [9:0] m362_64;
   assign m362_64 ={ {5{neg362[5]}} , neg362[5:1] };

   // m362_65 = W*in
   wire signed [9:0] m362_65;
   assign m362_65 =10'b0;

   // m362_66 = W*in
   wire signed [9:0] m362_66;
   assign m362_66 ={ {5{in362[5]}} , in362[5:1] };

   // m362_67 = W*in
   wire signed [9:0] m362_67;
   assign m362_67 =10'b0;

   // m362_68 = W*in
   wire signed [9:0] m362_68;
   assign m362_68 =10'b0;

   // m362_69 = W*in
   wire signed [9:0] m362_69;
   assign m362_69 =10'b0;

   // m362_70 = W*in
   wire signed [9:0] m362_70;
   assign m362_70 =10'b0;

   // m362_71 = W*in
   wire signed [9:0] m362_71;
   assign m362_71 =10'b0;

   // m362_72 = W*in
   wire signed [9:0] m362_72;
   assign m362_72 ={ {5{neg362[5]}} , neg362[5:1] };

   // m362_73 = W*in
   wire signed [9:0] m362_73;
   assign m362_73 =10'b0;

   // m362_74 = W*in
   wire signed [9:0] m362_74;
   assign m362_74 =10'b0;

   // m362_75 = W*in
   wire signed [9:0] m362_75;
   assign m362_75 =10'b0;

   // m362_76 = W*in
   wire signed [9:0] m362_76;
   assign m362_76 =10'b0;

   // m362_77 = W*in
   wire signed [9:0] m362_77;
   assign m362_77 =10'b0;

   // m362_78 = W*in
   wire signed [9:0] m362_78;
   assign m362_78 =10'b0;

   // m362_79 = W*in
   wire signed [9:0] m362_79;
   assign m362_79 =10'b0;

   // m362_80 = W*in
   wire signed [9:0] m362_80;
   assign m362_80 ={ {5{in362[5]}} , in362[5:1] };

   // m362_81 = W*in
   wire signed [9:0] m362_81;
   assign m362_81 ={ {5{neg362[5]}} , neg362[5:1] };

   // m362_82 = W*in
   wire signed [9:0] m362_82;
   assign m362_82 =10'b0;

   // m362_83 = W*in
   wire signed [9:0] m362_83;
   assign m362_83 =10'b0;

   // m362_84 = W*in
   wire signed [9:0] m362_84;
   assign m362_84 =10'b0;

   // m362_85 = W*in
   wire signed [9:0] m362_85;
   assign m362_85 =10'b0;

   // m362_86 = W*in
   wire signed [9:0] m362_86;
   assign m362_86 =10'b0;

   // m362_87 = W*in
   wire signed [9:0] m362_87;
   assign m362_87 =10'b0;

   // m362_88 = W*in
   wire signed [9:0] m362_88;
   assign m362_88 =10'b0;

   // m362_89 = W*in
   wire signed [9:0] m362_89;
   assign m362_89 =10'b0;

   // m362_90 = W*in
   wire signed [9:0] m362_90;
   assign m362_90 =10'b0;

   // m362_91 = W*in
   wire signed [9:0] m362_91;
   assign m362_91 =10'b0;

   // m362_92 = W*in
   wire signed [9:0] m362_92;
   assign m362_92 =10'b0;

   // m362_93 = W*in
   wire signed [9:0] m362_93;
   assign m362_93 =10'b0;

   // m362_94 = W*in
   wire signed [9:0] m362_94;
   assign m362_94 =10'b0;

   // m362_95 = W*in
   wire signed [9:0] m362_95;
   assign m362_95 =10'b0;

   // m362_96 = W*in
   wire signed [9:0] m362_96;
   assign m362_96 =10'b0;

   // m362_97 = W*in
   wire signed [9:0] m362_97;
   assign m362_97 =10'b0;

   // m362_98 = W*in
   wire signed [9:0] m362_98;
   assign m362_98 =10'b0;

   // m362_99 = W*in
   wire signed [9:0] m362_99;
   assign m362_99 =10'b0;

   // m362_100 = W*in
   wire signed [9:0] m362_100;
   assign m362_100 =10'b0;

   // m362_101 = W*in
   wire signed [9:0] m362_101;
   assign m362_101 =10'b0;

   // m362_102 = W*in
   wire signed [9:0] m362_102;
   assign m362_102 ={ {4{neg362[5]}} , neg362[5:0] };

   // m362_103 = W*in
   wire signed [9:0] m362_103;
   assign m362_103 =10'b0;

   // m362_104 = W*in
   wire signed [9:0] m362_104;
   assign m362_104 =10'b0;

   // m362_105 = W*in
   wire signed [9:0] m362_105;
   assign m362_105 =10'b0;

   // m362_106 = W*in
   wire signed [9:0] m362_106;
   assign m362_106 ={ {5{neg362[5]}} , neg362[5:1] };

   // m362_107 = W*in
   wire signed [9:0] m362_107;
   assign m362_107 =10'b0;

   // m362_108 = W*in
   wire signed [9:0] m362_108;
   assign m362_108 =10'b0;

   // m362_109 = W*in
   wire signed [9:0] m362_109;
   assign m362_109 =10'b0;

   // m362_110 = W*in
   wire signed [9:0] m362_110;
   assign m362_110 =10'b0;

   // m362_111 = W*in
   wire signed [9:0] m362_111;
   assign m362_111 =10'b0;

   // m362_112 = W*in
   wire signed [9:0] m362_112;
   assign m362_112 =10'b0;

   // m362_113 = W*in
   wire signed [9:0] m362_113;
   assign m362_113 =10'b0;

   // m362_114 = W*in
   wire signed [9:0] m362_114;
   assign m362_114 =10'b0;

   // m362_115 = W*in
   wire signed [9:0] m362_115;
   assign m362_115 =10'b0;

   // m362_116 = W*in
   wire signed [9:0] m362_116;
   assign m362_116 =10'b0;

   // m362_117 = W*in
   wire signed [9:0] m362_117;
   assign m362_117 =10'b0;

   // m363_1 = W*in
   wire signed [9:0] m363_1;
   assign m363_1 =10'b0;

   // m363_2 = W*in
   wire signed [9:0] m363_2;
   assign m363_2 ={ {4{in363[5]}} , in363[5:0] };

   // m363_3 = W*in
   wire signed [9:0] m363_3;
   assign m363_3 =10'b0;

   // m363_4 = W*in
   wire signed [9:0] m363_4;
   assign m363_4 =10'b0;

   // m363_5 = W*in
   wire signed [9:0] m363_5;
   assign m363_5 =10'b0;

   // m363_6 = W*in
   wire signed [9:0] m363_6;
   assign m363_6 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_7 = W*in
   wire signed [9:0] m363_7;
   assign m363_7 =10'b0;

   // m363_8 = W*in
   wire signed [9:0] m363_8;
   assign m363_8 =10'b0;

   // m363_9 = W*in
   wire signed [9:0] m363_9;
   assign m363_9 =10'b0;

   // m363_10 = W*in
   wire signed [9:0] m363_10;
   assign m363_10 =10'b0;

   // m363_11 = W*in
   wire signed [9:0] m363_11;
   assign m363_11 =10'b0;

   // m363_12 = W*in
   wire signed [9:0] m363_12;
   assign m363_12 ={ {4{in363[5]}} , in363[5:0] };

   // m363_13 = W*in
   wire signed [9:0] m363_13;
   assign m363_13 =10'b0;

   // m363_14 = W*in
   wire signed [9:0] m363_14;
   assign m363_14 =10'b0;

   // m363_15 = W*in
   wire signed [9:0] m363_15;
   assign m363_15 =10'b0;

   // m363_16 = W*in
   wire signed [9:0] m363_16;
   assign m363_16 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_17 = W*in
   wire signed [9:0] m363_17;
   assign m363_17 ={ {4{in363[5]}} , in363[5:0] };

   // m363_18 = W*in
   wire signed [9:0] m363_18;
   assign m363_18 =10'b0;

   // m363_19 = W*in
   wire signed [9:0] m363_19;
   assign m363_19 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_20 = W*in
   wire signed [9:0] m363_20;
   assign m363_20 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_21 = W*in
   wire signed [9:0] m363_21;
   assign m363_21 =10'b0;

   // m363_22 = W*in
   wire signed [9:0] m363_22;
   assign m363_22 =10'b0;

   // m363_23 = W*in
   wire signed [9:0] m363_23;
   assign m363_23 =10'b0;

   // m363_24 = W*in
   wire signed [9:0] m363_24;
   assign m363_24 =10'b0;

   // m363_25 = W*in
   wire signed [9:0] m363_25;
   assign m363_25 =10'b0;

   // m363_26 = W*in
   wire signed [9:0] m363_26;
   assign m363_26 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_27 = W*in
   wire signed [9:0] m363_27;
   assign m363_27 ={ {4{in363[5]}} , in363[5:0] };

   // m363_28 = W*in
   wire signed [9:0] m363_28;
   assign m363_28 =10'b0;

   // m363_29 = W*in
   wire signed [9:0] m363_29;
   assign m363_29 =10'b0;

   // m363_30 = W*in
   wire signed [9:0] m363_30;
   assign m363_30 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_31 = W*in
   wire signed [9:0] m363_31;
   assign m363_31 =10'b0;

   // m363_32 = W*in
   wire signed [9:0] m363_32;
   assign m363_32 =10'b0;

   // m363_33 = W*in
   wire signed [9:0] m363_33;
   assign m363_33 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_34 = W*in
   wire signed [9:0] m363_34;
   assign m363_34 =10'b0;

   // m363_35 = W*in
   wire signed [9:0] m363_35;
   assign m363_35 =10'b0;

   // m363_36 = W*in
   wire signed [9:0] m363_36;
   assign m363_36 =10'b0;

   // m363_37 = W*in
   wire signed [9:0] m363_37;
   assign m363_37 =10'b0;

   // m363_38 = W*in
   wire signed [9:0] m363_38;
   assign m363_38 =10'b0;

   // m363_39 = W*in
   wire signed [9:0] m363_39;
   assign m363_39 =10'b0;

   // m363_40 = W*in
   wire signed [9:0] m363_40;
   assign m363_40 =10'b0;

   // m363_41 = W*in
   wire signed [9:0] m363_41;
   assign m363_41 =10'b0;

   // m363_42 = W*in
   wire signed [9:0] m363_42;
   assign m363_42 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_43 = W*in
   wire signed [9:0] m363_43;
   assign m363_43 =10'b0;

   // m363_44 = W*in
   wire signed [9:0] m363_44;
   assign m363_44 =10'b0;

   // m363_45 = W*in
   wire signed [9:0] m363_45;
   assign m363_45 =10'b0;

   // m363_46 = W*in
   wire signed [9:0] m363_46;
   assign m363_46 =10'b0;

   // m363_47 = W*in
   wire signed [9:0] m363_47;
   assign m363_47 =10'b0;

   // m363_48 = W*in
   wire signed [9:0] m363_48;
   assign m363_48 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_49 = W*in
   wire signed [9:0] m363_49;
   assign m363_49 =10'b0;

   // m363_50 = W*in
   wire signed [9:0] m363_50;
   assign m363_50 =10'b0;

   // m363_51 = W*in
   wire signed [9:0] m363_51;
   assign m363_51 ={ {4{in363[5]}} , in363[5:0] };

   // m363_52 = W*in
   wire signed [9:0] m363_52;
   assign m363_52 ={ {4{in363[5]}} , in363[5:0] };

   // m363_53 = W*in
   wire signed [9:0] m363_53;
   assign m363_53 =10'b0;

   // m363_54 = W*in
   wire signed [9:0] m363_54;
   assign m363_54 =10'b0;

   // m363_55 = W*in
   wire signed [9:0] m363_55;
   assign m363_55 =10'b0;

   // m363_56 = W*in
   wire signed [9:0] m363_56;
   assign m363_56 =10'b0;

   // m363_57 = W*in
   wire signed [9:0] m363_57;
   assign m363_57 =10'b0;

   // m363_58 = W*in
   wire signed [9:0] m363_58;
   assign m363_58 =10'b0;

   // m363_59 = W*in
   wire signed [9:0] m363_59;
   assign m363_59 =10'b0;

   // m363_60 = W*in
   wire signed [9:0] m363_60;
   assign m363_60 ={ {4{in363[5]}} , in363[5:0] };

   // m363_61 = W*in
   wire signed [9:0] m363_61;
   assign m363_61 =10'b0;

   // m363_62 = W*in
   wire signed [9:0] m363_62;
   assign m363_62 =10'b0;

   // m363_63 = W*in
   wire signed [9:0] m363_63;
   assign m363_63 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_64 = W*in
   wire signed [9:0] m363_64;
   assign m363_64 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_65 = W*in
   wire signed [9:0] m363_65;
   assign m363_65 =10'b0;

   // m363_66 = W*in
   wire signed [9:0] m363_66;
   assign m363_66 =10'b0;

   // m363_67 = W*in
   wire signed [9:0] m363_67;
   assign m363_67 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_68 = W*in
   wire signed [9:0] m363_68;
   assign m363_68 ={ {4{in363[5]}} , in363[5:0] };

   // m363_69 = W*in
   wire signed [9:0] m363_69;
   assign m363_69 =10'b0;

   // m363_70 = W*in
   wire signed [9:0] m363_70;
   assign m363_70 =10'b0;

   // m363_71 = W*in
   wire signed [9:0] m363_71;
   assign m363_71 ={ {5{in363[5]}} , in363[5:1] };

   // m363_72 = W*in
   wire signed [9:0] m363_72;
   assign m363_72 =10'b0;

   // m363_73 = W*in
   wire signed [9:0] m363_73;
   assign m363_73 =10'b0;

   // m363_74 = W*in
   wire signed [9:0] m363_74;
   assign m363_74 =10'b0;

   // m363_75 = W*in
   wire signed [9:0] m363_75;
   assign m363_75 =10'b0;

   // m363_76 = W*in
   wire signed [9:0] m363_76;
   assign m363_76 =10'b0;

   // m363_77 = W*in
   wire signed [9:0] m363_77;
   assign m363_77 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_78 = W*in
   wire signed [9:0] m363_78;
   assign m363_78 =10'b0;

   // m363_79 = W*in
   wire signed [9:0] m363_79;
   assign m363_79 =10'b0;

   // m363_80 = W*in
   wire signed [9:0] m363_80;
   assign m363_80 ={ {5{in363[5]}} , in363[5:1] };

   // m363_81 = W*in
   wire signed [9:0] m363_81;
   assign m363_81 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_82 = W*in
   wire signed [9:0] m363_82;
   assign m363_82 =10'b0;

   // m363_83 = W*in
   wire signed [9:0] m363_83;
   assign m363_83 =10'b0;

   // m363_84 = W*in
   wire signed [9:0] m363_84;
   assign m363_84 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_85 = W*in
   wire signed [9:0] m363_85;
   assign m363_85 ={ {4{in363[5]}} , in363[5:0] };

   // m363_86 = W*in
   wire signed [9:0] m363_86;
   assign m363_86 =10'b0;

   // m363_87 = W*in
   wire signed [9:0] m363_87;
   assign m363_87 =10'b0;

   // m363_88 = W*in
   wire signed [9:0] m363_88;
   assign m363_88 =10'b0;

   // m363_89 = W*in
   wire signed [9:0] m363_89;
   assign m363_89 =10'b0;

   // m363_90 = W*in
   wire signed [9:0] m363_90;
   assign m363_90 =10'b0;

   // m363_91 = W*in
   wire signed [9:0] m363_91;
   assign m363_91 =10'b0;

   // m363_92 = W*in
   wire signed [9:0] m363_92;
   assign m363_92 =10'b0;

   // m363_93 = W*in
   wire signed [9:0] m363_93;
   assign m363_93 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_94 = W*in
   wire signed [9:0] m363_94;
   assign m363_94 =10'b0;

   // m363_95 = W*in
   wire signed [9:0] m363_95;
   assign m363_95 ={ {4{in363[5]}} , in363[5:0] };

   // m363_96 = W*in
   wire signed [9:0] m363_96;
   assign m363_96 =10'b0;

   // m363_97 = W*in
   wire signed [9:0] m363_97;
   assign m363_97 =10'b0;

   // m363_98 = W*in
   wire signed [9:0] m363_98;
   assign m363_98 =10'b0;

   // m363_99 = W*in
   wire signed [9:0] m363_99;
   assign m363_99 =10'b0;

   // m363_100 = W*in
   wire signed [9:0] m363_100;
   assign m363_100 =10'b0;

   // m363_101 = W*in
   wire signed [9:0] m363_101;
   assign m363_101 =10'b0;

   // m363_102 = W*in
   wire signed [9:0] m363_102;
   assign m363_102 ={ {4{neg363[5]}} , neg363[5:0] };

   // m363_103 = W*in
   wire signed [9:0] m363_103;
   assign m363_103 =10'b0;

   // m363_104 = W*in
   wire signed [9:0] m363_104;
   assign m363_104 ={ {4{in363[5]}} , in363[5:0] };

   // m363_105 = W*in
   wire signed [9:0] m363_105;
   assign m363_105 =10'b0;

   // m363_106 = W*in
   wire signed [9:0] m363_106;
   assign m363_106 ={ {5{neg363[5]}} , neg363[5:1] };

   // m363_107 = W*in
   wire signed [9:0] m363_107;
   assign m363_107 ={ {5{in363[5]}} , in363[5:1] };

   // m363_108 = W*in
   wire signed [9:0] m363_108;
   assign m363_108 =10'b0;

   // m363_109 = W*in
   wire signed [9:0] m363_109;
   assign m363_109 =10'b0;

   // m363_110 = W*in
   wire signed [9:0] m363_110;
   assign m363_110 =10'b0;

   // m363_111 = W*in
   wire signed [9:0] m363_111;
   assign m363_111 =10'b0;

   // m363_112 = W*in
   wire signed [9:0] m363_112;
   assign m363_112 =10'b0;

   // m363_113 = W*in
   wire signed [9:0] m363_113;
   assign m363_113 =10'b0;

   // m363_114 = W*in
   wire signed [9:0] m363_114;
   assign m363_114 =10'b0;

   // m363_115 = W*in
   wire signed [9:0] m363_115;
   assign m363_115 =10'b0;

   // m363_116 = W*in
   wire signed [9:0] m363_116;
   assign m363_116 =10'b0;

   // m363_117 = W*in
   wire signed [9:0] m363_117;
   assign m363_117 =10'b0;

   // m364_1 = W*in
   wire signed [9:0] m364_1;
   assign m364_1 =10'b0;

   // m364_2 = W*in
   wire signed [9:0] m364_2;
   assign m364_2 =10'b0;

   // m364_3 = W*in
   wire signed [9:0] m364_3;
   assign m364_3 =10'b0;

   // m364_4 = W*in
   wire signed [9:0] m364_4;
   assign m364_4 =10'b0;

   // m364_5 = W*in
   wire signed [9:0] m364_5;
   assign m364_5 =10'b0;

   // m364_6 = W*in
   wire signed [9:0] m364_6;
   assign m364_6 =10'b0;

   // m364_7 = W*in
   wire signed [9:0] m364_7;
   assign m364_7 =10'b0;

   // m364_8 = W*in
   wire signed [9:0] m364_8;
   assign m364_8 =10'b0;

   // m364_9 = W*in
   wire signed [9:0] m364_9;
   assign m364_9 =10'b0;

   // m364_10 = W*in
   wire signed [9:0] m364_10;
   assign m364_10 =10'b0;

   // m364_11 = W*in
   wire signed [9:0] m364_11;
   assign m364_11 =10'b0;

   // m364_12 = W*in
   wire signed [9:0] m364_12;
   assign m364_12 =10'b0;

   // m364_13 = W*in
   wire signed [9:0] m364_13;
   assign m364_13 ={ {4{in364[5]}} , in364[5:0] };

   // m364_14 = W*in
   wire signed [9:0] m364_14;
   assign m364_14 =10'b0;

   // m364_15 = W*in
   wire signed [9:0] m364_15;
   assign m364_15 ={ {4{in364[5]}} , in364[5:0] };

   // m364_16 = W*in
   wire signed [9:0] m364_16;
   assign m364_16 =10'b0;

   // m364_17 = W*in
   wire signed [9:0] m364_17;
   assign m364_17 ={ {5{in364[5]}} , in364[5:1] };

   // m364_18 = W*in
   wire signed [9:0] m364_18;
   assign m364_18 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_19 = W*in
   wire signed [9:0] m364_19;
   assign m364_19 =10'b0;

   // m364_20 = W*in
   wire signed [9:0] m364_20;
   assign m364_20 ={ {4{in364[5]}} , in364[5:0] };

   // m364_21 = W*in
   wire signed [9:0] m364_21;
   assign m364_21 =10'b0;

   // m364_22 = W*in
   wire signed [9:0] m364_22;
   assign m364_22 =10'b0;

   // m364_23 = W*in
   wire signed [9:0] m364_23;
   assign m364_23 =10'b0;

   // m364_24 = W*in
   wire signed [9:0] m364_24;
   assign m364_24 =10'b0;

   // m364_25 = W*in
   wire signed [9:0] m364_25;
   assign m364_25 ={ {5{in364[5]}} , in364[5:1] };

   // m364_26 = W*in
   wire signed [9:0] m364_26;
   assign m364_26 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_27 = W*in
   wire signed [9:0] m364_27;
   assign m364_27 =10'b0;

   // m364_28 = W*in
   wire signed [9:0] m364_28;
   assign m364_28 ={ {5{in364[5]}} , in364[5:1] };

   // m364_29 = W*in
   wire signed [9:0] m364_29;
   assign m364_29 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_30 = W*in
   wire signed [9:0] m364_30;
   assign m364_30 ={ {4{in364[5]}} , in364[5:0] };

   // m364_31 = W*in
   wire signed [9:0] m364_31;
   assign m364_31 =10'b0;

   // m364_32 = W*in
   wire signed [9:0] m364_32;
   assign m364_32 =10'b0;

   // m364_33 = W*in
   wire signed [9:0] m364_33;
   assign m364_33 =10'b0;

   // m364_34 = W*in
   wire signed [9:0] m364_34;
   assign m364_34 ={ {5{neg364[5]}} , neg364[5:1] };

   // m364_35 = W*in
   wire signed [9:0] m364_35;
   assign m364_35 ={ {4{in364[5]}} , in364[5:0] };

   // m364_36 = W*in
   wire signed [9:0] m364_36;
   assign m364_36 =10'b0;

   // m364_37 = W*in
   wire signed [9:0] m364_37;
   assign m364_37 ={ {4{in364[5]}} , in364[5:0] };

   // m364_38 = W*in
   wire signed [9:0] m364_38;
   assign m364_38 =10'b0;

   // m364_39 = W*in
   wire signed [9:0] m364_39;
   assign m364_39 =10'b0;

   // m364_40 = W*in
   wire signed [9:0] m364_40;
   assign m364_40 =10'b0;

   // m364_41 = W*in
   wire signed [9:0] m364_41;
   assign m364_41 ={ {4{in364[5]}} , in364[5:0] };

   // m364_42 = W*in
   wire signed [9:0] m364_42;
   assign m364_42 =10'b0;

   // m364_43 = W*in
   wire signed [9:0] m364_43;
   assign m364_43 =10'b0;

   // m364_44 = W*in
   wire signed [9:0] m364_44;
   assign m364_44 =10'b0;

   // m364_45 = W*in
   wire signed [9:0] m364_45;
   assign m364_45 =10'b0;

   // m364_46 = W*in
   wire signed [9:0] m364_46;
   assign m364_46 =10'b0;

   // m364_47 = W*in
   wire signed [9:0] m364_47;
   assign m364_47 =10'b0;

   // m364_48 = W*in
   wire signed [9:0] m364_48;
   assign m364_48 =10'b0;

   // m364_49 = W*in
   wire signed [9:0] m364_49;
   assign m364_49 =10'b0;

   // m364_50 = W*in
   wire signed [9:0] m364_50;
   assign m364_50 =10'b0;

   // m364_51 = W*in
   wire signed [9:0] m364_51;
   assign m364_51 =10'b0;

   // m364_52 = W*in
   wire signed [9:0] m364_52;
   assign m364_52 =10'b0;

   // m364_53 = W*in
   wire signed [9:0] m364_53;
   assign m364_53 =10'b0;

   // m364_54 = W*in
   wire signed [9:0] m364_54;
   assign m364_54 =10'b0;

   // m364_55 = W*in
   wire signed [9:0] m364_55;
   assign m364_55 =10'b0;

   // m364_56 = W*in
   wire signed [9:0] m364_56;
   assign m364_56 =10'b0;

   // m364_57 = W*in
   wire signed [9:0] m364_57;
   assign m364_57 =10'b0;

   // m364_58 = W*in
   wire signed [9:0] m364_58;
   assign m364_58 =10'b0;

   // m364_59 = W*in
   wire signed [9:0] m364_59;
   assign m364_59 =10'b0;

   // m364_60 = W*in
   wire signed [9:0] m364_60;
   assign m364_60 ={ {4{in364[5]}} , in364[5:0] };

   // m364_61 = W*in
   wire signed [9:0] m364_61;
   assign m364_61 ={ {4{in364[5]}} , in364[5:0] };

   // m364_62 = W*in
   wire signed [9:0] m364_62;
   assign m364_62 =10'b0;

   // m364_63 = W*in
   wire signed [9:0] m364_63;
   assign m364_63 =10'b0;

   // m364_64 = W*in
   wire signed [9:0] m364_64;
   assign m364_64 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_65 = W*in
   wire signed [9:0] m364_65;
   assign m364_65 ={ {5{neg364[5]}} , neg364[5:1] };

   // m364_66 = W*in
   wire signed [9:0] m364_66;
   assign m364_66 =10'b0;

   // m364_67 = W*in
   wire signed [9:0] m364_67;
   assign m364_67 =10'b0;

   // m364_68 = W*in
   wire signed [9:0] m364_68;
   assign m364_68 =10'b0;

   // m364_69 = W*in
   wire signed [9:0] m364_69;
   assign m364_69 =10'b0;

   // m364_70 = W*in
   wire signed [9:0] m364_70;
   assign m364_70 =10'b0;

   // m364_71 = W*in
   wire signed [9:0] m364_71;
   assign m364_71 =10'b0;

   // m364_72 = W*in
   wire signed [9:0] m364_72;
   assign m364_72 =10'b0;

   // m364_73 = W*in
   wire signed [9:0] m364_73;
   assign m364_73 =10'b0;

   // m364_74 = W*in
   wire signed [9:0] m364_74;
   assign m364_74 =10'b0;

   // m364_75 = W*in
   wire signed [9:0] m364_75;
   assign m364_75 =10'b0;

   // m364_76 = W*in
   wire signed [9:0] m364_76;
   assign m364_76 =10'b0;

   // m364_77 = W*in
   wire signed [9:0] m364_77;
   assign m364_77 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_78 = W*in
   wire signed [9:0] m364_78;
   assign m364_78 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_79 = W*in
   wire signed [9:0] m364_79;
   assign m364_79 ={ {4{in364[5]}} , in364[5:0] };

   // m364_80 = W*in
   wire signed [9:0] m364_80;
   assign m364_80 ={ {5{neg364[5]}} , neg364[5:1] };

   // m364_81 = W*in
   wire signed [9:0] m364_81;
   assign m364_81 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_82 = W*in
   wire signed [9:0] m364_82;
   assign m364_82 =10'b0;

   // m364_83 = W*in
   wire signed [9:0] m364_83;
   assign m364_83 ={ {5{in364[5]}} , in364[5:1] };

   // m364_84 = W*in
   wire signed [9:0] m364_84;
   assign m364_84 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_85 = W*in
   wire signed [9:0] m364_85;
   assign m364_85 ={ {4{in364[5]}} , in364[5:0] };

   // m364_86 = W*in
   wire signed [9:0] m364_86;
   assign m364_86 =10'b0;

   // m364_87 = W*in
   wire signed [9:0] m364_87;
   assign m364_87 =10'b0;

   // m364_88 = W*in
   wire signed [9:0] m364_88;
   assign m364_88 ={ {4{in364[5]}} , in364[5:0] };

   // m364_89 = W*in
   wire signed [9:0] m364_89;
   assign m364_89 ={ {4{in364[5]}} , in364[5:0] };

   // m364_90 = W*in
   wire signed [9:0] m364_90;
   assign m364_90 =10'b0;

   // m364_91 = W*in
   wire signed [9:0] m364_91;
   assign m364_91 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_92 = W*in
   wire signed [9:0] m364_92;
   assign m364_92 =10'b0;

   // m364_93 = W*in
   wire signed [9:0] m364_93;
   assign m364_93 =10'b0;

   // m364_94 = W*in
   wire signed [9:0] m364_94;
   assign m364_94 =10'b0;

   // m364_95 = W*in
   wire signed [9:0] m364_95;
   assign m364_95 ={ {4{in364[5]}} , in364[5:0] };

   // m364_96 = W*in
   wire signed [9:0] m364_96;
   assign m364_96 ={ {4{in364[5]}} , in364[5:0] };

   // m364_97 = W*in
   wire signed [9:0] m364_97;
   assign m364_97 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_98 = W*in
   wire signed [9:0] m364_98;
   assign m364_98 =10'b0;

   // m364_99 = W*in
   wire signed [9:0] m364_99;
   assign m364_99 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_100 = W*in
   wire signed [9:0] m364_100;
   assign m364_100 ={ {4{in364[5]}} , in364[5:0] };

   // m364_101 = W*in
   wire signed [9:0] m364_101;
   assign m364_101 =10'b0;

   // m364_102 = W*in
   wire signed [9:0] m364_102;
   assign m364_102 =10'b0;

   // m364_103 = W*in
   wire signed [9:0] m364_103;
   assign m364_103 =10'b0;

   // m364_104 = W*in
   wire signed [9:0] m364_104;
   assign m364_104 =10'b0;

   // m364_105 = W*in
   wire signed [9:0] m364_105;
   assign m364_105 =10'b0;

   // m364_106 = W*in
   wire signed [9:0] m364_106;
   assign m364_106 =10'b0;

   // m364_107 = W*in
   wire signed [9:0] m364_107;
   assign m364_107 =10'b0;

   // m364_108 = W*in
   wire signed [9:0] m364_108;
   assign m364_108 ={ {4{in364[5]}} , in364[5:0] };

   // m364_109 = W*in
   wire signed [9:0] m364_109;
   assign m364_109 ={ {3{in364[5]}} , in364 , {1{1'b0}} };

   // m364_110 = W*in
   wire signed [9:0] m364_110;
   assign m364_110 =10'b0;

   // m364_111 = W*in
   wire signed [9:0] m364_111;
   assign m364_111 ={ {4{neg364[5]}} , neg364[5:0] };

   // m364_112 = W*in
   wire signed [9:0] m364_112;
   assign m364_112 =10'b0;

   // m364_113 = W*in
   wire signed [9:0] m364_113;
   assign m364_113 =10'b0;

   // m364_114 = W*in
   wire signed [9:0] m364_114;
   assign m364_114 =10'b0;

   // m364_115 = W*in
   wire signed [9:0] m364_115;
   assign m364_115 ={ {5{in364[5]}} , in364[5:1] };

   // m364_116 = W*in
   wire signed [9:0] m364_116;
   assign m364_116 ={ {4{in364[5]}} , in364[5:0] };

   // m364_117 = W*in
   wire signed [9:0] m364_117;
   assign m364_117 ={ {4{in364[5]}} , in364[5:0] };

   // m365_1 = W*in
   wire signed [9:0] m365_1;
   assign m365_1 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_2 = W*in
   wire signed [9:0] m365_2;
   assign m365_2 =10'b0;

   // m365_3 = W*in
   wire signed [9:0] m365_3;
   assign m365_3 =10'b0;

   // m365_4 = W*in
   wire signed [9:0] m365_4;
   assign m365_4 =10'b0;

   // m365_5 = W*in
   wire signed [9:0] m365_5;
   assign m365_5 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_6 = W*in
   wire signed [9:0] m365_6;
   assign m365_6 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_7 = W*in
   wire signed [9:0] m365_7;
   assign m365_7 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_8 = W*in
   wire signed [9:0] m365_8;
   assign m365_8 =10'b0;

   // m365_9 = W*in
   wire signed [9:0] m365_9;
   assign m365_9 =10'b0;

   // m365_10 = W*in
   wire signed [9:0] m365_10;
   assign m365_10 =10'b0;

   // m365_11 = W*in
   wire signed [9:0] m365_11;
   assign m365_11 =10'b0;

   // m365_12 = W*in
   wire signed [9:0] m365_12;
   assign m365_12 =10'b0;

   // m365_13 = W*in
   wire signed [9:0] m365_13;
   assign m365_13 =10'b0;

   // m365_14 = W*in
   wire signed [9:0] m365_14;
   assign m365_14 =10'b0;

   // m365_15 = W*in
   wire signed [9:0] m365_15;
   assign m365_15 ={ {4{in365[5]}} , in365[5:0] };

   // m365_16 = W*in
   wire signed [9:0] m365_16;
   assign m365_16 =10'b0;

   // m365_17 = W*in
   wire signed [9:0] m365_17;
   assign m365_17 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_18 = W*in
   wire signed [9:0] m365_18;
   assign m365_18 =10'b0;

   // m365_19 = W*in
   wire signed [9:0] m365_19;
   assign m365_19 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_20 = W*in
   wire signed [9:0] m365_20;
   assign m365_20 =10'b0;

   // m365_21 = W*in
   wire signed [9:0] m365_21;
   assign m365_21 ={ {5{in365[5]}} , in365[5:1] };

   // m365_22 = W*in
   wire signed [9:0] m365_22;
   assign m365_22 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_23 = W*in
   wire signed [9:0] m365_23;
   assign m365_23 =10'b0;

   // m365_24 = W*in
   wire signed [9:0] m365_24;
   assign m365_24 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_25 = W*in
   wire signed [9:0] m365_25;
   assign m365_25 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_26 = W*in
   wire signed [9:0] m365_26;
   assign m365_26 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_27 = W*in
   wire signed [9:0] m365_27;
   assign m365_27 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_28 = W*in
   wire signed [9:0] m365_28;
   assign m365_28 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_29 = W*in
   wire signed [9:0] m365_29;
   assign m365_29 =10'b0;

   // m365_30 = W*in
   wire signed [9:0] m365_30;
   assign m365_30 ={ {3{in365[5]}} , in365 , {1{1'b0}} };

   // m365_31 = W*in
   wire signed [9:0] m365_31;
   assign m365_31 =10'b0;

   // m365_32 = W*in
   wire signed [9:0] m365_32;
   assign m365_32 =10'b0;

   // m365_33 = W*in
   wire signed [9:0] m365_33;
   assign m365_33 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_34 = W*in
   wire signed [9:0] m365_34;
   assign m365_34 =10'b0;

   // m365_35 = W*in
   wire signed [9:0] m365_35;
   assign m365_35 =10'b0;

   // m365_36 = W*in
   wire signed [9:0] m365_36;
   assign m365_36 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_37 = W*in
   wire signed [9:0] m365_37;
   assign m365_37 ={ {4{in365[5]}} , in365[5:0] };

   // m365_38 = W*in
   wire signed [9:0] m365_38;
   assign m365_38 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_39 = W*in
   wire signed [9:0] m365_39;
   assign m365_39 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_40 = W*in
   wire signed [9:0] m365_40;
   assign m365_40 =10'b0;

   // m365_41 = W*in
   wire signed [9:0] m365_41;
   assign m365_41 ={ {4{in365[5]}} , in365[5:0] };

   // m365_42 = W*in
   wire signed [9:0] m365_42;
   assign m365_42 =10'b0;

   // m365_43 = W*in
   wire signed [9:0] m365_43;
   assign m365_43 =10'b0;

   // m365_44 = W*in
   wire signed [9:0] m365_44;
   assign m365_44 =10'b0;

   // m365_45 = W*in
   wire signed [9:0] m365_45;
   assign m365_45 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_46 = W*in
   wire signed [9:0] m365_46;
   assign m365_46 =10'b0;

   // m365_47 = W*in
   wire signed [9:0] m365_47;
   assign m365_47 =10'b0;

   // m365_48 = W*in
   wire signed [9:0] m365_48;
   assign m365_48 =10'b0;

   // m365_49 = W*in
   wire signed [9:0] m365_49;
   assign m365_49 =10'b0;

   // m365_50 = W*in
   wire signed [9:0] m365_50;
   assign m365_50 ={ {4{in365[5]}} , in365[5:0] };

   // m365_51 = W*in
   wire signed [9:0] m365_51;
   assign m365_51 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_52 = W*in
   wire signed [9:0] m365_52;
   assign m365_52 =10'b0;

   // m365_53 = W*in
   wire signed [9:0] m365_53;
   assign m365_53 =10'b0;

   // m365_54 = W*in
   wire signed [9:0] m365_54;
   assign m365_54 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_55 = W*in
   wire signed [9:0] m365_55;
   assign m365_55 =10'b0;

   // m365_56 = W*in
   wire signed [9:0] m365_56;
   assign m365_56 =10'b0;

   // m365_57 = W*in
   wire signed [9:0] m365_57;
   assign m365_57 =10'b0;

   // m365_58 = W*in
   wire signed [9:0] m365_58;
   assign m365_58 =10'b0;

   // m365_59 = W*in
   wire signed [9:0] m365_59;
   assign m365_59 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_60 = W*in
   wire signed [9:0] m365_60;
   assign m365_60 =10'b0;

   // m365_61 = W*in
   wire signed [9:0] m365_61;
   assign m365_61 ={ {4{in365[5]}} , in365[5:0] };

   // m365_62 = W*in
   wire signed [9:0] m365_62;
   assign m365_62 =10'b0;

   // m365_63 = W*in
   wire signed [9:0] m365_63;
   assign m365_63 ={ {5{in365[5]}} , in365[5:1] };

   // m365_64 = W*in
   wire signed [9:0] m365_64;
   assign m365_64 =10'b0;

   // m365_65 = W*in
   wire signed [9:0] m365_65;
   assign m365_65 =10'b0;

   // m365_66 = W*in
   wire signed [9:0] m365_66;
   assign m365_66 ={ {4{in365[5]}} , in365[5:0] };

   // m365_67 = W*in
   wire signed [9:0] m365_67;
   assign m365_67 =10'b0;

   // m365_68 = W*in
   wire signed [9:0] m365_68;
   assign m365_68 =10'b0;

   // m365_69 = W*in
   wire signed [9:0] m365_69;
   assign m365_69 ={ {4{in365[5]}} , in365[5:0] };

   // m365_70 = W*in
   wire signed [9:0] m365_70;
   assign m365_70 ={ {4{in365[5]}} , in365[5:0] };

   // m365_71 = W*in
   wire signed [9:0] m365_71;
   assign m365_71 =10'b0;

   // m365_72 = W*in
   wire signed [9:0] m365_72;
   assign m365_72 ={ {4{in365[5]}} , in365[5:0] };

   // m365_73 = W*in
   wire signed [9:0] m365_73;
   assign m365_73 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_74 = W*in
   wire signed [9:0] m365_74;
   assign m365_74 =10'b0;

   // m365_75 = W*in
   wire signed [9:0] m365_75;
   assign m365_75 =10'b0;

   // m365_76 = W*in
   wire signed [9:0] m365_76;
   assign m365_76 =10'b0;

   // m365_77 = W*in
   wire signed [9:0] m365_77;
   assign m365_77 =10'b0;

   // m365_78 = W*in
   wire signed [9:0] m365_78;
   assign m365_78 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_79 = W*in
   wire signed [9:0] m365_79;
   assign m365_79 ={ {4{in365[5]}} , in365[5:0] };

   // m365_80 = W*in
   wire signed [9:0] m365_80;
   assign m365_80 =10'b0;

   // m365_81 = W*in
   wire signed [9:0] m365_81;
   assign m365_81 =10'b0;

   // m365_82 = W*in
   wire signed [9:0] m365_82;
   assign m365_82 ={ {4{in365[5]}} , in365[5:0] };

   // m365_83 = W*in
   wire signed [9:0] m365_83;
   assign m365_83 =10'b0;

   // m365_84 = W*in
   wire signed [9:0] m365_84;
   assign m365_84 =10'b0;

   // m365_85 = W*in
   wire signed [9:0] m365_85;
   assign m365_85 =10'b0;

   // m365_86 = W*in
   wire signed [9:0] m365_86;
   assign m365_86 ={ {4{in365[5]}} , in365[5:0] };

   // m365_87 = W*in
   wire signed [9:0] m365_87;
   assign m365_87 =10'b0;

   // m365_88 = W*in
   wire signed [9:0] m365_88;
   assign m365_88 ={ {3{in365[5]}} , in365 , {1{1'b0}} };

   // m365_89 = W*in
   wire signed [9:0] m365_89;
   assign m365_89 =10'b0;

   // m365_90 = W*in
   wire signed [9:0] m365_90;
   assign m365_90 =10'b0;

   // m365_91 = W*in
   wire signed [9:0] m365_91;
   assign m365_91 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_92 = W*in
   wire signed [9:0] m365_92;
   assign m365_92 ={ {3{in365[5]}} , in365 , {1{1'b0}} };

   // m365_93 = W*in
   wire signed [9:0] m365_93;
   assign m365_93 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_94 = W*in
   wire signed [9:0] m365_94;
   assign m365_94 ={ {4{in365[5]}} , in365[5:0] };

   // m365_95 = W*in
   wire signed [9:0] m365_95;
   assign m365_95 =10'b0;

   // m365_96 = W*in
   wire signed [9:0] m365_96;
   assign m365_96 ={ {4{in365[5]}} , in365[5:0] };

   // m365_97 = W*in
   wire signed [9:0] m365_97;
   assign m365_97 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_98 = W*in
   wire signed [9:0] m365_98;
   assign m365_98 =10'b0;

   // m365_99 = W*in
   wire signed [9:0] m365_99;
   assign m365_99 =10'b0;

   // m365_100 = W*in
   wire signed [9:0] m365_100;
   assign m365_100 ={ {4{in365[5]}} , in365[5:0] };

   // m365_101 = W*in
   wire signed [9:0] m365_101;
   assign m365_101 =10'b0;

   // m365_102 = W*in
   wire signed [9:0] m365_102;
   assign m365_102 =10'b0;

   // m365_103 = W*in
   wire signed [9:0] m365_103;
   assign m365_103 =10'b0;

   // m365_104 = W*in
   wire signed [9:0] m365_104;
   assign m365_104 =10'b0;

   // m365_105 = W*in
   wire signed [9:0] m365_105;
   assign m365_105 =10'b0;

   // m365_106 = W*in
   wire signed [9:0] m365_106;
   assign m365_106 =10'b0;

   // m365_107 = W*in
   wire signed [9:0] m365_107;
   assign m365_107 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_108 = W*in
   wire signed [9:0] m365_108;
   assign m365_108 ={ {4{in365[5]}} , in365[5:0] };

   // m365_109 = W*in
   wire signed [9:0] m365_109;
   assign m365_109 ={ {3{in365[5]}} , in365 , {1{1'b0}} };

   // m365_110 = W*in
   wire signed [9:0] m365_110;
   assign m365_110 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_111 = W*in
   wire signed [9:0] m365_111;
   assign m365_111 =10'b0;

   // m365_112 = W*in
   wire signed [9:0] m365_112;
   assign m365_112 =10'b0;

   // m365_113 = W*in
   wire signed [9:0] m365_113;
   assign m365_113 ={ {4{in365[5]}} , in365[5:0] };

   // m365_114 = W*in
   wire signed [9:0] m365_114;
   assign m365_114 ={ {4{neg365[5]}} , neg365[5:0] };

   // m365_115 = W*in
   wire signed [9:0] m365_115;
   assign m365_115 ={ {5{neg365[5]}} , neg365[5:1] };

   // m365_116 = W*in
   wire signed [9:0] m365_116;
   assign m365_116 ={ {4{in365[5]}} , in365[5:0] };

   // m365_117 = W*in
   wire signed [9:0] m365_117;
   assign m365_117 =10'b0;

   // m366_1 = W*in
   wire signed [9:0] m366_1;
   assign m366_1 =10'b0;

   // m366_2 = W*in
   wire signed [9:0] m366_2;
   assign m366_2 =10'b0;

   // m366_3 = W*in
   wire signed [9:0] m366_3;
   assign m366_3 =10'b0;

   // m366_4 = W*in
   wire signed [9:0] m366_4;
   assign m366_4 =10'b0;

   // m366_5 = W*in
   wire signed [9:0] m366_5;
   assign m366_5 =10'b0;

   // m366_6 = W*in
   wire signed [9:0] m366_6;
   assign m366_6 ={ {4{neg366[5]}} , neg366[5:0] };

   // m366_7 = W*in
   wire signed [9:0] m366_7;
   assign m366_7 =10'b0;

   // m366_8 = W*in
   wire signed [9:0] m366_8;
   assign m366_8 =10'b0;

   // m366_9 = W*in
   wire signed [9:0] m366_9;
   assign m366_9 =10'b0;

   // m366_10 = W*in
   wire signed [9:0] m366_10;
   assign m366_10 =10'b0;

   // m366_11 = W*in
   wire signed [9:0] m366_11;
   assign m366_11 =10'b0;

   // m366_12 = W*in
   wire signed [9:0] m366_12;
   assign m366_12 =10'b0;

   // m366_13 = W*in
   wire signed [9:0] m366_13;
   assign m366_13 =10'b0;

   // m366_14 = W*in
   wire signed [9:0] m366_14;
   assign m366_14 =10'b0;

   // m366_15 = W*in
   wire signed [9:0] m366_15;
   assign m366_15 =10'b0;

   // m366_16 = W*in
   wire signed [9:0] m366_16;
   assign m366_16 ={ {4{in366[5]}} , in366[5:0] };

   // m366_17 = W*in
   wire signed [9:0] m366_17;
   assign m366_17 ={ {4{neg366[5]}} , neg366[5:0] };

   // m366_18 = W*in
   wire signed [9:0] m366_18;
   assign m366_18 =10'b0;

   // m366_19 = W*in
   wire signed [9:0] m366_19;
   assign m366_19 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_20 = W*in
   wire signed [9:0] m366_20;
   assign m366_20 =10'b0;

   // m366_21 = W*in
   wire signed [9:0] m366_21;
   assign m366_21 ={ {4{in366[5]}} , in366[5:0] };

   // m366_22 = W*in
   wire signed [9:0] m366_22;
   assign m366_22 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_23 = W*in
   wire signed [9:0] m366_23;
   assign m366_23 =10'b0;

   // m366_24 = W*in
   wire signed [9:0] m366_24;
   assign m366_24 =10'b0;

   // m366_25 = W*in
   wire signed [9:0] m366_25;
   assign m366_25 =10'b0;

   // m366_26 = W*in
   wire signed [9:0] m366_26;
   assign m366_26 =10'b0;

   // m366_27 = W*in
   wire signed [9:0] m366_27;
   assign m366_27 ={ {4{neg366[5]}} , neg366[5:0] };

   // m366_28 = W*in
   wire signed [9:0] m366_28;
   assign m366_28 =10'b0;

   // m366_29 = W*in
   wire signed [9:0] m366_29;
   assign m366_29 =10'b0;

   // m366_30 = W*in
   wire signed [9:0] m366_30;
   assign m366_30 ={ {4{in366[5]}} , in366[5:0] };

   // m366_31 = W*in
   wire signed [9:0] m366_31;
   assign m366_31 =10'b0;

   // m366_32 = W*in
   wire signed [9:0] m366_32;
   assign m366_32 =10'b0;

   // m366_33 = W*in
   wire signed [9:0] m366_33;
   assign m366_33 =10'b0;

   // m366_34 = W*in
   wire signed [9:0] m366_34;
   assign m366_34 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_35 = W*in
   wire signed [9:0] m366_35;
   assign m366_35 =10'b0;

   // m366_36 = W*in
   wire signed [9:0] m366_36;
   assign m366_36 =10'b0;

   // m366_37 = W*in
   wire signed [9:0] m366_37;
   assign m366_37 ={ {4{in366[5]}} , in366[5:0] };

   // m366_38 = W*in
   wire signed [9:0] m366_38;
   assign m366_38 ={ {4{neg366[5]}} , neg366[5:0] };

   // m366_39 = W*in
   wire signed [9:0] m366_39;
   assign m366_39 =10'b0;

   // m366_40 = W*in
   wire signed [9:0] m366_40;
   assign m366_40 =10'b0;

   // m366_41 = W*in
   wire signed [9:0] m366_41;
   assign m366_41 ={ {4{in366[5]}} , in366[5:0] };

   // m366_42 = W*in
   wire signed [9:0] m366_42;
   assign m366_42 =10'b0;

   // m366_43 = W*in
   wire signed [9:0] m366_43;
   assign m366_43 =10'b0;

   // m366_44 = W*in
   wire signed [9:0] m366_44;
   assign m366_44 =10'b0;

   // m366_45 = W*in
   wire signed [9:0] m366_45;
   assign m366_45 =10'b0;

   // m366_46 = W*in
   wire signed [9:0] m366_46;
   assign m366_46 =10'b0;

   // m366_47 = W*in
   wire signed [9:0] m366_47;
   assign m366_47 =10'b0;

   // m366_48 = W*in
   wire signed [9:0] m366_48;
   assign m366_48 =10'b0;

   // m366_49 = W*in
   wire signed [9:0] m366_49;
   assign m366_49 =10'b0;

   // m366_50 = W*in
   wire signed [9:0] m366_50;
   assign m366_50 =10'b0;

   // m366_51 = W*in
   wire signed [9:0] m366_51;
   assign m366_51 =10'b0;

   // m366_52 = W*in
   wire signed [9:0] m366_52;
   assign m366_52 =10'b0;

   // m366_53 = W*in
   wire signed [9:0] m366_53;
   assign m366_53 =10'b0;

   // m366_54 = W*in
   wire signed [9:0] m366_54;
   assign m366_54 ={ {4{neg366[5]}} , neg366[5:0] };

   // m366_55 = W*in
   wire signed [9:0] m366_55;
   assign m366_55 =10'b0;

   // m366_56 = W*in
   wire signed [9:0] m366_56;
   assign m366_56 =10'b0;

   // m366_57 = W*in
   wire signed [9:0] m366_57;
   assign m366_57 =10'b0;

   // m366_58 = W*in
   wire signed [9:0] m366_58;
   assign m366_58 =10'b0;

   // m366_59 = W*in
   wire signed [9:0] m366_59;
   assign m366_59 =10'b0;

   // m366_60 = W*in
   wire signed [9:0] m366_60;
   assign m366_60 =10'b0;

   // m366_61 = W*in
   wire signed [9:0] m366_61;
   assign m366_61 ={ {4{in366[5]}} , in366[5:0] };

   // m366_62 = W*in
   wire signed [9:0] m366_62;
   assign m366_62 =10'b0;

   // m366_63 = W*in
   wire signed [9:0] m366_63;
   assign m366_63 =10'b0;

   // m366_64 = W*in
   wire signed [9:0] m366_64;
   assign m366_64 =10'b0;

   // m366_65 = W*in
   wire signed [9:0] m366_65;
   assign m366_65 ={ {5{in366[5]}} , in366[5:1] };

   // m366_66 = W*in
   wire signed [9:0] m366_66;
   assign m366_66 ={ {5{in366[5]}} , in366[5:1] };

   // m366_67 = W*in
   wire signed [9:0] m366_67;
   assign m366_67 ={ {4{neg366[5]}} , neg366[5:0] };

   // m366_68 = W*in
   wire signed [9:0] m366_68;
   assign m366_68 =10'b0;

   // m366_69 = W*in
   wire signed [9:0] m366_69;
   assign m366_69 ={ {4{in366[5]}} , in366[5:0] };

   // m366_70 = W*in
   wire signed [9:0] m366_70;
   assign m366_70 ={ {4{in366[5]}} , in366[5:0] };

   // m366_71 = W*in
   wire signed [9:0] m366_71;
   assign m366_71 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_72 = W*in
   wire signed [9:0] m366_72;
   assign m366_72 ={ {5{in366[5]}} , in366[5:1] };

   // m366_73 = W*in
   wire signed [9:0] m366_73;
   assign m366_73 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_74 = W*in
   wire signed [9:0] m366_74;
   assign m366_74 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_75 = W*in
   wire signed [9:0] m366_75;
   assign m366_75 =10'b0;

   // m366_76 = W*in
   wire signed [9:0] m366_76;
   assign m366_76 =10'b0;

   // m366_77 = W*in
   wire signed [9:0] m366_77;
   assign m366_77 =10'b0;

   // m366_78 = W*in
   wire signed [9:0] m366_78;
   assign m366_78 =10'b0;

   // m366_79 = W*in
   wire signed [9:0] m366_79;
   assign m366_79 =10'b0;

   // m366_80 = W*in
   wire signed [9:0] m366_80;
   assign m366_80 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_81 = W*in
   wire signed [9:0] m366_81;
   assign m366_81 =10'b0;

   // m366_82 = W*in
   wire signed [9:0] m366_82;
   assign m366_82 ={ {4{in366[5]}} , in366[5:0] };

   // m366_83 = W*in
   wire signed [9:0] m366_83;
   assign m366_83 =10'b0;

   // m366_84 = W*in
   wire signed [9:0] m366_84;
   assign m366_84 ={ {5{in366[5]}} , in366[5:1] };

   // m366_85 = W*in
   wire signed [9:0] m366_85;
   assign m366_85 =10'b0;

   // m366_86 = W*in
   wire signed [9:0] m366_86;
   assign m366_86 ={ {4{in366[5]}} , in366[5:0] };

   // m366_87 = W*in
   wire signed [9:0] m366_87;
   assign m366_87 =10'b0;

   // m366_88 = W*in
   wire signed [9:0] m366_88;
   assign m366_88 =10'b0;

   // m366_89 = W*in
   wire signed [9:0] m366_89;
   assign m366_89 =10'b0;

   // m366_90 = W*in
   wire signed [9:0] m366_90;
   assign m366_90 =10'b0;

   // m366_91 = W*in
   wire signed [9:0] m366_91;
   assign m366_91 =10'b0;

   // m366_92 = W*in
   wire signed [9:0] m366_92;
   assign m366_92 =10'b0;

   // m366_93 = W*in
   wire signed [9:0] m366_93;
   assign m366_93 =10'b0;

   // m366_94 = W*in
   wire signed [9:0] m366_94;
   assign m366_94 ={ {4{in366[5]}} , in366[5:0] };

   // m366_95 = W*in
   wire signed [9:0] m366_95;
   assign m366_95 =10'b0;

   // m366_96 = W*in
   wire signed [9:0] m366_96;
   assign m366_96 ={ {4{in366[5]}} , in366[5:0] };

   // m366_97 = W*in
   wire signed [9:0] m366_97;
   assign m366_97 =10'b0;

   // m366_98 = W*in
   wire signed [9:0] m366_98;
   assign m366_98 =10'b0;

   // m366_99 = W*in
   wire signed [9:0] m366_99;
   assign m366_99 =10'b0;

   // m366_100 = W*in
   wire signed [9:0] m366_100;
   assign m366_100 ={ {4{in366[5]}} , in366[5:0] };

   // m366_101 = W*in
   wire signed [9:0] m366_101;
   assign m366_101 =10'b0;

   // m366_102 = W*in
   wire signed [9:0] m366_102;
   assign m366_102 =10'b0;

   // m366_103 = W*in
   wire signed [9:0] m366_103;
   assign m366_103 =10'b0;

   // m366_104 = W*in
   wire signed [9:0] m366_104;
   assign m366_104 =10'b0;

   // m366_105 = W*in
   wire signed [9:0] m366_105;
   assign m366_105 =10'b0;

   // m366_106 = W*in
   wire signed [9:0] m366_106;
   assign m366_106 ={ {5{in366[5]}} , in366[5:1] };

   // m366_107 = W*in
   wire signed [9:0] m366_107;
   assign m366_107 ={ {5{neg366[5]}} , neg366[5:1] };

   // m366_108 = W*in
   wire signed [9:0] m366_108;
   assign m366_108 ={ {4{in366[5]}} , in366[5:0] };

   // m366_109 = W*in
   wire signed [9:0] m366_109;
   assign m366_109 =10'b0;

   // m366_110 = W*in
   wire signed [9:0] m366_110;
   assign m366_110 ={ {3{neg366[5]}} , neg366 , {1{1'b0}} };

   // m366_111 = W*in
   wire signed [9:0] m366_111;
   assign m366_111 =10'b0;

   // m366_112 = W*in
   wire signed [9:0] m366_112;
   assign m366_112 =10'b0;

   // m366_113 = W*in
   wire signed [9:0] m366_113;
   assign m366_113 =10'b0;

   // m366_114 = W*in
   wire signed [9:0] m366_114;
   assign m366_114 =10'b0;

   // m366_115 = W*in
   wire signed [9:0] m366_115;
   assign m366_115 =10'b0;

   // m366_116 = W*in
   wire signed [9:0] m366_116;
   assign m366_116 ={ {4{in366[5]}} , in366[5:0] };

   // m366_117 = W*in
   wire signed [9:0] m366_117;
   assign m366_117 =10'b0;

   // m367_1 = W*in
   wire signed [9:0] m367_1;
   assign m367_1 =10'b0;

   // m367_2 = W*in
   wire signed [9:0] m367_2;
   assign m367_2 =10'b0;

   // m367_3 = W*in
   wire signed [9:0] m367_3;
   assign m367_3 =10'b0;

   // m367_4 = W*in
   wire signed [9:0] m367_4;
   assign m367_4 =10'b0;

   // m367_5 = W*in
   wire signed [9:0] m367_5;
   assign m367_5 ={ {4{in367[5]}} , in367[5:0] };

   // m367_6 = W*in
   wire signed [9:0] m367_6;
   assign m367_6 =10'b0;

   // m367_7 = W*in
   wire signed [9:0] m367_7;
   assign m367_7 =10'b0;

   // m367_8 = W*in
   wire signed [9:0] m367_8;
   assign m367_8 =10'b0;

   // m367_9 = W*in
   wire signed [9:0] m367_9;
   assign m367_9 =10'b0;

   // m367_10 = W*in
   wire signed [9:0] m367_10;
   assign m367_10 =10'b0;

   // m367_11 = W*in
   wire signed [9:0] m367_11;
   assign m367_11 =10'b0;

   // m367_12 = W*in
   wire signed [9:0] m367_12;
   assign m367_12 =10'b0;

   // m367_13 = W*in
   wire signed [9:0] m367_13;
   assign m367_13 =10'b0;

   // m367_14 = W*in
   wire signed [9:0] m367_14;
   assign m367_14 =10'b0;

   // m367_15 = W*in
   wire signed [9:0] m367_15;
   assign m367_15 =10'b0;

   // m367_16 = W*in
   wire signed [9:0] m367_16;
   assign m367_16 =10'b0;

   // m367_17 = W*in
   wire signed [9:0] m367_17;
   assign m367_17 ={ {5{in367[5]}} , in367[5:1] };

   // m367_18 = W*in
   wire signed [9:0] m367_18;
   assign m367_18 ={ {4{neg367[5]}} , neg367[5:0] };

   // m367_19 = W*in
   wire signed [9:0] m367_19;
   assign m367_19 ={ {4{in367[5]}} , in367[5:0] };

   // m367_20 = W*in
   wire signed [9:0] m367_20;
   assign m367_20 ={ {5{neg367[5]}} , neg367[5:1] };

   // m367_21 = W*in
   wire signed [9:0] m367_21;
   assign m367_21 =10'b0;

   // m367_22 = W*in
   wire signed [9:0] m367_22;
   assign m367_22 =10'b0;

   // m367_23 = W*in
   wire signed [9:0] m367_23;
   assign m367_23 =10'b0;

   // m367_24 = W*in
   wire signed [9:0] m367_24;
   assign m367_24 =10'b0;

   // m367_25 = W*in
   wire signed [9:0] m367_25;
   assign m367_25 =10'b0;

   // m367_26 = W*in
   wire signed [9:0] m367_26;
   assign m367_26 ={ {5{neg367[5]}} , neg367[5:1] };

   // m367_27 = W*in
   wire signed [9:0] m367_27;
   assign m367_27 =10'b0;

   // m367_28 = W*in
   wire signed [9:0] m367_28;
   assign m367_28 =10'b0;

   // m367_29 = W*in
   wire signed [9:0] m367_29;
   assign m367_29 =10'b0;

   // m367_30 = W*in
   wire signed [9:0] m367_30;
   assign m367_30 =10'b0;

   // m367_31 = W*in
   wire signed [9:0] m367_31;
   assign m367_31 =10'b0;

   // m367_32 = W*in
   wire signed [9:0] m367_32;
   assign m367_32 =10'b0;

   // m367_33 = W*in
   wire signed [9:0] m367_33;
   assign m367_33 =10'b0;

   // m367_34 = W*in
   wire signed [9:0] m367_34;
   assign m367_34 ={ {5{neg367[5]}} , neg367[5:1] };

   // m367_35 = W*in
   wire signed [9:0] m367_35;
   assign m367_35 =10'b0;

   // m367_36 = W*in
   wire signed [9:0] m367_36;
   assign m367_36 =10'b0;

   // m367_37 = W*in
   wire signed [9:0] m367_37;
   assign m367_37 ={ {4{in367[5]}} , in367[5:0] };

   // m367_38 = W*in
   wire signed [9:0] m367_38;
   assign m367_38 =10'b0;

   // m367_39 = W*in
   wire signed [9:0] m367_39;
   assign m367_39 =10'b0;

   // m367_40 = W*in
   wire signed [9:0] m367_40;
   assign m367_40 =10'b0;

   // m367_41 = W*in
   wire signed [9:0] m367_41;
   assign m367_41 ={ {4{in367[5]}} , in367[5:0] };

   // m367_42 = W*in
   wire signed [9:0] m367_42;
   assign m367_42 ={ {4{neg367[5]}} , neg367[5:0] };

   // m367_43 = W*in
   wire signed [9:0] m367_43;
   assign m367_43 =10'b0;

   // m367_44 = W*in
   wire signed [9:0] m367_44;
   assign m367_44 =10'b0;

   // m367_45 = W*in
   wire signed [9:0] m367_45;
   assign m367_45 =10'b0;

   // m367_46 = W*in
   wire signed [9:0] m367_46;
   assign m367_46 =10'b0;

   // m367_47 = W*in
   wire signed [9:0] m367_47;
   assign m367_47 =10'b0;

   // m367_48 = W*in
   wire signed [9:0] m367_48;
   assign m367_48 =10'b0;

   // m367_49 = W*in
   wire signed [9:0] m367_49;
   assign m367_49 =10'b0;

   // m367_50 = W*in
   wire signed [9:0] m367_50;
   assign m367_50 =10'b0;

   // m367_51 = W*in
   wire signed [9:0] m367_51;
   assign m367_51 =10'b0;

   // m367_52 = W*in
   wire signed [9:0] m367_52;
   assign m367_52 =10'b0;

   // m367_53 = W*in
   wire signed [9:0] m367_53;
   assign m367_53 =10'b0;

   // m367_54 = W*in
   wire signed [9:0] m367_54;
   assign m367_54 =10'b0;

   // m367_55 = W*in
   wire signed [9:0] m367_55;
   assign m367_55 =10'b0;

   // m367_56 = W*in
   wire signed [9:0] m367_56;
   assign m367_56 =10'b0;

   // m367_57 = W*in
   wire signed [9:0] m367_57;
   assign m367_57 =10'b0;

   // m367_58 = W*in
   wire signed [9:0] m367_58;
   assign m367_58 =10'b0;

   // m367_59 = W*in
   wire signed [9:0] m367_59;
   assign m367_59 =10'b0;

   // m367_60 = W*in
   wire signed [9:0] m367_60;
   assign m367_60 =10'b0;

   // m367_61 = W*in
   wire signed [9:0] m367_61;
   assign m367_61 ={ {4{in367[5]}} , in367[5:0] };

   // m367_62 = W*in
   wire signed [9:0] m367_62;
   assign m367_62 =10'b0;

   // m367_63 = W*in
   wire signed [9:0] m367_63;
   assign m367_63 ={ {4{in367[5]}} , in367[5:0] };

   // m367_64 = W*in
   wire signed [9:0] m367_64;
   assign m367_64 ={ {4{neg367[5]}} , neg367[5:0] };

   // m367_65 = W*in
   wire signed [9:0] m367_65;
   assign m367_65 =10'b0;

   // m367_66 = W*in
   wire signed [9:0] m367_66;
   assign m367_66 =10'b0;

   // m367_67 = W*in
   wire signed [9:0] m367_67;
   assign m367_67 =10'b0;

   // m367_68 = W*in
   wire signed [9:0] m367_68;
   assign m367_68 =10'b0;

   // m367_69 = W*in
   wire signed [9:0] m367_69;
   assign m367_69 ={ {4{in367[5]}} , in367[5:0] };

   // m367_70 = W*in
   wire signed [9:0] m367_70;
   assign m367_70 =10'b0;

   // m367_71 = W*in
   wire signed [9:0] m367_71;
   assign m367_71 =10'b0;

   // m367_72 = W*in
   wire signed [9:0] m367_72;
   assign m367_72 =10'b0;

   // m367_73 = W*in
   wire signed [9:0] m367_73;
   assign m367_73 ={ {5{in367[5]}} , in367[5:1] };

   // m367_74 = W*in
   wire signed [9:0] m367_74;
   assign m367_74 ={ {4{neg367[5]}} , neg367[5:0] };

   // m367_75 = W*in
   wire signed [9:0] m367_75;
   assign m367_75 =10'b0;

   // m367_76 = W*in
   wire signed [9:0] m367_76;
   assign m367_76 ={ {4{neg367[5]}} , neg367[5:0] };

   // m367_77 = W*in
   wire signed [9:0] m367_77;
   assign m367_77 =10'b0;

   // m367_78 = W*in
   wire signed [9:0] m367_78;
   assign m367_78 =10'b0;

   // m367_79 = W*in
   wire signed [9:0] m367_79;
   assign m367_79 =10'b0;

   // m367_80 = W*in
   wire signed [9:0] m367_80;
   assign m367_80 ={ {5{in367[5]}} , in367[5:1] };

   // m367_81 = W*in
   wire signed [9:0] m367_81;
   assign m367_81 ={ {4{neg367[5]}} , neg367[5:0] };

   // m367_82 = W*in
   wire signed [9:0] m367_82;
   assign m367_82 ={ {4{in367[5]}} , in367[5:0] };

   // m367_83 = W*in
   wire signed [9:0] m367_83;
   assign m367_83 =10'b0;

   // m367_84 = W*in
   wire signed [9:0] m367_84;
   assign m367_84 =10'b0;

   // m367_85 = W*in
   wire signed [9:0] m367_85;
   assign m367_85 ={ {3{in367[5]}} , in367 , {1{1'b0}} };

   // m367_86 = W*in
   wire signed [9:0] m367_86;
   assign m367_86 =10'b0;

   // m367_87 = W*in
   wire signed [9:0] m367_87;
   assign m367_87 =10'b0;

   // m367_88 = W*in
   wire signed [9:0] m367_88;
   assign m367_88 =10'b0;

   // m367_89 = W*in
   wire signed [9:0] m367_89;
   assign m367_89 =10'b0;

   // m367_90 = W*in
   wire signed [9:0] m367_90;
   assign m367_90 =10'b0;

   // m367_91 = W*in
   wire signed [9:0] m367_91;
   assign m367_91 =10'b0;

   // m367_92 = W*in
   wire signed [9:0] m367_92;
   assign m367_92 =10'b0;

   // m367_93 = W*in
   wire signed [9:0] m367_93;
   assign m367_93 ={ {4{in367[5]}} , in367[5:0] };

   // m367_94 = W*in
   wire signed [9:0] m367_94;
   assign m367_94 =10'b0;

   // m367_95 = W*in
   wire signed [9:0] m367_95;
   assign m367_95 =10'b0;

   // m367_96 = W*in
   wire signed [9:0] m367_96;
   assign m367_96 =10'b0;

   // m367_97 = W*in
   wire signed [9:0] m367_97;
   assign m367_97 =10'b0;

   // m367_98 = W*in
   wire signed [9:0] m367_98;
   assign m367_98 =10'b0;

   // m367_99 = W*in
   wire signed [9:0] m367_99;
   assign m367_99 =10'b0;

   // m367_100 = W*in
   wire signed [9:0] m367_100;
   assign m367_100 =10'b0;

   // m367_101 = W*in
   wire signed [9:0] m367_101;
   assign m367_101 =10'b0;

   // m367_102 = W*in
   wire signed [9:0] m367_102;
   assign m367_102 =10'b0;

   // m367_103 = W*in
   wire signed [9:0] m367_103;
   assign m367_103 =10'b0;

   // m367_104 = W*in
   wire signed [9:0] m367_104;
   assign m367_104 =10'b0;

   // m367_105 = W*in
   wire signed [9:0] m367_105;
   assign m367_105 =10'b0;

   // m367_106 = W*in
   wire signed [9:0] m367_106;
   assign m367_106 ={ {5{neg367[5]}} , neg367[5:1] };

   // m367_107 = W*in
   wire signed [9:0] m367_107;
   assign m367_107 ={ {5{in367[5]}} , in367[5:1] };

   // m367_108 = W*in
   wire signed [9:0] m367_108;
   assign m367_108 =10'b0;

   // m367_109 = W*in
   wire signed [9:0] m367_109;
   assign m367_109 ={ {4{in367[5]}} , in367[5:0] };

   // m367_110 = W*in
   wire signed [9:0] m367_110;
   assign m367_110 =10'b0;

   // m367_111 = W*in
   wire signed [9:0] m367_111;
   assign m367_111 =10'b0;

   // m367_112 = W*in
   wire signed [9:0] m367_112;
   assign m367_112 =10'b0;

   // m367_113 = W*in
   wire signed [9:0] m367_113;
   assign m367_113 =10'b0;

   // m367_114 = W*in
   wire signed [9:0] m367_114;
   assign m367_114 =10'b0;

   // m367_115 = W*in
   wire signed [9:0] m367_115;
   assign m367_115 ={ {5{neg367[5]}} , neg367[5:1] };

   // m367_116 = W*in
   wire signed [9:0] m367_116;
   assign m367_116 ={ {4{in367[5]}} , in367[5:0] };

   // m367_117 = W*in
   wire signed [9:0] m367_117;
   assign m367_117 =10'b0;

   // m368_1 = W*in
   wire signed [9:0] m368_1;
   assign m368_1 =10'b0;

   // m368_2 = W*in
   wire signed [9:0] m368_2;
   assign m368_2 =10'b0;

   // m368_3 = W*in
   wire signed [9:0] m368_3;
   assign m368_3 ={ {4{in368[5]}} , in368[5:0] };

   // m368_4 = W*in
   wire signed [9:0] m368_4;
   assign m368_4 =10'b0;

   // m368_5 = W*in
   wire signed [9:0] m368_5;
   assign m368_5 =10'b0;

   // m368_6 = W*in
   wire signed [9:0] m368_6;
   assign m368_6 =10'b0;

   // m368_7 = W*in
   wire signed [9:0] m368_7;
   assign m368_7 =10'b0;

   // m368_8 = W*in
   wire signed [9:0] m368_8;
   assign m368_8 =10'b0;

   // m368_9 = W*in
   wire signed [9:0] m368_9;
   assign m368_9 =10'b0;

   // m368_10 = W*in
   wire signed [9:0] m368_10;
   assign m368_10 ={ {4{in368[5]}} , in368[5:0] };

   // m368_11 = W*in
   wire signed [9:0] m368_11;
   assign m368_11 ={ {4{in368[5]}} , in368[5:0] };

   // m368_12 = W*in
   wire signed [9:0] m368_12;
   assign m368_12 ={ {4{in368[5]}} , in368[5:0] };

   // m368_13 = W*in
   wire signed [9:0] m368_13;
   assign m368_13 =10'b0;

   // m368_14 = W*in
   wire signed [9:0] m368_14;
   assign m368_14 =10'b0;

   // m368_15 = W*in
   wire signed [9:0] m368_15;
   assign m368_15 =10'b0;

   // m368_16 = W*in
   wire signed [9:0] m368_16;
   assign m368_16 ={ {5{neg368[5]}} , neg368[5:1] };

   // m368_17 = W*in
   wire signed [9:0] m368_17;
   assign m368_17 ={ {4{in368[5]}} , in368[5:0] };

   // m368_18 = W*in
   wire signed [9:0] m368_18;
   assign m368_18 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_19 = W*in
   wire signed [9:0] m368_19;
   assign m368_19 ={ {4{in368[5]}} , in368[5:0] };

   // m368_20 = W*in
   wire signed [9:0] m368_20;
   assign m368_20 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_21 = W*in
   wire signed [9:0] m368_21;
   assign m368_21 ={ {4{in368[5]}} , in368[5:0] };

   // m368_22 = W*in
   wire signed [9:0] m368_22;
   assign m368_22 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_23 = W*in
   wire signed [9:0] m368_23;
   assign m368_23 =10'b0;

   // m368_24 = W*in
   wire signed [9:0] m368_24;
   assign m368_24 =10'b0;

   // m368_25 = W*in
   wire signed [9:0] m368_25;
   assign m368_25 ={ {5{in368[5]}} , in368[5:1] };

   // m368_26 = W*in
   wire signed [9:0] m368_26;
   assign m368_26 =10'b0;

   // m368_27 = W*in
   wire signed [9:0] m368_27;
   assign m368_27 =10'b0;

   // m368_28 = W*in
   wire signed [9:0] m368_28;
   assign m368_28 =10'b0;

   // m368_29 = W*in
   wire signed [9:0] m368_29;
   assign m368_29 ={ {4{in368[5]}} , in368[5:0] };

   // m368_30 = W*in
   wire signed [9:0] m368_30;
   assign m368_30 ={ {5{neg368[5]}} , neg368[5:1] };

   // m368_31 = W*in
   wire signed [9:0] m368_31;
   assign m368_31 =10'b0;

   // m368_32 = W*in
   wire signed [9:0] m368_32;
   assign m368_32 =10'b0;

   // m368_33 = W*in
   wire signed [9:0] m368_33;
   assign m368_33 =10'b0;

   // m368_34 = W*in
   wire signed [9:0] m368_34;
   assign m368_34 =10'b0;

   // m368_35 = W*in
   wire signed [9:0] m368_35;
   assign m368_35 ={ {5{neg368[5]}} , neg368[5:1] };

   // m368_36 = W*in
   wire signed [9:0] m368_36;
   assign m368_36 ={ {4{in368[5]}} , in368[5:0] };

   // m368_37 = W*in
   wire signed [9:0] m368_37;
   assign m368_37 ={ {3{in368[5]}} , in368 , {1{1'b0}} };

   // m368_38 = W*in
   wire signed [9:0] m368_38;
   assign m368_38 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_39 = W*in
   wire signed [9:0] m368_39;
   assign m368_39 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_40 = W*in
   wire signed [9:0] m368_40;
   assign m368_40 =10'b0;

   // m368_41 = W*in
   wire signed [9:0] m368_41;
   assign m368_41 ={ {4{in368[5]}} , in368[5:0] };

   // m368_42 = W*in
   wire signed [9:0] m368_42;
   assign m368_42 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_43 = W*in
   wire signed [9:0] m368_43;
   assign m368_43 =10'b0;

   // m368_44 = W*in
   wire signed [9:0] m368_44;
   assign m368_44 =10'b0;

   // m368_45 = W*in
   wire signed [9:0] m368_45;
   assign m368_45 =10'b0;

   // m368_46 = W*in
   wire signed [9:0] m368_46;
   assign m368_46 ={ {4{in368[5]}} , in368[5:0] };

   // m368_47 = W*in
   wire signed [9:0] m368_47;
   assign m368_47 =10'b0;

   // m368_48 = W*in
   wire signed [9:0] m368_48;
   assign m368_48 =10'b0;

   // m368_49 = W*in
   wire signed [9:0] m368_49;
   assign m368_49 =10'b0;

   // m368_50 = W*in
   wire signed [9:0] m368_50;
   assign m368_50 =10'b0;

   // m368_51 = W*in
   wire signed [9:0] m368_51;
   assign m368_51 =10'b0;

   // m368_52 = W*in
   wire signed [9:0] m368_52;
   assign m368_52 =10'b0;

   // m368_53 = W*in
   wire signed [9:0] m368_53;
   assign m368_53 ={ {4{in368[5]}} , in368[5:0] };

   // m368_54 = W*in
   wire signed [9:0] m368_54;
   assign m368_54 =10'b0;

   // m368_55 = W*in
   wire signed [9:0] m368_55;
   assign m368_55 =10'b0;

   // m368_56 = W*in
   wire signed [9:0] m368_56;
   assign m368_56 =10'b0;

   // m368_57 = W*in
   wire signed [9:0] m368_57;
   assign m368_57 =10'b0;

   // m368_58 = W*in
   wire signed [9:0] m368_58;
   assign m368_58 =10'b0;

   // m368_59 = W*in
   wire signed [9:0] m368_59;
   assign m368_59 =10'b0;

   // m368_60 = W*in
   wire signed [9:0] m368_60;
   assign m368_60 ={ {4{in368[5]}} , in368[5:0] };

   // m368_61 = W*in
   wire signed [9:0] m368_61;
   assign m368_61 =10'b0;

   // m368_62 = W*in
   wire signed [9:0] m368_62;
   assign m368_62 =10'b0;

   // m368_63 = W*in
   wire signed [9:0] m368_63;
   assign m368_63 =10'b0;

   // m368_64 = W*in
   wire signed [9:0] m368_64;
   assign m368_64 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_65 = W*in
   wire signed [9:0] m368_65;
   assign m368_65 =10'b0;

   // m368_66 = W*in
   wire signed [9:0] m368_66;
   assign m368_66 ={ {4{in368[5]}} , in368[5:0] };

   // m368_67 = W*in
   wire signed [9:0] m368_67;
   assign m368_67 ={ {4{in368[5]}} , in368[5:0] };

   // m368_68 = W*in
   wire signed [9:0] m368_68;
   assign m368_68 =10'b0;

   // m368_69 = W*in
   wire signed [9:0] m368_69;
   assign m368_69 =10'b0;

   // m368_70 = W*in
   wire signed [9:0] m368_70;
   assign m368_70 =10'b0;

   // m368_71 = W*in
   wire signed [9:0] m368_71;
   assign m368_71 =10'b0;

   // m368_72 = W*in
   wire signed [9:0] m368_72;
   assign m368_72 =10'b0;

   // m368_73 = W*in
   wire signed [9:0] m368_73;
   assign m368_73 =10'b0;

   // m368_74 = W*in
   wire signed [9:0] m368_74;
   assign m368_74 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_75 = W*in
   wire signed [9:0] m368_75;
   assign m368_75 =10'b0;

   // m368_76 = W*in
   wire signed [9:0] m368_76;
   assign m368_76 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_77 = W*in
   wire signed [9:0] m368_77;
   assign m368_77 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_78 = W*in
   wire signed [9:0] m368_78;
   assign m368_78 =10'b0;

   // m368_79 = W*in
   wire signed [9:0] m368_79;
   assign m368_79 ={ {4{in368[5]}} , in368[5:0] };

   // m368_80 = W*in
   wire signed [9:0] m368_80;
   assign m368_80 =10'b0;

   // m368_81 = W*in
   wire signed [9:0] m368_81;
   assign m368_81 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_82 = W*in
   wire signed [9:0] m368_82;
   assign m368_82 =10'b0;

   // m368_83 = W*in
   wire signed [9:0] m368_83;
   assign m368_83 =10'b0;

   // m368_84 = W*in
   wire signed [9:0] m368_84;
   assign m368_84 =10'b0;

   // m368_85 = W*in
   wire signed [9:0] m368_85;
   assign m368_85 ={ {3{in368[5]}} , in368 , {1{1'b0}} };

   // m368_86 = W*in
   wire signed [9:0] m368_86;
   assign m368_86 =10'b0;

   // m368_87 = W*in
   wire signed [9:0] m368_87;
   assign m368_87 =10'b0;

   // m368_88 = W*in
   wire signed [9:0] m368_88;
   assign m368_88 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_89 = W*in
   wire signed [9:0] m368_89;
   assign m368_89 =10'b0;

   // m368_90 = W*in
   wire signed [9:0] m368_90;
   assign m368_90 =10'b0;

   // m368_91 = W*in
   wire signed [9:0] m368_91;
   assign m368_91 =10'b0;

   // m368_92 = W*in
   wire signed [9:0] m368_92;
   assign m368_92 =10'b0;

   // m368_93 = W*in
   wire signed [9:0] m368_93;
   assign m368_93 ={ {4{in368[5]}} , in368[5:0] };

   // m368_94 = W*in
   wire signed [9:0] m368_94;
   assign m368_94 =10'b0;

   // m368_95 = W*in
   wire signed [9:0] m368_95;
   assign m368_95 ={ {4{in368[5]}} , in368[5:0] };

   // m368_96 = W*in
   wire signed [9:0] m368_96;
   assign m368_96 =10'b0;

   // m368_97 = W*in
   wire signed [9:0] m368_97;
   assign m368_97 =10'b0;

   // m368_98 = W*in
   wire signed [9:0] m368_98;
   assign m368_98 =10'b0;

   // m368_99 = W*in
   wire signed [9:0] m368_99;
   assign m368_99 =10'b0;

   // m368_100 = W*in
   wire signed [9:0] m368_100;
   assign m368_100 =10'b0;

   // m368_101 = W*in
   wire signed [9:0] m368_101;
   assign m368_101 =10'b0;

   // m368_102 = W*in
   wire signed [9:0] m368_102;
   assign m368_102 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_103 = W*in
   wire signed [9:0] m368_103;
   assign m368_103 ={ {4{in368[5]}} , in368[5:0] };

   // m368_104 = W*in
   wire signed [9:0] m368_104;
   assign m368_104 ={ {4{in368[5]}} , in368[5:0] };

   // m368_105 = W*in
   wire signed [9:0] m368_105;
   assign m368_105 =10'b0;

   // m368_106 = W*in
   wire signed [9:0] m368_106;
   assign m368_106 ={ {5{neg368[5]}} , neg368[5:1] };

   // m368_107 = W*in
   wire signed [9:0] m368_107;
   assign m368_107 ={ {4{in368[5]}} , in368[5:0] };

   // m368_108 = W*in
   wire signed [9:0] m368_108;
   assign m368_108 =10'b0;

   // m368_109 = W*in
   wire signed [9:0] m368_109;
   assign m368_109 =10'b0;

   // m368_110 = W*in
   wire signed [9:0] m368_110;
   assign m368_110 =10'b0;

   // m368_111 = W*in
   wire signed [9:0] m368_111;
   assign m368_111 =10'b0;

   // m368_112 = W*in
   wire signed [9:0] m368_112;
   assign m368_112 =10'b0;

   // m368_113 = W*in
   wire signed [9:0] m368_113;
   assign m368_113 ={ {4{neg368[5]}} , neg368[5:0] };

   // m368_114 = W*in
   wire signed [9:0] m368_114;
   assign m368_114 =10'b0;

   // m368_115 = W*in
   wire signed [9:0] m368_115;
   assign m368_115 ={ {5{neg368[5]}} , neg368[5:1] };

   // m368_116 = W*in
   wire signed [9:0] m368_116;
   assign m368_116 ={ {4{in368[5]}} , in368[5:0] };

   // m368_117 = W*in
   wire signed [9:0] m368_117;
   assign m368_117 ={ {4{neg368[5]}} , neg368[5:0] };

   // m369_1 = W*in
   wire signed [9:0] m369_1;
   assign m369_1 =10'b0;

   // m369_2 = W*in
   wire signed [9:0] m369_2;
   assign m369_2 =10'b0;

   // m369_3 = W*in
   wire signed [9:0] m369_3;
   assign m369_3 =10'b0;

   // m369_4 = W*in
   wire signed [9:0] m369_4;
   assign m369_4 =10'b0;

   // m369_5 = W*in
   wire signed [9:0] m369_5;
   assign m369_5 =10'b0;

   // m369_6 = W*in
   wire signed [9:0] m369_6;
   assign m369_6 =10'b0;

   // m369_7 = W*in
   wire signed [9:0] m369_7;
   assign m369_7 =10'b0;

   // m369_8 = W*in
   wire signed [9:0] m369_8;
   assign m369_8 =10'b0;

   // m369_9 = W*in
   wire signed [9:0] m369_9;
   assign m369_9 =10'b0;

   // m369_10 = W*in
   wire signed [9:0] m369_10;
   assign m369_10 ={ {4{in369[5]}} , in369[5:0] };

   // m369_11 = W*in
   wire signed [9:0] m369_11;
   assign m369_11 =10'b0;

   // m369_12 = W*in
   wire signed [9:0] m369_12;
   assign m369_12 =10'b0;

   // m369_13 = W*in
   wire signed [9:0] m369_13;
   assign m369_13 =10'b0;

   // m369_14 = W*in
   wire signed [9:0] m369_14;
   assign m369_14 =10'b0;

   // m369_15 = W*in
   wire signed [9:0] m369_15;
   assign m369_15 =10'b0;

   // m369_16 = W*in
   wire signed [9:0] m369_16;
   assign m369_16 ={ {5{neg369[5]}} , neg369[5:1] };

   // m369_17 = W*in
   wire signed [9:0] m369_17;
   assign m369_17 =10'b0;

   // m369_18 = W*in
   wire signed [9:0] m369_18;
   assign m369_18 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_19 = W*in
   wire signed [9:0] m369_19;
   assign m369_19 =10'b0;

   // m369_20 = W*in
   wire signed [9:0] m369_20;
   assign m369_20 ={ {4{in369[5]}} , in369[5:0] };

   // m369_21 = W*in
   wire signed [9:0] m369_21;
   assign m369_21 ={ {4{in369[5]}} , in369[5:0] };

   // m369_22 = W*in
   wire signed [9:0] m369_22;
   assign m369_22 =10'b0;

   // m369_23 = W*in
   wire signed [9:0] m369_23;
   assign m369_23 =10'b0;

   // m369_24 = W*in
   wire signed [9:0] m369_24;
   assign m369_24 =10'b0;

   // m369_25 = W*in
   wire signed [9:0] m369_25;
   assign m369_25 =10'b0;

   // m369_26 = W*in
   wire signed [9:0] m369_26;
   assign m369_26 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_27 = W*in
   wire signed [9:0] m369_27;
   assign m369_27 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_28 = W*in
   wire signed [9:0] m369_28;
   assign m369_28 ={ {5{neg369[5]}} , neg369[5:1] };

   // m369_29 = W*in
   wire signed [9:0] m369_29;
   assign m369_29 =10'b0;

   // m369_30 = W*in
   wire signed [9:0] m369_30;
   assign m369_30 =10'b0;

   // m369_31 = W*in
   wire signed [9:0] m369_31;
   assign m369_31 =10'b0;

   // m369_32 = W*in
   wire signed [9:0] m369_32;
   assign m369_32 =10'b0;

   // m369_33 = W*in
   wire signed [9:0] m369_33;
   assign m369_33 =10'b0;

   // m369_34 = W*in
   wire signed [9:0] m369_34;
   assign m369_34 =10'b0;

   // m369_35 = W*in
   wire signed [9:0] m369_35;
   assign m369_35 ={ {5{in369[5]}} , in369[5:1] };

   // m369_36 = W*in
   wire signed [9:0] m369_36;
   assign m369_36 =10'b0;

   // m369_37 = W*in
   wire signed [9:0] m369_37;
   assign m369_37 =10'b0;

   // m369_38 = W*in
   wire signed [9:0] m369_38;
   assign m369_38 =10'b0;

   // m369_39 = W*in
   wire signed [9:0] m369_39;
   assign m369_39 =10'b0;

   // m369_40 = W*in
   wire signed [9:0] m369_40;
   assign m369_40 =10'b0;

   // m369_41 = W*in
   wire signed [9:0] m369_41;
   assign m369_41 ={ {4{in369[5]}} , in369[5:0] };

   // m369_42 = W*in
   wire signed [9:0] m369_42;
   assign m369_42 =10'b0;

   // m369_43 = W*in
   wire signed [9:0] m369_43;
   assign m369_43 =10'b0;

   // m369_44 = W*in
   wire signed [9:0] m369_44;
   assign m369_44 =10'b0;

   // m369_45 = W*in
   wire signed [9:0] m369_45;
   assign m369_45 =10'b0;

   // m369_46 = W*in
   wire signed [9:0] m369_46;
   assign m369_46 =10'b0;

   // m369_47 = W*in
   wire signed [9:0] m369_47;
   assign m369_47 =10'b0;

   // m369_48 = W*in
   wire signed [9:0] m369_48;
   assign m369_48 =10'b0;

   // m369_49 = W*in
   wire signed [9:0] m369_49;
   assign m369_49 =10'b0;

   // m369_50 = W*in
   wire signed [9:0] m369_50;
   assign m369_50 =10'b0;

   // m369_51 = W*in
   wire signed [9:0] m369_51;
   assign m369_51 =10'b0;

   // m369_52 = W*in
   wire signed [9:0] m369_52;
   assign m369_52 =10'b0;

   // m369_53 = W*in
   wire signed [9:0] m369_53;
   assign m369_53 ={ {4{in369[5]}} , in369[5:0] };

   // m369_54 = W*in
   wire signed [9:0] m369_54;
   assign m369_54 =10'b0;

   // m369_55 = W*in
   wire signed [9:0] m369_55;
   assign m369_55 =10'b0;

   // m369_56 = W*in
   wire signed [9:0] m369_56;
   assign m369_56 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_57 = W*in
   wire signed [9:0] m369_57;
   assign m369_57 =10'b0;

   // m369_58 = W*in
   wire signed [9:0] m369_58;
   assign m369_58 =10'b0;

   // m369_59 = W*in
   wire signed [9:0] m369_59;
   assign m369_59 =10'b0;

   // m369_60 = W*in
   wire signed [9:0] m369_60;
   assign m369_60 =10'b0;

   // m369_61 = W*in
   wire signed [9:0] m369_61;
   assign m369_61 =10'b0;

   // m369_62 = W*in
   wire signed [9:0] m369_62;
   assign m369_62 =10'b0;

   // m369_63 = W*in
   wire signed [9:0] m369_63;
   assign m369_63 =10'b0;

   // m369_64 = W*in
   wire signed [9:0] m369_64;
   assign m369_64 =10'b0;

   // m369_65 = W*in
   wire signed [9:0] m369_65;
   assign m369_65 =10'b0;

   // m369_66 = W*in
   wire signed [9:0] m369_66;
   assign m369_66 =10'b0;

   // m369_67 = W*in
   wire signed [9:0] m369_67;
   assign m369_67 ={ {4{in369[5]}} , in369[5:0] };

   // m369_68 = W*in
   wire signed [9:0] m369_68;
   assign m369_68 =10'b0;

   // m369_69 = W*in
   wire signed [9:0] m369_69;
   assign m369_69 ={ {5{in369[5]}} , in369[5:1] };

   // m369_70 = W*in
   wire signed [9:0] m369_70;
   assign m369_70 =10'b0;

   // m369_71 = W*in
   wire signed [9:0] m369_71;
   assign m369_71 =10'b0;

   // m369_72 = W*in
   wire signed [9:0] m369_72;
   assign m369_72 ={ {4{in369[5]}} , in369[5:0] };

   // m369_73 = W*in
   wire signed [9:0] m369_73;
   assign m369_73 =10'b0;

   // m369_74 = W*in
   wire signed [9:0] m369_74;
   assign m369_74 =10'b0;

   // m369_75 = W*in
   wire signed [9:0] m369_75;
   assign m369_75 =10'b0;

   // m369_76 = W*in
   wire signed [9:0] m369_76;
   assign m369_76 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_77 = W*in
   wire signed [9:0] m369_77;
   assign m369_77 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_78 = W*in
   wire signed [9:0] m369_78;
   assign m369_78 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_79 = W*in
   wire signed [9:0] m369_79;
   assign m369_79 ={ {4{in369[5]}} , in369[5:0] };

   // m369_80 = W*in
   wire signed [9:0] m369_80;
   assign m369_80 ={ {5{neg369[5]}} , neg369[5:1] };

   // m369_81 = W*in
   wire signed [9:0] m369_81;
   assign m369_81 ={ {5{neg369[5]}} , neg369[5:1] };

   // m369_82 = W*in
   wire signed [9:0] m369_82;
   assign m369_82 =10'b0;

   // m369_83 = W*in
   wire signed [9:0] m369_83;
   assign m369_83 ={ {5{neg369[5]}} , neg369[5:1] };

   // m369_84 = W*in
   wire signed [9:0] m369_84;
   assign m369_84 ={ {5{in369[5]}} , in369[5:1] };

   // m369_85 = W*in
   wire signed [9:0] m369_85;
   assign m369_85 =10'b0;

   // m369_86 = W*in
   wire signed [9:0] m369_86;
   assign m369_86 =10'b0;

   // m369_87 = W*in
   wire signed [9:0] m369_87;
   assign m369_87 =10'b0;

   // m369_88 = W*in
   wire signed [9:0] m369_88;
   assign m369_88 =10'b0;

   // m369_89 = W*in
   wire signed [9:0] m369_89;
   assign m369_89 =10'b0;

   // m369_90 = W*in
   wire signed [9:0] m369_90;
   assign m369_90 =10'b0;

   // m369_91 = W*in
   wire signed [9:0] m369_91;
   assign m369_91 =10'b0;

   // m369_92 = W*in
   wire signed [9:0] m369_92;
   assign m369_92 =10'b0;

   // m369_93 = W*in
   wire signed [9:0] m369_93;
   assign m369_93 =10'b0;

   // m369_94 = W*in
   wire signed [9:0] m369_94;
   assign m369_94 =10'b0;

   // m369_95 = W*in
   wire signed [9:0] m369_95;
   assign m369_95 =10'b0;

   // m369_96 = W*in
   wire signed [9:0] m369_96;
   assign m369_96 =10'b0;

   // m369_97 = W*in
   wire signed [9:0] m369_97;
   assign m369_97 =10'b0;

   // m369_98 = W*in
   wire signed [9:0] m369_98;
   assign m369_98 ={ {4{neg369[5]}} , neg369[5:0] };

   // m369_99 = W*in
   wire signed [9:0] m369_99;
   assign m369_99 =10'b0;

   // m369_100 = W*in
   wire signed [9:0] m369_100;
   assign m369_100 =10'b0;

   // m369_101 = W*in
   wire signed [9:0] m369_101;
   assign m369_101 =10'b0;

   // m369_102 = W*in
   wire signed [9:0] m369_102;
   assign m369_102 =10'b0;

   // m369_103 = W*in
   wire signed [9:0] m369_103;
   assign m369_103 =10'b0;

   // m369_104 = W*in
   wire signed [9:0] m369_104;
   assign m369_104 =10'b0;

   // m369_105 = W*in
   wire signed [9:0] m369_105;
   assign m369_105 =10'b0;

   // m369_106 = W*in
   wire signed [9:0] m369_106;
   assign m369_106 =10'b0;

   // m369_107 = W*in
   wire signed [9:0] m369_107;
   assign m369_107 =10'b0;

   // m369_108 = W*in
   wire signed [9:0] m369_108;
   assign m369_108 ={ {4{in369[5]}} , in369[5:0] };

   // m369_109 = W*in
   wire signed [9:0] m369_109;
   assign m369_109 =10'b0;

   // m369_110 = W*in
   wire signed [9:0] m369_110;
   assign m369_110 =10'b0;

   // m369_111 = W*in
   wire signed [9:0] m369_111;
   assign m369_111 =10'b0;

   // m369_112 = W*in
   wire signed [9:0] m369_112;
   assign m369_112 =10'b0;

   // m369_113 = W*in
   wire signed [9:0] m369_113;
   assign m369_113 =10'b0;

   // m369_114 = W*in
   wire signed [9:0] m369_114;
   assign m369_114 =10'b0;

   // m369_115 = W*in
   wire signed [9:0] m369_115;
   assign m369_115 =10'b0;

   // m369_116 = W*in
   wire signed [9:0] m369_116;
   assign m369_116 ={ {4{in369[5]}} , in369[5:0] };

   // m369_117 = W*in
   wire signed [9:0] m369_117;
   assign m369_117 =10'b0;

   // m370_1 = W*in
   wire signed [9:0] m370_1;
   assign m370_1 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_2 = W*in
   wire signed [9:0] m370_2;
   assign m370_2 =10'b0;

   // m370_3 = W*in
   wire signed [9:0] m370_3;
   assign m370_3 =10'b0;

   // m370_4 = W*in
   wire signed [9:0] m370_4;
   assign m370_4 =10'b0;

   // m370_5 = W*in
   wire signed [9:0] m370_5;
   assign m370_5 =10'b0;

   // m370_6 = W*in
   wire signed [9:0] m370_6;
   assign m370_6 =10'b0;

   // m370_7 = W*in
   wire signed [9:0] m370_7;
   assign m370_7 =10'b0;

   // m370_8 = W*in
   wire signed [9:0] m370_8;
   assign m370_8 =10'b0;

   // m370_9 = W*in
   wire signed [9:0] m370_9;
   assign m370_9 =10'b0;

   // m370_10 = W*in
   wire signed [9:0] m370_10;
   assign m370_10 =10'b0;

   // m370_11 = W*in
   wire signed [9:0] m370_11;
   assign m370_11 =10'b0;

   // m370_12 = W*in
   wire signed [9:0] m370_12;
   assign m370_12 =10'b0;

   // m370_13 = W*in
   wire signed [9:0] m370_13;
   assign m370_13 =10'b0;

   // m370_14 = W*in
   wire signed [9:0] m370_14;
   assign m370_14 ={ {4{in370[5]}} , in370[5:0] };

   // m370_15 = W*in
   wire signed [9:0] m370_15;
   assign m370_15 =10'b0;

   // m370_16 = W*in
   wire signed [9:0] m370_16;
   assign m370_16 ={ {5{neg370[5]}} , neg370[5:1] };

   // m370_17 = W*in
   wire signed [9:0] m370_17;
   assign m370_17 ={ {5{neg370[5]}} , neg370[5:1] };

   // m370_18 = W*in
   wire signed [9:0] m370_18;
   assign m370_18 =10'b0;

   // m370_19 = W*in
   wire signed [9:0] m370_19;
   assign m370_19 =10'b0;

   // m370_20 = W*in
   wire signed [9:0] m370_20;
   assign m370_20 =10'b0;

   // m370_21 = W*in
   wire signed [9:0] m370_21;
   assign m370_21 ={ {4{in370[5]}} , in370[5:0] };

   // m370_22 = W*in
   wire signed [9:0] m370_22;
   assign m370_22 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_23 = W*in
   wire signed [9:0] m370_23;
   assign m370_23 =10'b0;

   // m370_24 = W*in
   wire signed [9:0] m370_24;
   assign m370_24 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_25 = W*in
   wire signed [9:0] m370_25;
   assign m370_25 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_26 = W*in
   wire signed [9:0] m370_26;
   assign m370_26 =10'b0;

   // m370_27 = W*in
   wire signed [9:0] m370_27;
   assign m370_27 ={ {5{neg370[5]}} , neg370[5:1] };

   // m370_28 = W*in
   wire signed [9:0] m370_28;
   assign m370_28 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_29 = W*in
   wire signed [9:0] m370_29;
   assign m370_29 ={ {4{in370[5]}} , in370[5:0] };

   // m370_30 = W*in
   wire signed [9:0] m370_30;
   assign m370_30 =10'b0;

   // m370_31 = W*in
   wire signed [9:0] m370_31;
   assign m370_31 =10'b0;

   // m370_32 = W*in
   wire signed [9:0] m370_32;
   assign m370_32 =10'b0;

   // m370_33 = W*in
   wire signed [9:0] m370_33;
   assign m370_33 =10'b0;

   // m370_34 = W*in
   wire signed [9:0] m370_34;
   assign m370_34 =10'b0;

   // m370_35 = W*in
   wire signed [9:0] m370_35;
   assign m370_35 =10'b0;

   // m370_36 = W*in
   wire signed [9:0] m370_36;
   assign m370_36 =10'b0;

   // m370_37 = W*in
   wire signed [9:0] m370_37;
   assign m370_37 =10'b0;

   // m370_38 = W*in
   wire signed [9:0] m370_38;
   assign m370_38 =10'b0;

   // m370_39 = W*in
   wire signed [9:0] m370_39;
   assign m370_39 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_40 = W*in
   wire signed [9:0] m370_40;
   assign m370_40 =10'b0;

   // m370_41 = W*in
   wire signed [9:0] m370_41;
   assign m370_41 =10'b0;

   // m370_42 = W*in
   wire signed [9:0] m370_42;
   assign m370_42 ={ {4{in370[5]}} , in370[5:0] };

   // m370_43 = W*in
   wire signed [9:0] m370_43;
   assign m370_43 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_44 = W*in
   wire signed [9:0] m370_44;
   assign m370_44 =10'b0;

   // m370_45 = W*in
   wire signed [9:0] m370_45;
   assign m370_45 =10'b0;

   // m370_46 = W*in
   wire signed [9:0] m370_46;
   assign m370_46 =10'b0;

   // m370_47 = W*in
   wire signed [9:0] m370_47;
   assign m370_47 =10'b0;

   // m370_48 = W*in
   wire signed [9:0] m370_48;
   assign m370_48 =10'b0;

   // m370_49 = W*in
   wire signed [9:0] m370_49;
   assign m370_49 =10'b0;

   // m370_50 = W*in
   wire signed [9:0] m370_50;
   assign m370_50 =10'b0;

   // m370_51 = W*in
   wire signed [9:0] m370_51;
   assign m370_51 =10'b0;

   // m370_52 = W*in
   wire signed [9:0] m370_52;
   assign m370_52 =10'b0;

   // m370_53 = W*in
   wire signed [9:0] m370_53;
   assign m370_53 ={ {4{in370[5]}} , in370[5:0] };

   // m370_54 = W*in
   wire signed [9:0] m370_54;
   assign m370_54 =10'b0;

   // m370_55 = W*in
   wire signed [9:0] m370_55;
   assign m370_55 =10'b0;

   // m370_56 = W*in
   wire signed [9:0] m370_56;
   assign m370_56 =10'b0;

   // m370_57 = W*in
   wire signed [9:0] m370_57;
   assign m370_57 =10'b0;

   // m370_58 = W*in
   wire signed [9:0] m370_58;
   assign m370_58 =10'b0;

   // m370_59 = W*in
   wire signed [9:0] m370_59;
   assign m370_59 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_60 = W*in
   wire signed [9:0] m370_60;
   assign m370_60 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_61 = W*in
   wire signed [9:0] m370_61;
   assign m370_61 =10'b0;

   // m370_62 = W*in
   wire signed [9:0] m370_62;
   assign m370_62 =10'b0;

   // m370_63 = W*in
   wire signed [9:0] m370_63;
   assign m370_63 ={ {5{in370[5]}} , in370[5:1] };

   // m370_64 = W*in
   wire signed [9:0] m370_64;
   assign m370_64 =10'b0;

   // m370_65 = W*in
   wire signed [9:0] m370_65;
   assign m370_65 ={ {5{in370[5]}} , in370[5:1] };

   // m370_66 = W*in
   wire signed [9:0] m370_66;
   assign m370_66 ={ {5{in370[5]}} , in370[5:1] };

   // m370_67 = W*in
   wire signed [9:0] m370_67;
   assign m370_67 =10'b0;

   // m370_68 = W*in
   wire signed [9:0] m370_68;
   assign m370_68 =10'b0;

   // m370_69 = W*in
   wire signed [9:0] m370_69;
   assign m370_69 ={ {4{in370[5]}} , in370[5:0] };

   // m370_70 = W*in
   wire signed [9:0] m370_70;
   assign m370_70 ={ {5{in370[5]}} , in370[5:1] };

   // m370_71 = W*in
   wire signed [9:0] m370_71;
   assign m370_71 =10'b0;

   // m370_72 = W*in
   wire signed [9:0] m370_72;
   assign m370_72 =10'b0;

   // m370_73 = W*in
   wire signed [9:0] m370_73;
   assign m370_73 =10'b0;

   // m370_74 = W*in
   wire signed [9:0] m370_74;
   assign m370_74 =10'b0;

   // m370_75 = W*in
   wire signed [9:0] m370_75;
   assign m370_75 =10'b0;

   // m370_76 = W*in
   wire signed [9:0] m370_76;
   assign m370_76 =10'b0;

   // m370_77 = W*in
   wire signed [9:0] m370_77;
   assign m370_77 ={ {4{in370[5]}} , in370[5:0] };

   // m370_78 = W*in
   wire signed [9:0] m370_78;
   assign m370_78 =10'b0;

   // m370_79 = W*in
   wire signed [9:0] m370_79;
   assign m370_79 =10'b0;

   // m370_80 = W*in
   wire signed [9:0] m370_80;
   assign m370_80 ={ {4{in370[5]}} , in370[5:0] };

   // m370_81 = W*in
   wire signed [9:0] m370_81;
   assign m370_81 =10'b0;

   // m370_82 = W*in
   wire signed [9:0] m370_82;
   assign m370_82 ={ {4{in370[5]}} , in370[5:0] };

   // m370_83 = W*in
   wire signed [9:0] m370_83;
   assign m370_83 =10'b0;

   // m370_84 = W*in
   wire signed [9:0] m370_84;
   assign m370_84 ={ {5{neg370[5]}} , neg370[5:1] };

   // m370_85 = W*in
   wire signed [9:0] m370_85;
   assign m370_85 ={ {4{in370[5]}} , in370[5:0] };

   // m370_86 = W*in
   wire signed [9:0] m370_86;
   assign m370_86 =10'b0;

   // m370_87 = W*in
   wire signed [9:0] m370_87;
   assign m370_87 =10'b0;

   // m370_88 = W*in
   wire signed [9:0] m370_88;
   assign m370_88 =10'b0;

   // m370_89 = W*in
   wire signed [9:0] m370_89;
   assign m370_89 =10'b0;

   // m370_90 = W*in
   wire signed [9:0] m370_90;
   assign m370_90 =10'b0;

   // m370_91 = W*in
   wire signed [9:0] m370_91;
   assign m370_91 =10'b0;

   // m370_92 = W*in
   wire signed [9:0] m370_92;
   assign m370_92 =10'b0;

   // m370_93 = W*in
   wire signed [9:0] m370_93;
   assign m370_93 ={ {4{in370[5]}} , in370[5:0] };

   // m370_94 = W*in
   wire signed [9:0] m370_94;
   assign m370_94 ={ {4{in370[5]}} , in370[5:0] };

   // m370_95 = W*in
   wire signed [9:0] m370_95;
   assign m370_95 =10'b0;

   // m370_96 = W*in
   wire signed [9:0] m370_96;
   assign m370_96 =10'b0;

   // m370_97 = W*in
   wire signed [9:0] m370_97;
   assign m370_97 =10'b0;

   // m370_98 = W*in
   wire signed [9:0] m370_98;
   assign m370_98 =10'b0;

   // m370_99 = W*in
   wire signed [9:0] m370_99;
   assign m370_99 =10'b0;

   // m370_100 = W*in
   wire signed [9:0] m370_100;
   assign m370_100 =10'b0;

   // m370_101 = W*in
   wire signed [9:0] m370_101;
   assign m370_101 =10'b0;

   // m370_102 = W*in
   wire signed [9:0] m370_102;
   assign m370_102 =10'b0;

   // m370_103 = W*in
   wire signed [9:0] m370_103;
   assign m370_103 =10'b0;

   // m370_104 = W*in
   wire signed [9:0] m370_104;
   assign m370_104 =10'b0;

   // m370_105 = W*in
   wire signed [9:0] m370_105;
   assign m370_105 =10'b0;

   // m370_106 = W*in
   wire signed [9:0] m370_106;
   assign m370_106 =10'b0;

   // m370_107 = W*in
   wire signed [9:0] m370_107;
   assign m370_107 ={ {5{neg370[5]}} , neg370[5:1] };

   // m370_108 = W*in
   wire signed [9:0] m370_108;
   assign m370_108 =10'b0;

   // m370_109 = W*in
   wire signed [9:0] m370_109;
   assign m370_109 =10'b0;

   // m370_110 = W*in
   wire signed [9:0] m370_110;
   assign m370_110 =10'b0;

   // m370_111 = W*in
   wire signed [9:0] m370_111;
   assign m370_111 =10'b0;

   // m370_112 = W*in
   wire signed [9:0] m370_112;
   assign m370_112 =10'b0;

   // m370_113 = W*in
   wire signed [9:0] m370_113;
   assign m370_113 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_114 = W*in
   wire signed [9:0] m370_114;
   assign m370_114 =10'b0;

   // m370_115 = W*in
   wire signed [9:0] m370_115;
   assign m370_115 ={ {4{neg370[5]}} , neg370[5:0] };

   // m370_116 = W*in
   wire signed [9:0] m370_116;
   assign m370_116 =10'b0;

   // m370_117 = W*in
   wire signed [9:0] m370_117;
   assign m370_117 ={ {4{neg370[5]}} , neg370[5:0] };

   // m371_1 = W*in
   wire signed [9:0] m371_1;
   assign m371_1 =10'b0;

   // m371_2 = W*in
   wire signed [9:0] m371_2;
   assign m371_2 =10'b0;

   // m371_3 = W*in
   wire signed [9:0] m371_3;
   assign m371_3 =10'b0;

   // m371_4 = W*in
   wire signed [9:0] m371_4;
   assign m371_4 =10'b0;

   // m371_5 = W*in
   wire signed [9:0] m371_5;
   assign m371_5 =10'b0;

   // m371_6 = W*in
   wire signed [9:0] m371_6;
   assign m371_6 =10'b0;

   // m371_7 = W*in
   wire signed [9:0] m371_7;
   assign m371_7 =10'b0;

   // m371_8 = W*in
   wire signed [9:0] m371_8;
   assign m371_8 =10'b0;

   // m371_9 = W*in
   wire signed [9:0] m371_9;
   assign m371_9 =10'b0;

   // m371_10 = W*in
   wire signed [9:0] m371_10;
   assign m371_10 =10'b0;

   // m371_11 = W*in
   wire signed [9:0] m371_11;
   assign m371_11 =10'b0;

   // m371_12 = W*in
   wire signed [9:0] m371_12;
   assign m371_12 =10'b0;

   // m371_13 = W*in
   wire signed [9:0] m371_13;
   assign m371_13 =10'b0;

   // m371_14 = W*in
   wire signed [9:0] m371_14;
   assign m371_14 =10'b0;

   // m371_15 = W*in
   wire signed [9:0] m371_15;
   assign m371_15 =10'b0;

   // m371_16 = W*in
   wire signed [9:0] m371_16;
   assign m371_16 =10'b0;

   // m371_17 = W*in
   wire signed [9:0] m371_17;
   assign m371_17 =10'b0;

   // m371_18 = W*in
   wire signed [9:0] m371_18;
   assign m371_18 =10'b0;

   // m371_19 = W*in
   wire signed [9:0] m371_19;
   assign m371_19 =10'b0;

   // m371_20 = W*in
   wire signed [9:0] m371_20;
   assign m371_20 ={ {5{neg371[5]}} , neg371[5:1] };

   // m371_21 = W*in
   wire signed [9:0] m371_21;
   assign m371_21 =10'b0;

   // m371_22 = W*in
   wire signed [9:0] m371_22;
   assign m371_22 =10'b0;

   // m371_23 = W*in
   wire signed [9:0] m371_23;
   assign m371_23 =10'b0;

   // m371_24 = W*in
   wire signed [9:0] m371_24;
   assign m371_24 =10'b0;

   // m371_25 = W*in
   wire signed [9:0] m371_25;
   assign m371_25 =10'b0;

   // m371_26 = W*in
   wire signed [9:0] m371_26;
   assign m371_26 =10'b0;

   // m371_27 = W*in
   wire signed [9:0] m371_27;
   assign m371_27 ={ {5{neg371[5]}} , neg371[5:1] };

   // m371_28 = W*in
   wire signed [9:0] m371_28;
   assign m371_28 =10'b0;

   // m371_29 = W*in
   wire signed [9:0] m371_29;
   assign m371_29 =10'b0;

   // m371_30 = W*in
   wire signed [9:0] m371_30;
   assign m371_30 =10'b0;

   // m371_31 = W*in
   wire signed [9:0] m371_31;
   assign m371_31 =10'b0;

   // m371_32 = W*in
   wire signed [9:0] m371_32;
   assign m371_32 =10'b0;

   // m371_33 = W*in
   wire signed [9:0] m371_33;
   assign m371_33 =10'b0;

   // m371_34 = W*in
   wire signed [9:0] m371_34;
   assign m371_34 ={ {5{neg371[5]}} , neg371[5:1] };

   // m371_35 = W*in
   wire signed [9:0] m371_35;
   assign m371_35 =10'b0;

   // m371_36 = W*in
   wire signed [9:0] m371_36;
   assign m371_36 =10'b0;

   // m371_37 = W*in
   wire signed [9:0] m371_37;
   assign m371_37 ={ {4{in371[5]}} , in371[5:0] };

   // m371_38 = W*in
   wire signed [9:0] m371_38;
   assign m371_38 =10'b0;

   // m371_39 = W*in
   wire signed [9:0] m371_39;
   assign m371_39 =10'b0;

   // m371_40 = W*in
   wire signed [9:0] m371_40;
   assign m371_40 =10'b0;

   // m371_41 = W*in
   wire signed [9:0] m371_41;
   assign m371_41 =10'b0;

   // m371_42 = W*in
   wire signed [9:0] m371_42;
   assign m371_42 =10'b0;

   // m371_43 = W*in
   wire signed [9:0] m371_43;
   assign m371_43 =10'b0;

   // m371_44 = W*in
   wire signed [9:0] m371_44;
   assign m371_44 =10'b0;

   // m371_45 = W*in
   wire signed [9:0] m371_45;
   assign m371_45 =10'b0;

   // m371_46 = W*in
   wire signed [9:0] m371_46;
   assign m371_46 =10'b0;

   // m371_47 = W*in
   wire signed [9:0] m371_47;
   assign m371_47 =10'b0;

   // m371_48 = W*in
   wire signed [9:0] m371_48;
   assign m371_48 =10'b0;

   // m371_49 = W*in
   wire signed [9:0] m371_49;
   assign m371_49 =10'b0;

   // m371_50 = W*in
   wire signed [9:0] m371_50;
   assign m371_50 =10'b0;

   // m371_51 = W*in
   wire signed [9:0] m371_51;
   assign m371_51 =10'b0;

   // m371_52 = W*in
   wire signed [9:0] m371_52;
   assign m371_52 =10'b0;

   // m371_53 = W*in
   wire signed [9:0] m371_53;
   assign m371_53 =10'b0;

   // m371_54 = W*in
   wire signed [9:0] m371_54;
   assign m371_54 =10'b0;

   // m371_55 = W*in
   wire signed [9:0] m371_55;
   assign m371_55 =10'b0;

   // m371_56 = W*in
   wire signed [9:0] m371_56;
   assign m371_56 =10'b0;

   // m371_57 = W*in
   wire signed [9:0] m371_57;
   assign m371_57 =10'b0;

   // m371_58 = W*in
   wire signed [9:0] m371_58;
   assign m371_58 =10'b0;

   // m371_59 = W*in
   wire signed [9:0] m371_59;
   assign m371_59 =10'b0;

   // m371_60 = W*in
   wire signed [9:0] m371_60;
   assign m371_60 =10'b0;

   // m371_61 = W*in
   wire signed [9:0] m371_61;
   assign m371_61 =10'b0;

   // m371_62 = W*in
   wire signed [9:0] m371_62;
   assign m371_62 =10'b0;

   // m371_63 = W*in
   wire signed [9:0] m371_63;
   assign m371_63 =10'b0;

   // m371_64 = W*in
   wire signed [9:0] m371_64;
   assign m371_64 ={ {5{neg371[5]}} , neg371[5:1] };

   // m371_65 = W*in
   wire signed [9:0] m371_65;
   assign m371_65 =10'b0;

   // m371_66 = W*in
   wire signed [9:0] m371_66;
   assign m371_66 ={ {5{in371[5]}} , in371[5:1] };

   // m371_67 = W*in
   wire signed [9:0] m371_67;
   assign m371_67 =10'b0;

   // m371_68 = W*in
   wire signed [9:0] m371_68;
   assign m371_68 =10'b0;

   // m371_69 = W*in
   wire signed [9:0] m371_69;
   assign m371_69 ={ {5{in371[5]}} , in371[5:1] };

   // m371_70 = W*in
   wire signed [9:0] m371_70;
   assign m371_70 =10'b0;

   // m371_71 = W*in
   wire signed [9:0] m371_71;
   assign m371_71 =10'b0;

   // m371_72 = W*in
   wire signed [9:0] m371_72;
   assign m371_72 =10'b0;

   // m371_73 = W*in
   wire signed [9:0] m371_73;
   assign m371_73 =10'b0;

   // m371_74 = W*in
   wire signed [9:0] m371_74;
   assign m371_74 =10'b0;

   // m371_75 = W*in
   wire signed [9:0] m371_75;
   assign m371_75 =10'b0;

   // m371_76 = W*in
   wire signed [9:0] m371_76;
   assign m371_76 =10'b0;

   // m371_77 = W*in
   wire signed [9:0] m371_77;
   assign m371_77 =10'b0;

   // m371_78 = W*in
   wire signed [9:0] m371_78;
   assign m371_78 =10'b0;

   // m371_79 = W*in
   wire signed [9:0] m371_79;
   assign m371_79 =10'b0;

   // m371_80 = W*in
   wire signed [9:0] m371_80;
   assign m371_80 =10'b0;

   // m371_81 = W*in
   wire signed [9:0] m371_81;
   assign m371_81 =10'b0;

   // m371_82 = W*in
   wire signed [9:0] m371_82;
   assign m371_82 =10'b0;

   // m371_83 = W*in
   wire signed [9:0] m371_83;
   assign m371_83 =10'b0;

   // m371_84 = W*in
   wire signed [9:0] m371_84;
   assign m371_84 =10'b0;

   // m371_85 = W*in
   wire signed [9:0] m371_85;
   assign m371_85 ={ {4{in371[5]}} , in371[5:0] };

   // m371_86 = W*in
   wire signed [9:0] m371_86;
   assign m371_86 =10'b0;

   // m371_87 = W*in
   wire signed [9:0] m371_87;
   assign m371_87 ={ {4{neg371[5]}} , neg371[5:0] };

   // m371_88 = W*in
   wire signed [9:0] m371_88;
   assign m371_88 =10'b0;

   // m371_89 = W*in
   wire signed [9:0] m371_89;
   assign m371_89 =10'b0;

   // m371_90 = W*in
   wire signed [9:0] m371_90;
   assign m371_90 =10'b0;

   // m371_91 = W*in
   wire signed [9:0] m371_91;
   assign m371_91 =10'b0;

   // m371_92 = W*in
   wire signed [9:0] m371_92;
   assign m371_92 =10'b0;

   // m371_93 = W*in
   wire signed [9:0] m371_93;
   assign m371_93 =10'b0;

   // m371_94 = W*in
   wire signed [9:0] m371_94;
   assign m371_94 =10'b0;

   // m371_95 = W*in
   wire signed [9:0] m371_95;
   assign m371_95 =10'b0;

   // m371_96 = W*in
   wire signed [9:0] m371_96;
   assign m371_96 =10'b0;

   // m371_97 = W*in
   wire signed [9:0] m371_97;
   assign m371_97 =10'b0;

   // m371_98 = W*in
   wire signed [9:0] m371_98;
   assign m371_98 =10'b0;

   // m371_99 = W*in
   wire signed [9:0] m371_99;
   assign m371_99 =10'b0;

   // m371_100 = W*in
   wire signed [9:0] m371_100;
   assign m371_100 =10'b0;

   // m371_101 = W*in
   wire signed [9:0] m371_101;
   assign m371_101 =10'b0;

   // m371_102 = W*in
   wire signed [9:0] m371_102;
   assign m371_102 =10'b0;

   // m371_103 = W*in
   wire signed [9:0] m371_103;
   assign m371_103 =10'b0;

   // m371_104 = W*in
   wire signed [9:0] m371_104;
   assign m371_104 =10'b0;

   // m371_105 = W*in
   wire signed [9:0] m371_105;
   assign m371_105 =10'b0;

   // m371_106 = W*in
   wire signed [9:0] m371_106;
   assign m371_106 =10'b0;

   // m371_107 = W*in
   wire signed [9:0] m371_107;
   assign m371_107 =10'b0;

   // m371_108 = W*in
   wire signed [9:0] m371_108;
   assign m371_108 =10'b0;

   // m371_109 = W*in
   wire signed [9:0] m371_109;
   assign m371_109 =10'b0;

   // m371_110 = W*in
   wire signed [9:0] m371_110;
   assign m371_110 =10'b0;

   // m371_111 = W*in
   wire signed [9:0] m371_111;
   assign m371_111 =10'b0;

   // m371_112 = W*in
   wire signed [9:0] m371_112;
   assign m371_112 =10'b0;

   // m371_113 = W*in
   wire signed [9:0] m371_113;
   assign m371_113 =10'b0;

   // m371_114 = W*in
   wire signed [9:0] m371_114;
   assign m371_114 =10'b0;

   // m371_115 = W*in
   wire signed [9:0] m371_115;
   assign m371_115 ={ {5{neg371[5]}} , neg371[5:1] };

   // m371_116 = W*in
   wire signed [9:0] m371_116;
   assign m371_116 =10'b0;

   // m371_117 = W*in
   wire signed [9:0] m371_117;
   assign m371_117 =10'b0;

   // m372_1 = W*in
   wire signed [9:0] m372_1;
   assign m372_1 =10'b0;

   // m372_2 = W*in
   wire signed [9:0] m372_2;
   assign m372_2 =10'b0;

   // m372_3 = W*in
   wire signed [9:0] m372_3;
   assign m372_3 =10'b0;

   // m372_4 = W*in
   wire signed [9:0] m372_4;
   assign m372_4 =10'b0;

   // m372_5 = W*in
   wire signed [9:0] m372_5;
   assign m372_5 =10'b0;

   // m372_6 = W*in
   wire signed [9:0] m372_6;
   assign m372_6 =10'b0;

   // m372_7 = W*in
   wire signed [9:0] m372_7;
   assign m372_7 =10'b0;

   // m372_8 = W*in
   wire signed [9:0] m372_8;
   assign m372_8 =10'b0;

   // m372_9 = W*in
   wire signed [9:0] m372_9;
   assign m372_9 =10'b0;

   // m372_10 = W*in
   wire signed [9:0] m372_10;
   assign m372_10 =10'b0;

   // m372_11 = W*in
   wire signed [9:0] m372_11;
   assign m372_11 =10'b0;

   // m372_12 = W*in
   wire signed [9:0] m372_12;
   assign m372_12 =10'b0;

   // m372_13 = W*in
   wire signed [9:0] m372_13;
   assign m372_13 =10'b0;

   // m372_14 = W*in
   wire signed [9:0] m372_14;
   assign m372_14 =10'b0;

   // m372_15 = W*in
   wire signed [9:0] m372_15;
   assign m372_15 =10'b0;

   // m372_16 = W*in
   wire signed [9:0] m372_16;
   assign m372_16 =10'b0;

   // m372_17 = W*in
   wire signed [9:0] m372_17;
   assign m372_17 ={ {5{in372[5]}} , in372[5:1] };

   // m372_18 = W*in
   wire signed [9:0] m372_18;
   assign m372_18 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_19 = W*in
   wire signed [9:0] m372_19;
   assign m372_19 =10'b0;

   // m372_20 = W*in
   wire signed [9:0] m372_20;
   assign m372_20 ={ {5{neg372[5]}} , neg372[5:1] };

   // m372_21 = W*in
   wire signed [9:0] m372_21;
   assign m372_21 =10'b0;

   // m372_22 = W*in
   wire signed [9:0] m372_22;
   assign m372_22 =10'b0;

   // m372_23 = W*in
   wire signed [9:0] m372_23;
   assign m372_23 ={ {4{in372[5]}} , in372[5:0] };

   // m372_24 = W*in
   wire signed [9:0] m372_24;
   assign m372_24 =10'b0;

   // m372_25 = W*in
   wire signed [9:0] m372_25;
   assign m372_25 =10'b0;

   // m372_26 = W*in
   wire signed [9:0] m372_26;
   assign m372_26 ={ {5{neg372[5]}} , neg372[5:1] };

   // m372_27 = W*in
   wire signed [9:0] m372_27;
   assign m372_27 =10'b0;

   // m372_28 = W*in
   wire signed [9:0] m372_28;
   assign m372_28 =10'b0;

   // m372_29 = W*in
   wire signed [9:0] m372_29;
   assign m372_29 =10'b0;

   // m372_30 = W*in
   wire signed [9:0] m372_30;
   assign m372_30 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_31 = W*in
   wire signed [9:0] m372_31;
   assign m372_31 =10'b0;

   // m372_32 = W*in
   wire signed [9:0] m372_32;
   assign m372_32 =10'b0;

   // m372_33 = W*in
   wire signed [9:0] m372_33;
   assign m372_33 =10'b0;

   // m372_34 = W*in
   wire signed [9:0] m372_34;
   assign m372_34 =10'b0;

   // m372_35 = W*in
   wire signed [9:0] m372_35;
   assign m372_35 ={ {5{neg372[5]}} , neg372[5:1] };

   // m372_36 = W*in
   wire signed [9:0] m372_36;
   assign m372_36 =10'b0;

   // m372_37 = W*in
   wire signed [9:0] m372_37;
   assign m372_37 =10'b0;

   // m372_38 = W*in
   wire signed [9:0] m372_38;
   assign m372_38 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_39 = W*in
   wire signed [9:0] m372_39;
   assign m372_39 =10'b0;

   // m372_40 = W*in
   wire signed [9:0] m372_40;
   assign m372_40 =10'b0;

   // m372_41 = W*in
   wire signed [9:0] m372_41;
   assign m372_41 =10'b0;

   // m372_42 = W*in
   wire signed [9:0] m372_42;
   assign m372_42 =10'b0;

   // m372_43 = W*in
   wire signed [9:0] m372_43;
   assign m372_43 =10'b0;

   // m372_44 = W*in
   wire signed [9:0] m372_44;
   assign m372_44 =10'b0;

   // m372_45 = W*in
   wire signed [9:0] m372_45;
   assign m372_45 ={ {4{in372[5]}} , in372[5:0] };

   // m372_46 = W*in
   wire signed [9:0] m372_46;
   assign m372_46 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_47 = W*in
   wire signed [9:0] m372_47;
   assign m372_47 =10'b0;

   // m372_48 = W*in
   wire signed [9:0] m372_48;
   assign m372_48 =10'b0;

   // m372_49 = W*in
   wire signed [9:0] m372_49;
   assign m372_49 =10'b0;

   // m372_50 = W*in
   wire signed [9:0] m372_50;
   assign m372_50 =10'b0;

   // m372_51 = W*in
   wire signed [9:0] m372_51;
   assign m372_51 =10'b0;

   // m372_52 = W*in
   wire signed [9:0] m372_52;
   assign m372_52 =10'b0;

   // m372_53 = W*in
   wire signed [9:0] m372_53;
   assign m372_53 =10'b0;

   // m372_54 = W*in
   wire signed [9:0] m372_54;
   assign m372_54 ={ {4{in372[5]}} , in372[5:0] };

   // m372_55 = W*in
   wire signed [9:0] m372_55;
   assign m372_55 =10'b0;

   // m372_56 = W*in
   wire signed [9:0] m372_56;
   assign m372_56 =10'b0;

   // m372_57 = W*in
   wire signed [9:0] m372_57;
   assign m372_57 =10'b0;

   // m372_58 = W*in
   wire signed [9:0] m372_58;
   assign m372_58 =10'b0;

   // m372_59 = W*in
   wire signed [9:0] m372_59;
   assign m372_59 =10'b0;

   // m372_60 = W*in
   wire signed [9:0] m372_60;
   assign m372_60 =10'b0;

   // m372_61 = W*in
   wire signed [9:0] m372_61;
   assign m372_61 =10'b0;

   // m372_62 = W*in
   wire signed [9:0] m372_62;
   assign m372_62 =10'b0;

   // m372_63 = W*in
   wire signed [9:0] m372_63;
   assign m372_63 =10'b0;

   // m372_64 = W*in
   wire signed [9:0] m372_64;
   assign m372_64 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_65 = W*in
   wire signed [9:0] m372_65;
   assign m372_65 =10'b0;

   // m372_66 = W*in
   wire signed [9:0] m372_66;
   assign m372_66 =10'b0;

   // m372_67 = W*in
   wire signed [9:0] m372_67;
   assign m372_67 =10'b0;

   // m372_68 = W*in
   wire signed [9:0] m372_68;
   assign m372_68 =10'b0;

   // m372_69 = W*in
   wire signed [9:0] m372_69;
   assign m372_69 ={ {4{in372[5]}} , in372[5:0] };

   // m372_70 = W*in
   wire signed [9:0] m372_70;
   assign m372_70 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_71 = W*in
   wire signed [9:0] m372_71;
   assign m372_71 =10'b0;

   // m372_72 = W*in
   wire signed [9:0] m372_72;
   assign m372_72 =10'b0;

   // m372_73 = W*in
   wire signed [9:0] m372_73;
   assign m372_73 ={ {4{in372[5]}} , in372[5:0] };

   // m372_74 = W*in
   wire signed [9:0] m372_74;
   assign m372_74 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_75 = W*in
   wire signed [9:0] m372_75;
   assign m372_75 =10'b0;

   // m372_76 = W*in
   wire signed [9:0] m372_76;
   assign m372_76 =10'b0;

   // m372_77 = W*in
   wire signed [9:0] m372_77;
   assign m372_77 =10'b0;

   // m372_78 = W*in
   wire signed [9:0] m372_78;
   assign m372_78 =10'b0;

   // m372_79 = W*in
   wire signed [9:0] m372_79;
   assign m372_79 =10'b0;

   // m372_80 = W*in
   wire signed [9:0] m372_80;
   assign m372_80 ={ {5{in372[5]}} , in372[5:1] };

   // m372_81 = W*in
   wire signed [9:0] m372_81;
   assign m372_81 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_82 = W*in
   wire signed [9:0] m372_82;
   assign m372_82 ={ {4{in372[5]}} , in372[5:0] };

   // m372_83 = W*in
   wire signed [9:0] m372_83;
   assign m372_83 ={ {5{in372[5]}} , in372[5:1] };

   // m372_84 = W*in
   wire signed [9:0] m372_84;
   assign m372_84 ={ {4{in372[5]}} , in372[5:0] };

   // m372_85 = W*in
   wire signed [9:0] m372_85;
   assign m372_85 =10'b0;

   // m372_86 = W*in
   wire signed [9:0] m372_86;
   assign m372_86 =10'b0;

   // m372_87 = W*in
   wire signed [9:0] m372_87;
   assign m372_87 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_88 = W*in
   wire signed [9:0] m372_88;
   assign m372_88 =10'b0;

   // m372_89 = W*in
   wire signed [9:0] m372_89;
   assign m372_89 =10'b0;

   // m372_90 = W*in
   wire signed [9:0] m372_90;
   assign m372_90 =10'b0;

   // m372_91 = W*in
   wire signed [9:0] m372_91;
   assign m372_91 =10'b0;

   // m372_92 = W*in
   wire signed [9:0] m372_92;
   assign m372_92 =10'b0;

   // m372_93 = W*in
   wire signed [9:0] m372_93;
   assign m372_93 ={ {4{in372[5]}} , in372[5:0] };

   // m372_94 = W*in
   wire signed [9:0] m372_94;
   assign m372_94 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_95 = W*in
   wire signed [9:0] m372_95;
   assign m372_95 ={ {4{in372[5]}} , in372[5:0] };

   // m372_96 = W*in
   wire signed [9:0] m372_96;
   assign m372_96 =10'b0;

   // m372_97 = W*in
   wire signed [9:0] m372_97;
   assign m372_97 =10'b0;

   // m372_98 = W*in
   wire signed [9:0] m372_98;
   assign m372_98 =10'b0;

   // m372_99 = W*in
   wire signed [9:0] m372_99;
   assign m372_99 ={ {4{neg372[5]}} , neg372[5:0] };

   // m372_100 = W*in
   wire signed [9:0] m372_100;
   assign m372_100 =10'b0;

   // m372_101 = W*in
   wire signed [9:0] m372_101;
   assign m372_101 =10'b0;

   // m372_102 = W*in
   wire signed [9:0] m372_102;
   assign m372_102 =10'b0;

   // m372_103 = W*in
   wire signed [9:0] m372_103;
   assign m372_103 =10'b0;

   // m372_104 = W*in
   wire signed [9:0] m372_104;
   assign m372_104 =10'b0;

   // m372_105 = W*in
   wire signed [9:0] m372_105;
   assign m372_105 =10'b0;

   // m372_106 = W*in
   wire signed [9:0] m372_106;
   assign m372_106 =10'b0;

   // m372_107 = W*in
   wire signed [9:0] m372_107;
   assign m372_107 ={ {5{in372[5]}} , in372[5:1] };

   // m372_108 = W*in
   wire signed [9:0] m372_108;
   assign m372_108 =10'b0;

   // m372_109 = W*in
   wire signed [9:0] m372_109;
   assign m372_109 =10'b0;

   // m372_110 = W*in
   wire signed [9:0] m372_110;
   assign m372_110 =10'b0;

   // m372_111 = W*in
   wire signed [9:0] m372_111;
   assign m372_111 =10'b0;

   // m372_112 = W*in
   wire signed [9:0] m372_112;
   assign m372_112 =10'b0;

   // m372_113 = W*in
   wire signed [9:0] m372_113;
   assign m372_113 =10'b0;

   // m372_114 = W*in
   wire signed [9:0] m372_114;
   assign m372_114 =10'b0;

   // m372_115 = W*in
   wire signed [9:0] m372_115;
   assign m372_115 ={ {5{neg372[5]}} , neg372[5:1] };

   // m372_116 = W*in
   wire signed [9:0] m372_116;
   assign m372_116 =10'b0;

   // m372_117 = W*in
   wire signed [9:0] m372_117;
   assign m372_117 =10'b0;

   // m373_1 = W*in
   wire signed [9:0] m373_1;
   assign m373_1 =10'b0;

   // m373_2 = W*in
   wire signed [9:0] m373_2;
   assign m373_2 =10'b0;

   // m373_3 = W*in
   wire signed [9:0] m373_3;
   assign m373_3 ={ {4{in373[5]}} , in373[5:0] };

   // m373_4 = W*in
   wire signed [9:0] m373_4;
   assign m373_4 =10'b0;

   // m373_5 = W*in
   wire signed [9:0] m373_5;
   assign m373_5 =10'b0;

   // m373_6 = W*in
   wire signed [9:0] m373_6;
   assign m373_6 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_7 = W*in
   wire signed [9:0] m373_7;
   assign m373_7 =10'b0;

   // m373_8 = W*in
   wire signed [9:0] m373_8;
   assign m373_8 =10'b0;

   // m373_9 = W*in
   wire signed [9:0] m373_9;
   assign m373_9 =10'b0;

   // m373_10 = W*in
   wire signed [9:0] m373_10;
   assign m373_10 ={ {4{in373[5]}} , in373[5:0] };

   // m373_11 = W*in
   wire signed [9:0] m373_11;
   assign m373_11 ={ {4{in373[5]}} , in373[5:0] };

   // m373_12 = W*in
   wire signed [9:0] m373_12;
   assign m373_12 =10'b0;

   // m373_13 = W*in
   wire signed [9:0] m373_13;
   assign m373_13 =10'b0;

   // m373_14 = W*in
   wire signed [9:0] m373_14;
   assign m373_14 =10'b0;

   // m373_15 = W*in
   wire signed [9:0] m373_15;
   assign m373_15 =10'b0;

   // m373_16 = W*in
   wire signed [9:0] m373_16;
   assign m373_16 =10'b0;

   // m373_17 = W*in
   wire signed [9:0] m373_17;
   assign m373_17 ={ {4{in373[5]}} , in373[5:0] };

   // m373_18 = W*in
   wire signed [9:0] m373_18;
   assign m373_18 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_19 = W*in
   wire signed [9:0] m373_19;
   assign m373_19 =10'b0;

   // m373_20 = W*in
   wire signed [9:0] m373_20;
   assign m373_20 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_21 = W*in
   wire signed [9:0] m373_21;
   assign m373_21 ={ {4{in373[5]}} , in373[5:0] };

   // m373_22 = W*in
   wire signed [9:0] m373_22;
   assign m373_22 =10'b0;

   // m373_23 = W*in
   wire signed [9:0] m373_23;
   assign m373_23 =10'b0;

   // m373_24 = W*in
   wire signed [9:0] m373_24;
   assign m373_24 =10'b0;

   // m373_25 = W*in
   wire signed [9:0] m373_25;
   assign m373_25 =10'b0;

   // m373_26 = W*in
   wire signed [9:0] m373_26;
   assign m373_26 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_27 = W*in
   wire signed [9:0] m373_27;
   assign m373_27 ={ {5{neg373[5]}} , neg373[5:1] };

   // m373_28 = W*in
   wire signed [9:0] m373_28;
   assign m373_28 =10'b0;

   // m373_29 = W*in
   wire signed [9:0] m373_29;
   assign m373_29 =10'b0;

   // m373_30 = W*in
   wire signed [9:0] m373_30;
   assign m373_30 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_31 = W*in
   wire signed [9:0] m373_31;
   assign m373_31 =10'b0;

   // m373_32 = W*in
   wire signed [9:0] m373_32;
   assign m373_32 =10'b0;

   // m373_33 = W*in
   wire signed [9:0] m373_33;
   assign m373_33 =10'b0;

   // m373_34 = W*in
   wire signed [9:0] m373_34;
   assign m373_34 =10'b0;

   // m373_35 = W*in
   wire signed [9:0] m373_35;
   assign m373_35 ={ {5{neg373[5]}} , neg373[5:1] };

   // m373_36 = W*in
   wire signed [9:0] m373_36;
   assign m373_36 =10'b0;

   // m373_37 = W*in
   wire signed [9:0] m373_37;
   assign m373_37 =10'b0;

   // m373_38 = W*in
   wire signed [9:0] m373_38;
   assign m373_38 =10'b0;

   // m373_39 = W*in
   wire signed [9:0] m373_39;
   assign m373_39 =10'b0;

   // m373_40 = W*in
   wire signed [9:0] m373_40;
   assign m373_40 =10'b0;

   // m373_41 = W*in
   wire signed [9:0] m373_41;
   assign m373_41 ={ {4{in373[5]}} , in373[5:0] };

   // m373_42 = W*in
   wire signed [9:0] m373_42;
   assign m373_42 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_43 = W*in
   wire signed [9:0] m373_43;
   assign m373_43 =10'b0;

   // m373_44 = W*in
   wire signed [9:0] m373_44;
   assign m373_44 =10'b0;

   // m373_45 = W*in
   wire signed [9:0] m373_45;
   assign m373_45 =10'b0;

   // m373_46 = W*in
   wire signed [9:0] m373_46;
   assign m373_46 =10'b0;

   // m373_47 = W*in
   wire signed [9:0] m373_47;
   assign m373_47 =10'b0;

   // m373_48 = W*in
   wire signed [9:0] m373_48;
   assign m373_48 =10'b0;

   // m373_49 = W*in
   wire signed [9:0] m373_49;
   assign m373_49 =10'b0;

   // m373_50 = W*in
   wire signed [9:0] m373_50;
   assign m373_50 =10'b0;

   // m373_51 = W*in
   wire signed [9:0] m373_51;
   assign m373_51 =10'b0;

   // m373_52 = W*in
   wire signed [9:0] m373_52;
   assign m373_52 =10'b0;

   // m373_53 = W*in
   wire signed [9:0] m373_53;
   assign m373_53 =10'b0;

   // m373_54 = W*in
   wire signed [9:0] m373_54;
   assign m373_54 =10'b0;

   // m373_55 = W*in
   wire signed [9:0] m373_55;
   assign m373_55 =10'b0;

   // m373_56 = W*in
   wire signed [9:0] m373_56;
   assign m373_56 =10'b0;

   // m373_57 = W*in
   wire signed [9:0] m373_57;
   assign m373_57 =10'b0;

   // m373_58 = W*in
   wire signed [9:0] m373_58;
   assign m373_58 =10'b0;

   // m373_59 = W*in
   wire signed [9:0] m373_59;
   assign m373_59 =10'b0;

   // m373_60 = W*in
   wire signed [9:0] m373_60;
   assign m373_60 =10'b0;

   // m373_61 = W*in
   wire signed [9:0] m373_61;
   assign m373_61 =10'b0;

   // m373_62 = W*in
   wire signed [9:0] m373_62;
   assign m373_62 =10'b0;

   // m373_63 = W*in
   wire signed [9:0] m373_63;
   assign m373_63 =10'b0;

   // m373_64 = W*in
   wire signed [9:0] m373_64;
   assign m373_64 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_65 = W*in
   wire signed [9:0] m373_65;
   assign m373_65 =10'b0;

   // m373_66 = W*in
   wire signed [9:0] m373_66;
   assign m373_66 =10'b0;

   // m373_67 = W*in
   wire signed [9:0] m373_67;
   assign m373_67 =10'b0;

   // m373_68 = W*in
   wire signed [9:0] m373_68;
   assign m373_68 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_69 = W*in
   wire signed [9:0] m373_69;
   assign m373_69 ={ {4{in373[5]}} , in373[5:0] };

   // m373_70 = W*in
   wire signed [9:0] m373_70;
   assign m373_70 =10'b0;

   // m373_71 = W*in
   wire signed [9:0] m373_71;
   assign m373_71 ={ {5{in373[5]}} , in373[5:1] };

   // m373_72 = W*in
   wire signed [9:0] m373_72;
   assign m373_72 =10'b0;

   // m373_73 = W*in
   wire signed [9:0] m373_73;
   assign m373_73 ={ {5{neg373[5]}} , neg373[5:1] };

   // m373_74 = W*in
   wire signed [9:0] m373_74;
   assign m373_74 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_75 = W*in
   wire signed [9:0] m373_75;
   assign m373_75 =10'b0;

   // m373_76 = W*in
   wire signed [9:0] m373_76;
   assign m373_76 =10'b0;

   // m373_77 = W*in
   wire signed [9:0] m373_77;
   assign m373_77 =10'b0;

   // m373_78 = W*in
   wire signed [9:0] m373_78;
   assign m373_78 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_79 = W*in
   wire signed [9:0] m373_79;
   assign m373_79 ={ {4{in373[5]}} , in373[5:0] };

   // m373_80 = W*in
   wire signed [9:0] m373_80;
   assign m373_80 =10'b0;

   // m373_81 = W*in
   wire signed [9:0] m373_81;
   assign m373_81 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_82 = W*in
   wire signed [9:0] m373_82;
   assign m373_82 ={ {3{in373[5]}} , in373 , {1{1'b0}} };

   // m373_83 = W*in
   wire signed [9:0] m373_83;
   assign m373_83 ={ {4{in373[5]}} , in373[5:0] };

   // m373_84 = W*in
   wire signed [9:0] m373_84;
   assign m373_84 ={ {5{in373[5]}} , in373[5:1] };

   // m373_85 = W*in
   wire signed [9:0] m373_85;
   assign m373_85 ={ {4{in373[5]}} , in373[5:0] };

   // m373_86 = W*in
   wire signed [9:0] m373_86;
   assign m373_86 =10'b0;

   // m373_87 = W*in
   wire signed [9:0] m373_87;
   assign m373_87 =10'b0;

   // m373_88 = W*in
   wire signed [9:0] m373_88;
   assign m373_88 =10'b0;

   // m373_89 = W*in
   wire signed [9:0] m373_89;
   assign m373_89 =10'b0;

   // m373_90 = W*in
   wire signed [9:0] m373_90;
   assign m373_90 =10'b0;

   // m373_91 = W*in
   wire signed [9:0] m373_91;
   assign m373_91 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_92 = W*in
   wire signed [9:0] m373_92;
   assign m373_92 =10'b0;

   // m373_93 = W*in
   wire signed [9:0] m373_93;
   assign m373_93 =10'b0;

   // m373_94 = W*in
   wire signed [9:0] m373_94;
   assign m373_94 ={ {4{neg373[5]}} , neg373[5:0] };

   // m373_95 = W*in
   wire signed [9:0] m373_95;
   assign m373_95 ={ {4{in373[5]}} , in373[5:0] };

   // m373_96 = W*in
   wire signed [9:0] m373_96;
   assign m373_96 =10'b0;

   // m373_97 = W*in
   wire signed [9:0] m373_97;
   assign m373_97 =10'b0;

   // m373_98 = W*in
   wire signed [9:0] m373_98;
   assign m373_98 =10'b0;

   // m373_99 = W*in
   wire signed [9:0] m373_99;
   assign m373_99 =10'b0;

   // m373_100 = W*in
   wire signed [9:0] m373_100;
   assign m373_100 =10'b0;

   // m373_101 = W*in
   wire signed [9:0] m373_101;
   assign m373_101 =10'b0;

   // m373_102 = W*in
   wire signed [9:0] m373_102;
   assign m373_102 =10'b0;

   // m373_103 = W*in
   wire signed [9:0] m373_103;
   assign m373_103 =10'b0;

   // m373_104 = W*in
   wire signed [9:0] m373_104;
   assign m373_104 =10'b0;

   // m373_105 = W*in
   wire signed [9:0] m373_105;
   assign m373_105 =10'b0;

   // m373_106 = W*in
   wire signed [9:0] m373_106;
   assign m373_106 ={ {5{neg373[5]}} , neg373[5:1] };

   // m373_107 = W*in
   wire signed [9:0] m373_107;
   assign m373_107 ={ {5{in373[5]}} , in373[5:1] };

   // m373_108 = W*in
   wire signed [9:0] m373_108;
   assign m373_108 ={ {4{in373[5]}} , in373[5:0] };

   // m373_109 = W*in
   wire signed [9:0] m373_109;
   assign m373_109 ={ {5{in373[5]}} , in373[5:1] };

   // m373_110 = W*in
   wire signed [9:0] m373_110;
   assign m373_110 ={ {4{in373[5]}} , in373[5:0] };

   // m373_111 = W*in
   wire signed [9:0] m373_111;
   assign m373_111 =10'b0;

   // m373_112 = W*in
   wire signed [9:0] m373_112;
   assign m373_112 =10'b0;

   // m373_113 = W*in
   wire signed [9:0] m373_113;
   assign m373_113 ={ {5{neg373[5]}} , neg373[5:1] };

   // m373_114 = W*in
   wire signed [9:0] m373_114;
   assign m373_114 =10'b0;

   // m373_115 = W*in
   wire signed [9:0] m373_115;
   assign m373_115 ={ {5{neg373[5]}} , neg373[5:1] };

   // m373_116 = W*in
   wire signed [9:0] m373_116;
   assign m373_116 =10'b0;

   // m373_117 = W*in
   wire signed [9:0] m373_117;
   assign m373_117 ={ {4{neg373[5]}} , neg373[5:0] };

   // m374_1 = W*in
   wire signed [9:0] m374_1;
   assign m374_1 =10'b0;

   // m374_2 = W*in
   wire signed [9:0] m374_2;
   assign m374_2 =10'b0;

   // m374_3 = W*in
   wire signed [9:0] m374_3;
   assign m374_3 =10'b0;

   // m374_4 = W*in
   wire signed [9:0] m374_4;
   assign m374_4 =10'b0;

   // m374_5 = W*in
   wire signed [9:0] m374_5;
   assign m374_5 =10'b0;

   // m374_6 = W*in
   wire signed [9:0] m374_6;
   assign m374_6 =10'b0;

   // m374_7 = W*in
   wire signed [9:0] m374_7;
   assign m374_7 =10'b0;

   // m374_8 = W*in
   wire signed [9:0] m374_8;
   assign m374_8 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_9 = W*in
   wire signed [9:0] m374_9;
   assign m374_9 =10'b0;

   // m374_10 = W*in
   wire signed [9:0] m374_10;
   assign m374_10 =10'b0;

   // m374_11 = W*in
   wire signed [9:0] m374_11;
   assign m374_11 ={ {4{in374[5]}} , in374[5:0] };

   // m374_12 = W*in
   wire signed [9:0] m374_12;
   assign m374_12 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_13 = W*in
   wire signed [9:0] m374_13;
   assign m374_13 =10'b0;

   // m374_14 = W*in
   wire signed [9:0] m374_14;
   assign m374_14 =10'b0;

   // m374_15 = W*in
   wire signed [9:0] m374_15;
   assign m374_15 =10'b0;

   // m374_16 = W*in
   wire signed [9:0] m374_16;
   assign m374_16 ={ {5{neg374[5]}} , neg374[5:1] };

   // m374_17 = W*in
   wire signed [9:0] m374_17;
   assign m374_17 ={ {5{in374[5]}} , in374[5:1] };

   // m374_18 = W*in
   wire signed [9:0] m374_18;
   assign m374_18 =10'b0;

   // m374_19 = W*in
   wire signed [9:0] m374_19;
   assign m374_19 =10'b0;

   // m374_20 = W*in
   wire signed [9:0] m374_20;
   assign m374_20 =10'b0;

   // m374_21 = W*in
   wire signed [9:0] m374_21;
   assign m374_21 =10'b0;

   // m374_22 = W*in
   wire signed [9:0] m374_22;
   assign m374_22 =10'b0;

   // m374_23 = W*in
   wire signed [9:0] m374_23;
   assign m374_23 =10'b0;

   // m374_24 = W*in
   wire signed [9:0] m374_24;
   assign m374_24 =10'b0;

   // m374_25 = W*in
   wire signed [9:0] m374_25;
   assign m374_25 ={ {5{neg374[5]}} , neg374[5:1] };

   // m374_26 = W*in
   wire signed [9:0] m374_26;
   assign m374_26 =10'b0;

   // m374_27 = W*in
   wire signed [9:0] m374_27;
   assign m374_27 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_28 = W*in
   wire signed [9:0] m374_28;
   assign m374_28 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_29 = W*in
   wire signed [9:0] m374_29;
   assign m374_29 =10'b0;

   // m374_30 = W*in
   wire signed [9:0] m374_30;
   assign m374_30 ={ {5{neg374[5]}} , neg374[5:1] };

   // m374_31 = W*in
   wire signed [9:0] m374_31;
   assign m374_31 =10'b0;

   // m374_32 = W*in
   wire signed [9:0] m374_32;
   assign m374_32 ={ {4{in374[5]}} , in374[5:0] };

   // m374_33 = W*in
   wire signed [9:0] m374_33;
   assign m374_33 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_34 = W*in
   wire signed [9:0] m374_34;
   assign m374_34 =10'b0;

   // m374_35 = W*in
   wire signed [9:0] m374_35;
   assign m374_35 =10'b0;

   // m374_36 = W*in
   wire signed [9:0] m374_36;
   assign m374_36 =10'b0;

   // m374_37 = W*in
   wire signed [9:0] m374_37;
   assign m374_37 =10'b0;

   // m374_38 = W*in
   wire signed [9:0] m374_38;
   assign m374_38 =10'b0;

   // m374_39 = W*in
   wire signed [9:0] m374_39;
   assign m374_39 =10'b0;

   // m374_40 = W*in
   wire signed [9:0] m374_40;
   assign m374_40 =10'b0;

   // m374_41 = W*in
   wire signed [9:0] m374_41;
   assign m374_41 =10'b0;

   // m374_42 = W*in
   wire signed [9:0] m374_42;
   assign m374_42 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_43 = W*in
   wire signed [9:0] m374_43;
   assign m374_43 =10'b0;

   // m374_44 = W*in
   wire signed [9:0] m374_44;
   assign m374_44 =10'b0;

   // m374_45 = W*in
   wire signed [9:0] m374_45;
   assign m374_45 =10'b0;

   // m374_46 = W*in
   wire signed [9:0] m374_46;
   assign m374_46 =10'b0;

   // m374_47 = W*in
   wire signed [9:0] m374_47;
   assign m374_47 =10'b0;

   // m374_48 = W*in
   wire signed [9:0] m374_48;
   assign m374_48 =10'b0;

   // m374_49 = W*in
   wire signed [9:0] m374_49;
   assign m374_49 ={ {4{in374[5]}} , in374[5:0] };

   // m374_50 = W*in
   wire signed [9:0] m374_50;
   assign m374_50 =10'b0;

   // m374_51 = W*in
   wire signed [9:0] m374_51;
   assign m374_51 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_52 = W*in
   wire signed [9:0] m374_52;
   assign m374_52 =10'b0;

   // m374_53 = W*in
   wire signed [9:0] m374_53;
   assign m374_53 =10'b0;

   // m374_54 = W*in
   wire signed [9:0] m374_54;
   assign m374_54 =10'b0;

   // m374_55 = W*in
   wire signed [9:0] m374_55;
   assign m374_55 =10'b0;

   // m374_56 = W*in
   wire signed [9:0] m374_56;
   assign m374_56 =10'b0;

   // m374_57 = W*in
   wire signed [9:0] m374_57;
   assign m374_57 ={ {4{in374[5]}} , in374[5:0] };

   // m374_58 = W*in
   wire signed [9:0] m374_58;
   assign m374_58 =10'b0;

   // m374_59 = W*in
   wire signed [9:0] m374_59;
   assign m374_59 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_60 = W*in
   wire signed [9:0] m374_60;
   assign m374_60 =10'b0;

   // m374_61 = W*in
   wire signed [9:0] m374_61;
   assign m374_61 ={ {5{in374[5]}} , in374[5:1] };

   // m374_62 = W*in
   wire signed [9:0] m374_62;
   assign m374_62 =10'b0;

   // m374_63 = W*in
   wire signed [9:0] m374_63;
   assign m374_63 ={ {4{in374[5]}} , in374[5:0] };

   // m374_64 = W*in
   wire signed [9:0] m374_64;
   assign m374_64 ={ {5{neg374[5]}} , neg374[5:1] };

   // m374_65 = W*in
   wire signed [9:0] m374_65;
   assign m374_65 ={ {5{neg374[5]}} , neg374[5:1] };

   // m374_66 = W*in
   wire signed [9:0] m374_66;
   assign m374_66 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_67 = W*in
   wire signed [9:0] m374_67;
   assign m374_67 =10'b0;

   // m374_68 = W*in
   wire signed [9:0] m374_68;
   assign m374_68 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_69 = W*in
   wire signed [9:0] m374_69;
   assign m374_69 ={ {4{in374[5]}} , in374[5:0] };

   // m374_70 = W*in
   wire signed [9:0] m374_70;
   assign m374_70 ={ {4{in374[5]}} , in374[5:0] };

   // m374_71 = W*in
   wire signed [9:0] m374_71;
   assign m374_71 ={ {5{in374[5]}} , in374[5:1] };

   // m374_72 = W*in
   wire signed [9:0] m374_72;
   assign m374_72 ={ {4{in374[5]}} , in374[5:0] };

   // m374_73 = W*in
   wire signed [9:0] m374_73;
   assign m374_73 =10'b0;

   // m374_74 = W*in
   wire signed [9:0] m374_74;
   assign m374_74 ={ {5{in374[5]}} , in374[5:1] };

   // m374_75 = W*in
   wire signed [9:0] m374_75;
   assign m374_75 =10'b0;

   // m374_76 = W*in
   wire signed [9:0] m374_76;
   assign m374_76 =10'b0;

   // m374_77 = W*in
   wire signed [9:0] m374_77;
   assign m374_77 =10'b0;

   // m374_78 = W*in
   wire signed [9:0] m374_78;
   assign m374_78 =10'b0;

   // m374_79 = W*in
   wire signed [9:0] m374_79;
   assign m374_79 =10'b0;

   // m374_80 = W*in
   wire signed [9:0] m374_80;
   assign m374_80 ={ {5{neg374[5]}} , neg374[5:1] };

   // m374_81 = W*in
   wire signed [9:0] m374_81;
   assign m374_81 =10'b0;

   // m374_82 = W*in
   wire signed [9:0] m374_82;
   assign m374_82 =10'b0;

   // m374_83 = W*in
   wire signed [9:0] m374_83;
   assign m374_83 ={ {5{in374[5]}} , in374[5:1] };

   // m374_84 = W*in
   wire signed [9:0] m374_84;
   assign m374_84 ={ {4{in374[5]}} , in374[5:0] };

   // m374_85 = W*in
   wire signed [9:0] m374_85;
   assign m374_85 =10'b0;

   // m374_86 = W*in
   wire signed [9:0] m374_86;
   assign m374_86 =10'b0;

   // m374_87 = W*in
   wire signed [9:0] m374_87;
   assign m374_87 ={ {4{in374[5]}} , in374[5:0] };

   // m374_88 = W*in
   wire signed [9:0] m374_88;
   assign m374_88 =10'b0;

   // m374_89 = W*in
   wire signed [9:0] m374_89;
   assign m374_89 =10'b0;

   // m374_90 = W*in
   wire signed [9:0] m374_90;
   assign m374_90 =10'b0;

   // m374_91 = W*in
   wire signed [9:0] m374_91;
   assign m374_91 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_92 = W*in
   wire signed [9:0] m374_92;
   assign m374_92 =10'b0;

   // m374_93 = W*in
   wire signed [9:0] m374_93;
   assign m374_93 ={ {5{in374[5]}} , in374[5:1] };

   // m374_94 = W*in
   wire signed [9:0] m374_94;
   assign m374_94 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_95 = W*in
   wire signed [9:0] m374_95;
   assign m374_95 ={ {4{in374[5]}} , in374[5:0] };

   // m374_96 = W*in
   wire signed [9:0] m374_96;
   assign m374_96 =10'b0;

   // m374_97 = W*in
   wire signed [9:0] m374_97;
   assign m374_97 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_98 = W*in
   wire signed [9:0] m374_98;
   assign m374_98 =10'b0;

   // m374_99 = W*in
   wire signed [9:0] m374_99;
   assign m374_99 =10'b0;

   // m374_100 = W*in
   wire signed [9:0] m374_100;
   assign m374_100 =10'b0;

   // m374_101 = W*in
   wire signed [9:0] m374_101;
   assign m374_101 =10'b0;

   // m374_102 = W*in
   wire signed [9:0] m374_102;
   assign m374_102 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_103 = W*in
   wire signed [9:0] m374_103;
   assign m374_103 =10'b0;

   // m374_104 = W*in
   wire signed [9:0] m374_104;
   assign m374_104 =10'b0;

   // m374_105 = W*in
   wire signed [9:0] m374_105;
   assign m374_105 =10'b0;

   // m374_106 = W*in
   wire signed [9:0] m374_106;
   assign m374_106 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_107 = W*in
   wire signed [9:0] m374_107;
   assign m374_107 ={ {4{in374[5]}} , in374[5:0] };

   // m374_108 = W*in
   wire signed [9:0] m374_108;
   assign m374_108 =10'b0;

   // m374_109 = W*in
   wire signed [9:0] m374_109;
   assign m374_109 =10'b0;

   // m374_110 = W*in
   wire signed [9:0] m374_110;
   assign m374_110 =10'b0;

   // m374_111 = W*in
   wire signed [9:0] m374_111;
   assign m374_111 =10'b0;

   // m374_112 = W*in
   wire signed [9:0] m374_112;
   assign m374_112 ={ {4{neg374[5]}} , neg374[5:0] };

   // m374_113 = W*in
   wire signed [9:0] m374_113;
   assign m374_113 =10'b0;

   // m374_114 = W*in
   wire signed [9:0] m374_114;
   assign m374_114 =10'b0;

   // m374_115 = W*in
   wire signed [9:0] m374_115;
   assign m374_115 =10'b0;

   // m374_116 = W*in
   wire signed [9:0] m374_116;
   assign m374_116 =10'b0;

   // m374_117 = W*in
   wire signed [9:0] m374_117;
   assign m374_117 =10'b0;

   // m375_1 = W*in
   wire signed [9:0] m375_1;
   assign m375_1 =10'b0;

   // m375_2 = W*in
   wire signed [9:0] m375_2;
   assign m375_2 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_3 = W*in
   wire signed [9:0] m375_3;
   assign m375_3 =10'b0;

   // m375_4 = W*in
   wire signed [9:0] m375_4;
   assign m375_4 =10'b0;

   // m375_5 = W*in
   wire signed [9:0] m375_5;
   assign m375_5 =10'b0;

   // m375_6 = W*in
   wire signed [9:0] m375_6;
   assign m375_6 =10'b0;

   // m375_7 = W*in
   wire signed [9:0] m375_7;
   assign m375_7 =10'b0;

   // m375_8 = W*in
   wire signed [9:0] m375_8;
   assign m375_8 =10'b0;

   // m375_9 = W*in
   wire signed [9:0] m375_9;
   assign m375_9 =10'b0;

   // m375_10 = W*in
   wire signed [9:0] m375_10;
   assign m375_10 =10'b0;

   // m375_11 = W*in
   wire signed [9:0] m375_11;
   assign m375_11 =10'b0;

   // m375_12 = W*in
   wire signed [9:0] m375_12;
   assign m375_12 =10'b0;

   // m375_13 = W*in
   wire signed [9:0] m375_13;
   assign m375_13 =10'b0;

   // m375_14 = W*in
   wire signed [9:0] m375_14;
   assign m375_14 =10'b0;

   // m375_15 = W*in
   wire signed [9:0] m375_15;
   assign m375_15 =10'b0;

   // m375_16 = W*in
   wire signed [9:0] m375_16;
   assign m375_16 ={ {5{neg375[5]}} , neg375[5:1] };

   // m375_17 = W*in
   wire signed [9:0] m375_17;
   assign m375_17 =10'b0;

   // m375_18 = W*in
   wire signed [9:0] m375_18;
   assign m375_18 =10'b0;

   // m375_19 = W*in
   wire signed [9:0] m375_19;
   assign m375_19 =10'b0;

   // m375_20 = W*in
   wire signed [9:0] m375_20;
   assign m375_20 =10'b0;

   // m375_21 = W*in
   wire signed [9:0] m375_21;
   assign m375_21 ={ {5{neg375[5]}} , neg375[5:1] };

   // m375_22 = W*in
   wire signed [9:0] m375_22;
   assign m375_22 =10'b0;

   // m375_23 = W*in
   wire signed [9:0] m375_23;
   assign m375_23 =10'b0;

   // m375_24 = W*in
   wire signed [9:0] m375_24;
   assign m375_24 =10'b0;

   // m375_25 = W*in
   wire signed [9:0] m375_25;
   assign m375_25 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_26 = W*in
   wire signed [9:0] m375_26;
   assign m375_26 =10'b0;

   // m375_27 = W*in
   wire signed [9:0] m375_27;
   assign m375_27 =10'b0;

   // m375_28 = W*in
   wire signed [9:0] m375_28;
   assign m375_28 =10'b0;

   // m375_29 = W*in
   wire signed [9:0] m375_29;
   assign m375_29 =10'b0;

   // m375_30 = W*in
   wire signed [9:0] m375_30;
   assign m375_30 =10'b0;

   // m375_31 = W*in
   wire signed [9:0] m375_31;
   assign m375_31 =10'b0;

   // m375_32 = W*in
   wire signed [9:0] m375_32;
   assign m375_32 =10'b0;

   // m375_33 = W*in
   wire signed [9:0] m375_33;
   assign m375_33 =10'b0;

   // m375_34 = W*in
   wire signed [9:0] m375_34;
   assign m375_34 =10'b0;

   // m375_35 = W*in
   wire signed [9:0] m375_35;
   assign m375_35 ={ {5{neg375[5]}} , neg375[5:1] };

   // m375_36 = W*in
   wire signed [9:0] m375_36;
   assign m375_36 =10'b0;

   // m375_37 = W*in
   wire signed [9:0] m375_37;
   assign m375_37 =10'b0;

   // m375_38 = W*in
   wire signed [9:0] m375_38;
   assign m375_38 =10'b0;

   // m375_39 = W*in
   wire signed [9:0] m375_39;
   assign m375_39 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_40 = W*in
   wire signed [9:0] m375_40;
   assign m375_40 =10'b0;

   // m375_41 = W*in
   wire signed [9:0] m375_41;
   assign m375_41 =10'b0;

   // m375_42 = W*in
   wire signed [9:0] m375_42;
   assign m375_42 ={ {4{in375[5]}} , in375[5:0] };

   // m375_43 = W*in
   wire signed [9:0] m375_43;
   assign m375_43 =10'b0;

   // m375_44 = W*in
   wire signed [9:0] m375_44;
   assign m375_44 =10'b0;

   // m375_45 = W*in
   wire signed [9:0] m375_45;
   assign m375_45 =10'b0;

   // m375_46 = W*in
   wire signed [9:0] m375_46;
   assign m375_46 =10'b0;

   // m375_47 = W*in
   wire signed [9:0] m375_47;
   assign m375_47 =10'b0;

   // m375_48 = W*in
   wire signed [9:0] m375_48;
   assign m375_48 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_49 = W*in
   wire signed [9:0] m375_49;
   assign m375_49 =10'b0;

   // m375_50 = W*in
   wire signed [9:0] m375_50;
   assign m375_50 =10'b0;

   // m375_51 = W*in
   wire signed [9:0] m375_51;
   assign m375_51 =10'b0;

   // m375_52 = W*in
   wire signed [9:0] m375_52;
   assign m375_52 =10'b0;

   // m375_53 = W*in
   wire signed [9:0] m375_53;
   assign m375_53 =10'b0;

   // m375_54 = W*in
   wire signed [9:0] m375_54;
   assign m375_54 =10'b0;

   // m375_55 = W*in
   wire signed [9:0] m375_55;
   assign m375_55 =10'b0;

   // m375_56 = W*in
   wire signed [9:0] m375_56;
   assign m375_56 =10'b0;

   // m375_57 = W*in
   wire signed [9:0] m375_57;
   assign m375_57 ={ {4{in375[5]}} , in375[5:0] };

   // m375_58 = W*in
   wire signed [9:0] m375_58;
   assign m375_58 =10'b0;

   // m375_59 = W*in
   wire signed [9:0] m375_59;
   assign m375_59 =10'b0;

   // m375_60 = W*in
   wire signed [9:0] m375_60;
   assign m375_60 =10'b0;

   // m375_61 = W*in
   wire signed [9:0] m375_61;
   assign m375_61 =10'b0;

   // m375_62 = W*in
   wire signed [9:0] m375_62;
   assign m375_62 =10'b0;

   // m375_63 = W*in
   wire signed [9:0] m375_63;
   assign m375_63 =10'b0;

   // m375_64 = W*in
   wire signed [9:0] m375_64;
   assign m375_64 ={ {4{in375[5]}} , in375[5:0] };

   // m375_65 = W*in
   wire signed [9:0] m375_65;
   assign m375_65 ={ {4{in375[5]}} , in375[5:0] };

   // m375_66 = W*in
   wire signed [9:0] m375_66;
   assign m375_66 ={ {4{in375[5]}} , in375[5:0] };

   // m375_67 = W*in
   wire signed [9:0] m375_67;
   assign m375_67 =10'b0;

   // m375_68 = W*in
   wire signed [9:0] m375_68;
   assign m375_68 =10'b0;

   // m375_69 = W*in
   wire signed [9:0] m375_69;
   assign m375_69 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_70 = W*in
   wire signed [9:0] m375_70;
   assign m375_70 =10'b0;

   // m375_71 = W*in
   wire signed [9:0] m375_71;
   assign m375_71 ={ {5{in375[5]}} , in375[5:1] };

   // m375_72 = W*in
   wire signed [9:0] m375_72;
   assign m375_72 ={ {5{neg375[5]}} , neg375[5:1] };

   // m375_73 = W*in
   wire signed [9:0] m375_73;
   assign m375_73 =10'b0;

   // m375_74 = W*in
   wire signed [9:0] m375_74;
   assign m375_74 =10'b0;

   // m375_75 = W*in
   wire signed [9:0] m375_75;
   assign m375_75 =10'b0;

   // m375_76 = W*in
   wire signed [9:0] m375_76;
   assign m375_76 =10'b0;

   // m375_77 = W*in
   wire signed [9:0] m375_77;
   assign m375_77 =10'b0;

   // m375_78 = W*in
   wire signed [9:0] m375_78;
   assign m375_78 =10'b0;

   // m375_79 = W*in
   wire signed [9:0] m375_79;
   assign m375_79 =10'b0;

   // m375_80 = W*in
   wire signed [9:0] m375_80;
   assign m375_80 =10'b0;

   // m375_81 = W*in
   wire signed [9:0] m375_81;
   assign m375_81 ={ {5{in375[5]}} , in375[5:1] };

   // m375_82 = W*in
   wire signed [9:0] m375_82;
   assign m375_82 =10'b0;

   // m375_83 = W*in
   wire signed [9:0] m375_83;
   assign m375_83 =10'b0;

   // m375_84 = W*in
   wire signed [9:0] m375_84;
   assign m375_84 =10'b0;

   // m375_85 = W*in
   wire signed [9:0] m375_85;
   assign m375_85 =10'b0;

   // m375_86 = W*in
   wire signed [9:0] m375_86;
   assign m375_86 =10'b0;

   // m375_87 = W*in
   wire signed [9:0] m375_87;
   assign m375_87 =10'b0;

   // m375_88 = W*in
   wire signed [9:0] m375_88;
   assign m375_88 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_89 = W*in
   wire signed [9:0] m375_89;
   assign m375_89 =10'b0;

   // m375_90 = W*in
   wire signed [9:0] m375_90;
   assign m375_90 =10'b0;

   // m375_91 = W*in
   wire signed [9:0] m375_91;
   assign m375_91 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_92 = W*in
   wire signed [9:0] m375_92;
   assign m375_92 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_93 = W*in
   wire signed [9:0] m375_93;
   assign m375_93 =10'b0;

   // m375_94 = W*in
   wire signed [9:0] m375_94;
   assign m375_94 =10'b0;

   // m375_95 = W*in
   wire signed [9:0] m375_95;
   assign m375_95 =10'b0;

   // m375_96 = W*in
   wire signed [9:0] m375_96;
   assign m375_96 =10'b0;

   // m375_97 = W*in
   wire signed [9:0] m375_97;
   assign m375_97 =10'b0;

   // m375_98 = W*in
   wire signed [9:0] m375_98;
   assign m375_98 =10'b0;

   // m375_99 = W*in
   wire signed [9:0] m375_99;
   assign m375_99 =10'b0;

   // m375_100 = W*in
   wire signed [9:0] m375_100;
   assign m375_100 ={ {4{in375[5]}} , in375[5:0] };

   // m375_101 = W*in
   wire signed [9:0] m375_101;
   assign m375_101 =10'b0;

   // m375_102 = W*in
   wire signed [9:0] m375_102;
   assign m375_102 =10'b0;

   // m375_103 = W*in
   wire signed [9:0] m375_103;
   assign m375_103 =10'b0;

   // m375_104 = W*in
   wire signed [9:0] m375_104;
   assign m375_104 =10'b0;

   // m375_105 = W*in
   wire signed [9:0] m375_105;
   assign m375_105 =10'b0;

   // m375_106 = W*in
   wire signed [9:0] m375_106;
   assign m375_106 =10'b0;

   // m375_107 = W*in
   wire signed [9:0] m375_107;
   assign m375_107 ={ {4{in375[5]}} , in375[5:0] };

   // m375_108 = W*in
   wire signed [9:0] m375_108;
   assign m375_108 =10'b0;

   // m375_109 = W*in
   wire signed [9:0] m375_109;
   assign m375_109 ={ {3{neg375[5]}} , neg375 , {1{1'b0}} };

   // m375_110 = W*in
   wire signed [9:0] m375_110;
   assign m375_110 ={ {4{in375[5]}} , in375[5:0] };

   // m375_111 = W*in
   wire signed [9:0] m375_111;
   assign m375_111 =10'b0;

   // m375_112 = W*in
   wire signed [9:0] m375_112;
   assign m375_112 =10'b0;

   // m375_113 = W*in
   wire signed [9:0] m375_113;
   assign m375_113 ={ {4{neg375[5]}} , neg375[5:0] };

   // m375_114 = W*in
   wire signed [9:0] m375_114;
   assign m375_114 =10'b0;

   // m375_115 = W*in
   wire signed [9:0] m375_115;
   assign m375_115 =10'b0;

   // m375_116 = W*in
   wire signed [9:0] m375_116;
   assign m375_116 =10'b0;

   // m375_117 = W*in
   wire signed [9:0] m375_117;
   assign m375_117 =10'b0;

   // m376_1 = W*in
   wire signed [9:0] m376_1;
   assign m376_1 =10'b0;

   // m376_2 = W*in
   wire signed [9:0] m376_2;
   assign m376_2 =10'b0;

   // m376_3 = W*in
   wire signed [9:0] m376_3;
   assign m376_3 =10'b0;

   // m376_4 = W*in
   wire signed [9:0] m376_4;
   assign m376_4 =10'b0;

   // m376_5 = W*in
   wire signed [9:0] m376_5;
   assign m376_5 =10'b0;

   // m376_6 = W*in
   wire signed [9:0] m376_6;
   assign m376_6 =10'b0;

   // m376_7 = W*in
   wire signed [9:0] m376_7;
   assign m376_7 =10'b0;

   // m376_8 = W*in
   wire signed [9:0] m376_8;
   assign m376_8 =10'b0;

   // m376_9 = W*in
   wire signed [9:0] m376_9;
   assign m376_9 =10'b0;

   // m376_10 = W*in
   wire signed [9:0] m376_10;
   assign m376_10 =10'b0;

   // m376_11 = W*in
   wire signed [9:0] m376_11;
   assign m376_11 =10'b0;

   // m376_12 = W*in
   wire signed [9:0] m376_12;
   assign m376_12 =10'b0;

   // m376_13 = W*in
   wire signed [9:0] m376_13;
   assign m376_13 =10'b0;

   // m376_14 = W*in
   wire signed [9:0] m376_14;
   assign m376_14 =10'b0;

   // m376_15 = W*in
   wire signed [9:0] m376_15;
   assign m376_15 =10'b0;

   // m376_16 = W*in
   wire signed [9:0] m376_16;
   assign m376_16 ={ {5{neg376[5]}} , neg376[5:1] };

   // m376_17 = W*in
   wire signed [9:0] m376_17;
   assign m376_17 =10'b0;

   // m376_18 = W*in
   wire signed [9:0] m376_18;
   assign m376_18 =10'b0;

   // m376_19 = W*in
   wire signed [9:0] m376_19;
   assign m376_19 =10'b0;

   // m376_20 = W*in
   wire signed [9:0] m376_20;
   assign m376_20 =10'b0;

   // m376_21 = W*in
   wire signed [9:0] m376_21;
   assign m376_21 ={ {5{neg376[5]}} , neg376[5:1] };

   // m376_22 = W*in
   wire signed [9:0] m376_22;
   assign m376_22 =10'b0;

   // m376_23 = W*in
   wire signed [9:0] m376_23;
   assign m376_23 =10'b0;

   // m376_24 = W*in
   wire signed [9:0] m376_24;
   assign m376_24 =10'b0;

   // m376_25 = W*in
   wire signed [9:0] m376_25;
   assign m376_25 =10'b0;

   // m376_26 = W*in
   wire signed [9:0] m376_26;
   assign m376_26 =10'b0;

   // m376_27 = W*in
   wire signed [9:0] m376_27;
   assign m376_27 =10'b0;

   // m376_28 = W*in
   wire signed [9:0] m376_28;
   assign m376_28 =10'b0;

   // m376_29 = W*in
   wire signed [9:0] m376_29;
   assign m376_29 =10'b0;

   // m376_30 = W*in
   wire signed [9:0] m376_30;
   assign m376_30 =10'b0;

   // m376_31 = W*in
   wire signed [9:0] m376_31;
   assign m376_31 =10'b0;

   // m376_32 = W*in
   wire signed [9:0] m376_32;
   assign m376_32 =10'b0;

   // m376_33 = W*in
   wire signed [9:0] m376_33;
   assign m376_33 =10'b0;

   // m376_34 = W*in
   wire signed [9:0] m376_34;
   assign m376_34 =10'b0;

   // m376_35 = W*in
   wire signed [9:0] m376_35;
   assign m376_35 =10'b0;

   // m376_36 = W*in
   wire signed [9:0] m376_36;
   assign m376_36 =10'b0;

   // m376_37 = W*in
   wire signed [9:0] m376_37;
   assign m376_37 =10'b0;

   // m376_38 = W*in
   wire signed [9:0] m376_38;
   assign m376_38 =10'b0;

   // m376_39 = W*in
   wire signed [9:0] m376_39;
   assign m376_39 =10'b0;

   // m376_40 = W*in
   wire signed [9:0] m376_40;
   assign m376_40 =10'b0;

   // m376_41 = W*in
   wire signed [9:0] m376_41;
   assign m376_41 =10'b0;

   // m376_42 = W*in
   wire signed [9:0] m376_42;
   assign m376_42 =10'b0;

   // m376_43 = W*in
   wire signed [9:0] m376_43;
   assign m376_43 =10'b0;

   // m376_44 = W*in
   wire signed [9:0] m376_44;
   assign m376_44 =10'b0;

   // m376_45 = W*in
   wire signed [9:0] m376_45;
   assign m376_45 =10'b0;

   // m376_46 = W*in
   wire signed [9:0] m376_46;
   assign m376_46 =10'b0;

   // m376_47 = W*in
   wire signed [9:0] m376_47;
   assign m376_47 =10'b0;

   // m376_48 = W*in
   wire signed [9:0] m376_48;
   assign m376_48 =10'b0;

   // m376_49 = W*in
   wire signed [9:0] m376_49;
   assign m376_49 =10'b0;

   // m376_50 = W*in
   wire signed [9:0] m376_50;
   assign m376_50 =10'b0;

   // m376_51 = W*in
   wire signed [9:0] m376_51;
   assign m376_51 =10'b0;

   // m376_52 = W*in
   wire signed [9:0] m376_52;
   assign m376_52 =10'b0;

   // m376_53 = W*in
   wire signed [9:0] m376_53;
   assign m376_53 =10'b0;

   // m376_54 = W*in
   wire signed [9:0] m376_54;
   assign m376_54 =10'b0;

   // m376_55 = W*in
   wire signed [9:0] m376_55;
   assign m376_55 =10'b0;

   // m376_56 = W*in
   wire signed [9:0] m376_56;
   assign m376_56 =10'b0;

   // m376_57 = W*in
   wire signed [9:0] m376_57;
   assign m376_57 =10'b0;

   // m376_58 = W*in
   wire signed [9:0] m376_58;
   assign m376_58 =10'b0;

   // m376_59 = W*in
   wire signed [9:0] m376_59;
   assign m376_59 =10'b0;

   // m376_60 = W*in
   wire signed [9:0] m376_60;
   assign m376_60 =10'b0;

   // m376_61 = W*in
   wire signed [9:0] m376_61;
   assign m376_61 =10'b0;

   // m376_62 = W*in
   wire signed [9:0] m376_62;
   assign m376_62 =10'b0;

   // m376_63 = W*in
   wire signed [9:0] m376_63;
   assign m376_63 ={ {5{neg376[5]}} , neg376[5:1] };

   // m376_64 = W*in
   wire signed [9:0] m376_64;
   assign m376_64 ={ {5{in376[5]}} , in376[5:1] };

   // m376_65 = W*in
   wire signed [9:0] m376_65;
   assign m376_65 =10'b0;

   // m376_66 = W*in
   wire signed [9:0] m376_66;
   assign m376_66 =10'b0;

   // m376_67 = W*in
   wire signed [9:0] m376_67;
   assign m376_67 =10'b0;

   // m376_68 = W*in
   wire signed [9:0] m376_68;
   assign m376_68 =10'b0;

   // m376_69 = W*in
   wire signed [9:0] m376_69;
   assign m376_69 ={ {4{neg376[5]}} , neg376[5:0] };

   // m376_70 = W*in
   wire signed [9:0] m376_70;
   assign m376_70 =10'b0;

   // m376_71 = W*in
   wire signed [9:0] m376_71;
   assign m376_71 =10'b0;

   // m376_72 = W*in
   wire signed [9:0] m376_72;
   assign m376_72 ={ {5{neg376[5]}} , neg376[5:1] };

   // m376_73 = W*in
   wire signed [9:0] m376_73;
   assign m376_73 ={ {5{in376[5]}} , in376[5:1] };

   // m376_74 = W*in
   wire signed [9:0] m376_74;
   assign m376_74 ={ {5{neg376[5]}} , neg376[5:1] };

   // m376_75 = W*in
   wire signed [9:0] m376_75;
   assign m376_75 =10'b0;

   // m376_76 = W*in
   wire signed [9:0] m376_76;
   assign m376_76 =10'b0;

   // m376_77 = W*in
   wire signed [9:0] m376_77;
   assign m376_77 =10'b0;

   // m376_78 = W*in
   wire signed [9:0] m376_78;
   assign m376_78 =10'b0;

   // m376_79 = W*in
   wire signed [9:0] m376_79;
   assign m376_79 =10'b0;

   // m376_80 = W*in
   wire signed [9:0] m376_80;
   assign m376_80 =10'b0;

   // m376_81 = W*in
   wire signed [9:0] m376_81;
   assign m376_81 =10'b0;

   // m376_82 = W*in
   wire signed [9:0] m376_82;
   assign m376_82 =10'b0;

   // m376_83 = W*in
   wire signed [9:0] m376_83;
   assign m376_83 =10'b0;

   // m376_84 = W*in
   wire signed [9:0] m376_84;
   assign m376_84 =10'b0;

   // m376_85 = W*in
   wire signed [9:0] m376_85;
   assign m376_85 =10'b0;

   // m376_86 = W*in
   wire signed [9:0] m376_86;
   assign m376_86 =10'b0;

   // m376_87 = W*in
   wire signed [9:0] m376_87;
   assign m376_87 =10'b0;

   // m376_88 = W*in
   wire signed [9:0] m376_88;
   assign m376_88 =10'b0;

   // m376_89 = W*in
   wire signed [9:0] m376_89;
   assign m376_89 =10'b0;

   // m376_90 = W*in
   wire signed [9:0] m376_90;
   assign m376_90 =10'b0;

   // m376_91 = W*in
   wire signed [9:0] m376_91;
   assign m376_91 ={ {4{neg376[5]}} , neg376[5:0] };

   // m376_92 = W*in
   wire signed [9:0] m376_92;
   assign m376_92 =10'b0;

   // m376_93 = W*in
   wire signed [9:0] m376_93;
   assign m376_93 =10'b0;

   // m376_94 = W*in
   wire signed [9:0] m376_94;
   assign m376_94 =10'b0;

   // m376_95 = W*in
   wire signed [9:0] m376_95;
   assign m376_95 =10'b0;

   // m376_96 = W*in
   wire signed [9:0] m376_96;
   assign m376_96 =10'b0;

   // m376_97 = W*in
   wire signed [9:0] m376_97;
   assign m376_97 =10'b0;

   // m376_98 = W*in
   wire signed [9:0] m376_98;
   assign m376_98 =10'b0;

   // m376_99 = W*in
   wire signed [9:0] m376_99;
   assign m376_99 =10'b0;

   // m376_100 = W*in
   wire signed [9:0] m376_100;
   assign m376_100 =10'b0;

   // m376_101 = W*in
   wire signed [9:0] m376_101;
   assign m376_101 =10'b0;

   // m376_102 = W*in
   wire signed [9:0] m376_102;
   assign m376_102 =10'b0;

   // m376_103 = W*in
   wire signed [9:0] m376_103;
   assign m376_103 =10'b0;

   // m376_104 = W*in
   wire signed [9:0] m376_104;
   assign m376_104 =10'b0;

   // m376_105 = W*in
   wire signed [9:0] m376_105;
   assign m376_105 =10'b0;

   // m376_106 = W*in
   wire signed [9:0] m376_106;
   assign m376_106 =10'b0;

   // m376_107 = W*in
   wire signed [9:0] m376_107;
   assign m376_107 ={ {5{in376[5]}} , in376[5:1] };

   // m376_108 = W*in
   wire signed [9:0] m376_108;
   assign m376_108 =10'b0;

   // m376_109 = W*in
   wire signed [9:0] m376_109;
   assign m376_109 =10'b0;

   // m376_110 = W*in
   wire signed [9:0] m376_110;
   assign m376_110 =10'b0;

   // m376_111 = W*in
   wire signed [9:0] m376_111;
   assign m376_111 =10'b0;

   // m376_112 = W*in
   wire signed [9:0] m376_112;
   assign m376_112 =10'b0;

   // m376_113 = W*in
   wire signed [9:0] m376_113;
   assign m376_113 =10'b0;

   // m376_114 = W*in
   wire signed [9:0] m376_114;
   assign m376_114 =10'b0;

   // m376_115 = W*in
   wire signed [9:0] m376_115;
   assign m376_115 =10'b0;

   // m376_116 = W*in
   wire signed [9:0] m376_116;
   assign m376_116 =10'b0;

   // m376_117 = W*in
   wire signed [9:0] m376_117;
   assign m376_117 =10'b0;

   // m377_1 = W*in
   wire signed [9:0] m377_1;
   assign m377_1 =10'b0;

   // m377_2 = W*in
   wire signed [9:0] m377_2;
   assign m377_2 =10'b0;

   // m377_3 = W*in
   wire signed [9:0] m377_3;
   assign m377_3 =10'b0;

   // m377_4 = W*in
   wire signed [9:0] m377_4;
   assign m377_4 =10'b0;

   // m377_5 = W*in
   wire signed [9:0] m377_5;
   assign m377_5 ={ {4{in377[5]}} , in377[5:0] };

   // m377_6 = W*in
   wire signed [9:0] m377_6;
   assign m377_6 =10'b0;

   // m377_7 = W*in
   wire signed [9:0] m377_7;
   assign m377_7 =10'b0;

   // m377_8 = W*in
   wire signed [9:0] m377_8;
   assign m377_8 =10'b0;

   // m377_9 = W*in
   wire signed [9:0] m377_9;
   assign m377_9 =10'b0;

   // m377_10 = W*in
   wire signed [9:0] m377_10;
   assign m377_10 =10'b0;

   // m377_11 = W*in
   wire signed [9:0] m377_11;
   assign m377_11 =10'b0;

   // m377_12 = W*in
   wire signed [9:0] m377_12;
   assign m377_12 =10'b0;

   // m377_13 = W*in
   wire signed [9:0] m377_13;
   assign m377_13 =10'b0;

   // m377_14 = W*in
   wire signed [9:0] m377_14;
   assign m377_14 =10'b0;

   // m377_15 = W*in
   wire signed [9:0] m377_15;
   assign m377_15 =10'b0;

   // m377_16 = W*in
   wire signed [9:0] m377_16;
   assign m377_16 =10'b0;

   // m377_17 = W*in
   wire signed [9:0] m377_17;
   assign m377_17 =10'b0;

   // m377_18 = W*in
   wire signed [9:0] m377_18;
   assign m377_18 ={ {4{neg377[5]}} , neg377[5:0] };

   // m377_19 = W*in
   wire signed [9:0] m377_19;
   assign m377_19 ={ {5{in377[5]}} , in377[5:1] };

   // m377_20 = W*in
   wire signed [9:0] m377_20;
   assign m377_20 ={ {4{neg377[5]}} , neg377[5:0] };

   // m377_21 = W*in
   wire signed [9:0] m377_21;
   assign m377_21 ={ {5{in377[5]}} , in377[5:1] };

   // m377_22 = W*in
   wire signed [9:0] m377_22;
   assign m377_22 =10'b0;

   // m377_23 = W*in
   wire signed [9:0] m377_23;
   assign m377_23 =10'b0;

   // m377_24 = W*in
   wire signed [9:0] m377_24;
   assign m377_24 =10'b0;

   // m377_25 = W*in
   wire signed [9:0] m377_25;
   assign m377_25 =10'b0;

   // m377_26 = W*in
   wire signed [9:0] m377_26;
   assign m377_26 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_27 = W*in
   wire signed [9:0] m377_27;
   assign m377_27 =10'b0;

   // m377_28 = W*in
   wire signed [9:0] m377_28;
   assign m377_28 =10'b0;

   // m377_29 = W*in
   wire signed [9:0] m377_29;
   assign m377_29 ={ {4{in377[5]}} , in377[5:0] };

   // m377_30 = W*in
   wire signed [9:0] m377_30;
   assign m377_30 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_31 = W*in
   wire signed [9:0] m377_31;
   assign m377_31 =10'b0;

   // m377_32 = W*in
   wire signed [9:0] m377_32;
   assign m377_32 =10'b0;

   // m377_33 = W*in
   wire signed [9:0] m377_33;
   assign m377_33 =10'b0;

   // m377_34 = W*in
   wire signed [9:0] m377_34;
   assign m377_34 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_35 = W*in
   wire signed [9:0] m377_35;
   assign m377_35 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_36 = W*in
   wire signed [9:0] m377_36;
   assign m377_36 =10'b0;

   // m377_37 = W*in
   wire signed [9:0] m377_37;
   assign m377_37 =10'b0;

   // m377_38 = W*in
   wire signed [9:0] m377_38;
   assign m377_38 =10'b0;

   // m377_39 = W*in
   wire signed [9:0] m377_39;
   assign m377_39 =10'b0;

   // m377_40 = W*in
   wire signed [9:0] m377_40;
   assign m377_40 =10'b0;

   // m377_41 = W*in
   wire signed [9:0] m377_41;
   assign m377_41 =10'b0;

   // m377_42 = W*in
   wire signed [9:0] m377_42;
   assign m377_42 =10'b0;

   // m377_43 = W*in
   wire signed [9:0] m377_43;
   assign m377_43 =10'b0;

   // m377_44 = W*in
   wire signed [9:0] m377_44;
   assign m377_44 ={ {4{in377[5]}} , in377[5:0] };

   // m377_45 = W*in
   wire signed [9:0] m377_45;
   assign m377_45 =10'b0;

   // m377_46 = W*in
   wire signed [9:0] m377_46;
   assign m377_46 =10'b0;

   // m377_47 = W*in
   wire signed [9:0] m377_47;
   assign m377_47 =10'b0;

   // m377_48 = W*in
   wire signed [9:0] m377_48;
   assign m377_48 =10'b0;

   // m377_49 = W*in
   wire signed [9:0] m377_49;
   assign m377_49 =10'b0;

   // m377_50 = W*in
   wire signed [9:0] m377_50;
   assign m377_50 =10'b0;

   // m377_51 = W*in
   wire signed [9:0] m377_51;
   assign m377_51 =10'b0;

   // m377_52 = W*in
   wire signed [9:0] m377_52;
   assign m377_52 =10'b0;

   // m377_53 = W*in
   wire signed [9:0] m377_53;
   assign m377_53 =10'b0;

   // m377_54 = W*in
   wire signed [9:0] m377_54;
   assign m377_54 ={ {4{in377[5]}} , in377[5:0] };

   // m377_55 = W*in
   wire signed [9:0] m377_55;
   assign m377_55 =10'b0;

   // m377_56 = W*in
   wire signed [9:0] m377_56;
   assign m377_56 =10'b0;

   // m377_57 = W*in
   wire signed [9:0] m377_57;
   assign m377_57 =10'b0;

   // m377_58 = W*in
   wire signed [9:0] m377_58;
   assign m377_58 =10'b0;

   // m377_59 = W*in
   wire signed [9:0] m377_59;
   assign m377_59 =10'b0;

   // m377_60 = W*in
   wire signed [9:0] m377_60;
   assign m377_60 =10'b0;

   // m377_61 = W*in
   wire signed [9:0] m377_61;
   assign m377_61 =10'b0;

   // m377_62 = W*in
   wire signed [9:0] m377_62;
   assign m377_62 =10'b0;

   // m377_63 = W*in
   wire signed [9:0] m377_63;
   assign m377_63 ={ {5{in377[5]}} , in377[5:1] };

   // m377_64 = W*in
   wire signed [9:0] m377_64;
   assign m377_64 ={ {4{neg377[5]}} , neg377[5:0] };

   // m377_65 = W*in
   wire signed [9:0] m377_65;
   assign m377_65 =10'b0;

   // m377_66 = W*in
   wire signed [9:0] m377_66;
   assign m377_66 =10'b0;

   // m377_67 = W*in
   wire signed [9:0] m377_67;
   assign m377_67 =10'b0;

   // m377_68 = W*in
   wire signed [9:0] m377_68;
   assign m377_68 ={ {4{neg377[5]}} , neg377[5:0] };

   // m377_69 = W*in
   wire signed [9:0] m377_69;
   assign m377_69 ={ {4{in377[5]}} , in377[5:0] };

   // m377_70 = W*in
   wire signed [9:0] m377_70;
   assign m377_70 =10'b0;

   // m377_71 = W*in
   wire signed [9:0] m377_71;
   assign m377_71 =10'b0;

   // m377_72 = W*in
   wire signed [9:0] m377_72;
   assign m377_72 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_73 = W*in
   wire signed [9:0] m377_73;
   assign m377_73 =10'b0;

   // m377_74 = W*in
   wire signed [9:0] m377_74;
   assign m377_74 ={ {4{neg377[5]}} , neg377[5:0] };

   // m377_75 = W*in
   wire signed [9:0] m377_75;
   assign m377_75 =10'b0;

   // m377_76 = W*in
   wire signed [9:0] m377_76;
   assign m377_76 =10'b0;

   // m377_77 = W*in
   wire signed [9:0] m377_77;
   assign m377_77 =10'b0;

   // m377_78 = W*in
   wire signed [9:0] m377_78;
   assign m377_78 =10'b0;

   // m377_79 = W*in
   wire signed [9:0] m377_79;
   assign m377_79 =10'b0;

   // m377_80 = W*in
   wire signed [9:0] m377_80;
   assign m377_80 =10'b0;

   // m377_81 = W*in
   wire signed [9:0] m377_81;
   assign m377_81 ={ {4{neg377[5]}} , neg377[5:0] };

   // m377_82 = W*in
   wire signed [9:0] m377_82;
   assign m377_82 ={ {4{in377[5]}} , in377[5:0] };

   // m377_83 = W*in
   wire signed [9:0] m377_83;
   assign m377_83 ={ {5{in377[5]}} , in377[5:1] };

   // m377_84 = W*in
   wire signed [9:0] m377_84;
   assign m377_84 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_85 = W*in
   wire signed [9:0] m377_85;
   assign m377_85 ={ {4{in377[5]}} , in377[5:0] };

   // m377_86 = W*in
   wire signed [9:0] m377_86;
   assign m377_86 =10'b0;

   // m377_87 = W*in
   wire signed [9:0] m377_87;
   assign m377_87 =10'b0;

   // m377_88 = W*in
   wire signed [9:0] m377_88;
   assign m377_88 =10'b0;

   // m377_89 = W*in
   wire signed [9:0] m377_89;
   assign m377_89 =10'b0;

   // m377_90 = W*in
   wire signed [9:0] m377_90;
   assign m377_90 =10'b0;

   // m377_91 = W*in
   wire signed [9:0] m377_91;
   assign m377_91 =10'b0;

   // m377_92 = W*in
   wire signed [9:0] m377_92;
   assign m377_92 =10'b0;

   // m377_93 = W*in
   wire signed [9:0] m377_93;
   assign m377_93 ={ {4{in377[5]}} , in377[5:0] };

   // m377_94 = W*in
   wire signed [9:0] m377_94;
   assign m377_94 =10'b0;

   // m377_95 = W*in
   wire signed [9:0] m377_95;
   assign m377_95 ={ {4{in377[5]}} , in377[5:0] };

   // m377_96 = W*in
   wire signed [9:0] m377_96;
   assign m377_96 =10'b0;

   // m377_97 = W*in
   wire signed [9:0] m377_97;
   assign m377_97 =10'b0;

   // m377_98 = W*in
   wire signed [9:0] m377_98;
   assign m377_98 =10'b0;

   // m377_99 = W*in
   wire signed [9:0] m377_99;
   assign m377_99 =10'b0;

   // m377_100 = W*in
   wire signed [9:0] m377_100;
   assign m377_100 =10'b0;

   // m377_101 = W*in
   wire signed [9:0] m377_101;
   assign m377_101 =10'b0;

   // m377_102 = W*in
   wire signed [9:0] m377_102;
   assign m377_102 =10'b0;

   // m377_103 = W*in
   wire signed [9:0] m377_103;
   assign m377_103 =10'b0;

   // m377_104 = W*in
   wire signed [9:0] m377_104;
   assign m377_104 =10'b0;

   // m377_105 = W*in
   wire signed [9:0] m377_105;
   assign m377_105 =10'b0;

   // m377_106 = W*in
   wire signed [9:0] m377_106;
   assign m377_106 =10'b0;

   // m377_107 = W*in
   wire signed [9:0] m377_107;
   assign m377_107 ={ {5{in377[5]}} , in377[5:1] };

   // m377_108 = W*in
   wire signed [9:0] m377_108;
   assign m377_108 =10'b0;

   // m377_109 = W*in
   wire signed [9:0] m377_109;
   assign m377_109 =10'b0;

   // m377_110 = W*in
   wire signed [9:0] m377_110;
   assign m377_110 =10'b0;

   // m377_111 = W*in
   wire signed [9:0] m377_111;
   assign m377_111 =10'b0;

   // m377_112 = W*in
   wire signed [9:0] m377_112;
   assign m377_112 =10'b0;

   // m377_113 = W*in
   wire signed [9:0] m377_113;
   assign m377_113 =10'b0;

   // m377_114 = W*in
   wire signed [9:0] m377_114;
   assign m377_114 =10'b0;

   // m377_115 = W*in
   wire signed [9:0] m377_115;
   assign m377_115 ={ {5{neg377[5]}} , neg377[5:1] };

   // m377_116 = W*in
   wire signed [9:0] m377_116;
   assign m377_116 =10'b0;

   // m377_117 = W*in
   wire signed [9:0] m377_117;
   assign m377_117 =10'b0;

   // m378_1 = W*in
   wire signed [9:0] m378_1;
   assign m378_1 =10'b0;

   // m378_2 = W*in
   wire signed [9:0] m378_2;
   assign m378_2 ={ {3{neg378[5]}} , neg378 , {1{1'b0}} };

   // m378_3 = W*in
   wire signed [9:0] m378_3;
   assign m378_3 =10'b0;

   // m378_4 = W*in
   wire signed [9:0] m378_4;
   assign m378_4 =10'b0;

   // m378_5 = W*in
   wire signed [9:0] m378_5;
   assign m378_5 =10'b0;

   // m378_6 = W*in
   wire signed [9:0] m378_6;
   assign m378_6 ={ {4{in378[5]}} , in378[5:0] };

   // m378_7 = W*in
   wire signed [9:0] m378_7;
   assign m378_7 =10'b0;

   // m378_8 = W*in
   wire signed [9:0] m378_8;
   assign m378_8 ={ {3{neg378[5]}} , neg378 , {1{1'b0}} };

   // m378_9 = W*in
   wire signed [9:0] m378_9;
   assign m378_9 =10'b0;

   // m378_10 = W*in
   wire signed [9:0] m378_10;
   assign m378_10 =10'b0;

   // m378_11 = W*in
   wire signed [9:0] m378_11;
   assign m378_11 ={ {4{in378[5]}} , in378[5:0] };

   // m378_12 = W*in
   wire signed [9:0] m378_12;
   assign m378_12 =10'b0;

   // m378_13 = W*in
   wire signed [9:0] m378_13;
   assign m378_13 =10'b0;

   // m378_14 = W*in
   wire signed [9:0] m378_14;
   assign m378_14 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_15 = W*in
   wire signed [9:0] m378_15;
   assign m378_15 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_16 = W*in
   wire signed [9:0] m378_16;
   assign m378_16 =10'b0;

   // m378_17 = W*in
   wire signed [9:0] m378_17;
   assign m378_17 =10'b0;

   // m378_18 = W*in
   wire signed [9:0] m378_18;
   assign m378_18 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_19 = W*in
   wire signed [9:0] m378_19;
   assign m378_19 =10'b0;

   // m378_20 = W*in
   wire signed [9:0] m378_20;
   assign m378_20 =10'b0;

   // m378_21 = W*in
   wire signed [9:0] m378_21;
   assign m378_21 ={ {5{in378[5]}} , in378[5:1] };

   // m378_22 = W*in
   wire signed [9:0] m378_22;
   assign m378_22 =10'b0;

   // m378_23 = W*in
   wire signed [9:0] m378_23;
   assign m378_23 =10'b0;

   // m378_24 = W*in
   wire signed [9:0] m378_24;
   assign m378_24 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_25 = W*in
   wire signed [9:0] m378_25;
   assign m378_25 =10'b0;

   // m378_26 = W*in
   wire signed [9:0] m378_26;
   assign m378_26 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_27 = W*in
   wire signed [9:0] m378_27;
   assign m378_27 =10'b0;

   // m378_28 = W*in
   wire signed [9:0] m378_28;
   assign m378_28 =10'b0;

   // m378_29 = W*in
   wire signed [9:0] m378_29;
   assign m378_29 =10'b0;

   // m378_30 = W*in
   wire signed [9:0] m378_30;
   assign m378_30 =10'b0;

   // m378_31 = W*in
   wire signed [9:0] m378_31;
   assign m378_31 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_32 = W*in
   wire signed [9:0] m378_32;
   assign m378_32 =10'b0;

   // m378_33 = W*in
   wire signed [9:0] m378_33;
   assign m378_33 =10'b0;

   // m378_34 = W*in
   wire signed [9:0] m378_34;
   assign m378_34 =10'b0;

   // m378_35 = W*in
   wire signed [9:0] m378_35;
   assign m378_35 =10'b0;

   // m378_36 = W*in
   wire signed [9:0] m378_36;
   assign m378_36 =10'b0;

   // m378_37 = W*in
   wire signed [9:0] m378_37;
   assign m378_37 =10'b0;

   // m378_38 = W*in
   wire signed [9:0] m378_38;
   assign m378_38 =10'b0;

   // m378_39 = W*in
   wire signed [9:0] m378_39;
   assign m378_39 =10'b0;

   // m378_40 = W*in
   wire signed [9:0] m378_40;
   assign m378_40 =10'b0;

   // m378_41 = W*in
   wire signed [9:0] m378_41;
   assign m378_41 ={ {4{in378[5]}} , in378[5:0] };

   // m378_42 = W*in
   wire signed [9:0] m378_42;
   assign m378_42 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_43 = W*in
   wire signed [9:0] m378_43;
   assign m378_43 =10'b0;

   // m378_44 = W*in
   wire signed [9:0] m378_44;
   assign m378_44 ={ {4{in378[5]}} , in378[5:0] };

   // m378_45 = W*in
   wire signed [9:0] m378_45;
   assign m378_45 =10'b0;

   // m378_46 = W*in
   wire signed [9:0] m378_46;
   assign m378_46 =10'b0;

   // m378_47 = W*in
   wire signed [9:0] m378_47;
   assign m378_47 =10'b0;

   // m378_48 = W*in
   wire signed [9:0] m378_48;
   assign m378_48 =10'b0;

   // m378_49 = W*in
   wire signed [9:0] m378_49;
   assign m378_49 =10'b0;

   // m378_50 = W*in
   wire signed [9:0] m378_50;
   assign m378_50 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_51 = W*in
   wire signed [9:0] m378_51;
   assign m378_51 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_52 = W*in
   wire signed [9:0] m378_52;
   assign m378_52 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_53 = W*in
   wire signed [9:0] m378_53;
   assign m378_53 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_54 = W*in
   wire signed [9:0] m378_54;
   assign m378_54 ={ {4{in378[5]}} , in378[5:0] };

   // m378_55 = W*in
   wire signed [9:0] m378_55;
   assign m378_55 =10'b0;

   // m378_56 = W*in
   wire signed [9:0] m378_56;
   assign m378_56 =10'b0;

   // m378_57 = W*in
   wire signed [9:0] m378_57;
   assign m378_57 ={ {4{in378[5]}} , in378[5:0] };

   // m378_58 = W*in
   wire signed [9:0] m378_58;
   assign m378_58 =10'b0;

   // m378_59 = W*in
   wire signed [9:0] m378_59;
   assign m378_59 =10'b0;

   // m378_60 = W*in
   wire signed [9:0] m378_60;
   assign m378_60 ={ {4{in378[5]}} , in378[5:0] };

   // m378_61 = W*in
   wire signed [9:0] m378_61;
   assign m378_61 ={ {4{in378[5]}} , in378[5:0] };

   // m378_62 = W*in
   wire signed [9:0] m378_62;
   assign m378_62 =10'b0;

   // m378_63 = W*in
   wire signed [9:0] m378_63;
   assign m378_63 ={ {4{in378[5]}} , in378[5:0] };

   // m378_64 = W*in
   wire signed [9:0] m378_64;
   assign m378_64 =10'b0;

   // m378_65 = W*in
   wire signed [9:0] m378_65;
   assign m378_65 =10'b0;

   // m378_66 = W*in
   wire signed [9:0] m378_66;
   assign m378_66 ={ {5{in378[5]}} , in378[5:1] };

   // m378_67 = W*in
   wire signed [9:0] m378_67;
   assign m378_67 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_68 = W*in
   wire signed [9:0] m378_68;
   assign m378_68 ={ {3{neg378[5]}} , neg378 , {1{1'b0}} };

   // m378_69 = W*in
   wire signed [9:0] m378_69;
   assign m378_69 ={ {4{in378[5]}} , in378[5:0] };

   // m378_70 = W*in
   wire signed [9:0] m378_70;
   assign m378_70 ={ {5{in378[5]}} , in378[5:1] };

   // m378_71 = W*in
   wire signed [9:0] m378_71;
   assign m378_71 =10'b0;

   // m378_72 = W*in
   wire signed [9:0] m378_72;
   assign m378_72 =10'b0;

   // m378_73 = W*in
   wire signed [9:0] m378_73;
   assign m378_73 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_74 = W*in
   wire signed [9:0] m378_74;
   assign m378_74 =10'b0;

   // m378_75 = W*in
   wire signed [9:0] m378_75;
   assign m378_75 =10'b0;

   // m378_76 = W*in
   wire signed [9:0] m378_76;
   assign m378_76 =10'b0;

   // m378_77 = W*in
   wire signed [9:0] m378_77;
   assign m378_77 ={ {4{in378[5]}} , in378[5:0] };

   // m378_78 = W*in
   wire signed [9:0] m378_78;
   assign m378_78 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_79 = W*in
   wire signed [9:0] m378_79;
   assign m378_79 =10'b0;

   // m378_80 = W*in
   wire signed [9:0] m378_80;
   assign m378_80 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_81 = W*in
   wire signed [9:0] m378_81;
   assign m378_81 =10'b0;

   // m378_82 = W*in
   wire signed [9:0] m378_82;
   assign m378_82 =10'b0;

   // m378_83 = W*in
   wire signed [9:0] m378_83;
   assign m378_83 =10'b0;

   // m378_84 = W*in
   wire signed [9:0] m378_84;
   assign m378_84 =10'b0;

   // m378_85 = W*in
   wire signed [9:0] m378_85;
   assign m378_85 =10'b0;

   // m378_86 = W*in
   wire signed [9:0] m378_86;
   assign m378_86 =10'b0;

   // m378_87 = W*in
   wire signed [9:0] m378_87;
   assign m378_87 =10'b0;

   // m378_88 = W*in
   wire signed [9:0] m378_88;
   assign m378_88 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_89 = W*in
   wire signed [9:0] m378_89;
   assign m378_89 =10'b0;

   // m378_90 = W*in
   wire signed [9:0] m378_90;
   assign m378_90 ={ {3{neg378[5]}} , neg378 , {1{1'b0}} };

   // m378_91 = W*in
   wire signed [9:0] m378_91;
   assign m378_91 =10'b0;

   // m378_92 = W*in
   wire signed [9:0] m378_92;
   assign m378_92 =10'b0;

   // m378_93 = W*in
   wire signed [9:0] m378_93;
   assign m378_93 =10'b0;

   // m378_94 = W*in
   wire signed [9:0] m378_94;
   assign m378_94 =10'b0;

   // m378_95 = W*in
   wire signed [9:0] m378_95;
   assign m378_95 ={ {4{in378[5]}} , in378[5:0] };

   // m378_96 = W*in
   wire signed [9:0] m378_96;
   assign m378_96 =10'b0;

   // m378_97 = W*in
   wire signed [9:0] m378_97;
   assign m378_97 =10'b0;

   // m378_98 = W*in
   wire signed [9:0] m378_98;
   assign m378_98 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_99 = W*in
   wire signed [9:0] m378_99;
   assign m378_99 ={ {4{in378[5]}} , in378[5:0] };

   // m378_100 = W*in
   wire signed [9:0] m378_100;
   assign m378_100 =10'b0;

   // m378_101 = W*in
   wire signed [9:0] m378_101;
   assign m378_101 ={ {5{in378[5]}} , in378[5:1] };

   // m378_102 = W*in
   wire signed [9:0] m378_102;
   assign m378_102 =10'b0;

   // m378_103 = W*in
   wire signed [9:0] m378_103;
   assign m378_103 =10'b0;

   // m378_104 = W*in
   wire signed [9:0] m378_104;
   assign m378_104 =10'b0;

   // m378_105 = W*in
   wire signed [9:0] m378_105;
   assign m378_105 ={ {4{neg378[5]}} , neg378[5:0] };

   // m378_106 = W*in
   wire signed [9:0] m378_106;
   assign m378_106 =10'b0;

   // m378_107 = W*in
   wire signed [9:0] m378_107;
   assign m378_107 =10'b0;

   // m378_108 = W*in
   wire signed [9:0] m378_108;
   assign m378_108 =10'b0;

   // m378_109 = W*in
   wire signed [9:0] m378_109;
   assign m378_109 =10'b0;

   // m378_110 = W*in
   wire signed [9:0] m378_110;
   assign m378_110 ={ {4{in378[5]}} , in378[5:0] };

   // m378_111 = W*in
   wire signed [9:0] m378_111;
   assign m378_111 =10'b0;

   // m378_112 = W*in
   wire signed [9:0] m378_112;
   assign m378_112 =10'b0;

   // m378_113 = W*in
   wire signed [9:0] m378_113;
   assign m378_113 =10'b0;

   // m378_114 = W*in
   wire signed [9:0] m378_114;
   assign m378_114 =10'b0;

   // m378_115 = W*in
   wire signed [9:0] m378_115;
   assign m378_115 =10'b0;

   // m378_116 = W*in
   wire signed [9:0] m378_116;
   assign m378_116 =10'b0;

   // m378_117 = W*in
   wire signed [9:0] m378_117;
   assign m378_117 =10'b0;

   // m379_1 = W*in
   wire signed [9:0] m379_1;
   assign m379_1 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_2 = W*in
   wire signed [9:0] m379_2;
   assign m379_2 ={ {3{neg379[5]}} , neg379 , {1{1'b0}} };

   // m379_3 = W*in
   wire signed [9:0] m379_3;
   assign m379_3 =10'b0;

   // m379_4 = W*in
   wire signed [9:0] m379_4;
   assign m379_4 =10'b0;

   // m379_5 = W*in
   wire signed [9:0] m379_5;
   assign m379_5 =10'b0;

   // m379_6 = W*in
   wire signed [9:0] m379_6;
   assign m379_6 =10'b0;

   // m379_7 = W*in
   wire signed [9:0] m379_7;
   assign m379_7 =10'b0;

   // m379_8 = W*in
   wire signed [9:0] m379_8;
   assign m379_8 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_9 = W*in
   wire signed [9:0] m379_9;
   assign m379_9 =10'b0;

   // m379_10 = W*in
   wire signed [9:0] m379_10;
   assign m379_10 =10'b0;

   // m379_11 = W*in
   wire signed [9:0] m379_11;
   assign m379_11 =10'b0;

   // m379_12 = W*in
   wire signed [9:0] m379_12;
   assign m379_12 =10'b0;

   // m379_13 = W*in
   wire signed [9:0] m379_13;
   assign m379_13 =10'b0;

   // m379_14 = W*in
   wire signed [9:0] m379_14;
   assign m379_14 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_15 = W*in
   wire signed [9:0] m379_15;
   assign m379_15 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_16 = W*in
   wire signed [9:0] m379_16;
   assign m379_16 =10'b0;

   // m379_17 = W*in
   wire signed [9:0] m379_17;
   assign m379_17 ={ {4{in379[5]}} , in379[5:0] };

   // m379_18 = W*in
   wire signed [9:0] m379_18;
   assign m379_18 =10'b0;

   // m379_19 = W*in
   wire signed [9:0] m379_19;
   assign m379_19 =10'b0;

   // m379_20 = W*in
   wire signed [9:0] m379_20;
   assign m379_20 ={ {4{in379[5]}} , in379[5:0] };

   // m379_21 = W*in
   wire signed [9:0] m379_21;
   assign m379_21 =10'b0;

   // m379_22 = W*in
   wire signed [9:0] m379_22;
   assign m379_22 =10'b0;

   // m379_23 = W*in
   wire signed [9:0] m379_23;
   assign m379_23 =10'b0;

   // m379_24 = W*in
   wire signed [9:0] m379_24;
   assign m379_24 =10'b0;

   // m379_25 = W*in
   wire signed [9:0] m379_25;
   assign m379_25 =10'b0;

   // m379_26 = W*in
   wire signed [9:0] m379_26;
   assign m379_26 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_27 = W*in
   wire signed [9:0] m379_27;
   assign m379_27 =10'b0;

   // m379_28 = W*in
   wire signed [9:0] m379_28;
   assign m379_28 =10'b0;

   // m379_29 = W*in
   wire signed [9:0] m379_29;
   assign m379_29 =10'b0;

   // m379_30 = W*in
   wire signed [9:0] m379_30;
   assign m379_30 ={ {4{in379[5]}} , in379[5:0] };

   // m379_31 = W*in
   wire signed [9:0] m379_31;
   assign m379_31 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_32 = W*in
   wire signed [9:0] m379_32;
   assign m379_32 =10'b0;

   // m379_33 = W*in
   wire signed [9:0] m379_33;
   assign m379_33 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_34 = W*in
   wire signed [9:0] m379_34;
   assign m379_34 =10'b0;

   // m379_35 = W*in
   wire signed [9:0] m379_35;
   assign m379_35 ={ {4{in379[5]}} , in379[5:0] };

   // m379_36 = W*in
   wire signed [9:0] m379_36;
   assign m379_36 =10'b0;

   // m379_37 = W*in
   wire signed [9:0] m379_37;
   assign m379_37 =10'b0;

   // m379_38 = W*in
   wire signed [9:0] m379_38;
   assign m379_38 ={ {4{in379[5]}} , in379[5:0] };

   // m379_39 = W*in
   wire signed [9:0] m379_39;
   assign m379_39 =10'b0;

   // m379_40 = W*in
   wire signed [9:0] m379_40;
   assign m379_40 =10'b0;

   // m379_41 = W*in
   wire signed [9:0] m379_41;
   assign m379_41 =10'b0;

   // m379_42 = W*in
   wire signed [9:0] m379_42;
   assign m379_42 =10'b0;

   // m379_43 = W*in
   wire signed [9:0] m379_43;
   assign m379_43 =10'b0;

   // m379_44 = W*in
   wire signed [9:0] m379_44;
   assign m379_44 ={ {4{in379[5]}} , in379[5:0] };

   // m379_45 = W*in
   wire signed [9:0] m379_45;
   assign m379_45 =10'b0;

   // m379_46 = W*in
   wire signed [9:0] m379_46;
   assign m379_46 =10'b0;

   // m379_47 = W*in
   wire signed [9:0] m379_47;
   assign m379_47 =10'b0;

   // m379_48 = W*in
   wire signed [9:0] m379_48;
   assign m379_48 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_49 = W*in
   wire signed [9:0] m379_49;
   assign m379_49 =10'b0;

   // m379_50 = W*in
   wire signed [9:0] m379_50;
   assign m379_50 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_51 = W*in
   wire signed [9:0] m379_51;
   assign m379_51 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_52 = W*in
   wire signed [9:0] m379_52;
   assign m379_52 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_53 = W*in
   wire signed [9:0] m379_53;
   assign m379_53 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_54 = W*in
   wire signed [9:0] m379_54;
   assign m379_54 =10'b0;

   // m379_55 = W*in
   wire signed [9:0] m379_55;
   assign m379_55 =10'b0;

   // m379_56 = W*in
   wire signed [9:0] m379_56;
   assign m379_56 =10'b0;

   // m379_57 = W*in
   wire signed [9:0] m379_57;
   assign m379_57 ={ {4{in379[5]}} , in379[5:0] };

   // m379_58 = W*in
   wire signed [9:0] m379_58;
   assign m379_58 =10'b0;

   // m379_59 = W*in
   wire signed [9:0] m379_59;
   assign m379_59 =10'b0;

   // m379_60 = W*in
   wire signed [9:0] m379_60;
   assign m379_60 ={ {4{in379[5]}} , in379[5:0] };

   // m379_61 = W*in
   wire signed [9:0] m379_61;
   assign m379_61 ={ {4{in379[5]}} , in379[5:0] };

   // m379_62 = W*in
   wire signed [9:0] m379_62;
   assign m379_62 =10'b0;

   // m379_63 = W*in
   wire signed [9:0] m379_63;
   assign m379_63 =10'b0;

   // m379_64 = W*in
   wire signed [9:0] m379_64;
   assign m379_64 ={ {4{in379[5]}} , in379[5:0] };

   // m379_65 = W*in
   wire signed [9:0] m379_65;
   assign m379_65 ={ {5{neg379[5]}} , neg379[5:1] };

   // m379_66 = W*in
   wire signed [9:0] m379_66;
   assign m379_66 ={ {4{in379[5]}} , in379[5:0] };

   // m379_67 = W*in
   wire signed [9:0] m379_67;
   assign m379_67 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_68 = W*in
   wire signed [9:0] m379_68;
   assign m379_68 ={ {3{neg379[5]}} , neg379 , {1{1'b0}} };

   // m379_69 = W*in
   wire signed [9:0] m379_69;
   assign m379_69 =10'b0;

   // m379_70 = W*in
   wire signed [9:0] m379_70;
   assign m379_70 =10'b0;

   // m379_71 = W*in
   wire signed [9:0] m379_71;
   assign m379_71 ={ {5{in379[5]}} , in379[5:1] };

   // m379_72 = W*in
   wire signed [9:0] m379_72;
   assign m379_72 ={ {5{neg379[5]}} , neg379[5:1] };

   // m379_73 = W*in
   wire signed [9:0] m379_73;
   assign m379_73 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_74 = W*in
   wire signed [9:0] m379_74;
   assign m379_74 ={ {4{in379[5]}} , in379[5:0] };

   // m379_75 = W*in
   wire signed [9:0] m379_75;
   assign m379_75 =10'b0;

   // m379_76 = W*in
   wire signed [9:0] m379_76;
   assign m379_76 =10'b0;

   // m379_77 = W*in
   wire signed [9:0] m379_77;
   assign m379_77 =10'b0;

   // m379_78 = W*in
   wire signed [9:0] m379_78;
   assign m379_78 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_79 = W*in
   wire signed [9:0] m379_79;
   assign m379_79 ={ {4{in379[5]}} , in379[5:0] };

   // m379_80 = W*in
   wire signed [9:0] m379_80;
   assign m379_80 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_81 = W*in
   wire signed [9:0] m379_81;
   assign m379_81 ={ {4{in379[5]}} , in379[5:0] };

   // m379_82 = W*in
   wire signed [9:0] m379_82;
   assign m379_82 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_83 = W*in
   wire signed [9:0] m379_83;
   assign m379_83 =10'b0;

   // m379_84 = W*in
   wire signed [9:0] m379_84;
   assign m379_84 ={ {5{neg379[5]}} , neg379[5:1] };

   // m379_85 = W*in
   wire signed [9:0] m379_85;
   assign m379_85 =10'b0;

   // m379_86 = W*in
   wire signed [9:0] m379_86;
   assign m379_86 =10'b0;

   // m379_87 = W*in
   wire signed [9:0] m379_87;
   assign m379_87 =10'b0;

   // m379_88 = W*in
   wire signed [9:0] m379_88;
   assign m379_88 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_89 = W*in
   wire signed [9:0] m379_89;
   assign m379_89 =10'b0;

   // m379_90 = W*in
   wire signed [9:0] m379_90;
   assign m379_90 ={ {3{neg379[5]}} , neg379 , {1{1'b0}} };

   // m379_91 = W*in
   wire signed [9:0] m379_91;
   assign m379_91 ={ {5{in379[5]}} , in379[5:1] };

   // m379_92 = W*in
   wire signed [9:0] m379_92;
   assign m379_92 =10'b0;

   // m379_93 = W*in
   wire signed [9:0] m379_93;
   assign m379_93 =10'b0;

   // m379_94 = W*in
   wire signed [9:0] m379_94;
   assign m379_94 =10'b0;

   // m379_95 = W*in
   wire signed [9:0] m379_95;
   assign m379_95 =10'b0;

   // m379_96 = W*in
   wire signed [9:0] m379_96;
   assign m379_96 =10'b0;

   // m379_97 = W*in
   wire signed [9:0] m379_97;
   assign m379_97 =10'b0;

   // m379_98 = W*in
   wire signed [9:0] m379_98;
   assign m379_98 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_99 = W*in
   wire signed [9:0] m379_99;
   assign m379_99 ={ {4{in379[5]}} , in379[5:0] };

   // m379_100 = W*in
   wire signed [9:0] m379_100;
   assign m379_100 ={ {4{in379[5]}} , in379[5:0] };

   // m379_101 = W*in
   wire signed [9:0] m379_101;
   assign m379_101 ={ {4{in379[5]}} , in379[5:0] };

   // m379_102 = W*in
   wire signed [9:0] m379_102;
   assign m379_102 =10'b0;

   // m379_103 = W*in
   wire signed [9:0] m379_103;
   assign m379_103 =10'b0;

   // m379_104 = W*in
   wire signed [9:0] m379_104;
   assign m379_104 =10'b0;

   // m379_105 = W*in
   wire signed [9:0] m379_105;
   assign m379_105 =10'b0;

   // m379_106 = W*in
   wire signed [9:0] m379_106;
   assign m379_106 =10'b0;

   // m379_107 = W*in
   wire signed [9:0] m379_107;
   assign m379_107 ={ {4{neg379[5]}} , neg379[5:0] };

   // m379_108 = W*in
   wire signed [9:0] m379_108;
   assign m379_108 =10'b0;

   // m379_109 = W*in
   wire signed [9:0] m379_109;
   assign m379_109 =10'b0;

   // m379_110 = W*in
   wire signed [9:0] m379_110;
   assign m379_110 ={ {4{in379[5]}} , in379[5:0] };

   // m379_111 = W*in
   wire signed [9:0] m379_111;
   assign m379_111 ={ {5{neg379[5]}} , neg379[5:1] };

   // m379_112 = W*in
   wire signed [9:0] m379_112;
   assign m379_112 =10'b0;

   // m379_113 = W*in
   wire signed [9:0] m379_113;
   assign m379_113 ={ {5{neg379[5]}} , neg379[5:1] };

   // m379_114 = W*in
   wire signed [9:0] m379_114;
   assign m379_114 ={ {4{in379[5]}} , in379[5:0] };

   // m379_115 = W*in
   wire signed [9:0] m379_115;
   assign m379_115 =10'b0;

   // m379_116 = W*in
   wire signed [9:0] m379_116;
   assign m379_116 =10'b0;

   // m379_117 = W*in
   wire signed [9:0] m379_117;
   assign m379_117 ={ {4{in379[5]}} , in379[5:0] };

   // m380_1 = W*in
   wire signed [9:0] m380_1;
   assign m380_1 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_2 = W*in
   wire signed [9:0] m380_2;
   assign m380_2 =10'b0;

   // m380_3 = W*in
   wire signed [9:0] m380_3;
   assign m380_3 =10'b0;

   // m380_4 = W*in
   wire signed [9:0] m380_4;
   assign m380_4 =10'b0;

   // m380_5 = W*in
   wire signed [9:0] m380_5;
   assign m380_5 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_6 = W*in
   wire signed [9:0] m380_6;
   assign m380_6 ={ {4{in380[5]}} , in380[5:0] };

   // m380_7 = W*in
   wire signed [9:0] m380_7;
   assign m380_7 =10'b0;

   // m380_8 = W*in
   wire signed [9:0] m380_8;
   assign m380_8 =10'b0;

   // m380_9 = W*in
   wire signed [9:0] m380_9;
   assign m380_9 =10'b0;

   // m380_10 = W*in
   wire signed [9:0] m380_10;
   assign m380_10 ={ {4{in380[5]}} , in380[5:0] };

   // m380_11 = W*in
   wire signed [9:0] m380_11;
   assign m380_11 =10'b0;

   // m380_12 = W*in
   wire signed [9:0] m380_12;
   assign m380_12 =10'b0;

   // m380_13 = W*in
   wire signed [9:0] m380_13;
   assign m380_13 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_14 = W*in
   wire signed [9:0] m380_14;
   assign m380_14 =10'b0;

   // m380_15 = W*in
   wire signed [9:0] m380_15;
   assign m380_15 =10'b0;

   // m380_16 = W*in
   wire signed [9:0] m380_16;
   assign m380_16 =10'b0;

   // m380_17 = W*in
   wire signed [9:0] m380_17;
   assign m380_17 =10'b0;

   // m380_18 = W*in
   wire signed [9:0] m380_18;
   assign m380_18 =10'b0;

   // m380_19 = W*in
   wire signed [9:0] m380_19;
   assign m380_19 =10'b0;

   // m380_20 = W*in
   wire signed [9:0] m380_20;
   assign m380_20 =10'b0;

   // m380_21 = W*in
   wire signed [9:0] m380_21;
   assign m380_21 =10'b0;

   // m380_22 = W*in
   wire signed [9:0] m380_22;
   assign m380_22 =10'b0;

   // m380_23 = W*in
   wire signed [9:0] m380_23;
   assign m380_23 =10'b0;

   // m380_24 = W*in
   wire signed [9:0] m380_24;
   assign m380_24 =10'b0;

   // m380_25 = W*in
   wire signed [9:0] m380_25;
   assign m380_25 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_26 = W*in
   wire signed [9:0] m380_26;
   assign m380_26 =10'b0;

   // m380_27 = W*in
   wire signed [9:0] m380_27;
   assign m380_27 =10'b0;

   // m380_28 = W*in
   wire signed [9:0] m380_28;
   assign m380_28 ={ {5{neg380[5]}} , neg380[5:1] };

   // m380_29 = W*in
   wire signed [9:0] m380_29;
   assign m380_29 =10'b0;

   // m380_30 = W*in
   wire signed [9:0] m380_30;
   assign m380_30 ={ {5{in380[5]}} , in380[5:1] };

   // m380_31 = W*in
   wire signed [9:0] m380_31;
   assign m380_31 =10'b0;

   // m380_32 = W*in
   wire signed [9:0] m380_32;
   assign m380_32 =10'b0;

   // m380_33 = W*in
   wire signed [9:0] m380_33;
   assign m380_33 =10'b0;

   // m380_34 = W*in
   wire signed [9:0] m380_34;
   assign m380_34 =10'b0;

   // m380_35 = W*in
   wire signed [9:0] m380_35;
   assign m380_35 ={ {4{in380[5]}} , in380[5:0] };

   // m380_36 = W*in
   wire signed [9:0] m380_36;
   assign m380_36 =10'b0;

   // m380_37 = W*in
   wire signed [9:0] m380_37;
   assign m380_37 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_38 = W*in
   wire signed [9:0] m380_38;
   assign m380_38 ={ {4{in380[5]}} , in380[5:0] };

   // m380_39 = W*in
   wire signed [9:0] m380_39;
   assign m380_39 =10'b0;

   // m380_40 = W*in
   wire signed [9:0] m380_40;
   assign m380_40 =10'b0;

   // m380_41 = W*in
   wire signed [9:0] m380_41;
   assign m380_41 =10'b0;

   // m380_42 = W*in
   wire signed [9:0] m380_42;
   assign m380_42 =10'b0;

   // m380_43 = W*in
   wire signed [9:0] m380_43;
   assign m380_43 =10'b0;

   // m380_44 = W*in
   wire signed [9:0] m380_44;
   assign m380_44 =10'b0;

   // m380_45 = W*in
   wire signed [9:0] m380_45;
   assign m380_45 =10'b0;

   // m380_46 = W*in
   wire signed [9:0] m380_46;
   assign m380_46 =10'b0;

   // m380_47 = W*in
   wire signed [9:0] m380_47;
   assign m380_47 =10'b0;

   // m380_48 = W*in
   wire signed [9:0] m380_48;
   assign m380_48 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_49 = W*in
   wire signed [9:0] m380_49;
   assign m380_49 =10'b0;

   // m380_50 = W*in
   wire signed [9:0] m380_50;
   assign m380_50 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_51 = W*in
   wire signed [9:0] m380_51;
   assign m380_51 =10'b0;

   // m380_52 = W*in
   wire signed [9:0] m380_52;
   assign m380_52 =10'b0;

   // m380_53 = W*in
   wire signed [9:0] m380_53;
   assign m380_53 =10'b0;

   // m380_54 = W*in
   wire signed [9:0] m380_54;
   assign m380_54 =10'b0;

   // m380_55 = W*in
   wire signed [9:0] m380_55;
   assign m380_55 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_56 = W*in
   wire signed [9:0] m380_56;
   assign m380_56 =10'b0;

   // m380_57 = W*in
   wire signed [9:0] m380_57;
   assign m380_57 ={ {4{in380[5]}} , in380[5:0] };

   // m380_58 = W*in
   wire signed [9:0] m380_58;
   assign m380_58 =10'b0;

   // m380_59 = W*in
   wire signed [9:0] m380_59;
   assign m380_59 =10'b0;

   // m380_60 = W*in
   wire signed [9:0] m380_60;
   assign m380_60 =10'b0;

   // m380_61 = W*in
   wire signed [9:0] m380_61;
   assign m380_61 ={ {4{in380[5]}} , in380[5:0] };

   // m380_62 = W*in
   wire signed [9:0] m380_62;
   assign m380_62 =10'b0;

   // m380_63 = W*in
   wire signed [9:0] m380_63;
   assign m380_63 ={ {5{neg380[5]}} , neg380[5:1] };

   // m380_64 = W*in
   wire signed [9:0] m380_64;
   assign m380_64 ={ {4{in380[5]}} , in380[5:0] };

   // m380_65 = W*in
   wire signed [9:0] m380_65;
   assign m380_65 =10'b0;

   // m380_66 = W*in
   wire signed [9:0] m380_66;
   assign m380_66 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_67 = W*in
   wire signed [9:0] m380_67;
   assign m380_67 =10'b0;

   // m380_68 = W*in
   wire signed [9:0] m380_68;
   assign m380_68 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_69 = W*in
   wire signed [9:0] m380_69;
   assign m380_69 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_70 = W*in
   wire signed [9:0] m380_70;
   assign m380_70 =10'b0;

   // m380_71 = W*in
   wire signed [9:0] m380_71;
   assign m380_71 =10'b0;

   // m380_72 = W*in
   wire signed [9:0] m380_72;
   assign m380_72 =10'b0;

   // m380_73 = W*in
   wire signed [9:0] m380_73;
   assign m380_73 ={ {5{neg380[5]}} , neg380[5:1] };

   // m380_74 = W*in
   wire signed [9:0] m380_74;
   assign m380_74 ={ {4{in380[5]}} , in380[5:0] };

   // m380_75 = W*in
   wire signed [9:0] m380_75;
   assign m380_75 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_76 = W*in
   wire signed [9:0] m380_76;
   assign m380_76 =10'b0;

   // m380_77 = W*in
   wire signed [9:0] m380_77;
   assign m380_77 =10'b0;

   // m380_78 = W*in
   wire signed [9:0] m380_78;
   assign m380_78 =10'b0;

   // m380_79 = W*in
   wire signed [9:0] m380_79;
   assign m380_79 =10'b0;

   // m380_80 = W*in
   wire signed [9:0] m380_80;
   assign m380_80 =10'b0;

   // m380_81 = W*in
   wire signed [9:0] m380_81;
   assign m380_81 ={ {4{in380[5]}} , in380[5:0] };

   // m380_82 = W*in
   wire signed [9:0] m380_82;
   assign m380_82 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_83 = W*in
   wire signed [9:0] m380_83;
   assign m380_83 =10'b0;

   // m380_84 = W*in
   wire signed [9:0] m380_84;
   assign m380_84 =10'b0;

   // m380_85 = W*in
   wire signed [9:0] m380_85;
   assign m380_85 =10'b0;

   // m380_86 = W*in
   wire signed [9:0] m380_86;
   assign m380_86 =10'b0;

   // m380_87 = W*in
   wire signed [9:0] m380_87;
   assign m380_87 =10'b0;

   // m380_88 = W*in
   wire signed [9:0] m380_88;
   assign m380_88 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_89 = W*in
   wire signed [9:0] m380_89;
   assign m380_89 =10'b0;

   // m380_90 = W*in
   wire signed [9:0] m380_90;
   assign m380_90 =10'b0;

   // m380_91 = W*in
   wire signed [9:0] m380_91;
   assign m380_91 =10'b0;

   // m380_92 = W*in
   wire signed [9:0] m380_92;
   assign m380_92 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_93 = W*in
   wire signed [9:0] m380_93;
   assign m380_93 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_94 = W*in
   wire signed [9:0] m380_94;
   assign m380_94 =10'b0;

   // m380_95 = W*in
   wire signed [9:0] m380_95;
   assign m380_95 =10'b0;

   // m380_96 = W*in
   wire signed [9:0] m380_96;
   assign m380_96 ={ {4{neg380[5]}} , neg380[5:0] };

   // m380_97 = W*in
   wire signed [9:0] m380_97;
   assign m380_97 =10'b0;

   // m380_98 = W*in
   wire signed [9:0] m380_98;
   assign m380_98 =10'b0;

   // m380_99 = W*in
   wire signed [9:0] m380_99;
   assign m380_99 =10'b0;

   // m380_100 = W*in
   wire signed [9:0] m380_100;
   assign m380_100 =10'b0;

   // m380_101 = W*in
   wire signed [9:0] m380_101;
   assign m380_101 =10'b0;

   // m380_102 = W*in
   wire signed [9:0] m380_102;
   assign m380_102 =10'b0;

   // m380_103 = W*in
   wire signed [9:0] m380_103;
   assign m380_103 =10'b0;

   // m380_104 = W*in
   wire signed [9:0] m380_104;
   assign m380_104 =10'b0;

   // m380_105 = W*in
   wire signed [9:0] m380_105;
   assign m380_105 =10'b0;

   // m380_106 = W*in
   wire signed [9:0] m380_106;
   assign m380_106 =10'b0;

   // m380_107 = W*in
   wire signed [9:0] m380_107;
   assign m380_107 =10'b0;

   // m380_108 = W*in
   wire signed [9:0] m380_108;
   assign m380_108 =10'b0;

   // m380_109 = W*in
   wire signed [9:0] m380_109;
   assign m380_109 =10'b0;

   // m380_110 = W*in
   wire signed [9:0] m380_110;
   assign m380_110 =10'b0;

   // m380_111 = W*in
   wire signed [9:0] m380_111;
   assign m380_111 ={ {5{neg380[5]}} , neg380[5:1] };

   // m380_112 = W*in
   wire signed [9:0] m380_112;
   assign m380_112 =10'b0;

   // m380_113 = W*in
   wire signed [9:0] m380_113;
   assign m380_113 =10'b0;

   // m380_114 = W*in
   wire signed [9:0] m380_114;
   assign m380_114 =10'b0;

   // m380_115 = W*in
   wire signed [9:0] m380_115;
   assign m380_115 ={ {4{in380[5]}} , in380[5:0] };

   // m380_116 = W*in
   wire signed [9:0] m380_116;
   assign m380_116 =10'b0;

   // m380_117 = W*in
   wire signed [9:0] m380_117;
   assign m380_117 =10'b0;

   // m381_1 = W*in
   wire signed [9:0] m381_1;
   assign m381_1 =10'b0;

   // m381_2 = W*in
   wire signed [9:0] m381_2;
   assign m381_2 =10'b0;

   // m381_3 = W*in
   wire signed [9:0] m381_3;
   assign m381_3 =10'b0;

   // m381_4 = W*in
   wire signed [9:0] m381_4;
   assign m381_4 =10'b0;

   // m381_5 = W*in
   wire signed [9:0] m381_5;
   assign m381_5 =10'b0;

   // m381_6 = W*in
   wire signed [9:0] m381_6;
   assign m381_6 =10'b0;

   // m381_7 = W*in
   wire signed [9:0] m381_7;
   assign m381_7 =10'b0;

   // m381_8 = W*in
   wire signed [9:0] m381_8;
   assign m381_8 =10'b0;

   // m381_9 = W*in
   wire signed [9:0] m381_9;
   assign m381_9 =10'b0;

   // m381_10 = W*in
   wire signed [9:0] m381_10;
   assign m381_10 =10'b0;

   // m381_11 = W*in
   wire signed [9:0] m381_11;
   assign m381_11 =10'b0;

   // m381_12 = W*in
   wire signed [9:0] m381_12;
   assign m381_12 =10'b0;

   // m381_13 = W*in
   wire signed [9:0] m381_13;
   assign m381_13 =10'b0;

   // m381_14 = W*in
   wire signed [9:0] m381_14;
   assign m381_14 =10'b0;

   // m381_15 = W*in
   wire signed [9:0] m381_15;
   assign m381_15 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_16 = W*in
   wire signed [9:0] m381_16;
   assign m381_16 =10'b0;

   // m381_17 = W*in
   wire signed [9:0] m381_17;
   assign m381_17 =10'b0;

   // m381_18 = W*in
   wire signed [9:0] m381_18;
   assign m381_18 =10'b0;

   // m381_19 = W*in
   wire signed [9:0] m381_19;
   assign m381_19 ={ {5{neg381[5]}} , neg381[5:1] };

   // m381_20 = W*in
   wire signed [9:0] m381_20;
   assign m381_20 =10'b0;

   // m381_21 = W*in
   wire signed [9:0] m381_21;
   assign m381_21 =10'b0;

   // m381_22 = W*in
   wire signed [9:0] m381_22;
   assign m381_22 =10'b0;

   // m381_23 = W*in
   wire signed [9:0] m381_23;
   assign m381_23 =10'b0;

   // m381_24 = W*in
   wire signed [9:0] m381_24;
   assign m381_24 =10'b0;

   // m381_25 = W*in
   wire signed [9:0] m381_25;
   assign m381_25 =10'b0;

   // m381_26 = W*in
   wire signed [9:0] m381_26;
   assign m381_26 =10'b0;

   // m381_27 = W*in
   wire signed [9:0] m381_27;
   assign m381_27 ={ {4{in381[5]}} , in381[5:0] };

   // m381_28 = W*in
   wire signed [9:0] m381_28;
   assign m381_28 ={ {5{in381[5]}} , in381[5:1] };

   // m381_29 = W*in
   wire signed [9:0] m381_29;
   assign m381_29 =10'b0;

   // m381_30 = W*in
   wire signed [9:0] m381_30;
   assign m381_30 =10'b0;

   // m381_31 = W*in
   wire signed [9:0] m381_31;
   assign m381_31 =10'b0;

   // m381_32 = W*in
   wire signed [9:0] m381_32;
   assign m381_32 =10'b0;

   // m381_33 = W*in
   wire signed [9:0] m381_33;
   assign m381_33 =10'b0;

   // m381_34 = W*in
   wire signed [9:0] m381_34;
   assign m381_34 =10'b0;

   // m381_35 = W*in
   wire signed [9:0] m381_35;
   assign m381_35 ={ {4{in381[5]}} , in381[5:0] };

   // m381_36 = W*in
   wire signed [9:0] m381_36;
   assign m381_36 =10'b0;

   // m381_37 = W*in
   wire signed [9:0] m381_37;
   assign m381_37 =10'b0;

   // m381_38 = W*in
   wire signed [9:0] m381_38;
   assign m381_38 =10'b0;

   // m381_39 = W*in
   wire signed [9:0] m381_39;
   assign m381_39 ={ {4{in381[5]}} , in381[5:0] };

   // m381_40 = W*in
   wire signed [9:0] m381_40;
   assign m381_40 =10'b0;

   // m381_41 = W*in
   wire signed [9:0] m381_41;
   assign m381_41 =10'b0;

   // m381_42 = W*in
   wire signed [9:0] m381_42;
   assign m381_42 =10'b0;

   // m381_43 = W*in
   wire signed [9:0] m381_43;
   assign m381_43 =10'b0;

   // m381_44 = W*in
   wire signed [9:0] m381_44;
   assign m381_44 =10'b0;

   // m381_45 = W*in
   wire signed [9:0] m381_45;
   assign m381_45 =10'b0;

   // m381_46 = W*in
   wire signed [9:0] m381_46;
   assign m381_46 =10'b0;

   // m381_47 = W*in
   wire signed [9:0] m381_47;
   assign m381_47 =10'b0;

   // m381_48 = W*in
   wire signed [9:0] m381_48;
   assign m381_48 =10'b0;

   // m381_49 = W*in
   wire signed [9:0] m381_49;
   assign m381_49 =10'b0;

   // m381_50 = W*in
   wire signed [9:0] m381_50;
   assign m381_50 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_51 = W*in
   wire signed [9:0] m381_51;
   assign m381_51 =10'b0;

   // m381_52 = W*in
   wire signed [9:0] m381_52;
   assign m381_52 =10'b0;

   // m381_53 = W*in
   wire signed [9:0] m381_53;
   assign m381_53 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_54 = W*in
   wire signed [9:0] m381_54;
   assign m381_54 =10'b0;

   // m381_55 = W*in
   wire signed [9:0] m381_55;
   assign m381_55 =10'b0;

   // m381_56 = W*in
   wire signed [9:0] m381_56;
   assign m381_56 =10'b0;

   // m381_57 = W*in
   wire signed [9:0] m381_57;
   assign m381_57 ={ {4{in381[5]}} , in381[5:0] };

   // m381_58 = W*in
   wire signed [9:0] m381_58;
   assign m381_58 =10'b0;

   // m381_59 = W*in
   wire signed [9:0] m381_59;
   assign m381_59 =10'b0;

   // m381_60 = W*in
   wire signed [9:0] m381_60;
   assign m381_60 ={ {4{in381[5]}} , in381[5:0] };

   // m381_61 = W*in
   wire signed [9:0] m381_61;
   assign m381_61 ={ {4{in381[5]}} , in381[5:0] };

   // m381_62 = W*in
   wire signed [9:0] m381_62;
   assign m381_62 =10'b0;

   // m381_63 = W*in
   wire signed [9:0] m381_63;
   assign m381_63 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_64 = W*in
   wire signed [9:0] m381_64;
   assign m381_64 =10'b0;

   // m381_65 = W*in
   wire signed [9:0] m381_65;
   assign m381_65 ={ {5{neg381[5]}} , neg381[5:1] };

   // m381_66 = W*in
   wire signed [9:0] m381_66;
   assign m381_66 =10'b0;

   // m381_67 = W*in
   wire signed [9:0] m381_67;
   assign m381_67 =10'b0;

   // m381_68 = W*in
   wire signed [9:0] m381_68;
   assign m381_68 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_69 = W*in
   wire signed [9:0] m381_69;
   assign m381_69 ={ {5{neg381[5]}} , neg381[5:1] };

   // m381_70 = W*in
   wire signed [9:0] m381_70;
   assign m381_70 =10'b0;

   // m381_71 = W*in
   wire signed [9:0] m381_71;
   assign m381_71 =10'b0;

   // m381_72 = W*in
   wire signed [9:0] m381_72;
   assign m381_72 ={ {5{neg381[5]}} , neg381[5:1] };

   // m381_73 = W*in
   wire signed [9:0] m381_73;
   assign m381_73 =10'b0;

   // m381_74 = W*in
   wire signed [9:0] m381_74;
   assign m381_74 =10'b0;

   // m381_75 = W*in
   wire signed [9:0] m381_75;
   assign m381_75 =10'b0;

   // m381_76 = W*in
   wire signed [9:0] m381_76;
   assign m381_76 =10'b0;

   // m381_77 = W*in
   wire signed [9:0] m381_77;
   assign m381_77 =10'b0;

   // m381_78 = W*in
   wire signed [9:0] m381_78;
   assign m381_78 =10'b0;

   // m381_79 = W*in
   wire signed [9:0] m381_79;
   assign m381_79 =10'b0;

   // m381_80 = W*in
   wire signed [9:0] m381_80;
   assign m381_80 =10'b0;

   // m381_81 = W*in
   wire signed [9:0] m381_81;
   assign m381_81 ={ {5{neg381[5]}} , neg381[5:1] };

   // m381_82 = W*in
   wire signed [9:0] m381_82;
   assign m381_82 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_83 = W*in
   wire signed [9:0] m381_83;
   assign m381_83 =10'b0;

   // m381_84 = W*in
   wire signed [9:0] m381_84;
   assign m381_84 =10'b0;

   // m381_85 = W*in
   wire signed [9:0] m381_85;
   assign m381_85 =10'b0;

   // m381_86 = W*in
   wire signed [9:0] m381_86;
   assign m381_86 =10'b0;

   // m381_87 = W*in
   wire signed [9:0] m381_87;
   assign m381_87 =10'b0;

   // m381_88 = W*in
   wire signed [9:0] m381_88;
   assign m381_88 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_89 = W*in
   wire signed [9:0] m381_89;
   assign m381_89 =10'b0;

   // m381_90 = W*in
   wire signed [9:0] m381_90;
   assign m381_90 =10'b0;

   // m381_91 = W*in
   wire signed [9:0] m381_91;
   assign m381_91 =10'b0;

   // m381_92 = W*in
   wire signed [9:0] m381_92;
   assign m381_92 ={ {4{neg381[5]}} , neg381[5:0] };

   // m381_93 = W*in
   wire signed [9:0] m381_93;
   assign m381_93 =10'b0;

   // m381_94 = W*in
   wire signed [9:0] m381_94;
   assign m381_94 =10'b0;

   // m381_95 = W*in
   wire signed [9:0] m381_95;
   assign m381_95 =10'b0;

   // m381_96 = W*in
   wire signed [9:0] m381_96;
   assign m381_96 =10'b0;

   // m381_97 = W*in
   wire signed [9:0] m381_97;
   assign m381_97 =10'b0;

   // m381_98 = W*in
   wire signed [9:0] m381_98;
   assign m381_98 =10'b0;

   // m381_99 = W*in
   wire signed [9:0] m381_99;
   assign m381_99 =10'b0;

   // m381_100 = W*in
   wire signed [9:0] m381_100;
   assign m381_100 =10'b0;

   // m381_101 = W*in
   wire signed [9:0] m381_101;
   assign m381_101 =10'b0;

   // m381_102 = W*in
   wire signed [9:0] m381_102;
   assign m381_102 =10'b0;

   // m381_103 = W*in
   wire signed [9:0] m381_103;
   assign m381_103 =10'b0;

   // m381_104 = W*in
   wire signed [9:0] m381_104;
   assign m381_104 =10'b0;

   // m381_105 = W*in
   wire signed [9:0] m381_105;
   assign m381_105 =10'b0;

   // m381_106 = W*in
   wire signed [9:0] m381_106;
   assign m381_106 =10'b0;

   // m381_107 = W*in
   wire signed [9:0] m381_107;
   assign m381_107 ={ {4{in381[5]}} , in381[5:0] };

   // m381_108 = W*in
   wire signed [9:0] m381_108;
   assign m381_108 =10'b0;

   // m381_109 = W*in
   wire signed [9:0] m381_109;
   assign m381_109 =10'b0;

   // m381_110 = W*in
   wire signed [9:0] m381_110;
   assign m381_110 =10'b0;

   // m381_111 = W*in
   wire signed [9:0] m381_111;
   assign m381_111 =10'b0;

   // m381_112 = W*in
   wire signed [9:0] m381_112;
   assign m381_112 =10'b0;

   // m381_113 = W*in
   wire signed [9:0] m381_113;
   assign m381_113 =10'b0;

   // m381_114 = W*in
   wire signed [9:0] m381_114;
   assign m381_114 =10'b0;

   // m381_115 = W*in
   wire signed [9:0] m381_115;
   assign m381_115 =10'b0;

   // m381_116 = W*in
   wire signed [9:0] m381_116;
   assign m381_116 =10'b0;

   // m381_117 = W*in
   wire signed [9:0] m381_117;
   assign m381_117 ={ {4{in381[5]}} , in381[5:0] };

   //Perceptron Adders
   always @(posedge clk) out1 <= m1_1+m2_1+m3_1+m4_1+m5_1+m6_1+m7_1+m8_1+m9_1+m10_1+m11_1+m12_1+m13_1+m14_1+m15_1+m16_1+m17_1+m18_1+m19_1+m20_1+m21_1+m22_1+m23_1+m24_1+m25_1+m26_1+m27_1+m28_1+m29_1+m30_1+m31_1+m32_1+m33_1+m34_1+m35_1+m36_1+m37_1+m38_1+m39_1+m40_1+m41_1+m42_1+m43_1+m44_1+m45_1+m46_1+m47_1+m48_1+m49_1+m50_1+m51_1+m52_1+m53_1+m54_1+m55_1+m56_1+m57_1+m58_1+m59_1+m60_1+m61_1+m62_1+m63_1+m64_1+m65_1+m66_1+m67_1+m68_1+m69_1+m70_1+m71_1+m72_1+m73_1+m74_1+m75_1+m76_1+m77_1+m78_1+m79_1+m80_1+m81_1+m82_1+m83_1+m84_1+m85_1+m86_1+m87_1+m88_1+m89_1+m90_1+m91_1+m92_1+m93_1+m94_1+m95_1+m96_1+m97_1+m98_1+m99_1+m100_1+m101_1+m102_1+m103_1+m104_1+m105_1+m106_1+m107_1+m108_1+m109_1+m110_1+m111_1+m112_1+m113_1+m114_1+m115_1+m116_1+m117_1+m118_1+m119_1+m120_1+m121_1+m122_1+m123_1+m124_1+m125_1+m126_1+m127_1+m128_1+m129_1+m130_1+m131_1+m132_1+m133_1+m134_1+m135_1+m136_1+m137_1+m138_1+m139_1+m140_1+m141_1+m142_1+m143_1+m144_1+m145_1+m146_1+m147_1+m148_1+m149_1+m150_1+m151_1+m152_1+m153_1+m154_1+m155_1+m156_1+m157_1+m158_1+m159_1+m160_1+m161_1+m162_1+m163_1+m164_1+m165_1+m166_1+m167_1+m168_1+m169_1+m170_1+m171_1+m172_1+m173_1+m174_1+m175_1+m176_1+m177_1+m178_1+m179_1+m180_1+m181_1+m182_1+m183_1+m184_1+m185_1+m186_1+m187_1+m188_1+m189_1+m190_1+m191_1+m192_1+m193_1+m194_1+m195_1+m196_1+m197_1+m198_1+m199_1+m200_1+m201_1+m202_1+m203_1+m204_1+m205_1+m206_1+m207_1+m208_1+m209_1+m210_1+m211_1+m212_1+m213_1+m214_1+m215_1+m216_1+m217_1+m218_1+m219_1+m220_1+m221_1+m222_1+m223_1+m224_1+m225_1+m226_1+m227_1+m228_1+m229_1+m230_1+m231_1+m232_1+m233_1+m234_1+m235_1+m236_1+m237_1+m238_1+m239_1+m240_1+m241_1+m242_1+m243_1+m244_1+m245_1+m246_1+m247_1+m248_1+m249_1+m250_1+m251_1+m252_1+m253_1+m254_1+m255_1+m256_1+m257_1+m258_1+m259_1+m260_1+m261_1+m262_1+m263_1+m264_1+m265_1+m266_1+m267_1+m268_1+m269_1+m270_1+m271_1+m272_1+m273_1+m274_1+m275_1+m276_1+m277_1+m278_1+m279_1+m280_1+m281_1+m282_1+m283_1+m284_1+m285_1+m286_1+m287_1+m288_1+m289_1+m290_1+m291_1+m292_1+m293_1+m294_1+m295_1+m296_1+m297_1+m298_1+m299_1+m300_1+m301_1+m302_1+m303_1+m304_1+m305_1+m306_1+m307_1+m308_1+m309_1+m310_1+m311_1+m312_1+m313_1+m314_1+m315_1+m316_1+m317_1+m318_1+m319_1+m320_1+m321_1+m322_1+m323_1+m324_1+m325_1+m326_1+m327_1+m328_1+m329_1+m330_1+m331_1+m332_1+m333_1+m334_1+m335_1+m336_1+m337_1+m338_1+m339_1+m340_1+m341_1+m342_1+m343_1+m344_1+m345_1+m346_1+m347_1+m348_1+m349_1+m350_1+m351_1+m352_1+m353_1+m354_1+m355_1+m356_1+m357_1+m358_1+m359_1+m360_1+m361_1+m362_1+m363_1+m364_1+m365_1+m366_1+m367_1+m368_1+m369_1+m370_1+m371_1+m372_1+m373_1+m374_1+m375_1+m376_1+m377_1+m378_1+m379_1+m380_1+m381_1+b1;
   always @(posedge clk) out2 <= m1_2+m2_2+m3_2+m4_2+m5_2+m6_2+m7_2+m8_2+m9_2+m10_2+m11_2+m12_2+m13_2+m14_2+m15_2+m16_2+m17_2+m18_2+m19_2+m20_2+m21_2+m22_2+m23_2+m24_2+m25_2+m26_2+m27_2+m28_2+m29_2+m30_2+m31_2+m32_2+m33_2+m34_2+m35_2+m36_2+m37_2+m38_2+m39_2+m40_2+m41_2+m42_2+m43_2+m44_2+m45_2+m46_2+m47_2+m48_2+m49_2+m50_2+m51_2+m52_2+m53_2+m54_2+m55_2+m56_2+m57_2+m58_2+m59_2+m60_2+m61_2+m62_2+m63_2+m64_2+m65_2+m66_2+m67_2+m68_2+m69_2+m70_2+m71_2+m72_2+m73_2+m74_2+m75_2+m76_2+m77_2+m78_2+m79_2+m80_2+m81_2+m82_2+m83_2+m84_2+m85_2+m86_2+m87_2+m88_2+m89_2+m90_2+m91_2+m92_2+m93_2+m94_2+m95_2+m96_2+m97_2+m98_2+m99_2+m100_2+m101_2+m102_2+m103_2+m104_2+m105_2+m106_2+m107_2+m108_2+m109_2+m110_2+m111_2+m112_2+m113_2+m114_2+m115_2+m116_2+m117_2+m118_2+m119_2+m120_2+m121_2+m122_2+m123_2+m124_2+m125_2+m126_2+m127_2+m128_2+m129_2+m130_2+m131_2+m132_2+m133_2+m134_2+m135_2+m136_2+m137_2+m138_2+m139_2+m140_2+m141_2+m142_2+m143_2+m144_2+m145_2+m146_2+m147_2+m148_2+m149_2+m150_2+m151_2+m152_2+m153_2+m154_2+m155_2+m156_2+m157_2+m158_2+m159_2+m160_2+m161_2+m162_2+m163_2+m164_2+m165_2+m166_2+m167_2+m168_2+m169_2+m170_2+m171_2+m172_2+m173_2+m174_2+m175_2+m176_2+m177_2+m178_2+m179_2+m180_2+m181_2+m182_2+m183_2+m184_2+m185_2+m186_2+m187_2+m188_2+m189_2+m190_2+m191_2+m192_2+m193_2+m194_2+m195_2+m196_2+m197_2+m198_2+m199_2+m200_2+m201_2+m202_2+m203_2+m204_2+m205_2+m206_2+m207_2+m208_2+m209_2+m210_2+m211_2+m212_2+m213_2+m214_2+m215_2+m216_2+m217_2+m218_2+m219_2+m220_2+m221_2+m222_2+m223_2+m224_2+m225_2+m226_2+m227_2+m228_2+m229_2+m230_2+m231_2+m232_2+m233_2+m234_2+m235_2+m236_2+m237_2+m238_2+m239_2+m240_2+m241_2+m242_2+m243_2+m244_2+m245_2+m246_2+m247_2+m248_2+m249_2+m250_2+m251_2+m252_2+m253_2+m254_2+m255_2+m256_2+m257_2+m258_2+m259_2+m260_2+m261_2+m262_2+m263_2+m264_2+m265_2+m266_2+m267_2+m268_2+m269_2+m270_2+m271_2+m272_2+m273_2+m274_2+m275_2+m276_2+m277_2+m278_2+m279_2+m280_2+m281_2+m282_2+m283_2+m284_2+m285_2+m286_2+m287_2+m288_2+m289_2+m290_2+m291_2+m292_2+m293_2+m294_2+m295_2+m296_2+m297_2+m298_2+m299_2+m300_2+m301_2+m302_2+m303_2+m304_2+m305_2+m306_2+m307_2+m308_2+m309_2+m310_2+m311_2+m312_2+m313_2+m314_2+m315_2+m316_2+m317_2+m318_2+m319_2+m320_2+m321_2+m322_2+m323_2+m324_2+m325_2+m326_2+m327_2+m328_2+m329_2+m330_2+m331_2+m332_2+m333_2+m334_2+m335_2+m336_2+m337_2+m338_2+m339_2+m340_2+m341_2+m342_2+m343_2+m344_2+m345_2+m346_2+m347_2+m348_2+m349_2+m350_2+m351_2+m352_2+m353_2+m354_2+m355_2+m356_2+m357_2+m358_2+m359_2+m360_2+m361_2+m362_2+m363_2+m364_2+m365_2+m366_2+m367_2+m368_2+m369_2+m370_2+m371_2+m372_2+m373_2+m374_2+m375_2+m376_2+m377_2+m378_2+m379_2+m380_2+m381_2+b2;
   always @(posedge clk) out3 <= m1_3+m2_3+m3_3+m4_3+m5_3+m6_3+m7_3+m8_3+m9_3+m10_3+m11_3+m12_3+m13_3+m14_3+m15_3+m16_3+m17_3+m18_3+m19_3+m20_3+m21_3+m22_3+m23_3+m24_3+m25_3+m26_3+m27_3+m28_3+m29_3+m30_3+m31_3+m32_3+m33_3+m34_3+m35_3+m36_3+m37_3+m38_3+m39_3+m40_3+m41_3+m42_3+m43_3+m44_3+m45_3+m46_3+m47_3+m48_3+m49_3+m50_3+m51_3+m52_3+m53_3+m54_3+m55_3+m56_3+m57_3+m58_3+m59_3+m60_3+m61_3+m62_3+m63_3+m64_3+m65_3+m66_3+m67_3+m68_3+m69_3+m70_3+m71_3+m72_3+m73_3+m74_3+m75_3+m76_3+m77_3+m78_3+m79_3+m80_3+m81_3+m82_3+m83_3+m84_3+m85_3+m86_3+m87_3+m88_3+m89_3+m90_3+m91_3+m92_3+m93_3+m94_3+m95_3+m96_3+m97_3+m98_3+m99_3+m100_3+m101_3+m102_3+m103_3+m104_3+m105_3+m106_3+m107_3+m108_3+m109_3+m110_3+m111_3+m112_3+m113_3+m114_3+m115_3+m116_3+m117_3+m118_3+m119_3+m120_3+m121_3+m122_3+m123_3+m124_3+m125_3+m126_3+m127_3+m128_3+m129_3+m130_3+m131_3+m132_3+m133_3+m134_3+m135_3+m136_3+m137_3+m138_3+m139_3+m140_3+m141_3+m142_3+m143_3+m144_3+m145_3+m146_3+m147_3+m148_3+m149_3+m150_3+m151_3+m152_3+m153_3+m154_3+m155_3+m156_3+m157_3+m158_3+m159_3+m160_3+m161_3+m162_3+m163_3+m164_3+m165_3+m166_3+m167_3+m168_3+m169_3+m170_3+m171_3+m172_3+m173_3+m174_3+m175_3+m176_3+m177_3+m178_3+m179_3+m180_3+m181_3+m182_3+m183_3+m184_3+m185_3+m186_3+m187_3+m188_3+m189_3+m190_3+m191_3+m192_3+m193_3+m194_3+m195_3+m196_3+m197_3+m198_3+m199_3+m200_3+m201_3+m202_3+m203_3+m204_3+m205_3+m206_3+m207_3+m208_3+m209_3+m210_3+m211_3+m212_3+m213_3+m214_3+m215_3+m216_3+m217_3+m218_3+m219_3+m220_3+m221_3+m222_3+m223_3+m224_3+m225_3+m226_3+m227_3+m228_3+m229_3+m230_3+m231_3+m232_3+m233_3+m234_3+m235_3+m236_3+m237_3+m238_3+m239_3+m240_3+m241_3+m242_3+m243_3+m244_3+m245_3+m246_3+m247_3+m248_3+m249_3+m250_3+m251_3+m252_3+m253_3+m254_3+m255_3+m256_3+m257_3+m258_3+m259_3+m260_3+m261_3+m262_3+m263_3+m264_3+m265_3+m266_3+m267_3+m268_3+m269_3+m270_3+m271_3+m272_3+m273_3+m274_3+m275_3+m276_3+m277_3+m278_3+m279_3+m280_3+m281_3+m282_3+m283_3+m284_3+m285_3+m286_3+m287_3+m288_3+m289_3+m290_3+m291_3+m292_3+m293_3+m294_3+m295_3+m296_3+m297_3+m298_3+m299_3+m300_3+m301_3+m302_3+m303_3+m304_3+m305_3+m306_3+m307_3+m308_3+m309_3+m310_3+m311_3+m312_3+m313_3+m314_3+m315_3+m316_3+m317_3+m318_3+m319_3+m320_3+m321_3+m322_3+m323_3+m324_3+m325_3+m326_3+m327_3+m328_3+m329_3+m330_3+m331_3+m332_3+m333_3+m334_3+m335_3+m336_3+m337_3+m338_3+m339_3+m340_3+m341_3+m342_3+m343_3+m344_3+m345_3+m346_3+m347_3+m348_3+m349_3+m350_3+m351_3+m352_3+m353_3+m354_3+m355_3+m356_3+m357_3+m358_3+m359_3+m360_3+m361_3+m362_3+m363_3+m364_3+m365_3+m366_3+m367_3+m368_3+m369_3+m370_3+m371_3+m372_3+m373_3+m374_3+m375_3+m376_3+m377_3+m378_3+m379_3+m380_3+m381_3+b3;
   always @(posedge clk) out4 <= m1_4+m2_4+m3_4+m4_4+m5_4+m6_4+m7_4+m8_4+m9_4+m10_4+m11_4+m12_4+m13_4+m14_4+m15_4+m16_4+m17_4+m18_4+m19_4+m20_4+m21_4+m22_4+m23_4+m24_4+m25_4+m26_4+m27_4+m28_4+m29_4+m30_4+m31_4+m32_4+m33_4+m34_4+m35_4+m36_4+m37_4+m38_4+m39_4+m40_4+m41_4+m42_4+m43_4+m44_4+m45_4+m46_4+m47_4+m48_4+m49_4+m50_4+m51_4+m52_4+m53_4+m54_4+m55_4+m56_4+m57_4+m58_4+m59_4+m60_4+m61_4+m62_4+m63_4+m64_4+m65_4+m66_4+m67_4+m68_4+m69_4+m70_4+m71_4+m72_4+m73_4+m74_4+m75_4+m76_4+m77_4+m78_4+m79_4+m80_4+m81_4+m82_4+m83_4+m84_4+m85_4+m86_4+m87_4+m88_4+m89_4+m90_4+m91_4+m92_4+m93_4+m94_4+m95_4+m96_4+m97_4+m98_4+m99_4+m100_4+m101_4+m102_4+m103_4+m104_4+m105_4+m106_4+m107_4+m108_4+m109_4+m110_4+m111_4+m112_4+m113_4+m114_4+m115_4+m116_4+m117_4+m118_4+m119_4+m120_4+m121_4+m122_4+m123_4+m124_4+m125_4+m126_4+m127_4+m128_4+m129_4+m130_4+m131_4+m132_4+m133_4+m134_4+m135_4+m136_4+m137_4+m138_4+m139_4+m140_4+m141_4+m142_4+m143_4+m144_4+m145_4+m146_4+m147_4+m148_4+m149_4+m150_4+m151_4+m152_4+m153_4+m154_4+m155_4+m156_4+m157_4+m158_4+m159_4+m160_4+m161_4+m162_4+m163_4+m164_4+m165_4+m166_4+m167_4+m168_4+m169_4+m170_4+m171_4+m172_4+m173_4+m174_4+m175_4+m176_4+m177_4+m178_4+m179_4+m180_4+m181_4+m182_4+m183_4+m184_4+m185_4+m186_4+m187_4+m188_4+m189_4+m190_4+m191_4+m192_4+m193_4+m194_4+m195_4+m196_4+m197_4+m198_4+m199_4+m200_4+m201_4+m202_4+m203_4+m204_4+m205_4+m206_4+m207_4+m208_4+m209_4+m210_4+m211_4+m212_4+m213_4+m214_4+m215_4+m216_4+m217_4+m218_4+m219_4+m220_4+m221_4+m222_4+m223_4+m224_4+m225_4+m226_4+m227_4+m228_4+m229_4+m230_4+m231_4+m232_4+m233_4+m234_4+m235_4+m236_4+m237_4+m238_4+m239_4+m240_4+m241_4+m242_4+m243_4+m244_4+m245_4+m246_4+m247_4+m248_4+m249_4+m250_4+m251_4+m252_4+m253_4+m254_4+m255_4+m256_4+m257_4+m258_4+m259_4+m260_4+m261_4+m262_4+m263_4+m264_4+m265_4+m266_4+m267_4+m268_4+m269_4+m270_4+m271_4+m272_4+m273_4+m274_4+m275_4+m276_4+m277_4+m278_4+m279_4+m280_4+m281_4+m282_4+m283_4+m284_4+m285_4+m286_4+m287_4+m288_4+m289_4+m290_4+m291_4+m292_4+m293_4+m294_4+m295_4+m296_4+m297_4+m298_4+m299_4+m300_4+m301_4+m302_4+m303_4+m304_4+m305_4+m306_4+m307_4+m308_4+m309_4+m310_4+m311_4+m312_4+m313_4+m314_4+m315_4+m316_4+m317_4+m318_4+m319_4+m320_4+m321_4+m322_4+m323_4+m324_4+m325_4+m326_4+m327_4+m328_4+m329_4+m330_4+m331_4+m332_4+m333_4+m334_4+m335_4+m336_4+m337_4+m338_4+m339_4+m340_4+m341_4+m342_4+m343_4+m344_4+m345_4+m346_4+m347_4+m348_4+m349_4+m350_4+m351_4+m352_4+m353_4+m354_4+m355_4+m356_4+m357_4+m358_4+m359_4+m360_4+m361_4+m362_4+m363_4+m364_4+m365_4+m366_4+m367_4+m368_4+m369_4+m370_4+m371_4+m372_4+m373_4+m374_4+m375_4+m376_4+m377_4+m378_4+m379_4+m380_4+m381_4+b4;
   always @(posedge clk) out5 <= m1_5+m2_5+m3_5+m4_5+m5_5+m6_5+m7_5+m8_5+m9_5+m10_5+m11_5+m12_5+m13_5+m14_5+m15_5+m16_5+m17_5+m18_5+m19_5+m20_5+m21_5+m22_5+m23_5+m24_5+m25_5+m26_5+m27_5+m28_5+m29_5+m30_5+m31_5+m32_5+m33_5+m34_5+m35_5+m36_5+m37_5+m38_5+m39_5+m40_5+m41_5+m42_5+m43_5+m44_5+m45_5+m46_5+m47_5+m48_5+m49_5+m50_5+m51_5+m52_5+m53_5+m54_5+m55_5+m56_5+m57_5+m58_5+m59_5+m60_5+m61_5+m62_5+m63_5+m64_5+m65_5+m66_5+m67_5+m68_5+m69_5+m70_5+m71_5+m72_5+m73_5+m74_5+m75_5+m76_5+m77_5+m78_5+m79_5+m80_5+m81_5+m82_5+m83_5+m84_5+m85_5+m86_5+m87_5+m88_5+m89_5+m90_5+m91_5+m92_5+m93_5+m94_5+m95_5+m96_5+m97_5+m98_5+m99_5+m100_5+m101_5+m102_5+m103_5+m104_5+m105_5+m106_5+m107_5+m108_5+m109_5+m110_5+m111_5+m112_5+m113_5+m114_5+m115_5+m116_5+m117_5+m118_5+m119_5+m120_5+m121_5+m122_5+m123_5+m124_5+m125_5+m126_5+m127_5+m128_5+m129_5+m130_5+m131_5+m132_5+m133_5+m134_5+m135_5+m136_5+m137_5+m138_5+m139_5+m140_5+m141_5+m142_5+m143_5+m144_5+m145_5+m146_5+m147_5+m148_5+m149_5+m150_5+m151_5+m152_5+m153_5+m154_5+m155_5+m156_5+m157_5+m158_5+m159_5+m160_5+m161_5+m162_5+m163_5+m164_5+m165_5+m166_5+m167_5+m168_5+m169_5+m170_5+m171_5+m172_5+m173_5+m174_5+m175_5+m176_5+m177_5+m178_5+m179_5+m180_5+m181_5+m182_5+m183_5+m184_5+m185_5+m186_5+m187_5+m188_5+m189_5+m190_5+m191_5+m192_5+m193_5+m194_5+m195_5+m196_5+m197_5+m198_5+m199_5+m200_5+m201_5+m202_5+m203_5+m204_5+m205_5+m206_5+m207_5+m208_5+m209_5+m210_5+m211_5+m212_5+m213_5+m214_5+m215_5+m216_5+m217_5+m218_5+m219_5+m220_5+m221_5+m222_5+m223_5+m224_5+m225_5+m226_5+m227_5+m228_5+m229_5+m230_5+m231_5+m232_5+m233_5+m234_5+m235_5+m236_5+m237_5+m238_5+m239_5+m240_5+m241_5+m242_5+m243_5+m244_5+m245_5+m246_5+m247_5+m248_5+m249_5+m250_5+m251_5+m252_5+m253_5+m254_5+m255_5+m256_5+m257_5+m258_5+m259_5+m260_5+m261_5+m262_5+m263_5+m264_5+m265_5+m266_5+m267_5+m268_5+m269_5+m270_5+m271_5+m272_5+m273_5+m274_5+m275_5+m276_5+m277_5+m278_5+m279_5+m280_5+m281_5+m282_5+m283_5+m284_5+m285_5+m286_5+m287_5+m288_5+m289_5+m290_5+m291_5+m292_5+m293_5+m294_5+m295_5+m296_5+m297_5+m298_5+m299_5+m300_5+m301_5+m302_5+m303_5+m304_5+m305_5+m306_5+m307_5+m308_5+m309_5+m310_5+m311_5+m312_5+m313_5+m314_5+m315_5+m316_5+m317_5+m318_5+m319_5+m320_5+m321_5+m322_5+m323_5+m324_5+m325_5+m326_5+m327_5+m328_5+m329_5+m330_5+m331_5+m332_5+m333_5+m334_5+m335_5+m336_5+m337_5+m338_5+m339_5+m340_5+m341_5+m342_5+m343_5+m344_5+m345_5+m346_5+m347_5+m348_5+m349_5+m350_5+m351_5+m352_5+m353_5+m354_5+m355_5+m356_5+m357_5+m358_5+m359_5+m360_5+m361_5+m362_5+m363_5+m364_5+m365_5+m366_5+m367_5+m368_5+m369_5+m370_5+m371_5+m372_5+m373_5+m374_5+m375_5+m376_5+m377_5+m378_5+m379_5+m380_5+m381_5+b5;
   always @(posedge clk) out6 <= m1_6+m2_6+m3_6+m4_6+m5_6+m6_6+m7_6+m8_6+m9_6+m10_6+m11_6+m12_6+m13_6+m14_6+m15_6+m16_6+m17_6+m18_6+m19_6+m20_6+m21_6+m22_6+m23_6+m24_6+m25_6+m26_6+m27_6+m28_6+m29_6+m30_6+m31_6+m32_6+m33_6+m34_6+m35_6+m36_6+m37_6+m38_6+m39_6+m40_6+m41_6+m42_6+m43_6+m44_6+m45_6+m46_6+m47_6+m48_6+m49_6+m50_6+m51_6+m52_6+m53_6+m54_6+m55_6+m56_6+m57_6+m58_6+m59_6+m60_6+m61_6+m62_6+m63_6+m64_6+m65_6+m66_6+m67_6+m68_6+m69_6+m70_6+m71_6+m72_6+m73_6+m74_6+m75_6+m76_6+m77_6+m78_6+m79_6+m80_6+m81_6+m82_6+m83_6+m84_6+m85_6+m86_6+m87_6+m88_6+m89_6+m90_6+m91_6+m92_6+m93_6+m94_6+m95_6+m96_6+m97_6+m98_6+m99_6+m100_6+m101_6+m102_6+m103_6+m104_6+m105_6+m106_6+m107_6+m108_6+m109_6+m110_6+m111_6+m112_6+m113_6+m114_6+m115_6+m116_6+m117_6+m118_6+m119_6+m120_6+m121_6+m122_6+m123_6+m124_6+m125_6+m126_6+m127_6+m128_6+m129_6+m130_6+m131_6+m132_6+m133_6+m134_6+m135_6+m136_6+m137_6+m138_6+m139_6+m140_6+m141_6+m142_6+m143_6+m144_6+m145_6+m146_6+m147_6+m148_6+m149_6+m150_6+m151_6+m152_6+m153_6+m154_6+m155_6+m156_6+m157_6+m158_6+m159_6+m160_6+m161_6+m162_6+m163_6+m164_6+m165_6+m166_6+m167_6+m168_6+m169_6+m170_6+m171_6+m172_6+m173_6+m174_6+m175_6+m176_6+m177_6+m178_6+m179_6+m180_6+m181_6+m182_6+m183_6+m184_6+m185_6+m186_6+m187_6+m188_6+m189_6+m190_6+m191_6+m192_6+m193_6+m194_6+m195_6+m196_6+m197_6+m198_6+m199_6+m200_6+m201_6+m202_6+m203_6+m204_6+m205_6+m206_6+m207_6+m208_6+m209_6+m210_6+m211_6+m212_6+m213_6+m214_6+m215_6+m216_6+m217_6+m218_6+m219_6+m220_6+m221_6+m222_6+m223_6+m224_6+m225_6+m226_6+m227_6+m228_6+m229_6+m230_6+m231_6+m232_6+m233_6+m234_6+m235_6+m236_6+m237_6+m238_6+m239_6+m240_6+m241_6+m242_6+m243_6+m244_6+m245_6+m246_6+m247_6+m248_6+m249_6+m250_6+m251_6+m252_6+m253_6+m254_6+m255_6+m256_6+m257_6+m258_6+m259_6+m260_6+m261_6+m262_6+m263_6+m264_6+m265_6+m266_6+m267_6+m268_6+m269_6+m270_6+m271_6+m272_6+m273_6+m274_6+m275_6+m276_6+m277_6+m278_6+m279_6+m280_6+m281_6+m282_6+m283_6+m284_6+m285_6+m286_6+m287_6+m288_6+m289_6+m290_6+m291_6+m292_6+m293_6+m294_6+m295_6+m296_6+m297_6+m298_6+m299_6+m300_6+m301_6+m302_6+m303_6+m304_6+m305_6+m306_6+m307_6+m308_6+m309_6+m310_6+m311_6+m312_6+m313_6+m314_6+m315_6+m316_6+m317_6+m318_6+m319_6+m320_6+m321_6+m322_6+m323_6+m324_6+m325_6+m326_6+m327_6+m328_6+m329_6+m330_6+m331_6+m332_6+m333_6+m334_6+m335_6+m336_6+m337_6+m338_6+m339_6+m340_6+m341_6+m342_6+m343_6+m344_6+m345_6+m346_6+m347_6+m348_6+m349_6+m350_6+m351_6+m352_6+m353_6+m354_6+m355_6+m356_6+m357_6+m358_6+m359_6+m360_6+m361_6+m362_6+m363_6+m364_6+m365_6+m366_6+m367_6+m368_6+m369_6+m370_6+m371_6+m372_6+m373_6+m374_6+m375_6+m376_6+m377_6+m378_6+m379_6+m380_6+m381_6+b6;
   always @(posedge clk) out7 <= m1_7+m2_7+m3_7+m4_7+m5_7+m6_7+m7_7+m8_7+m9_7+m10_7+m11_7+m12_7+m13_7+m14_7+m15_7+m16_7+m17_7+m18_7+m19_7+m20_7+m21_7+m22_7+m23_7+m24_7+m25_7+m26_7+m27_7+m28_7+m29_7+m30_7+m31_7+m32_7+m33_7+m34_7+m35_7+m36_7+m37_7+m38_7+m39_7+m40_7+m41_7+m42_7+m43_7+m44_7+m45_7+m46_7+m47_7+m48_7+m49_7+m50_7+m51_7+m52_7+m53_7+m54_7+m55_7+m56_7+m57_7+m58_7+m59_7+m60_7+m61_7+m62_7+m63_7+m64_7+m65_7+m66_7+m67_7+m68_7+m69_7+m70_7+m71_7+m72_7+m73_7+m74_7+m75_7+m76_7+m77_7+m78_7+m79_7+m80_7+m81_7+m82_7+m83_7+m84_7+m85_7+m86_7+m87_7+m88_7+m89_7+m90_7+m91_7+m92_7+m93_7+m94_7+m95_7+m96_7+m97_7+m98_7+m99_7+m100_7+m101_7+m102_7+m103_7+m104_7+m105_7+m106_7+m107_7+m108_7+m109_7+m110_7+m111_7+m112_7+m113_7+m114_7+m115_7+m116_7+m117_7+m118_7+m119_7+m120_7+m121_7+m122_7+m123_7+m124_7+m125_7+m126_7+m127_7+m128_7+m129_7+m130_7+m131_7+m132_7+m133_7+m134_7+m135_7+m136_7+m137_7+m138_7+m139_7+m140_7+m141_7+m142_7+m143_7+m144_7+m145_7+m146_7+m147_7+m148_7+m149_7+m150_7+m151_7+m152_7+m153_7+m154_7+m155_7+m156_7+m157_7+m158_7+m159_7+m160_7+m161_7+m162_7+m163_7+m164_7+m165_7+m166_7+m167_7+m168_7+m169_7+m170_7+m171_7+m172_7+m173_7+m174_7+m175_7+m176_7+m177_7+m178_7+m179_7+m180_7+m181_7+m182_7+m183_7+m184_7+m185_7+m186_7+m187_7+m188_7+m189_7+m190_7+m191_7+m192_7+m193_7+m194_7+m195_7+m196_7+m197_7+m198_7+m199_7+m200_7+m201_7+m202_7+m203_7+m204_7+m205_7+m206_7+m207_7+m208_7+m209_7+m210_7+m211_7+m212_7+m213_7+m214_7+m215_7+m216_7+m217_7+m218_7+m219_7+m220_7+m221_7+m222_7+m223_7+m224_7+m225_7+m226_7+m227_7+m228_7+m229_7+m230_7+m231_7+m232_7+m233_7+m234_7+m235_7+m236_7+m237_7+m238_7+m239_7+m240_7+m241_7+m242_7+m243_7+m244_7+m245_7+m246_7+m247_7+m248_7+m249_7+m250_7+m251_7+m252_7+m253_7+m254_7+m255_7+m256_7+m257_7+m258_7+m259_7+m260_7+m261_7+m262_7+m263_7+m264_7+m265_7+m266_7+m267_7+m268_7+m269_7+m270_7+m271_7+m272_7+m273_7+m274_7+m275_7+m276_7+m277_7+m278_7+m279_7+m280_7+m281_7+m282_7+m283_7+m284_7+m285_7+m286_7+m287_7+m288_7+m289_7+m290_7+m291_7+m292_7+m293_7+m294_7+m295_7+m296_7+m297_7+m298_7+m299_7+m300_7+m301_7+m302_7+m303_7+m304_7+m305_7+m306_7+m307_7+m308_7+m309_7+m310_7+m311_7+m312_7+m313_7+m314_7+m315_7+m316_7+m317_7+m318_7+m319_7+m320_7+m321_7+m322_7+m323_7+m324_7+m325_7+m326_7+m327_7+m328_7+m329_7+m330_7+m331_7+m332_7+m333_7+m334_7+m335_7+m336_7+m337_7+m338_7+m339_7+m340_7+m341_7+m342_7+m343_7+m344_7+m345_7+m346_7+m347_7+m348_7+m349_7+m350_7+m351_7+m352_7+m353_7+m354_7+m355_7+m356_7+m357_7+m358_7+m359_7+m360_7+m361_7+m362_7+m363_7+m364_7+m365_7+m366_7+m367_7+m368_7+m369_7+m370_7+m371_7+m372_7+m373_7+m374_7+m375_7+m376_7+m377_7+m378_7+m379_7+m380_7+m381_7+b7;
   always @(posedge clk) out8 <= m1_8+m2_8+m3_8+m4_8+m5_8+m6_8+m7_8+m8_8+m9_8+m10_8+m11_8+m12_8+m13_8+m14_8+m15_8+m16_8+m17_8+m18_8+m19_8+m20_8+m21_8+m22_8+m23_8+m24_8+m25_8+m26_8+m27_8+m28_8+m29_8+m30_8+m31_8+m32_8+m33_8+m34_8+m35_8+m36_8+m37_8+m38_8+m39_8+m40_8+m41_8+m42_8+m43_8+m44_8+m45_8+m46_8+m47_8+m48_8+m49_8+m50_8+m51_8+m52_8+m53_8+m54_8+m55_8+m56_8+m57_8+m58_8+m59_8+m60_8+m61_8+m62_8+m63_8+m64_8+m65_8+m66_8+m67_8+m68_8+m69_8+m70_8+m71_8+m72_8+m73_8+m74_8+m75_8+m76_8+m77_8+m78_8+m79_8+m80_8+m81_8+m82_8+m83_8+m84_8+m85_8+m86_8+m87_8+m88_8+m89_8+m90_8+m91_8+m92_8+m93_8+m94_8+m95_8+m96_8+m97_8+m98_8+m99_8+m100_8+m101_8+m102_8+m103_8+m104_8+m105_8+m106_8+m107_8+m108_8+m109_8+m110_8+m111_8+m112_8+m113_8+m114_8+m115_8+m116_8+m117_8+m118_8+m119_8+m120_8+m121_8+m122_8+m123_8+m124_8+m125_8+m126_8+m127_8+m128_8+m129_8+m130_8+m131_8+m132_8+m133_8+m134_8+m135_8+m136_8+m137_8+m138_8+m139_8+m140_8+m141_8+m142_8+m143_8+m144_8+m145_8+m146_8+m147_8+m148_8+m149_8+m150_8+m151_8+m152_8+m153_8+m154_8+m155_8+m156_8+m157_8+m158_8+m159_8+m160_8+m161_8+m162_8+m163_8+m164_8+m165_8+m166_8+m167_8+m168_8+m169_8+m170_8+m171_8+m172_8+m173_8+m174_8+m175_8+m176_8+m177_8+m178_8+m179_8+m180_8+m181_8+m182_8+m183_8+m184_8+m185_8+m186_8+m187_8+m188_8+m189_8+m190_8+m191_8+m192_8+m193_8+m194_8+m195_8+m196_8+m197_8+m198_8+m199_8+m200_8+m201_8+m202_8+m203_8+m204_8+m205_8+m206_8+m207_8+m208_8+m209_8+m210_8+m211_8+m212_8+m213_8+m214_8+m215_8+m216_8+m217_8+m218_8+m219_8+m220_8+m221_8+m222_8+m223_8+m224_8+m225_8+m226_8+m227_8+m228_8+m229_8+m230_8+m231_8+m232_8+m233_8+m234_8+m235_8+m236_8+m237_8+m238_8+m239_8+m240_8+m241_8+m242_8+m243_8+m244_8+m245_8+m246_8+m247_8+m248_8+m249_8+m250_8+m251_8+m252_8+m253_8+m254_8+m255_8+m256_8+m257_8+m258_8+m259_8+m260_8+m261_8+m262_8+m263_8+m264_8+m265_8+m266_8+m267_8+m268_8+m269_8+m270_8+m271_8+m272_8+m273_8+m274_8+m275_8+m276_8+m277_8+m278_8+m279_8+m280_8+m281_8+m282_8+m283_8+m284_8+m285_8+m286_8+m287_8+m288_8+m289_8+m290_8+m291_8+m292_8+m293_8+m294_8+m295_8+m296_8+m297_8+m298_8+m299_8+m300_8+m301_8+m302_8+m303_8+m304_8+m305_8+m306_8+m307_8+m308_8+m309_8+m310_8+m311_8+m312_8+m313_8+m314_8+m315_8+m316_8+m317_8+m318_8+m319_8+m320_8+m321_8+m322_8+m323_8+m324_8+m325_8+m326_8+m327_8+m328_8+m329_8+m330_8+m331_8+m332_8+m333_8+m334_8+m335_8+m336_8+m337_8+m338_8+m339_8+m340_8+m341_8+m342_8+m343_8+m344_8+m345_8+m346_8+m347_8+m348_8+m349_8+m350_8+m351_8+m352_8+m353_8+m354_8+m355_8+m356_8+m357_8+m358_8+m359_8+m360_8+m361_8+m362_8+m363_8+m364_8+m365_8+m366_8+m367_8+m368_8+m369_8+m370_8+m371_8+m372_8+m373_8+m374_8+m375_8+m376_8+m377_8+m378_8+m379_8+m380_8+m381_8+b8;
   always @(posedge clk) out9 <= m1_9+m2_9+m3_9+m4_9+m5_9+m6_9+m7_9+m8_9+m9_9+m10_9+m11_9+m12_9+m13_9+m14_9+m15_9+m16_9+m17_9+m18_9+m19_9+m20_9+m21_9+m22_9+m23_9+m24_9+m25_9+m26_9+m27_9+m28_9+m29_9+m30_9+m31_9+m32_9+m33_9+m34_9+m35_9+m36_9+m37_9+m38_9+m39_9+m40_9+m41_9+m42_9+m43_9+m44_9+m45_9+m46_9+m47_9+m48_9+m49_9+m50_9+m51_9+m52_9+m53_9+m54_9+m55_9+m56_9+m57_9+m58_9+m59_9+m60_9+m61_9+m62_9+m63_9+m64_9+m65_9+m66_9+m67_9+m68_9+m69_9+m70_9+m71_9+m72_9+m73_9+m74_9+m75_9+m76_9+m77_9+m78_9+m79_9+m80_9+m81_9+m82_9+m83_9+m84_9+m85_9+m86_9+m87_9+m88_9+m89_9+m90_9+m91_9+m92_9+m93_9+m94_9+m95_9+m96_9+m97_9+m98_9+m99_9+m100_9+m101_9+m102_9+m103_9+m104_9+m105_9+m106_9+m107_9+m108_9+m109_9+m110_9+m111_9+m112_9+m113_9+m114_9+m115_9+m116_9+m117_9+m118_9+m119_9+m120_9+m121_9+m122_9+m123_9+m124_9+m125_9+m126_9+m127_9+m128_9+m129_9+m130_9+m131_9+m132_9+m133_9+m134_9+m135_9+m136_9+m137_9+m138_9+m139_9+m140_9+m141_9+m142_9+m143_9+m144_9+m145_9+m146_9+m147_9+m148_9+m149_9+m150_9+m151_9+m152_9+m153_9+m154_9+m155_9+m156_9+m157_9+m158_9+m159_9+m160_9+m161_9+m162_9+m163_9+m164_9+m165_9+m166_9+m167_9+m168_9+m169_9+m170_9+m171_9+m172_9+m173_9+m174_9+m175_9+m176_9+m177_9+m178_9+m179_9+m180_9+m181_9+m182_9+m183_9+m184_9+m185_9+m186_9+m187_9+m188_9+m189_9+m190_9+m191_9+m192_9+m193_9+m194_9+m195_9+m196_9+m197_9+m198_9+m199_9+m200_9+m201_9+m202_9+m203_9+m204_9+m205_9+m206_9+m207_9+m208_9+m209_9+m210_9+m211_9+m212_9+m213_9+m214_9+m215_9+m216_9+m217_9+m218_9+m219_9+m220_9+m221_9+m222_9+m223_9+m224_9+m225_9+m226_9+m227_9+m228_9+m229_9+m230_9+m231_9+m232_9+m233_9+m234_9+m235_9+m236_9+m237_9+m238_9+m239_9+m240_9+m241_9+m242_9+m243_9+m244_9+m245_9+m246_9+m247_9+m248_9+m249_9+m250_9+m251_9+m252_9+m253_9+m254_9+m255_9+m256_9+m257_9+m258_9+m259_9+m260_9+m261_9+m262_9+m263_9+m264_9+m265_9+m266_9+m267_9+m268_9+m269_9+m270_9+m271_9+m272_9+m273_9+m274_9+m275_9+m276_9+m277_9+m278_9+m279_9+m280_9+m281_9+m282_9+m283_9+m284_9+m285_9+m286_9+m287_9+m288_9+m289_9+m290_9+m291_9+m292_9+m293_9+m294_9+m295_9+m296_9+m297_9+m298_9+m299_9+m300_9+m301_9+m302_9+m303_9+m304_9+m305_9+m306_9+m307_9+m308_9+m309_9+m310_9+m311_9+m312_9+m313_9+m314_9+m315_9+m316_9+m317_9+m318_9+m319_9+m320_9+m321_9+m322_9+m323_9+m324_9+m325_9+m326_9+m327_9+m328_9+m329_9+m330_9+m331_9+m332_9+m333_9+m334_9+m335_9+m336_9+m337_9+m338_9+m339_9+m340_9+m341_9+m342_9+m343_9+m344_9+m345_9+m346_9+m347_9+m348_9+m349_9+m350_9+m351_9+m352_9+m353_9+m354_9+m355_9+m356_9+m357_9+m358_9+m359_9+m360_9+m361_9+m362_9+m363_9+m364_9+m365_9+m366_9+m367_9+m368_9+m369_9+m370_9+m371_9+m372_9+m373_9+m374_9+m375_9+m376_9+m377_9+m378_9+m379_9+m380_9+m381_9+b9;
   always @(posedge clk) out10 <= m1_10+m2_10+m3_10+m4_10+m5_10+m6_10+m7_10+m8_10+m9_10+m10_10+m11_10+m12_10+m13_10+m14_10+m15_10+m16_10+m17_10+m18_10+m19_10+m20_10+m21_10+m22_10+m23_10+m24_10+m25_10+m26_10+m27_10+m28_10+m29_10+m30_10+m31_10+m32_10+m33_10+m34_10+m35_10+m36_10+m37_10+m38_10+m39_10+m40_10+m41_10+m42_10+m43_10+m44_10+m45_10+m46_10+m47_10+m48_10+m49_10+m50_10+m51_10+m52_10+m53_10+m54_10+m55_10+m56_10+m57_10+m58_10+m59_10+m60_10+m61_10+m62_10+m63_10+m64_10+m65_10+m66_10+m67_10+m68_10+m69_10+m70_10+m71_10+m72_10+m73_10+m74_10+m75_10+m76_10+m77_10+m78_10+m79_10+m80_10+m81_10+m82_10+m83_10+m84_10+m85_10+m86_10+m87_10+m88_10+m89_10+m90_10+m91_10+m92_10+m93_10+m94_10+m95_10+m96_10+m97_10+m98_10+m99_10+m100_10+m101_10+m102_10+m103_10+m104_10+m105_10+m106_10+m107_10+m108_10+m109_10+m110_10+m111_10+m112_10+m113_10+m114_10+m115_10+m116_10+m117_10+m118_10+m119_10+m120_10+m121_10+m122_10+m123_10+m124_10+m125_10+m126_10+m127_10+m128_10+m129_10+m130_10+m131_10+m132_10+m133_10+m134_10+m135_10+m136_10+m137_10+m138_10+m139_10+m140_10+m141_10+m142_10+m143_10+m144_10+m145_10+m146_10+m147_10+m148_10+m149_10+m150_10+m151_10+m152_10+m153_10+m154_10+m155_10+m156_10+m157_10+m158_10+m159_10+m160_10+m161_10+m162_10+m163_10+m164_10+m165_10+m166_10+m167_10+m168_10+m169_10+m170_10+m171_10+m172_10+m173_10+m174_10+m175_10+m176_10+m177_10+m178_10+m179_10+m180_10+m181_10+m182_10+m183_10+m184_10+m185_10+m186_10+m187_10+m188_10+m189_10+m190_10+m191_10+m192_10+m193_10+m194_10+m195_10+m196_10+m197_10+m198_10+m199_10+m200_10+m201_10+m202_10+m203_10+m204_10+m205_10+m206_10+m207_10+m208_10+m209_10+m210_10+m211_10+m212_10+m213_10+m214_10+m215_10+m216_10+m217_10+m218_10+m219_10+m220_10+m221_10+m222_10+m223_10+m224_10+m225_10+m226_10+m227_10+m228_10+m229_10+m230_10+m231_10+m232_10+m233_10+m234_10+m235_10+m236_10+m237_10+m238_10+m239_10+m240_10+m241_10+m242_10+m243_10+m244_10+m245_10+m246_10+m247_10+m248_10+m249_10+m250_10+m251_10+m252_10+m253_10+m254_10+m255_10+m256_10+m257_10+m258_10+m259_10+m260_10+m261_10+m262_10+m263_10+m264_10+m265_10+m266_10+m267_10+m268_10+m269_10+m270_10+m271_10+m272_10+m273_10+m274_10+m275_10+m276_10+m277_10+m278_10+m279_10+m280_10+m281_10+m282_10+m283_10+m284_10+m285_10+m286_10+m287_10+m288_10+m289_10+m290_10+m291_10+m292_10+m293_10+m294_10+m295_10+m296_10+m297_10+m298_10+m299_10+m300_10+m301_10+m302_10+m303_10+m304_10+m305_10+m306_10+m307_10+m308_10+m309_10+m310_10+m311_10+m312_10+m313_10+m314_10+m315_10+m316_10+m317_10+m318_10+m319_10+m320_10+m321_10+m322_10+m323_10+m324_10+m325_10+m326_10+m327_10+m328_10+m329_10+m330_10+m331_10+m332_10+m333_10+m334_10+m335_10+m336_10+m337_10+m338_10+m339_10+m340_10+m341_10+m342_10+m343_10+m344_10+m345_10+m346_10+m347_10+m348_10+m349_10+m350_10+m351_10+m352_10+m353_10+m354_10+m355_10+m356_10+m357_10+m358_10+m359_10+m360_10+m361_10+m362_10+m363_10+m364_10+m365_10+m366_10+m367_10+m368_10+m369_10+m370_10+m371_10+m372_10+m373_10+m374_10+m375_10+m376_10+m377_10+m378_10+m379_10+m380_10+m381_10+b10;
   always @(posedge clk) out11 <= m1_11+m2_11+m3_11+m4_11+m5_11+m6_11+m7_11+m8_11+m9_11+m10_11+m11_11+m12_11+m13_11+m14_11+m15_11+m16_11+m17_11+m18_11+m19_11+m20_11+m21_11+m22_11+m23_11+m24_11+m25_11+m26_11+m27_11+m28_11+m29_11+m30_11+m31_11+m32_11+m33_11+m34_11+m35_11+m36_11+m37_11+m38_11+m39_11+m40_11+m41_11+m42_11+m43_11+m44_11+m45_11+m46_11+m47_11+m48_11+m49_11+m50_11+m51_11+m52_11+m53_11+m54_11+m55_11+m56_11+m57_11+m58_11+m59_11+m60_11+m61_11+m62_11+m63_11+m64_11+m65_11+m66_11+m67_11+m68_11+m69_11+m70_11+m71_11+m72_11+m73_11+m74_11+m75_11+m76_11+m77_11+m78_11+m79_11+m80_11+m81_11+m82_11+m83_11+m84_11+m85_11+m86_11+m87_11+m88_11+m89_11+m90_11+m91_11+m92_11+m93_11+m94_11+m95_11+m96_11+m97_11+m98_11+m99_11+m100_11+m101_11+m102_11+m103_11+m104_11+m105_11+m106_11+m107_11+m108_11+m109_11+m110_11+m111_11+m112_11+m113_11+m114_11+m115_11+m116_11+m117_11+m118_11+m119_11+m120_11+m121_11+m122_11+m123_11+m124_11+m125_11+m126_11+m127_11+m128_11+m129_11+m130_11+m131_11+m132_11+m133_11+m134_11+m135_11+m136_11+m137_11+m138_11+m139_11+m140_11+m141_11+m142_11+m143_11+m144_11+m145_11+m146_11+m147_11+m148_11+m149_11+m150_11+m151_11+m152_11+m153_11+m154_11+m155_11+m156_11+m157_11+m158_11+m159_11+m160_11+m161_11+m162_11+m163_11+m164_11+m165_11+m166_11+m167_11+m168_11+m169_11+m170_11+m171_11+m172_11+m173_11+m174_11+m175_11+m176_11+m177_11+m178_11+m179_11+m180_11+m181_11+m182_11+m183_11+m184_11+m185_11+m186_11+m187_11+m188_11+m189_11+m190_11+m191_11+m192_11+m193_11+m194_11+m195_11+m196_11+m197_11+m198_11+m199_11+m200_11+m201_11+m202_11+m203_11+m204_11+m205_11+m206_11+m207_11+m208_11+m209_11+m210_11+m211_11+m212_11+m213_11+m214_11+m215_11+m216_11+m217_11+m218_11+m219_11+m220_11+m221_11+m222_11+m223_11+m224_11+m225_11+m226_11+m227_11+m228_11+m229_11+m230_11+m231_11+m232_11+m233_11+m234_11+m235_11+m236_11+m237_11+m238_11+m239_11+m240_11+m241_11+m242_11+m243_11+m244_11+m245_11+m246_11+m247_11+m248_11+m249_11+m250_11+m251_11+m252_11+m253_11+m254_11+m255_11+m256_11+m257_11+m258_11+m259_11+m260_11+m261_11+m262_11+m263_11+m264_11+m265_11+m266_11+m267_11+m268_11+m269_11+m270_11+m271_11+m272_11+m273_11+m274_11+m275_11+m276_11+m277_11+m278_11+m279_11+m280_11+m281_11+m282_11+m283_11+m284_11+m285_11+m286_11+m287_11+m288_11+m289_11+m290_11+m291_11+m292_11+m293_11+m294_11+m295_11+m296_11+m297_11+m298_11+m299_11+m300_11+m301_11+m302_11+m303_11+m304_11+m305_11+m306_11+m307_11+m308_11+m309_11+m310_11+m311_11+m312_11+m313_11+m314_11+m315_11+m316_11+m317_11+m318_11+m319_11+m320_11+m321_11+m322_11+m323_11+m324_11+m325_11+m326_11+m327_11+m328_11+m329_11+m330_11+m331_11+m332_11+m333_11+m334_11+m335_11+m336_11+m337_11+m338_11+m339_11+m340_11+m341_11+m342_11+m343_11+m344_11+m345_11+m346_11+m347_11+m348_11+m349_11+m350_11+m351_11+m352_11+m353_11+m354_11+m355_11+m356_11+m357_11+m358_11+m359_11+m360_11+m361_11+m362_11+m363_11+m364_11+m365_11+m366_11+m367_11+m368_11+m369_11+m370_11+m371_11+m372_11+m373_11+m374_11+m375_11+m376_11+m377_11+m378_11+m379_11+m380_11+m381_11+b11;
   always @(posedge clk) out12 <= m1_12+m2_12+m3_12+m4_12+m5_12+m6_12+m7_12+m8_12+m9_12+m10_12+m11_12+m12_12+m13_12+m14_12+m15_12+m16_12+m17_12+m18_12+m19_12+m20_12+m21_12+m22_12+m23_12+m24_12+m25_12+m26_12+m27_12+m28_12+m29_12+m30_12+m31_12+m32_12+m33_12+m34_12+m35_12+m36_12+m37_12+m38_12+m39_12+m40_12+m41_12+m42_12+m43_12+m44_12+m45_12+m46_12+m47_12+m48_12+m49_12+m50_12+m51_12+m52_12+m53_12+m54_12+m55_12+m56_12+m57_12+m58_12+m59_12+m60_12+m61_12+m62_12+m63_12+m64_12+m65_12+m66_12+m67_12+m68_12+m69_12+m70_12+m71_12+m72_12+m73_12+m74_12+m75_12+m76_12+m77_12+m78_12+m79_12+m80_12+m81_12+m82_12+m83_12+m84_12+m85_12+m86_12+m87_12+m88_12+m89_12+m90_12+m91_12+m92_12+m93_12+m94_12+m95_12+m96_12+m97_12+m98_12+m99_12+m100_12+m101_12+m102_12+m103_12+m104_12+m105_12+m106_12+m107_12+m108_12+m109_12+m110_12+m111_12+m112_12+m113_12+m114_12+m115_12+m116_12+m117_12+m118_12+m119_12+m120_12+m121_12+m122_12+m123_12+m124_12+m125_12+m126_12+m127_12+m128_12+m129_12+m130_12+m131_12+m132_12+m133_12+m134_12+m135_12+m136_12+m137_12+m138_12+m139_12+m140_12+m141_12+m142_12+m143_12+m144_12+m145_12+m146_12+m147_12+m148_12+m149_12+m150_12+m151_12+m152_12+m153_12+m154_12+m155_12+m156_12+m157_12+m158_12+m159_12+m160_12+m161_12+m162_12+m163_12+m164_12+m165_12+m166_12+m167_12+m168_12+m169_12+m170_12+m171_12+m172_12+m173_12+m174_12+m175_12+m176_12+m177_12+m178_12+m179_12+m180_12+m181_12+m182_12+m183_12+m184_12+m185_12+m186_12+m187_12+m188_12+m189_12+m190_12+m191_12+m192_12+m193_12+m194_12+m195_12+m196_12+m197_12+m198_12+m199_12+m200_12+m201_12+m202_12+m203_12+m204_12+m205_12+m206_12+m207_12+m208_12+m209_12+m210_12+m211_12+m212_12+m213_12+m214_12+m215_12+m216_12+m217_12+m218_12+m219_12+m220_12+m221_12+m222_12+m223_12+m224_12+m225_12+m226_12+m227_12+m228_12+m229_12+m230_12+m231_12+m232_12+m233_12+m234_12+m235_12+m236_12+m237_12+m238_12+m239_12+m240_12+m241_12+m242_12+m243_12+m244_12+m245_12+m246_12+m247_12+m248_12+m249_12+m250_12+m251_12+m252_12+m253_12+m254_12+m255_12+m256_12+m257_12+m258_12+m259_12+m260_12+m261_12+m262_12+m263_12+m264_12+m265_12+m266_12+m267_12+m268_12+m269_12+m270_12+m271_12+m272_12+m273_12+m274_12+m275_12+m276_12+m277_12+m278_12+m279_12+m280_12+m281_12+m282_12+m283_12+m284_12+m285_12+m286_12+m287_12+m288_12+m289_12+m290_12+m291_12+m292_12+m293_12+m294_12+m295_12+m296_12+m297_12+m298_12+m299_12+m300_12+m301_12+m302_12+m303_12+m304_12+m305_12+m306_12+m307_12+m308_12+m309_12+m310_12+m311_12+m312_12+m313_12+m314_12+m315_12+m316_12+m317_12+m318_12+m319_12+m320_12+m321_12+m322_12+m323_12+m324_12+m325_12+m326_12+m327_12+m328_12+m329_12+m330_12+m331_12+m332_12+m333_12+m334_12+m335_12+m336_12+m337_12+m338_12+m339_12+m340_12+m341_12+m342_12+m343_12+m344_12+m345_12+m346_12+m347_12+m348_12+m349_12+m350_12+m351_12+m352_12+m353_12+m354_12+m355_12+m356_12+m357_12+m358_12+m359_12+m360_12+m361_12+m362_12+m363_12+m364_12+m365_12+m366_12+m367_12+m368_12+m369_12+m370_12+m371_12+m372_12+m373_12+m374_12+m375_12+m376_12+m377_12+m378_12+m379_12+m380_12+m381_12+b12;
   always @(posedge clk) out13 <= m1_13+m2_13+m3_13+m4_13+m5_13+m6_13+m7_13+m8_13+m9_13+m10_13+m11_13+m12_13+m13_13+m14_13+m15_13+m16_13+m17_13+m18_13+m19_13+m20_13+m21_13+m22_13+m23_13+m24_13+m25_13+m26_13+m27_13+m28_13+m29_13+m30_13+m31_13+m32_13+m33_13+m34_13+m35_13+m36_13+m37_13+m38_13+m39_13+m40_13+m41_13+m42_13+m43_13+m44_13+m45_13+m46_13+m47_13+m48_13+m49_13+m50_13+m51_13+m52_13+m53_13+m54_13+m55_13+m56_13+m57_13+m58_13+m59_13+m60_13+m61_13+m62_13+m63_13+m64_13+m65_13+m66_13+m67_13+m68_13+m69_13+m70_13+m71_13+m72_13+m73_13+m74_13+m75_13+m76_13+m77_13+m78_13+m79_13+m80_13+m81_13+m82_13+m83_13+m84_13+m85_13+m86_13+m87_13+m88_13+m89_13+m90_13+m91_13+m92_13+m93_13+m94_13+m95_13+m96_13+m97_13+m98_13+m99_13+m100_13+m101_13+m102_13+m103_13+m104_13+m105_13+m106_13+m107_13+m108_13+m109_13+m110_13+m111_13+m112_13+m113_13+m114_13+m115_13+m116_13+m117_13+m118_13+m119_13+m120_13+m121_13+m122_13+m123_13+m124_13+m125_13+m126_13+m127_13+m128_13+m129_13+m130_13+m131_13+m132_13+m133_13+m134_13+m135_13+m136_13+m137_13+m138_13+m139_13+m140_13+m141_13+m142_13+m143_13+m144_13+m145_13+m146_13+m147_13+m148_13+m149_13+m150_13+m151_13+m152_13+m153_13+m154_13+m155_13+m156_13+m157_13+m158_13+m159_13+m160_13+m161_13+m162_13+m163_13+m164_13+m165_13+m166_13+m167_13+m168_13+m169_13+m170_13+m171_13+m172_13+m173_13+m174_13+m175_13+m176_13+m177_13+m178_13+m179_13+m180_13+m181_13+m182_13+m183_13+m184_13+m185_13+m186_13+m187_13+m188_13+m189_13+m190_13+m191_13+m192_13+m193_13+m194_13+m195_13+m196_13+m197_13+m198_13+m199_13+m200_13+m201_13+m202_13+m203_13+m204_13+m205_13+m206_13+m207_13+m208_13+m209_13+m210_13+m211_13+m212_13+m213_13+m214_13+m215_13+m216_13+m217_13+m218_13+m219_13+m220_13+m221_13+m222_13+m223_13+m224_13+m225_13+m226_13+m227_13+m228_13+m229_13+m230_13+m231_13+m232_13+m233_13+m234_13+m235_13+m236_13+m237_13+m238_13+m239_13+m240_13+m241_13+m242_13+m243_13+m244_13+m245_13+m246_13+m247_13+m248_13+m249_13+m250_13+m251_13+m252_13+m253_13+m254_13+m255_13+m256_13+m257_13+m258_13+m259_13+m260_13+m261_13+m262_13+m263_13+m264_13+m265_13+m266_13+m267_13+m268_13+m269_13+m270_13+m271_13+m272_13+m273_13+m274_13+m275_13+m276_13+m277_13+m278_13+m279_13+m280_13+m281_13+m282_13+m283_13+m284_13+m285_13+m286_13+m287_13+m288_13+m289_13+m290_13+m291_13+m292_13+m293_13+m294_13+m295_13+m296_13+m297_13+m298_13+m299_13+m300_13+m301_13+m302_13+m303_13+m304_13+m305_13+m306_13+m307_13+m308_13+m309_13+m310_13+m311_13+m312_13+m313_13+m314_13+m315_13+m316_13+m317_13+m318_13+m319_13+m320_13+m321_13+m322_13+m323_13+m324_13+m325_13+m326_13+m327_13+m328_13+m329_13+m330_13+m331_13+m332_13+m333_13+m334_13+m335_13+m336_13+m337_13+m338_13+m339_13+m340_13+m341_13+m342_13+m343_13+m344_13+m345_13+m346_13+m347_13+m348_13+m349_13+m350_13+m351_13+m352_13+m353_13+m354_13+m355_13+m356_13+m357_13+m358_13+m359_13+m360_13+m361_13+m362_13+m363_13+m364_13+m365_13+m366_13+m367_13+m368_13+m369_13+m370_13+m371_13+m372_13+m373_13+m374_13+m375_13+m376_13+m377_13+m378_13+m379_13+m380_13+m381_13+b13;
   always @(posedge clk) out14 <= m1_14+m2_14+m3_14+m4_14+m5_14+m6_14+m7_14+m8_14+m9_14+m10_14+m11_14+m12_14+m13_14+m14_14+m15_14+m16_14+m17_14+m18_14+m19_14+m20_14+m21_14+m22_14+m23_14+m24_14+m25_14+m26_14+m27_14+m28_14+m29_14+m30_14+m31_14+m32_14+m33_14+m34_14+m35_14+m36_14+m37_14+m38_14+m39_14+m40_14+m41_14+m42_14+m43_14+m44_14+m45_14+m46_14+m47_14+m48_14+m49_14+m50_14+m51_14+m52_14+m53_14+m54_14+m55_14+m56_14+m57_14+m58_14+m59_14+m60_14+m61_14+m62_14+m63_14+m64_14+m65_14+m66_14+m67_14+m68_14+m69_14+m70_14+m71_14+m72_14+m73_14+m74_14+m75_14+m76_14+m77_14+m78_14+m79_14+m80_14+m81_14+m82_14+m83_14+m84_14+m85_14+m86_14+m87_14+m88_14+m89_14+m90_14+m91_14+m92_14+m93_14+m94_14+m95_14+m96_14+m97_14+m98_14+m99_14+m100_14+m101_14+m102_14+m103_14+m104_14+m105_14+m106_14+m107_14+m108_14+m109_14+m110_14+m111_14+m112_14+m113_14+m114_14+m115_14+m116_14+m117_14+m118_14+m119_14+m120_14+m121_14+m122_14+m123_14+m124_14+m125_14+m126_14+m127_14+m128_14+m129_14+m130_14+m131_14+m132_14+m133_14+m134_14+m135_14+m136_14+m137_14+m138_14+m139_14+m140_14+m141_14+m142_14+m143_14+m144_14+m145_14+m146_14+m147_14+m148_14+m149_14+m150_14+m151_14+m152_14+m153_14+m154_14+m155_14+m156_14+m157_14+m158_14+m159_14+m160_14+m161_14+m162_14+m163_14+m164_14+m165_14+m166_14+m167_14+m168_14+m169_14+m170_14+m171_14+m172_14+m173_14+m174_14+m175_14+m176_14+m177_14+m178_14+m179_14+m180_14+m181_14+m182_14+m183_14+m184_14+m185_14+m186_14+m187_14+m188_14+m189_14+m190_14+m191_14+m192_14+m193_14+m194_14+m195_14+m196_14+m197_14+m198_14+m199_14+m200_14+m201_14+m202_14+m203_14+m204_14+m205_14+m206_14+m207_14+m208_14+m209_14+m210_14+m211_14+m212_14+m213_14+m214_14+m215_14+m216_14+m217_14+m218_14+m219_14+m220_14+m221_14+m222_14+m223_14+m224_14+m225_14+m226_14+m227_14+m228_14+m229_14+m230_14+m231_14+m232_14+m233_14+m234_14+m235_14+m236_14+m237_14+m238_14+m239_14+m240_14+m241_14+m242_14+m243_14+m244_14+m245_14+m246_14+m247_14+m248_14+m249_14+m250_14+m251_14+m252_14+m253_14+m254_14+m255_14+m256_14+m257_14+m258_14+m259_14+m260_14+m261_14+m262_14+m263_14+m264_14+m265_14+m266_14+m267_14+m268_14+m269_14+m270_14+m271_14+m272_14+m273_14+m274_14+m275_14+m276_14+m277_14+m278_14+m279_14+m280_14+m281_14+m282_14+m283_14+m284_14+m285_14+m286_14+m287_14+m288_14+m289_14+m290_14+m291_14+m292_14+m293_14+m294_14+m295_14+m296_14+m297_14+m298_14+m299_14+m300_14+m301_14+m302_14+m303_14+m304_14+m305_14+m306_14+m307_14+m308_14+m309_14+m310_14+m311_14+m312_14+m313_14+m314_14+m315_14+m316_14+m317_14+m318_14+m319_14+m320_14+m321_14+m322_14+m323_14+m324_14+m325_14+m326_14+m327_14+m328_14+m329_14+m330_14+m331_14+m332_14+m333_14+m334_14+m335_14+m336_14+m337_14+m338_14+m339_14+m340_14+m341_14+m342_14+m343_14+m344_14+m345_14+m346_14+m347_14+m348_14+m349_14+m350_14+m351_14+m352_14+m353_14+m354_14+m355_14+m356_14+m357_14+m358_14+m359_14+m360_14+m361_14+m362_14+m363_14+m364_14+m365_14+m366_14+m367_14+m368_14+m369_14+m370_14+m371_14+m372_14+m373_14+m374_14+m375_14+m376_14+m377_14+m378_14+m379_14+m380_14+m381_14+b14;
   always @(posedge clk) out15 <= m1_15+m2_15+m3_15+m4_15+m5_15+m6_15+m7_15+m8_15+m9_15+m10_15+m11_15+m12_15+m13_15+m14_15+m15_15+m16_15+m17_15+m18_15+m19_15+m20_15+m21_15+m22_15+m23_15+m24_15+m25_15+m26_15+m27_15+m28_15+m29_15+m30_15+m31_15+m32_15+m33_15+m34_15+m35_15+m36_15+m37_15+m38_15+m39_15+m40_15+m41_15+m42_15+m43_15+m44_15+m45_15+m46_15+m47_15+m48_15+m49_15+m50_15+m51_15+m52_15+m53_15+m54_15+m55_15+m56_15+m57_15+m58_15+m59_15+m60_15+m61_15+m62_15+m63_15+m64_15+m65_15+m66_15+m67_15+m68_15+m69_15+m70_15+m71_15+m72_15+m73_15+m74_15+m75_15+m76_15+m77_15+m78_15+m79_15+m80_15+m81_15+m82_15+m83_15+m84_15+m85_15+m86_15+m87_15+m88_15+m89_15+m90_15+m91_15+m92_15+m93_15+m94_15+m95_15+m96_15+m97_15+m98_15+m99_15+m100_15+m101_15+m102_15+m103_15+m104_15+m105_15+m106_15+m107_15+m108_15+m109_15+m110_15+m111_15+m112_15+m113_15+m114_15+m115_15+m116_15+m117_15+m118_15+m119_15+m120_15+m121_15+m122_15+m123_15+m124_15+m125_15+m126_15+m127_15+m128_15+m129_15+m130_15+m131_15+m132_15+m133_15+m134_15+m135_15+m136_15+m137_15+m138_15+m139_15+m140_15+m141_15+m142_15+m143_15+m144_15+m145_15+m146_15+m147_15+m148_15+m149_15+m150_15+m151_15+m152_15+m153_15+m154_15+m155_15+m156_15+m157_15+m158_15+m159_15+m160_15+m161_15+m162_15+m163_15+m164_15+m165_15+m166_15+m167_15+m168_15+m169_15+m170_15+m171_15+m172_15+m173_15+m174_15+m175_15+m176_15+m177_15+m178_15+m179_15+m180_15+m181_15+m182_15+m183_15+m184_15+m185_15+m186_15+m187_15+m188_15+m189_15+m190_15+m191_15+m192_15+m193_15+m194_15+m195_15+m196_15+m197_15+m198_15+m199_15+m200_15+m201_15+m202_15+m203_15+m204_15+m205_15+m206_15+m207_15+m208_15+m209_15+m210_15+m211_15+m212_15+m213_15+m214_15+m215_15+m216_15+m217_15+m218_15+m219_15+m220_15+m221_15+m222_15+m223_15+m224_15+m225_15+m226_15+m227_15+m228_15+m229_15+m230_15+m231_15+m232_15+m233_15+m234_15+m235_15+m236_15+m237_15+m238_15+m239_15+m240_15+m241_15+m242_15+m243_15+m244_15+m245_15+m246_15+m247_15+m248_15+m249_15+m250_15+m251_15+m252_15+m253_15+m254_15+m255_15+m256_15+m257_15+m258_15+m259_15+m260_15+m261_15+m262_15+m263_15+m264_15+m265_15+m266_15+m267_15+m268_15+m269_15+m270_15+m271_15+m272_15+m273_15+m274_15+m275_15+m276_15+m277_15+m278_15+m279_15+m280_15+m281_15+m282_15+m283_15+m284_15+m285_15+m286_15+m287_15+m288_15+m289_15+m290_15+m291_15+m292_15+m293_15+m294_15+m295_15+m296_15+m297_15+m298_15+m299_15+m300_15+m301_15+m302_15+m303_15+m304_15+m305_15+m306_15+m307_15+m308_15+m309_15+m310_15+m311_15+m312_15+m313_15+m314_15+m315_15+m316_15+m317_15+m318_15+m319_15+m320_15+m321_15+m322_15+m323_15+m324_15+m325_15+m326_15+m327_15+m328_15+m329_15+m330_15+m331_15+m332_15+m333_15+m334_15+m335_15+m336_15+m337_15+m338_15+m339_15+m340_15+m341_15+m342_15+m343_15+m344_15+m345_15+m346_15+m347_15+m348_15+m349_15+m350_15+m351_15+m352_15+m353_15+m354_15+m355_15+m356_15+m357_15+m358_15+m359_15+m360_15+m361_15+m362_15+m363_15+m364_15+m365_15+m366_15+m367_15+m368_15+m369_15+m370_15+m371_15+m372_15+m373_15+m374_15+m375_15+m376_15+m377_15+m378_15+m379_15+m380_15+m381_15+b15;
   always @(posedge clk) out16 <= m1_16+m2_16+m3_16+m4_16+m5_16+m6_16+m7_16+m8_16+m9_16+m10_16+m11_16+m12_16+m13_16+m14_16+m15_16+m16_16+m17_16+m18_16+m19_16+m20_16+m21_16+m22_16+m23_16+m24_16+m25_16+m26_16+m27_16+m28_16+m29_16+m30_16+m31_16+m32_16+m33_16+m34_16+m35_16+m36_16+m37_16+m38_16+m39_16+m40_16+m41_16+m42_16+m43_16+m44_16+m45_16+m46_16+m47_16+m48_16+m49_16+m50_16+m51_16+m52_16+m53_16+m54_16+m55_16+m56_16+m57_16+m58_16+m59_16+m60_16+m61_16+m62_16+m63_16+m64_16+m65_16+m66_16+m67_16+m68_16+m69_16+m70_16+m71_16+m72_16+m73_16+m74_16+m75_16+m76_16+m77_16+m78_16+m79_16+m80_16+m81_16+m82_16+m83_16+m84_16+m85_16+m86_16+m87_16+m88_16+m89_16+m90_16+m91_16+m92_16+m93_16+m94_16+m95_16+m96_16+m97_16+m98_16+m99_16+m100_16+m101_16+m102_16+m103_16+m104_16+m105_16+m106_16+m107_16+m108_16+m109_16+m110_16+m111_16+m112_16+m113_16+m114_16+m115_16+m116_16+m117_16+m118_16+m119_16+m120_16+m121_16+m122_16+m123_16+m124_16+m125_16+m126_16+m127_16+m128_16+m129_16+m130_16+m131_16+m132_16+m133_16+m134_16+m135_16+m136_16+m137_16+m138_16+m139_16+m140_16+m141_16+m142_16+m143_16+m144_16+m145_16+m146_16+m147_16+m148_16+m149_16+m150_16+m151_16+m152_16+m153_16+m154_16+m155_16+m156_16+m157_16+m158_16+m159_16+m160_16+m161_16+m162_16+m163_16+m164_16+m165_16+m166_16+m167_16+m168_16+m169_16+m170_16+m171_16+m172_16+m173_16+m174_16+m175_16+m176_16+m177_16+m178_16+m179_16+m180_16+m181_16+m182_16+m183_16+m184_16+m185_16+m186_16+m187_16+m188_16+m189_16+m190_16+m191_16+m192_16+m193_16+m194_16+m195_16+m196_16+m197_16+m198_16+m199_16+m200_16+m201_16+m202_16+m203_16+m204_16+m205_16+m206_16+m207_16+m208_16+m209_16+m210_16+m211_16+m212_16+m213_16+m214_16+m215_16+m216_16+m217_16+m218_16+m219_16+m220_16+m221_16+m222_16+m223_16+m224_16+m225_16+m226_16+m227_16+m228_16+m229_16+m230_16+m231_16+m232_16+m233_16+m234_16+m235_16+m236_16+m237_16+m238_16+m239_16+m240_16+m241_16+m242_16+m243_16+m244_16+m245_16+m246_16+m247_16+m248_16+m249_16+m250_16+m251_16+m252_16+m253_16+m254_16+m255_16+m256_16+m257_16+m258_16+m259_16+m260_16+m261_16+m262_16+m263_16+m264_16+m265_16+m266_16+m267_16+m268_16+m269_16+m270_16+m271_16+m272_16+m273_16+m274_16+m275_16+m276_16+m277_16+m278_16+m279_16+m280_16+m281_16+m282_16+m283_16+m284_16+m285_16+m286_16+m287_16+m288_16+m289_16+m290_16+m291_16+m292_16+m293_16+m294_16+m295_16+m296_16+m297_16+m298_16+m299_16+m300_16+m301_16+m302_16+m303_16+m304_16+m305_16+m306_16+m307_16+m308_16+m309_16+m310_16+m311_16+m312_16+m313_16+m314_16+m315_16+m316_16+m317_16+m318_16+m319_16+m320_16+m321_16+m322_16+m323_16+m324_16+m325_16+m326_16+m327_16+m328_16+m329_16+m330_16+m331_16+m332_16+m333_16+m334_16+m335_16+m336_16+m337_16+m338_16+m339_16+m340_16+m341_16+m342_16+m343_16+m344_16+m345_16+m346_16+m347_16+m348_16+m349_16+m350_16+m351_16+m352_16+m353_16+m354_16+m355_16+m356_16+m357_16+m358_16+m359_16+m360_16+m361_16+m362_16+m363_16+m364_16+m365_16+m366_16+m367_16+m368_16+m369_16+m370_16+m371_16+m372_16+m373_16+m374_16+m375_16+m376_16+m377_16+m378_16+m379_16+m380_16+m381_16+b16;
   always @(posedge clk) out17 <= m1_17+m2_17+m3_17+m4_17+m5_17+m6_17+m7_17+m8_17+m9_17+m10_17+m11_17+m12_17+m13_17+m14_17+m15_17+m16_17+m17_17+m18_17+m19_17+m20_17+m21_17+m22_17+m23_17+m24_17+m25_17+m26_17+m27_17+m28_17+m29_17+m30_17+m31_17+m32_17+m33_17+m34_17+m35_17+m36_17+m37_17+m38_17+m39_17+m40_17+m41_17+m42_17+m43_17+m44_17+m45_17+m46_17+m47_17+m48_17+m49_17+m50_17+m51_17+m52_17+m53_17+m54_17+m55_17+m56_17+m57_17+m58_17+m59_17+m60_17+m61_17+m62_17+m63_17+m64_17+m65_17+m66_17+m67_17+m68_17+m69_17+m70_17+m71_17+m72_17+m73_17+m74_17+m75_17+m76_17+m77_17+m78_17+m79_17+m80_17+m81_17+m82_17+m83_17+m84_17+m85_17+m86_17+m87_17+m88_17+m89_17+m90_17+m91_17+m92_17+m93_17+m94_17+m95_17+m96_17+m97_17+m98_17+m99_17+m100_17+m101_17+m102_17+m103_17+m104_17+m105_17+m106_17+m107_17+m108_17+m109_17+m110_17+m111_17+m112_17+m113_17+m114_17+m115_17+m116_17+m117_17+m118_17+m119_17+m120_17+m121_17+m122_17+m123_17+m124_17+m125_17+m126_17+m127_17+m128_17+m129_17+m130_17+m131_17+m132_17+m133_17+m134_17+m135_17+m136_17+m137_17+m138_17+m139_17+m140_17+m141_17+m142_17+m143_17+m144_17+m145_17+m146_17+m147_17+m148_17+m149_17+m150_17+m151_17+m152_17+m153_17+m154_17+m155_17+m156_17+m157_17+m158_17+m159_17+m160_17+m161_17+m162_17+m163_17+m164_17+m165_17+m166_17+m167_17+m168_17+m169_17+m170_17+m171_17+m172_17+m173_17+m174_17+m175_17+m176_17+m177_17+m178_17+m179_17+m180_17+m181_17+m182_17+m183_17+m184_17+m185_17+m186_17+m187_17+m188_17+m189_17+m190_17+m191_17+m192_17+m193_17+m194_17+m195_17+m196_17+m197_17+m198_17+m199_17+m200_17+m201_17+m202_17+m203_17+m204_17+m205_17+m206_17+m207_17+m208_17+m209_17+m210_17+m211_17+m212_17+m213_17+m214_17+m215_17+m216_17+m217_17+m218_17+m219_17+m220_17+m221_17+m222_17+m223_17+m224_17+m225_17+m226_17+m227_17+m228_17+m229_17+m230_17+m231_17+m232_17+m233_17+m234_17+m235_17+m236_17+m237_17+m238_17+m239_17+m240_17+m241_17+m242_17+m243_17+m244_17+m245_17+m246_17+m247_17+m248_17+m249_17+m250_17+m251_17+m252_17+m253_17+m254_17+m255_17+m256_17+m257_17+m258_17+m259_17+m260_17+m261_17+m262_17+m263_17+m264_17+m265_17+m266_17+m267_17+m268_17+m269_17+m270_17+m271_17+m272_17+m273_17+m274_17+m275_17+m276_17+m277_17+m278_17+m279_17+m280_17+m281_17+m282_17+m283_17+m284_17+m285_17+m286_17+m287_17+m288_17+m289_17+m290_17+m291_17+m292_17+m293_17+m294_17+m295_17+m296_17+m297_17+m298_17+m299_17+m300_17+m301_17+m302_17+m303_17+m304_17+m305_17+m306_17+m307_17+m308_17+m309_17+m310_17+m311_17+m312_17+m313_17+m314_17+m315_17+m316_17+m317_17+m318_17+m319_17+m320_17+m321_17+m322_17+m323_17+m324_17+m325_17+m326_17+m327_17+m328_17+m329_17+m330_17+m331_17+m332_17+m333_17+m334_17+m335_17+m336_17+m337_17+m338_17+m339_17+m340_17+m341_17+m342_17+m343_17+m344_17+m345_17+m346_17+m347_17+m348_17+m349_17+m350_17+m351_17+m352_17+m353_17+m354_17+m355_17+m356_17+m357_17+m358_17+m359_17+m360_17+m361_17+m362_17+m363_17+m364_17+m365_17+m366_17+m367_17+m368_17+m369_17+m370_17+m371_17+m372_17+m373_17+m374_17+m375_17+m376_17+m377_17+m378_17+m379_17+m380_17+m381_17+b17;
   always @(posedge clk) out18 <= m1_18+m2_18+m3_18+m4_18+m5_18+m6_18+m7_18+m8_18+m9_18+m10_18+m11_18+m12_18+m13_18+m14_18+m15_18+m16_18+m17_18+m18_18+m19_18+m20_18+m21_18+m22_18+m23_18+m24_18+m25_18+m26_18+m27_18+m28_18+m29_18+m30_18+m31_18+m32_18+m33_18+m34_18+m35_18+m36_18+m37_18+m38_18+m39_18+m40_18+m41_18+m42_18+m43_18+m44_18+m45_18+m46_18+m47_18+m48_18+m49_18+m50_18+m51_18+m52_18+m53_18+m54_18+m55_18+m56_18+m57_18+m58_18+m59_18+m60_18+m61_18+m62_18+m63_18+m64_18+m65_18+m66_18+m67_18+m68_18+m69_18+m70_18+m71_18+m72_18+m73_18+m74_18+m75_18+m76_18+m77_18+m78_18+m79_18+m80_18+m81_18+m82_18+m83_18+m84_18+m85_18+m86_18+m87_18+m88_18+m89_18+m90_18+m91_18+m92_18+m93_18+m94_18+m95_18+m96_18+m97_18+m98_18+m99_18+m100_18+m101_18+m102_18+m103_18+m104_18+m105_18+m106_18+m107_18+m108_18+m109_18+m110_18+m111_18+m112_18+m113_18+m114_18+m115_18+m116_18+m117_18+m118_18+m119_18+m120_18+m121_18+m122_18+m123_18+m124_18+m125_18+m126_18+m127_18+m128_18+m129_18+m130_18+m131_18+m132_18+m133_18+m134_18+m135_18+m136_18+m137_18+m138_18+m139_18+m140_18+m141_18+m142_18+m143_18+m144_18+m145_18+m146_18+m147_18+m148_18+m149_18+m150_18+m151_18+m152_18+m153_18+m154_18+m155_18+m156_18+m157_18+m158_18+m159_18+m160_18+m161_18+m162_18+m163_18+m164_18+m165_18+m166_18+m167_18+m168_18+m169_18+m170_18+m171_18+m172_18+m173_18+m174_18+m175_18+m176_18+m177_18+m178_18+m179_18+m180_18+m181_18+m182_18+m183_18+m184_18+m185_18+m186_18+m187_18+m188_18+m189_18+m190_18+m191_18+m192_18+m193_18+m194_18+m195_18+m196_18+m197_18+m198_18+m199_18+m200_18+m201_18+m202_18+m203_18+m204_18+m205_18+m206_18+m207_18+m208_18+m209_18+m210_18+m211_18+m212_18+m213_18+m214_18+m215_18+m216_18+m217_18+m218_18+m219_18+m220_18+m221_18+m222_18+m223_18+m224_18+m225_18+m226_18+m227_18+m228_18+m229_18+m230_18+m231_18+m232_18+m233_18+m234_18+m235_18+m236_18+m237_18+m238_18+m239_18+m240_18+m241_18+m242_18+m243_18+m244_18+m245_18+m246_18+m247_18+m248_18+m249_18+m250_18+m251_18+m252_18+m253_18+m254_18+m255_18+m256_18+m257_18+m258_18+m259_18+m260_18+m261_18+m262_18+m263_18+m264_18+m265_18+m266_18+m267_18+m268_18+m269_18+m270_18+m271_18+m272_18+m273_18+m274_18+m275_18+m276_18+m277_18+m278_18+m279_18+m280_18+m281_18+m282_18+m283_18+m284_18+m285_18+m286_18+m287_18+m288_18+m289_18+m290_18+m291_18+m292_18+m293_18+m294_18+m295_18+m296_18+m297_18+m298_18+m299_18+m300_18+m301_18+m302_18+m303_18+m304_18+m305_18+m306_18+m307_18+m308_18+m309_18+m310_18+m311_18+m312_18+m313_18+m314_18+m315_18+m316_18+m317_18+m318_18+m319_18+m320_18+m321_18+m322_18+m323_18+m324_18+m325_18+m326_18+m327_18+m328_18+m329_18+m330_18+m331_18+m332_18+m333_18+m334_18+m335_18+m336_18+m337_18+m338_18+m339_18+m340_18+m341_18+m342_18+m343_18+m344_18+m345_18+m346_18+m347_18+m348_18+m349_18+m350_18+m351_18+m352_18+m353_18+m354_18+m355_18+m356_18+m357_18+m358_18+m359_18+m360_18+m361_18+m362_18+m363_18+m364_18+m365_18+m366_18+m367_18+m368_18+m369_18+m370_18+m371_18+m372_18+m373_18+m374_18+m375_18+m376_18+m377_18+m378_18+m379_18+m380_18+m381_18+b18;
   always @(posedge clk) out19 <= m1_19+m2_19+m3_19+m4_19+m5_19+m6_19+m7_19+m8_19+m9_19+m10_19+m11_19+m12_19+m13_19+m14_19+m15_19+m16_19+m17_19+m18_19+m19_19+m20_19+m21_19+m22_19+m23_19+m24_19+m25_19+m26_19+m27_19+m28_19+m29_19+m30_19+m31_19+m32_19+m33_19+m34_19+m35_19+m36_19+m37_19+m38_19+m39_19+m40_19+m41_19+m42_19+m43_19+m44_19+m45_19+m46_19+m47_19+m48_19+m49_19+m50_19+m51_19+m52_19+m53_19+m54_19+m55_19+m56_19+m57_19+m58_19+m59_19+m60_19+m61_19+m62_19+m63_19+m64_19+m65_19+m66_19+m67_19+m68_19+m69_19+m70_19+m71_19+m72_19+m73_19+m74_19+m75_19+m76_19+m77_19+m78_19+m79_19+m80_19+m81_19+m82_19+m83_19+m84_19+m85_19+m86_19+m87_19+m88_19+m89_19+m90_19+m91_19+m92_19+m93_19+m94_19+m95_19+m96_19+m97_19+m98_19+m99_19+m100_19+m101_19+m102_19+m103_19+m104_19+m105_19+m106_19+m107_19+m108_19+m109_19+m110_19+m111_19+m112_19+m113_19+m114_19+m115_19+m116_19+m117_19+m118_19+m119_19+m120_19+m121_19+m122_19+m123_19+m124_19+m125_19+m126_19+m127_19+m128_19+m129_19+m130_19+m131_19+m132_19+m133_19+m134_19+m135_19+m136_19+m137_19+m138_19+m139_19+m140_19+m141_19+m142_19+m143_19+m144_19+m145_19+m146_19+m147_19+m148_19+m149_19+m150_19+m151_19+m152_19+m153_19+m154_19+m155_19+m156_19+m157_19+m158_19+m159_19+m160_19+m161_19+m162_19+m163_19+m164_19+m165_19+m166_19+m167_19+m168_19+m169_19+m170_19+m171_19+m172_19+m173_19+m174_19+m175_19+m176_19+m177_19+m178_19+m179_19+m180_19+m181_19+m182_19+m183_19+m184_19+m185_19+m186_19+m187_19+m188_19+m189_19+m190_19+m191_19+m192_19+m193_19+m194_19+m195_19+m196_19+m197_19+m198_19+m199_19+m200_19+m201_19+m202_19+m203_19+m204_19+m205_19+m206_19+m207_19+m208_19+m209_19+m210_19+m211_19+m212_19+m213_19+m214_19+m215_19+m216_19+m217_19+m218_19+m219_19+m220_19+m221_19+m222_19+m223_19+m224_19+m225_19+m226_19+m227_19+m228_19+m229_19+m230_19+m231_19+m232_19+m233_19+m234_19+m235_19+m236_19+m237_19+m238_19+m239_19+m240_19+m241_19+m242_19+m243_19+m244_19+m245_19+m246_19+m247_19+m248_19+m249_19+m250_19+m251_19+m252_19+m253_19+m254_19+m255_19+m256_19+m257_19+m258_19+m259_19+m260_19+m261_19+m262_19+m263_19+m264_19+m265_19+m266_19+m267_19+m268_19+m269_19+m270_19+m271_19+m272_19+m273_19+m274_19+m275_19+m276_19+m277_19+m278_19+m279_19+m280_19+m281_19+m282_19+m283_19+m284_19+m285_19+m286_19+m287_19+m288_19+m289_19+m290_19+m291_19+m292_19+m293_19+m294_19+m295_19+m296_19+m297_19+m298_19+m299_19+m300_19+m301_19+m302_19+m303_19+m304_19+m305_19+m306_19+m307_19+m308_19+m309_19+m310_19+m311_19+m312_19+m313_19+m314_19+m315_19+m316_19+m317_19+m318_19+m319_19+m320_19+m321_19+m322_19+m323_19+m324_19+m325_19+m326_19+m327_19+m328_19+m329_19+m330_19+m331_19+m332_19+m333_19+m334_19+m335_19+m336_19+m337_19+m338_19+m339_19+m340_19+m341_19+m342_19+m343_19+m344_19+m345_19+m346_19+m347_19+m348_19+m349_19+m350_19+m351_19+m352_19+m353_19+m354_19+m355_19+m356_19+m357_19+m358_19+m359_19+m360_19+m361_19+m362_19+m363_19+m364_19+m365_19+m366_19+m367_19+m368_19+m369_19+m370_19+m371_19+m372_19+m373_19+m374_19+m375_19+m376_19+m377_19+m378_19+m379_19+m380_19+m381_19+b19;
   always @(posedge clk) out20 <= m1_20+m2_20+m3_20+m4_20+m5_20+m6_20+m7_20+m8_20+m9_20+m10_20+m11_20+m12_20+m13_20+m14_20+m15_20+m16_20+m17_20+m18_20+m19_20+m20_20+m21_20+m22_20+m23_20+m24_20+m25_20+m26_20+m27_20+m28_20+m29_20+m30_20+m31_20+m32_20+m33_20+m34_20+m35_20+m36_20+m37_20+m38_20+m39_20+m40_20+m41_20+m42_20+m43_20+m44_20+m45_20+m46_20+m47_20+m48_20+m49_20+m50_20+m51_20+m52_20+m53_20+m54_20+m55_20+m56_20+m57_20+m58_20+m59_20+m60_20+m61_20+m62_20+m63_20+m64_20+m65_20+m66_20+m67_20+m68_20+m69_20+m70_20+m71_20+m72_20+m73_20+m74_20+m75_20+m76_20+m77_20+m78_20+m79_20+m80_20+m81_20+m82_20+m83_20+m84_20+m85_20+m86_20+m87_20+m88_20+m89_20+m90_20+m91_20+m92_20+m93_20+m94_20+m95_20+m96_20+m97_20+m98_20+m99_20+m100_20+m101_20+m102_20+m103_20+m104_20+m105_20+m106_20+m107_20+m108_20+m109_20+m110_20+m111_20+m112_20+m113_20+m114_20+m115_20+m116_20+m117_20+m118_20+m119_20+m120_20+m121_20+m122_20+m123_20+m124_20+m125_20+m126_20+m127_20+m128_20+m129_20+m130_20+m131_20+m132_20+m133_20+m134_20+m135_20+m136_20+m137_20+m138_20+m139_20+m140_20+m141_20+m142_20+m143_20+m144_20+m145_20+m146_20+m147_20+m148_20+m149_20+m150_20+m151_20+m152_20+m153_20+m154_20+m155_20+m156_20+m157_20+m158_20+m159_20+m160_20+m161_20+m162_20+m163_20+m164_20+m165_20+m166_20+m167_20+m168_20+m169_20+m170_20+m171_20+m172_20+m173_20+m174_20+m175_20+m176_20+m177_20+m178_20+m179_20+m180_20+m181_20+m182_20+m183_20+m184_20+m185_20+m186_20+m187_20+m188_20+m189_20+m190_20+m191_20+m192_20+m193_20+m194_20+m195_20+m196_20+m197_20+m198_20+m199_20+m200_20+m201_20+m202_20+m203_20+m204_20+m205_20+m206_20+m207_20+m208_20+m209_20+m210_20+m211_20+m212_20+m213_20+m214_20+m215_20+m216_20+m217_20+m218_20+m219_20+m220_20+m221_20+m222_20+m223_20+m224_20+m225_20+m226_20+m227_20+m228_20+m229_20+m230_20+m231_20+m232_20+m233_20+m234_20+m235_20+m236_20+m237_20+m238_20+m239_20+m240_20+m241_20+m242_20+m243_20+m244_20+m245_20+m246_20+m247_20+m248_20+m249_20+m250_20+m251_20+m252_20+m253_20+m254_20+m255_20+m256_20+m257_20+m258_20+m259_20+m260_20+m261_20+m262_20+m263_20+m264_20+m265_20+m266_20+m267_20+m268_20+m269_20+m270_20+m271_20+m272_20+m273_20+m274_20+m275_20+m276_20+m277_20+m278_20+m279_20+m280_20+m281_20+m282_20+m283_20+m284_20+m285_20+m286_20+m287_20+m288_20+m289_20+m290_20+m291_20+m292_20+m293_20+m294_20+m295_20+m296_20+m297_20+m298_20+m299_20+m300_20+m301_20+m302_20+m303_20+m304_20+m305_20+m306_20+m307_20+m308_20+m309_20+m310_20+m311_20+m312_20+m313_20+m314_20+m315_20+m316_20+m317_20+m318_20+m319_20+m320_20+m321_20+m322_20+m323_20+m324_20+m325_20+m326_20+m327_20+m328_20+m329_20+m330_20+m331_20+m332_20+m333_20+m334_20+m335_20+m336_20+m337_20+m338_20+m339_20+m340_20+m341_20+m342_20+m343_20+m344_20+m345_20+m346_20+m347_20+m348_20+m349_20+m350_20+m351_20+m352_20+m353_20+m354_20+m355_20+m356_20+m357_20+m358_20+m359_20+m360_20+m361_20+m362_20+m363_20+m364_20+m365_20+m366_20+m367_20+m368_20+m369_20+m370_20+m371_20+m372_20+m373_20+m374_20+m375_20+m376_20+m377_20+m378_20+m379_20+m380_20+m381_20+b20;
   always @(posedge clk) out21 <= m1_21+m2_21+m3_21+m4_21+m5_21+m6_21+m7_21+m8_21+m9_21+m10_21+m11_21+m12_21+m13_21+m14_21+m15_21+m16_21+m17_21+m18_21+m19_21+m20_21+m21_21+m22_21+m23_21+m24_21+m25_21+m26_21+m27_21+m28_21+m29_21+m30_21+m31_21+m32_21+m33_21+m34_21+m35_21+m36_21+m37_21+m38_21+m39_21+m40_21+m41_21+m42_21+m43_21+m44_21+m45_21+m46_21+m47_21+m48_21+m49_21+m50_21+m51_21+m52_21+m53_21+m54_21+m55_21+m56_21+m57_21+m58_21+m59_21+m60_21+m61_21+m62_21+m63_21+m64_21+m65_21+m66_21+m67_21+m68_21+m69_21+m70_21+m71_21+m72_21+m73_21+m74_21+m75_21+m76_21+m77_21+m78_21+m79_21+m80_21+m81_21+m82_21+m83_21+m84_21+m85_21+m86_21+m87_21+m88_21+m89_21+m90_21+m91_21+m92_21+m93_21+m94_21+m95_21+m96_21+m97_21+m98_21+m99_21+m100_21+m101_21+m102_21+m103_21+m104_21+m105_21+m106_21+m107_21+m108_21+m109_21+m110_21+m111_21+m112_21+m113_21+m114_21+m115_21+m116_21+m117_21+m118_21+m119_21+m120_21+m121_21+m122_21+m123_21+m124_21+m125_21+m126_21+m127_21+m128_21+m129_21+m130_21+m131_21+m132_21+m133_21+m134_21+m135_21+m136_21+m137_21+m138_21+m139_21+m140_21+m141_21+m142_21+m143_21+m144_21+m145_21+m146_21+m147_21+m148_21+m149_21+m150_21+m151_21+m152_21+m153_21+m154_21+m155_21+m156_21+m157_21+m158_21+m159_21+m160_21+m161_21+m162_21+m163_21+m164_21+m165_21+m166_21+m167_21+m168_21+m169_21+m170_21+m171_21+m172_21+m173_21+m174_21+m175_21+m176_21+m177_21+m178_21+m179_21+m180_21+m181_21+m182_21+m183_21+m184_21+m185_21+m186_21+m187_21+m188_21+m189_21+m190_21+m191_21+m192_21+m193_21+m194_21+m195_21+m196_21+m197_21+m198_21+m199_21+m200_21+m201_21+m202_21+m203_21+m204_21+m205_21+m206_21+m207_21+m208_21+m209_21+m210_21+m211_21+m212_21+m213_21+m214_21+m215_21+m216_21+m217_21+m218_21+m219_21+m220_21+m221_21+m222_21+m223_21+m224_21+m225_21+m226_21+m227_21+m228_21+m229_21+m230_21+m231_21+m232_21+m233_21+m234_21+m235_21+m236_21+m237_21+m238_21+m239_21+m240_21+m241_21+m242_21+m243_21+m244_21+m245_21+m246_21+m247_21+m248_21+m249_21+m250_21+m251_21+m252_21+m253_21+m254_21+m255_21+m256_21+m257_21+m258_21+m259_21+m260_21+m261_21+m262_21+m263_21+m264_21+m265_21+m266_21+m267_21+m268_21+m269_21+m270_21+m271_21+m272_21+m273_21+m274_21+m275_21+m276_21+m277_21+m278_21+m279_21+m280_21+m281_21+m282_21+m283_21+m284_21+m285_21+m286_21+m287_21+m288_21+m289_21+m290_21+m291_21+m292_21+m293_21+m294_21+m295_21+m296_21+m297_21+m298_21+m299_21+m300_21+m301_21+m302_21+m303_21+m304_21+m305_21+m306_21+m307_21+m308_21+m309_21+m310_21+m311_21+m312_21+m313_21+m314_21+m315_21+m316_21+m317_21+m318_21+m319_21+m320_21+m321_21+m322_21+m323_21+m324_21+m325_21+m326_21+m327_21+m328_21+m329_21+m330_21+m331_21+m332_21+m333_21+m334_21+m335_21+m336_21+m337_21+m338_21+m339_21+m340_21+m341_21+m342_21+m343_21+m344_21+m345_21+m346_21+m347_21+m348_21+m349_21+m350_21+m351_21+m352_21+m353_21+m354_21+m355_21+m356_21+m357_21+m358_21+m359_21+m360_21+m361_21+m362_21+m363_21+m364_21+m365_21+m366_21+m367_21+m368_21+m369_21+m370_21+m371_21+m372_21+m373_21+m374_21+m375_21+m376_21+m377_21+m378_21+m379_21+m380_21+m381_21+b21;
   always @(posedge clk) out22 <= m1_22+m2_22+m3_22+m4_22+m5_22+m6_22+m7_22+m8_22+m9_22+m10_22+m11_22+m12_22+m13_22+m14_22+m15_22+m16_22+m17_22+m18_22+m19_22+m20_22+m21_22+m22_22+m23_22+m24_22+m25_22+m26_22+m27_22+m28_22+m29_22+m30_22+m31_22+m32_22+m33_22+m34_22+m35_22+m36_22+m37_22+m38_22+m39_22+m40_22+m41_22+m42_22+m43_22+m44_22+m45_22+m46_22+m47_22+m48_22+m49_22+m50_22+m51_22+m52_22+m53_22+m54_22+m55_22+m56_22+m57_22+m58_22+m59_22+m60_22+m61_22+m62_22+m63_22+m64_22+m65_22+m66_22+m67_22+m68_22+m69_22+m70_22+m71_22+m72_22+m73_22+m74_22+m75_22+m76_22+m77_22+m78_22+m79_22+m80_22+m81_22+m82_22+m83_22+m84_22+m85_22+m86_22+m87_22+m88_22+m89_22+m90_22+m91_22+m92_22+m93_22+m94_22+m95_22+m96_22+m97_22+m98_22+m99_22+m100_22+m101_22+m102_22+m103_22+m104_22+m105_22+m106_22+m107_22+m108_22+m109_22+m110_22+m111_22+m112_22+m113_22+m114_22+m115_22+m116_22+m117_22+m118_22+m119_22+m120_22+m121_22+m122_22+m123_22+m124_22+m125_22+m126_22+m127_22+m128_22+m129_22+m130_22+m131_22+m132_22+m133_22+m134_22+m135_22+m136_22+m137_22+m138_22+m139_22+m140_22+m141_22+m142_22+m143_22+m144_22+m145_22+m146_22+m147_22+m148_22+m149_22+m150_22+m151_22+m152_22+m153_22+m154_22+m155_22+m156_22+m157_22+m158_22+m159_22+m160_22+m161_22+m162_22+m163_22+m164_22+m165_22+m166_22+m167_22+m168_22+m169_22+m170_22+m171_22+m172_22+m173_22+m174_22+m175_22+m176_22+m177_22+m178_22+m179_22+m180_22+m181_22+m182_22+m183_22+m184_22+m185_22+m186_22+m187_22+m188_22+m189_22+m190_22+m191_22+m192_22+m193_22+m194_22+m195_22+m196_22+m197_22+m198_22+m199_22+m200_22+m201_22+m202_22+m203_22+m204_22+m205_22+m206_22+m207_22+m208_22+m209_22+m210_22+m211_22+m212_22+m213_22+m214_22+m215_22+m216_22+m217_22+m218_22+m219_22+m220_22+m221_22+m222_22+m223_22+m224_22+m225_22+m226_22+m227_22+m228_22+m229_22+m230_22+m231_22+m232_22+m233_22+m234_22+m235_22+m236_22+m237_22+m238_22+m239_22+m240_22+m241_22+m242_22+m243_22+m244_22+m245_22+m246_22+m247_22+m248_22+m249_22+m250_22+m251_22+m252_22+m253_22+m254_22+m255_22+m256_22+m257_22+m258_22+m259_22+m260_22+m261_22+m262_22+m263_22+m264_22+m265_22+m266_22+m267_22+m268_22+m269_22+m270_22+m271_22+m272_22+m273_22+m274_22+m275_22+m276_22+m277_22+m278_22+m279_22+m280_22+m281_22+m282_22+m283_22+m284_22+m285_22+m286_22+m287_22+m288_22+m289_22+m290_22+m291_22+m292_22+m293_22+m294_22+m295_22+m296_22+m297_22+m298_22+m299_22+m300_22+m301_22+m302_22+m303_22+m304_22+m305_22+m306_22+m307_22+m308_22+m309_22+m310_22+m311_22+m312_22+m313_22+m314_22+m315_22+m316_22+m317_22+m318_22+m319_22+m320_22+m321_22+m322_22+m323_22+m324_22+m325_22+m326_22+m327_22+m328_22+m329_22+m330_22+m331_22+m332_22+m333_22+m334_22+m335_22+m336_22+m337_22+m338_22+m339_22+m340_22+m341_22+m342_22+m343_22+m344_22+m345_22+m346_22+m347_22+m348_22+m349_22+m350_22+m351_22+m352_22+m353_22+m354_22+m355_22+m356_22+m357_22+m358_22+m359_22+m360_22+m361_22+m362_22+m363_22+m364_22+m365_22+m366_22+m367_22+m368_22+m369_22+m370_22+m371_22+m372_22+m373_22+m374_22+m375_22+m376_22+m377_22+m378_22+m379_22+m380_22+m381_22+b22;
   always @(posedge clk) out23 <= m1_23+m2_23+m3_23+m4_23+m5_23+m6_23+m7_23+m8_23+m9_23+m10_23+m11_23+m12_23+m13_23+m14_23+m15_23+m16_23+m17_23+m18_23+m19_23+m20_23+m21_23+m22_23+m23_23+m24_23+m25_23+m26_23+m27_23+m28_23+m29_23+m30_23+m31_23+m32_23+m33_23+m34_23+m35_23+m36_23+m37_23+m38_23+m39_23+m40_23+m41_23+m42_23+m43_23+m44_23+m45_23+m46_23+m47_23+m48_23+m49_23+m50_23+m51_23+m52_23+m53_23+m54_23+m55_23+m56_23+m57_23+m58_23+m59_23+m60_23+m61_23+m62_23+m63_23+m64_23+m65_23+m66_23+m67_23+m68_23+m69_23+m70_23+m71_23+m72_23+m73_23+m74_23+m75_23+m76_23+m77_23+m78_23+m79_23+m80_23+m81_23+m82_23+m83_23+m84_23+m85_23+m86_23+m87_23+m88_23+m89_23+m90_23+m91_23+m92_23+m93_23+m94_23+m95_23+m96_23+m97_23+m98_23+m99_23+m100_23+m101_23+m102_23+m103_23+m104_23+m105_23+m106_23+m107_23+m108_23+m109_23+m110_23+m111_23+m112_23+m113_23+m114_23+m115_23+m116_23+m117_23+m118_23+m119_23+m120_23+m121_23+m122_23+m123_23+m124_23+m125_23+m126_23+m127_23+m128_23+m129_23+m130_23+m131_23+m132_23+m133_23+m134_23+m135_23+m136_23+m137_23+m138_23+m139_23+m140_23+m141_23+m142_23+m143_23+m144_23+m145_23+m146_23+m147_23+m148_23+m149_23+m150_23+m151_23+m152_23+m153_23+m154_23+m155_23+m156_23+m157_23+m158_23+m159_23+m160_23+m161_23+m162_23+m163_23+m164_23+m165_23+m166_23+m167_23+m168_23+m169_23+m170_23+m171_23+m172_23+m173_23+m174_23+m175_23+m176_23+m177_23+m178_23+m179_23+m180_23+m181_23+m182_23+m183_23+m184_23+m185_23+m186_23+m187_23+m188_23+m189_23+m190_23+m191_23+m192_23+m193_23+m194_23+m195_23+m196_23+m197_23+m198_23+m199_23+m200_23+m201_23+m202_23+m203_23+m204_23+m205_23+m206_23+m207_23+m208_23+m209_23+m210_23+m211_23+m212_23+m213_23+m214_23+m215_23+m216_23+m217_23+m218_23+m219_23+m220_23+m221_23+m222_23+m223_23+m224_23+m225_23+m226_23+m227_23+m228_23+m229_23+m230_23+m231_23+m232_23+m233_23+m234_23+m235_23+m236_23+m237_23+m238_23+m239_23+m240_23+m241_23+m242_23+m243_23+m244_23+m245_23+m246_23+m247_23+m248_23+m249_23+m250_23+m251_23+m252_23+m253_23+m254_23+m255_23+m256_23+m257_23+m258_23+m259_23+m260_23+m261_23+m262_23+m263_23+m264_23+m265_23+m266_23+m267_23+m268_23+m269_23+m270_23+m271_23+m272_23+m273_23+m274_23+m275_23+m276_23+m277_23+m278_23+m279_23+m280_23+m281_23+m282_23+m283_23+m284_23+m285_23+m286_23+m287_23+m288_23+m289_23+m290_23+m291_23+m292_23+m293_23+m294_23+m295_23+m296_23+m297_23+m298_23+m299_23+m300_23+m301_23+m302_23+m303_23+m304_23+m305_23+m306_23+m307_23+m308_23+m309_23+m310_23+m311_23+m312_23+m313_23+m314_23+m315_23+m316_23+m317_23+m318_23+m319_23+m320_23+m321_23+m322_23+m323_23+m324_23+m325_23+m326_23+m327_23+m328_23+m329_23+m330_23+m331_23+m332_23+m333_23+m334_23+m335_23+m336_23+m337_23+m338_23+m339_23+m340_23+m341_23+m342_23+m343_23+m344_23+m345_23+m346_23+m347_23+m348_23+m349_23+m350_23+m351_23+m352_23+m353_23+m354_23+m355_23+m356_23+m357_23+m358_23+m359_23+m360_23+m361_23+m362_23+m363_23+m364_23+m365_23+m366_23+m367_23+m368_23+m369_23+m370_23+m371_23+m372_23+m373_23+m374_23+m375_23+m376_23+m377_23+m378_23+m379_23+m380_23+m381_23+b23;
   always @(posedge clk) out24 <= m1_24+m2_24+m3_24+m4_24+m5_24+m6_24+m7_24+m8_24+m9_24+m10_24+m11_24+m12_24+m13_24+m14_24+m15_24+m16_24+m17_24+m18_24+m19_24+m20_24+m21_24+m22_24+m23_24+m24_24+m25_24+m26_24+m27_24+m28_24+m29_24+m30_24+m31_24+m32_24+m33_24+m34_24+m35_24+m36_24+m37_24+m38_24+m39_24+m40_24+m41_24+m42_24+m43_24+m44_24+m45_24+m46_24+m47_24+m48_24+m49_24+m50_24+m51_24+m52_24+m53_24+m54_24+m55_24+m56_24+m57_24+m58_24+m59_24+m60_24+m61_24+m62_24+m63_24+m64_24+m65_24+m66_24+m67_24+m68_24+m69_24+m70_24+m71_24+m72_24+m73_24+m74_24+m75_24+m76_24+m77_24+m78_24+m79_24+m80_24+m81_24+m82_24+m83_24+m84_24+m85_24+m86_24+m87_24+m88_24+m89_24+m90_24+m91_24+m92_24+m93_24+m94_24+m95_24+m96_24+m97_24+m98_24+m99_24+m100_24+m101_24+m102_24+m103_24+m104_24+m105_24+m106_24+m107_24+m108_24+m109_24+m110_24+m111_24+m112_24+m113_24+m114_24+m115_24+m116_24+m117_24+m118_24+m119_24+m120_24+m121_24+m122_24+m123_24+m124_24+m125_24+m126_24+m127_24+m128_24+m129_24+m130_24+m131_24+m132_24+m133_24+m134_24+m135_24+m136_24+m137_24+m138_24+m139_24+m140_24+m141_24+m142_24+m143_24+m144_24+m145_24+m146_24+m147_24+m148_24+m149_24+m150_24+m151_24+m152_24+m153_24+m154_24+m155_24+m156_24+m157_24+m158_24+m159_24+m160_24+m161_24+m162_24+m163_24+m164_24+m165_24+m166_24+m167_24+m168_24+m169_24+m170_24+m171_24+m172_24+m173_24+m174_24+m175_24+m176_24+m177_24+m178_24+m179_24+m180_24+m181_24+m182_24+m183_24+m184_24+m185_24+m186_24+m187_24+m188_24+m189_24+m190_24+m191_24+m192_24+m193_24+m194_24+m195_24+m196_24+m197_24+m198_24+m199_24+m200_24+m201_24+m202_24+m203_24+m204_24+m205_24+m206_24+m207_24+m208_24+m209_24+m210_24+m211_24+m212_24+m213_24+m214_24+m215_24+m216_24+m217_24+m218_24+m219_24+m220_24+m221_24+m222_24+m223_24+m224_24+m225_24+m226_24+m227_24+m228_24+m229_24+m230_24+m231_24+m232_24+m233_24+m234_24+m235_24+m236_24+m237_24+m238_24+m239_24+m240_24+m241_24+m242_24+m243_24+m244_24+m245_24+m246_24+m247_24+m248_24+m249_24+m250_24+m251_24+m252_24+m253_24+m254_24+m255_24+m256_24+m257_24+m258_24+m259_24+m260_24+m261_24+m262_24+m263_24+m264_24+m265_24+m266_24+m267_24+m268_24+m269_24+m270_24+m271_24+m272_24+m273_24+m274_24+m275_24+m276_24+m277_24+m278_24+m279_24+m280_24+m281_24+m282_24+m283_24+m284_24+m285_24+m286_24+m287_24+m288_24+m289_24+m290_24+m291_24+m292_24+m293_24+m294_24+m295_24+m296_24+m297_24+m298_24+m299_24+m300_24+m301_24+m302_24+m303_24+m304_24+m305_24+m306_24+m307_24+m308_24+m309_24+m310_24+m311_24+m312_24+m313_24+m314_24+m315_24+m316_24+m317_24+m318_24+m319_24+m320_24+m321_24+m322_24+m323_24+m324_24+m325_24+m326_24+m327_24+m328_24+m329_24+m330_24+m331_24+m332_24+m333_24+m334_24+m335_24+m336_24+m337_24+m338_24+m339_24+m340_24+m341_24+m342_24+m343_24+m344_24+m345_24+m346_24+m347_24+m348_24+m349_24+m350_24+m351_24+m352_24+m353_24+m354_24+m355_24+m356_24+m357_24+m358_24+m359_24+m360_24+m361_24+m362_24+m363_24+m364_24+m365_24+m366_24+m367_24+m368_24+m369_24+m370_24+m371_24+m372_24+m373_24+m374_24+m375_24+m376_24+m377_24+m378_24+m379_24+m380_24+m381_24+b24;
   always @(posedge clk) out25 <= m1_25+m2_25+m3_25+m4_25+m5_25+m6_25+m7_25+m8_25+m9_25+m10_25+m11_25+m12_25+m13_25+m14_25+m15_25+m16_25+m17_25+m18_25+m19_25+m20_25+m21_25+m22_25+m23_25+m24_25+m25_25+m26_25+m27_25+m28_25+m29_25+m30_25+m31_25+m32_25+m33_25+m34_25+m35_25+m36_25+m37_25+m38_25+m39_25+m40_25+m41_25+m42_25+m43_25+m44_25+m45_25+m46_25+m47_25+m48_25+m49_25+m50_25+m51_25+m52_25+m53_25+m54_25+m55_25+m56_25+m57_25+m58_25+m59_25+m60_25+m61_25+m62_25+m63_25+m64_25+m65_25+m66_25+m67_25+m68_25+m69_25+m70_25+m71_25+m72_25+m73_25+m74_25+m75_25+m76_25+m77_25+m78_25+m79_25+m80_25+m81_25+m82_25+m83_25+m84_25+m85_25+m86_25+m87_25+m88_25+m89_25+m90_25+m91_25+m92_25+m93_25+m94_25+m95_25+m96_25+m97_25+m98_25+m99_25+m100_25+m101_25+m102_25+m103_25+m104_25+m105_25+m106_25+m107_25+m108_25+m109_25+m110_25+m111_25+m112_25+m113_25+m114_25+m115_25+m116_25+m117_25+m118_25+m119_25+m120_25+m121_25+m122_25+m123_25+m124_25+m125_25+m126_25+m127_25+m128_25+m129_25+m130_25+m131_25+m132_25+m133_25+m134_25+m135_25+m136_25+m137_25+m138_25+m139_25+m140_25+m141_25+m142_25+m143_25+m144_25+m145_25+m146_25+m147_25+m148_25+m149_25+m150_25+m151_25+m152_25+m153_25+m154_25+m155_25+m156_25+m157_25+m158_25+m159_25+m160_25+m161_25+m162_25+m163_25+m164_25+m165_25+m166_25+m167_25+m168_25+m169_25+m170_25+m171_25+m172_25+m173_25+m174_25+m175_25+m176_25+m177_25+m178_25+m179_25+m180_25+m181_25+m182_25+m183_25+m184_25+m185_25+m186_25+m187_25+m188_25+m189_25+m190_25+m191_25+m192_25+m193_25+m194_25+m195_25+m196_25+m197_25+m198_25+m199_25+m200_25+m201_25+m202_25+m203_25+m204_25+m205_25+m206_25+m207_25+m208_25+m209_25+m210_25+m211_25+m212_25+m213_25+m214_25+m215_25+m216_25+m217_25+m218_25+m219_25+m220_25+m221_25+m222_25+m223_25+m224_25+m225_25+m226_25+m227_25+m228_25+m229_25+m230_25+m231_25+m232_25+m233_25+m234_25+m235_25+m236_25+m237_25+m238_25+m239_25+m240_25+m241_25+m242_25+m243_25+m244_25+m245_25+m246_25+m247_25+m248_25+m249_25+m250_25+m251_25+m252_25+m253_25+m254_25+m255_25+m256_25+m257_25+m258_25+m259_25+m260_25+m261_25+m262_25+m263_25+m264_25+m265_25+m266_25+m267_25+m268_25+m269_25+m270_25+m271_25+m272_25+m273_25+m274_25+m275_25+m276_25+m277_25+m278_25+m279_25+m280_25+m281_25+m282_25+m283_25+m284_25+m285_25+m286_25+m287_25+m288_25+m289_25+m290_25+m291_25+m292_25+m293_25+m294_25+m295_25+m296_25+m297_25+m298_25+m299_25+m300_25+m301_25+m302_25+m303_25+m304_25+m305_25+m306_25+m307_25+m308_25+m309_25+m310_25+m311_25+m312_25+m313_25+m314_25+m315_25+m316_25+m317_25+m318_25+m319_25+m320_25+m321_25+m322_25+m323_25+m324_25+m325_25+m326_25+m327_25+m328_25+m329_25+m330_25+m331_25+m332_25+m333_25+m334_25+m335_25+m336_25+m337_25+m338_25+m339_25+m340_25+m341_25+m342_25+m343_25+m344_25+m345_25+m346_25+m347_25+m348_25+m349_25+m350_25+m351_25+m352_25+m353_25+m354_25+m355_25+m356_25+m357_25+m358_25+m359_25+m360_25+m361_25+m362_25+m363_25+m364_25+m365_25+m366_25+m367_25+m368_25+m369_25+m370_25+m371_25+m372_25+m373_25+m374_25+m375_25+m376_25+m377_25+m378_25+m379_25+m380_25+m381_25+b25;
   always @(posedge clk) out26 <= m1_26+m2_26+m3_26+m4_26+m5_26+m6_26+m7_26+m8_26+m9_26+m10_26+m11_26+m12_26+m13_26+m14_26+m15_26+m16_26+m17_26+m18_26+m19_26+m20_26+m21_26+m22_26+m23_26+m24_26+m25_26+m26_26+m27_26+m28_26+m29_26+m30_26+m31_26+m32_26+m33_26+m34_26+m35_26+m36_26+m37_26+m38_26+m39_26+m40_26+m41_26+m42_26+m43_26+m44_26+m45_26+m46_26+m47_26+m48_26+m49_26+m50_26+m51_26+m52_26+m53_26+m54_26+m55_26+m56_26+m57_26+m58_26+m59_26+m60_26+m61_26+m62_26+m63_26+m64_26+m65_26+m66_26+m67_26+m68_26+m69_26+m70_26+m71_26+m72_26+m73_26+m74_26+m75_26+m76_26+m77_26+m78_26+m79_26+m80_26+m81_26+m82_26+m83_26+m84_26+m85_26+m86_26+m87_26+m88_26+m89_26+m90_26+m91_26+m92_26+m93_26+m94_26+m95_26+m96_26+m97_26+m98_26+m99_26+m100_26+m101_26+m102_26+m103_26+m104_26+m105_26+m106_26+m107_26+m108_26+m109_26+m110_26+m111_26+m112_26+m113_26+m114_26+m115_26+m116_26+m117_26+m118_26+m119_26+m120_26+m121_26+m122_26+m123_26+m124_26+m125_26+m126_26+m127_26+m128_26+m129_26+m130_26+m131_26+m132_26+m133_26+m134_26+m135_26+m136_26+m137_26+m138_26+m139_26+m140_26+m141_26+m142_26+m143_26+m144_26+m145_26+m146_26+m147_26+m148_26+m149_26+m150_26+m151_26+m152_26+m153_26+m154_26+m155_26+m156_26+m157_26+m158_26+m159_26+m160_26+m161_26+m162_26+m163_26+m164_26+m165_26+m166_26+m167_26+m168_26+m169_26+m170_26+m171_26+m172_26+m173_26+m174_26+m175_26+m176_26+m177_26+m178_26+m179_26+m180_26+m181_26+m182_26+m183_26+m184_26+m185_26+m186_26+m187_26+m188_26+m189_26+m190_26+m191_26+m192_26+m193_26+m194_26+m195_26+m196_26+m197_26+m198_26+m199_26+m200_26+m201_26+m202_26+m203_26+m204_26+m205_26+m206_26+m207_26+m208_26+m209_26+m210_26+m211_26+m212_26+m213_26+m214_26+m215_26+m216_26+m217_26+m218_26+m219_26+m220_26+m221_26+m222_26+m223_26+m224_26+m225_26+m226_26+m227_26+m228_26+m229_26+m230_26+m231_26+m232_26+m233_26+m234_26+m235_26+m236_26+m237_26+m238_26+m239_26+m240_26+m241_26+m242_26+m243_26+m244_26+m245_26+m246_26+m247_26+m248_26+m249_26+m250_26+m251_26+m252_26+m253_26+m254_26+m255_26+m256_26+m257_26+m258_26+m259_26+m260_26+m261_26+m262_26+m263_26+m264_26+m265_26+m266_26+m267_26+m268_26+m269_26+m270_26+m271_26+m272_26+m273_26+m274_26+m275_26+m276_26+m277_26+m278_26+m279_26+m280_26+m281_26+m282_26+m283_26+m284_26+m285_26+m286_26+m287_26+m288_26+m289_26+m290_26+m291_26+m292_26+m293_26+m294_26+m295_26+m296_26+m297_26+m298_26+m299_26+m300_26+m301_26+m302_26+m303_26+m304_26+m305_26+m306_26+m307_26+m308_26+m309_26+m310_26+m311_26+m312_26+m313_26+m314_26+m315_26+m316_26+m317_26+m318_26+m319_26+m320_26+m321_26+m322_26+m323_26+m324_26+m325_26+m326_26+m327_26+m328_26+m329_26+m330_26+m331_26+m332_26+m333_26+m334_26+m335_26+m336_26+m337_26+m338_26+m339_26+m340_26+m341_26+m342_26+m343_26+m344_26+m345_26+m346_26+m347_26+m348_26+m349_26+m350_26+m351_26+m352_26+m353_26+m354_26+m355_26+m356_26+m357_26+m358_26+m359_26+m360_26+m361_26+m362_26+m363_26+m364_26+m365_26+m366_26+m367_26+m368_26+m369_26+m370_26+m371_26+m372_26+m373_26+m374_26+m375_26+m376_26+m377_26+m378_26+m379_26+m380_26+m381_26+b26;
   always @(posedge clk) out27 <= m1_27+m2_27+m3_27+m4_27+m5_27+m6_27+m7_27+m8_27+m9_27+m10_27+m11_27+m12_27+m13_27+m14_27+m15_27+m16_27+m17_27+m18_27+m19_27+m20_27+m21_27+m22_27+m23_27+m24_27+m25_27+m26_27+m27_27+m28_27+m29_27+m30_27+m31_27+m32_27+m33_27+m34_27+m35_27+m36_27+m37_27+m38_27+m39_27+m40_27+m41_27+m42_27+m43_27+m44_27+m45_27+m46_27+m47_27+m48_27+m49_27+m50_27+m51_27+m52_27+m53_27+m54_27+m55_27+m56_27+m57_27+m58_27+m59_27+m60_27+m61_27+m62_27+m63_27+m64_27+m65_27+m66_27+m67_27+m68_27+m69_27+m70_27+m71_27+m72_27+m73_27+m74_27+m75_27+m76_27+m77_27+m78_27+m79_27+m80_27+m81_27+m82_27+m83_27+m84_27+m85_27+m86_27+m87_27+m88_27+m89_27+m90_27+m91_27+m92_27+m93_27+m94_27+m95_27+m96_27+m97_27+m98_27+m99_27+m100_27+m101_27+m102_27+m103_27+m104_27+m105_27+m106_27+m107_27+m108_27+m109_27+m110_27+m111_27+m112_27+m113_27+m114_27+m115_27+m116_27+m117_27+m118_27+m119_27+m120_27+m121_27+m122_27+m123_27+m124_27+m125_27+m126_27+m127_27+m128_27+m129_27+m130_27+m131_27+m132_27+m133_27+m134_27+m135_27+m136_27+m137_27+m138_27+m139_27+m140_27+m141_27+m142_27+m143_27+m144_27+m145_27+m146_27+m147_27+m148_27+m149_27+m150_27+m151_27+m152_27+m153_27+m154_27+m155_27+m156_27+m157_27+m158_27+m159_27+m160_27+m161_27+m162_27+m163_27+m164_27+m165_27+m166_27+m167_27+m168_27+m169_27+m170_27+m171_27+m172_27+m173_27+m174_27+m175_27+m176_27+m177_27+m178_27+m179_27+m180_27+m181_27+m182_27+m183_27+m184_27+m185_27+m186_27+m187_27+m188_27+m189_27+m190_27+m191_27+m192_27+m193_27+m194_27+m195_27+m196_27+m197_27+m198_27+m199_27+m200_27+m201_27+m202_27+m203_27+m204_27+m205_27+m206_27+m207_27+m208_27+m209_27+m210_27+m211_27+m212_27+m213_27+m214_27+m215_27+m216_27+m217_27+m218_27+m219_27+m220_27+m221_27+m222_27+m223_27+m224_27+m225_27+m226_27+m227_27+m228_27+m229_27+m230_27+m231_27+m232_27+m233_27+m234_27+m235_27+m236_27+m237_27+m238_27+m239_27+m240_27+m241_27+m242_27+m243_27+m244_27+m245_27+m246_27+m247_27+m248_27+m249_27+m250_27+m251_27+m252_27+m253_27+m254_27+m255_27+m256_27+m257_27+m258_27+m259_27+m260_27+m261_27+m262_27+m263_27+m264_27+m265_27+m266_27+m267_27+m268_27+m269_27+m270_27+m271_27+m272_27+m273_27+m274_27+m275_27+m276_27+m277_27+m278_27+m279_27+m280_27+m281_27+m282_27+m283_27+m284_27+m285_27+m286_27+m287_27+m288_27+m289_27+m290_27+m291_27+m292_27+m293_27+m294_27+m295_27+m296_27+m297_27+m298_27+m299_27+m300_27+m301_27+m302_27+m303_27+m304_27+m305_27+m306_27+m307_27+m308_27+m309_27+m310_27+m311_27+m312_27+m313_27+m314_27+m315_27+m316_27+m317_27+m318_27+m319_27+m320_27+m321_27+m322_27+m323_27+m324_27+m325_27+m326_27+m327_27+m328_27+m329_27+m330_27+m331_27+m332_27+m333_27+m334_27+m335_27+m336_27+m337_27+m338_27+m339_27+m340_27+m341_27+m342_27+m343_27+m344_27+m345_27+m346_27+m347_27+m348_27+m349_27+m350_27+m351_27+m352_27+m353_27+m354_27+m355_27+m356_27+m357_27+m358_27+m359_27+m360_27+m361_27+m362_27+m363_27+m364_27+m365_27+m366_27+m367_27+m368_27+m369_27+m370_27+m371_27+m372_27+m373_27+m374_27+m375_27+m376_27+m377_27+m378_27+m379_27+m380_27+m381_27+b27;
   always @(posedge clk) out28 <= m1_28+m2_28+m3_28+m4_28+m5_28+m6_28+m7_28+m8_28+m9_28+m10_28+m11_28+m12_28+m13_28+m14_28+m15_28+m16_28+m17_28+m18_28+m19_28+m20_28+m21_28+m22_28+m23_28+m24_28+m25_28+m26_28+m27_28+m28_28+m29_28+m30_28+m31_28+m32_28+m33_28+m34_28+m35_28+m36_28+m37_28+m38_28+m39_28+m40_28+m41_28+m42_28+m43_28+m44_28+m45_28+m46_28+m47_28+m48_28+m49_28+m50_28+m51_28+m52_28+m53_28+m54_28+m55_28+m56_28+m57_28+m58_28+m59_28+m60_28+m61_28+m62_28+m63_28+m64_28+m65_28+m66_28+m67_28+m68_28+m69_28+m70_28+m71_28+m72_28+m73_28+m74_28+m75_28+m76_28+m77_28+m78_28+m79_28+m80_28+m81_28+m82_28+m83_28+m84_28+m85_28+m86_28+m87_28+m88_28+m89_28+m90_28+m91_28+m92_28+m93_28+m94_28+m95_28+m96_28+m97_28+m98_28+m99_28+m100_28+m101_28+m102_28+m103_28+m104_28+m105_28+m106_28+m107_28+m108_28+m109_28+m110_28+m111_28+m112_28+m113_28+m114_28+m115_28+m116_28+m117_28+m118_28+m119_28+m120_28+m121_28+m122_28+m123_28+m124_28+m125_28+m126_28+m127_28+m128_28+m129_28+m130_28+m131_28+m132_28+m133_28+m134_28+m135_28+m136_28+m137_28+m138_28+m139_28+m140_28+m141_28+m142_28+m143_28+m144_28+m145_28+m146_28+m147_28+m148_28+m149_28+m150_28+m151_28+m152_28+m153_28+m154_28+m155_28+m156_28+m157_28+m158_28+m159_28+m160_28+m161_28+m162_28+m163_28+m164_28+m165_28+m166_28+m167_28+m168_28+m169_28+m170_28+m171_28+m172_28+m173_28+m174_28+m175_28+m176_28+m177_28+m178_28+m179_28+m180_28+m181_28+m182_28+m183_28+m184_28+m185_28+m186_28+m187_28+m188_28+m189_28+m190_28+m191_28+m192_28+m193_28+m194_28+m195_28+m196_28+m197_28+m198_28+m199_28+m200_28+m201_28+m202_28+m203_28+m204_28+m205_28+m206_28+m207_28+m208_28+m209_28+m210_28+m211_28+m212_28+m213_28+m214_28+m215_28+m216_28+m217_28+m218_28+m219_28+m220_28+m221_28+m222_28+m223_28+m224_28+m225_28+m226_28+m227_28+m228_28+m229_28+m230_28+m231_28+m232_28+m233_28+m234_28+m235_28+m236_28+m237_28+m238_28+m239_28+m240_28+m241_28+m242_28+m243_28+m244_28+m245_28+m246_28+m247_28+m248_28+m249_28+m250_28+m251_28+m252_28+m253_28+m254_28+m255_28+m256_28+m257_28+m258_28+m259_28+m260_28+m261_28+m262_28+m263_28+m264_28+m265_28+m266_28+m267_28+m268_28+m269_28+m270_28+m271_28+m272_28+m273_28+m274_28+m275_28+m276_28+m277_28+m278_28+m279_28+m280_28+m281_28+m282_28+m283_28+m284_28+m285_28+m286_28+m287_28+m288_28+m289_28+m290_28+m291_28+m292_28+m293_28+m294_28+m295_28+m296_28+m297_28+m298_28+m299_28+m300_28+m301_28+m302_28+m303_28+m304_28+m305_28+m306_28+m307_28+m308_28+m309_28+m310_28+m311_28+m312_28+m313_28+m314_28+m315_28+m316_28+m317_28+m318_28+m319_28+m320_28+m321_28+m322_28+m323_28+m324_28+m325_28+m326_28+m327_28+m328_28+m329_28+m330_28+m331_28+m332_28+m333_28+m334_28+m335_28+m336_28+m337_28+m338_28+m339_28+m340_28+m341_28+m342_28+m343_28+m344_28+m345_28+m346_28+m347_28+m348_28+m349_28+m350_28+m351_28+m352_28+m353_28+m354_28+m355_28+m356_28+m357_28+m358_28+m359_28+m360_28+m361_28+m362_28+m363_28+m364_28+m365_28+m366_28+m367_28+m368_28+m369_28+m370_28+m371_28+m372_28+m373_28+m374_28+m375_28+m376_28+m377_28+m378_28+m379_28+m380_28+m381_28+b28;
   always @(posedge clk) out29 <= m1_29+m2_29+m3_29+m4_29+m5_29+m6_29+m7_29+m8_29+m9_29+m10_29+m11_29+m12_29+m13_29+m14_29+m15_29+m16_29+m17_29+m18_29+m19_29+m20_29+m21_29+m22_29+m23_29+m24_29+m25_29+m26_29+m27_29+m28_29+m29_29+m30_29+m31_29+m32_29+m33_29+m34_29+m35_29+m36_29+m37_29+m38_29+m39_29+m40_29+m41_29+m42_29+m43_29+m44_29+m45_29+m46_29+m47_29+m48_29+m49_29+m50_29+m51_29+m52_29+m53_29+m54_29+m55_29+m56_29+m57_29+m58_29+m59_29+m60_29+m61_29+m62_29+m63_29+m64_29+m65_29+m66_29+m67_29+m68_29+m69_29+m70_29+m71_29+m72_29+m73_29+m74_29+m75_29+m76_29+m77_29+m78_29+m79_29+m80_29+m81_29+m82_29+m83_29+m84_29+m85_29+m86_29+m87_29+m88_29+m89_29+m90_29+m91_29+m92_29+m93_29+m94_29+m95_29+m96_29+m97_29+m98_29+m99_29+m100_29+m101_29+m102_29+m103_29+m104_29+m105_29+m106_29+m107_29+m108_29+m109_29+m110_29+m111_29+m112_29+m113_29+m114_29+m115_29+m116_29+m117_29+m118_29+m119_29+m120_29+m121_29+m122_29+m123_29+m124_29+m125_29+m126_29+m127_29+m128_29+m129_29+m130_29+m131_29+m132_29+m133_29+m134_29+m135_29+m136_29+m137_29+m138_29+m139_29+m140_29+m141_29+m142_29+m143_29+m144_29+m145_29+m146_29+m147_29+m148_29+m149_29+m150_29+m151_29+m152_29+m153_29+m154_29+m155_29+m156_29+m157_29+m158_29+m159_29+m160_29+m161_29+m162_29+m163_29+m164_29+m165_29+m166_29+m167_29+m168_29+m169_29+m170_29+m171_29+m172_29+m173_29+m174_29+m175_29+m176_29+m177_29+m178_29+m179_29+m180_29+m181_29+m182_29+m183_29+m184_29+m185_29+m186_29+m187_29+m188_29+m189_29+m190_29+m191_29+m192_29+m193_29+m194_29+m195_29+m196_29+m197_29+m198_29+m199_29+m200_29+m201_29+m202_29+m203_29+m204_29+m205_29+m206_29+m207_29+m208_29+m209_29+m210_29+m211_29+m212_29+m213_29+m214_29+m215_29+m216_29+m217_29+m218_29+m219_29+m220_29+m221_29+m222_29+m223_29+m224_29+m225_29+m226_29+m227_29+m228_29+m229_29+m230_29+m231_29+m232_29+m233_29+m234_29+m235_29+m236_29+m237_29+m238_29+m239_29+m240_29+m241_29+m242_29+m243_29+m244_29+m245_29+m246_29+m247_29+m248_29+m249_29+m250_29+m251_29+m252_29+m253_29+m254_29+m255_29+m256_29+m257_29+m258_29+m259_29+m260_29+m261_29+m262_29+m263_29+m264_29+m265_29+m266_29+m267_29+m268_29+m269_29+m270_29+m271_29+m272_29+m273_29+m274_29+m275_29+m276_29+m277_29+m278_29+m279_29+m280_29+m281_29+m282_29+m283_29+m284_29+m285_29+m286_29+m287_29+m288_29+m289_29+m290_29+m291_29+m292_29+m293_29+m294_29+m295_29+m296_29+m297_29+m298_29+m299_29+m300_29+m301_29+m302_29+m303_29+m304_29+m305_29+m306_29+m307_29+m308_29+m309_29+m310_29+m311_29+m312_29+m313_29+m314_29+m315_29+m316_29+m317_29+m318_29+m319_29+m320_29+m321_29+m322_29+m323_29+m324_29+m325_29+m326_29+m327_29+m328_29+m329_29+m330_29+m331_29+m332_29+m333_29+m334_29+m335_29+m336_29+m337_29+m338_29+m339_29+m340_29+m341_29+m342_29+m343_29+m344_29+m345_29+m346_29+m347_29+m348_29+m349_29+m350_29+m351_29+m352_29+m353_29+m354_29+m355_29+m356_29+m357_29+m358_29+m359_29+m360_29+m361_29+m362_29+m363_29+m364_29+m365_29+m366_29+m367_29+m368_29+m369_29+m370_29+m371_29+m372_29+m373_29+m374_29+m375_29+m376_29+m377_29+m378_29+m379_29+m380_29+m381_29+b29;
   always @(posedge clk) out30 <= m1_30+m2_30+m3_30+m4_30+m5_30+m6_30+m7_30+m8_30+m9_30+m10_30+m11_30+m12_30+m13_30+m14_30+m15_30+m16_30+m17_30+m18_30+m19_30+m20_30+m21_30+m22_30+m23_30+m24_30+m25_30+m26_30+m27_30+m28_30+m29_30+m30_30+m31_30+m32_30+m33_30+m34_30+m35_30+m36_30+m37_30+m38_30+m39_30+m40_30+m41_30+m42_30+m43_30+m44_30+m45_30+m46_30+m47_30+m48_30+m49_30+m50_30+m51_30+m52_30+m53_30+m54_30+m55_30+m56_30+m57_30+m58_30+m59_30+m60_30+m61_30+m62_30+m63_30+m64_30+m65_30+m66_30+m67_30+m68_30+m69_30+m70_30+m71_30+m72_30+m73_30+m74_30+m75_30+m76_30+m77_30+m78_30+m79_30+m80_30+m81_30+m82_30+m83_30+m84_30+m85_30+m86_30+m87_30+m88_30+m89_30+m90_30+m91_30+m92_30+m93_30+m94_30+m95_30+m96_30+m97_30+m98_30+m99_30+m100_30+m101_30+m102_30+m103_30+m104_30+m105_30+m106_30+m107_30+m108_30+m109_30+m110_30+m111_30+m112_30+m113_30+m114_30+m115_30+m116_30+m117_30+m118_30+m119_30+m120_30+m121_30+m122_30+m123_30+m124_30+m125_30+m126_30+m127_30+m128_30+m129_30+m130_30+m131_30+m132_30+m133_30+m134_30+m135_30+m136_30+m137_30+m138_30+m139_30+m140_30+m141_30+m142_30+m143_30+m144_30+m145_30+m146_30+m147_30+m148_30+m149_30+m150_30+m151_30+m152_30+m153_30+m154_30+m155_30+m156_30+m157_30+m158_30+m159_30+m160_30+m161_30+m162_30+m163_30+m164_30+m165_30+m166_30+m167_30+m168_30+m169_30+m170_30+m171_30+m172_30+m173_30+m174_30+m175_30+m176_30+m177_30+m178_30+m179_30+m180_30+m181_30+m182_30+m183_30+m184_30+m185_30+m186_30+m187_30+m188_30+m189_30+m190_30+m191_30+m192_30+m193_30+m194_30+m195_30+m196_30+m197_30+m198_30+m199_30+m200_30+m201_30+m202_30+m203_30+m204_30+m205_30+m206_30+m207_30+m208_30+m209_30+m210_30+m211_30+m212_30+m213_30+m214_30+m215_30+m216_30+m217_30+m218_30+m219_30+m220_30+m221_30+m222_30+m223_30+m224_30+m225_30+m226_30+m227_30+m228_30+m229_30+m230_30+m231_30+m232_30+m233_30+m234_30+m235_30+m236_30+m237_30+m238_30+m239_30+m240_30+m241_30+m242_30+m243_30+m244_30+m245_30+m246_30+m247_30+m248_30+m249_30+m250_30+m251_30+m252_30+m253_30+m254_30+m255_30+m256_30+m257_30+m258_30+m259_30+m260_30+m261_30+m262_30+m263_30+m264_30+m265_30+m266_30+m267_30+m268_30+m269_30+m270_30+m271_30+m272_30+m273_30+m274_30+m275_30+m276_30+m277_30+m278_30+m279_30+m280_30+m281_30+m282_30+m283_30+m284_30+m285_30+m286_30+m287_30+m288_30+m289_30+m290_30+m291_30+m292_30+m293_30+m294_30+m295_30+m296_30+m297_30+m298_30+m299_30+m300_30+m301_30+m302_30+m303_30+m304_30+m305_30+m306_30+m307_30+m308_30+m309_30+m310_30+m311_30+m312_30+m313_30+m314_30+m315_30+m316_30+m317_30+m318_30+m319_30+m320_30+m321_30+m322_30+m323_30+m324_30+m325_30+m326_30+m327_30+m328_30+m329_30+m330_30+m331_30+m332_30+m333_30+m334_30+m335_30+m336_30+m337_30+m338_30+m339_30+m340_30+m341_30+m342_30+m343_30+m344_30+m345_30+m346_30+m347_30+m348_30+m349_30+m350_30+m351_30+m352_30+m353_30+m354_30+m355_30+m356_30+m357_30+m358_30+m359_30+m360_30+m361_30+m362_30+m363_30+m364_30+m365_30+m366_30+m367_30+m368_30+m369_30+m370_30+m371_30+m372_30+m373_30+m374_30+m375_30+m376_30+m377_30+m378_30+m379_30+m380_30+m381_30+b30;
   always @(posedge clk) out31 <= m1_31+m2_31+m3_31+m4_31+m5_31+m6_31+m7_31+m8_31+m9_31+m10_31+m11_31+m12_31+m13_31+m14_31+m15_31+m16_31+m17_31+m18_31+m19_31+m20_31+m21_31+m22_31+m23_31+m24_31+m25_31+m26_31+m27_31+m28_31+m29_31+m30_31+m31_31+m32_31+m33_31+m34_31+m35_31+m36_31+m37_31+m38_31+m39_31+m40_31+m41_31+m42_31+m43_31+m44_31+m45_31+m46_31+m47_31+m48_31+m49_31+m50_31+m51_31+m52_31+m53_31+m54_31+m55_31+m56_31+m57_31+m58_31+m59_31+m60_31+m61_31+m62_31+m63_31+m64_31+m65_31+m66_31+m67_31+m68_31+m69_31+m70_31+m71_31+m72_31+m73_31+m74_31+m75_31+m76_31+m77_31+m78_31+m79_31+m80_31+m81_31+m82_31+m83_31+m84_31+m85_31+m86_31+m87_31+m88_31+m89_31+m90_31+m91_31+m92_31+m93_31+m94_31+m95_31+m96_31+m97_31+m98_31+m99_31+m100_31+m101_31+m102_31+m103_31+m104_31+m105_31+m106_31+m107_31+m108_31+m109_31+m110_31+m111_31+m112_31+m113_31+m114_31+m115_31+m116_31+m117_31+m118_31+m119_31+m120_31+m121_31+m122_31+m123_31+m124_31+m125_31+m126_31+m127_31+m128_31+m129_31+m130_31+m131_31+m132_31+m133_31+m134_31+m135_31+m136_31+m137_31+m138_31+m139_31+m140_31+m141_31+m142_31+m143_31+m144_31+m145_31+m146_31+m147_31+m148_31+m149_31+m150_31+m151_31+m152_31+m153_31+m154_31+m155_31+m156_31+m157_31+m158_31+m159_31+m160_31+m161_31+m162_31+m163_31+m164_31+m165_31+m166_31+m167_31+m168_31+m169_31+m170_31+m171_31+m172_31+m173_31+m174_31+m175_31+m176_31+m177_31+m178_31+m179_31+m180_31+m181_31+m182_31+m183_31+m184_31+m185_31+m186_31+m187_31+m188_31+m189_31+m190_31+m191_31+m192_31+m193_31+m194_31+m195_31+m196_31+m197_31+m198_31+m199_31+m200_31+m201_31+m202_31+m203_31+m204_31+m205_31+m206_31+m207_31+m208_31+m209_31+m210_31+m211_31+m212_31+m213_31+m214_31+m215_31+m216_31+m217_31+m218_31+m219_31+m220_31+m221_31+m222_31+m223_31+m224_31+m225_31+m226_31+m227_31+m228_31+m229_31+m230_31+m231_31+m232_31+m233_31+m234_31+m235_31+m236_31+m237_31+m238_31+m239_31+m240_31+m241_31+m242_31+m243_31+m244_31+m245_31+m246_31+m247_31+m248_31+m249_31+m250_31+m251_31+m252_31+m253_31+m254_31+m255_31+m256_31+m257_31+m258_31+m259_31+m260_31+m261_31+m262_31+m263_31+m264_31+m265_31+m266_31+m267_31+m268_31+m269_31+m270_31+m271_31+m272_31+m273_31+m274_31+m275_31+m276_31+m277_31+m278_31+m279_31+m280_31+m281_31+m282_31+m283_31+m284_31+m285_31+m286_31+m287_31+m288_31+m289_31+m290_31+m291_31+m292_31+m293_31+m294_31+m295_31+m296_31+m297_31+m298_31+m299_31+m300_31+m301_31+m302_31+m303_31+m304_31+m305_31+m306_31+m307_31+m308_31+m309_31+m310_31+m311_31+m312_31+m313_31+m314_31+m315_31+m316_31+m317_31+m318_31+m319_31+m320_31+m321_31+m322_31+m323_31+m324_31+m325_31+m326_31+m327_31+m328_31+m329_31+m330_31+m331_31+m332_31+m333_31+m334_31+m335_31+m336_31+m337_31+m338_31+m339_31+m340_31+m341_31+m342_31+m343_31+m344_31+m345_31+m346_31+m347_31+m348_31+m349_31+m350_31+m351_31+m352_31+m353_31+m354_31+m355_31+m356_31+m357_31+m358_31+m359_31+m360_31+m361_31+m362_31+m363_31+m364_31+m365_31+m366_31+m367_31+m368_31+m369_31+m370_31+m371_31+m372_31+m373_31+m374_31+m375_31+m376_31+m377_31+m378_31+m379_31+m380_31+m381_31+b31;
   always @(posedge clk) out32 <= m1_32+m2_32+m3_32+m4_32+m5_32+m6_32+m7_32+m8_32+m9_32+m10_32+m11_32+m12_32+m13_32+m14_32+m15_32+m16_32+m17_32+m18_32+m19_32+m20_32+m21_32+m22_32+m23_32+m24_32+m25_32+m26_32+m27_32+m28_32+m29_32+m30_32+m31_32+m32_32+m33_32+m34_32+m35_32+m36_32+m37_32+m38_32+m39_32+m40_32+m41_32+m42_32+m43_32+m44_32+m45_32+m46_32+m47_32+m48_32+m49_32+m50_32+m51_32+m52_32+m53_32+m54_32+m55_32+m56_32+m57_32+m58_32+m59_32+m60_32+m61_32+m62_32+m63_32+m64_32+m65_32+m66_32+m67_32+m68_32+m69_32+m70_32+m71_32+m72_32+m73_32+m74_32+m75_32+m76_32+m77_32+m78_32+m79_32+m80_32+m81_32+m82_32+m83_32+m84_32+m85_32+m86_32+m87_32+m88_32+m89_32+m90_32+m91_32+m92_32+m93_32+m94_32+m95_32+m96_32+m97_32+m98_32+m99_32+m100_32+m101_32+m102_32+m103_32+m104_32+m105_32+m106_32+m107_32+m108_32+m109_32+m110_32+m111_32+m112_32+m113_32+m114_32+m115_32+m116_32+m117_32+m118_32+m119_32+m120_32+m121_32+m122_32+m123_32+m124_32+m125_32+m126_32+m127_32+m128_32+m129_32+m130_32+m131_32+m132_32+m133_32+m134_32+m135_32+m136_32+m137_32+m138_32+m139_32+m140_32+m141_32+m142_32+m143_32+m144_32+m145_32+m146_32+m147_32+m148_32+m149_32+m150_32+m151_32+m152_32+m153_32+m154_32+m155_32+m156_32+m157_32+m158_32+m159_32+m160_32+m161_32+m162_32+m163_32+m164_32+m165_32+m166_32+m167_32+m168_32+m169_32+m170_32+m171_32+m172_32+m173_32+m174_32+m175_32+m176_32+m177_32+m178_32+m179_32+m180_32+m181_32+m182_32+m183_32+m184_32+m185_32+m186_32+m187_32+m188_32+m189_32+m190_32+m191_32+m192_32+m193_32+m194_32+m195_32+m196_32+m197_32+m198_32+m199_32+m200_32+m201_32+m202_32+m203_32+m204_32+m205_32+m206_32+m207_32+m208_32+m209_32+m210_32+m211_32+m212_32+m213_32+m214_32+m215_32+m216_32+m217_32+m218_32+m219_32+m220_32+m221_32+m222_32+m223_32+m224_32+m225_32+m226_32+m227_32+m228_32+m229_32+m230_32+m231_32+m232_32+m233_32+m234_32+m235_32+m236_32+m237_32+m238_32+m239_32+m240_32+m241_32+m242_32+m243_32+m244_32+m245_32+m246_32+m247_32+m248_32+m249_32+m250_32+m251_32+m252_32+m253_32+m254_32+m255_32+m256_32+m257_32+m258_32+m259_32+m260_32+m261_32+m262_32+m263_32+m264_32+m265_32+m266_32+m267_32+m268_32+m269_32+m270_32+m271_32+m272_32+m273_32+m274_32+m275_32+m276_32+m277_32+m278_32+m279_32+m280_32+m281_32+m282_32+m283_32+m284_32+m285_32+m286_32+m287_32+m288_32+m289_32+m290_32+m291_32+m292_32+m293_32+m294_32+m295_32+m296_32+m297_32+m298_32+m299_32+m300_32+m301_32+m302_32+m303_32+m304_32+m305_32+m306_32+m307_32+m308_32+m309_32+m310_32+m311_32+m312_32+m313_32+m314_32+m315_32+m316_32+m317_32+m318_32+m319_32+m320_32+m321_32+m322_32+m323_32+m324_32+m325_32+m326_32+m327_32+m328_32+m329_32+m330_32+m331_32+m332_32+m333_32+m334_32+m335_32+m336_32+m337_32+m338_32+m339_32+m340_32+m341_32+m342_32+m343_32+m344_32+m345_32+m346_32+m347_32+m348_32+m349_32+m350_32+m351_32+m352_32+m353_32+m354_32+m355_32+m356_32+m357_32+m358_32+m359_32+m360_32+m361_32+m362_32+m363_32+m364_32+m365_32+m366_32+m367_32+m368_32+m369_32+m370_32+m371_32+m372_32+m373_32+m374_32+m375_32+m376_32+m377_32+m378_32+m379_32+m380_32+m381_32+b32;
   always @(posedge clk) out33 <= m1_33+m2_33+m3_33+m4_33+m5_33+m6_33+m7_33+m8_33+m9_33+m10_33+m11_33+m12_33+m13_33+m14_33+m15_33+m16_33+m17_33+m18_33+m19_33+m20_33+m21_33+m22_33+m23_33+m24_33+m25_33+m26_33+m27_33+m28_33+m29_33+m30_33+m31_33+m32_33+m33_33+m34_33+m35_33+m36_33+m37_33+m38_33+m39_33+m40_33+m41_33+m42_33+m43_33+m44_33+m45_33+m46_33+m47_33+m48_33+m49_33+m50_33+m51_33+m52_33+m53_33+m54_33+m55_33+m56_33+m57_33+m58_33+m59_33+m60_33+m61_33+m62_33+m63_33+m64_33+m65_33+m66_33+m67_33+m68_33+m69_33+m70_33+m71_33+m72_33+m73_33+m74_33+m75_33+m76_33+m77_33+m78_33+m79_33+m80_33+m81_33+m82_33+m83_33+m84_33+m85_33+m86_33+m87_33+m88_33+m89_33+m90_33+m91_33+m92_33+m93_33+m94_33+m95_33+m96_33+m97_33+m98_33+m99_33+m100_33+m101_33+m102_33+m103_33+m104_33+m105_33+m106_33+m107_33+m108_33+m109_33+m110_33+m111_33+m112_33+m113_33+m114_33+m115_33+m116_33+m117_33+m118_33+m119_33+m120_33+m121_33+m122_33+m123_33+m124_33+m125_33+m126_33+m127_33+m128_33+m129_33+m130_33+m131_33+m132_33+m133_33+m134_33+m135_33+m136_33+m137_33+m138_33+m139_33+m140_33+m141_33+m142_33+m143_33+m144_33+m145_33+m146_33+m147_33+m148_33+m149_33+m150_33+m151_33+m152_33+m153_33+m154_33+m155_33+m156_33+m157_33+m158_33+m159_33+m160_33+m161_33+m162_33+m163_33+m164_33+m165_33+m166_33+m167_33+m168_33+m169_33+m170_33+m171_33+m172_33+m173_33+m174_33+m175_33+m176_33+m177_33+m178_33+m179_33+m180_33+m181_33+m182_33+m183_33+m184_33+m185_33+m186_33+m187_33+m188_33+m189_33+m190_33+m191_33+m192_33+m193_33+m194_33+m195_33+m196_33+m197_33+m198_33+m199_33+m200_33+m201_33+m202_33+m203_33+m204_33+m205_33+m206_33+m207_33+m208_33+m209_33+m210_33+m211_33+m212_33+m213_33+m214_33+m215_33+m216_33+m217_33+m218_33+m219_33+m220_33+m221_33+m222_33+m223_33+m224_33+m225_33+m226_33+m227_33+m228_33+m229_33+m230_33+m231_33+m232_33+m233_33+m234_33+m235_33+m236_33+m237_33+m238_33+m239_33+m240_33+m241_33+m242_33+m243_33+m244_33+m245_33+m246_33+m247_33+m248_33+m249_33+m250_33+m251_33+m252_33+m253_33+m254_33+m255_33+m256_33+m257_33+m258_33+m259_33+m260_33+m261_33+m262_33+m263_33+m264_33+m265_33+m266_33+m267_33+m268_33+m269_33+m270_33+m271_33+m272_33+m273_33+m274_33+m275_33+m276_33+m277_33+m278_33+m279_33+m280_33+m281_33+m282_33+m283_33+m284_33+m285_33+m286_33+m287_33+m288_33+m289_33+m290_33+m291_33+m292_33+m293_33+m294_33+m295_33+m296_33+m297_33+m298_33+m299_33+m300_33+m301_33+m302_33+m303_33+m304_33+m305_33+m306_33+m307_33+m308_33+m309_33+m310_33+m311_33+m312_33+m313_33+m314_33+m315_33+m316_33+m317_33+m318_33+m319_33+m320_33+m321_33+m322_33+m323_33+m324_33+m325_33+m326_33+m327_33+m328_33+m329_33+m330_33+m331_33+m332_33+m333_33+m334_33+m335_33+m336_33+m337_33+m338_33+m339_33+m340_33+m341_33+m342_33+m343_33+m344_33+m345_33+m346_33+m347_33+m348_33+m349_33+m350_33+m351_33+m352_33+m353_33+m354_33+m355_33+m356_33+m357_33+m358_33+m359_33+m360_33+m361_33+m362_33+m363_33+m364_33+m365_33+m366_33+m367_33+m368_33+m369_33+m370_33+m371_33+m372_33+m373_33+m374_33+m375_33+m376_33+m377_33+m378_33+m379_33+m380_33+m381_33+b33;
   always @(posedge clk) out34 <= m1_34+m2_34+m3_34+m4_34+m5_34+m6_34+m7_34+m8_34+m9_34+m10_34+m11_34+m12_34+m13_34+m14_34+m15_34+m16_34+m17_34+m18_34+m19_34+m20_34+m21_34+m22_34+m23_34+m24_34+m25_34+m26_34+m27_34+m28_34+m29_34+m30_34+m31_34+m32_34+m33_34+m34_34+m35_34+m36_34+m37_34+m38_34+m39_34+m40_34+m41_34+m42_34+m43_34+m44_34+m45_34+m46_34+m47_34+m48_34+m49_34+m50_34+m51_34+m52_34+m53_34+m54_34+m55_34+m56_34+m57_34+m58_34+m59_34+m60_34+m61_34+m62_34+m63_34+m64_34+m65_34+m66_34+m67_34+m68_34+m69_34+m70_34+m71_34+m72_34+m73_34+m74_34+m75_34+m76_34+m77_34+m78_34+m79_34+m80_34+m81_34+m82_34+m83_34+m84_34+m85_34+m86_34+m87_34+m88_34+m89_34+m90_34+m91_34+m92_34+m93_34+m94_34+m95_34+m96_34+m97_34+m98_34+m99_34+m100_34+m101_34+m102_34+m103_34+m104_34+m105_34+m106_34+m107_34+m108_34+m109_34+m110_34+m111_34+m112_34+m113_34+m114_34+m115_34+m116_34+m117_34+m118_34+m119_34+m120_34+m121_34+m122_34+m123_34+m124_34+m125_34+m126_34+m127_34+m128_34+m129_34+m130_34+m131_34+m132_34+m133_34+m134_34+m135_34+m136_34+m137_34+m138_34+m139_34+m140_34+m141_34+m142_34+m143_34+m144_34+m145_34+m146_34+m147_34+m148_34+m149_34+m150_34+m151_34+m152_34+m153_34+m154_34+m155_34+m156_34+m157_34+m158_34+m159_34+m160_34+m161_34+m162_34+m163_34+m164_34+m165_34+m166_34+m167_34+m168_34+m169_34+m170_34+m171_34+m172_34+m173_34+m174_34+m175_34+m176_34+m177_34+m178_34+m179_34+m180_34+m181_34+m182_34+m183_34+m184_34+m185_34+m186_34+m187_34+m188_34+m189_34+m190_34+m191_34+m192_34+m193_34+m194_34+m195_34+m196_34+m197_34+m198_34+m199_34+m200_34+m201_34+m202_34+m203_34+m204_34+m205_34+m206_34+m207_34+m208_34+m209_34+m210_34+m211_34+m212_34+m213_34+m214_34+m215_34+m216_34+m217_34+m218_34+m219_34+m220_34+m221_34+m222_34+m223_34+m224_34+m225_34+m226_34+m227_34+m228_34+m229_34+m230_34+m231_34+m232_34+m233_34+m234_34+m235_34+m236_34+m237_34+m238_34+m239_34+m240_34+m241_34+m242_34+m243_34+m244_34+m245_34+m246_34+m247_34+m248_34+m249_34+m250_34+m251_34+m252_34+m253_34+m254_34+m255_34+m256_34+m257_34+m258_34+m259_34+m260_34+m261_34+m262_34+m263_34+m264_34+m265_34+m266_34+m267_34+m268_34+m269_34+m270_34+m271_34+m272_34+m273_34+m274_34+m275_34+m276_34+m277_34+m278_34+m279_34+m280_34+m281_34+m282_34+m283_34+m284_34+m285_34+m286_34+m287_34+m288_34+m289_34+m290_34+m291_34+m292_34+m293_34+m294_34+m295_34+m296_34+m297_34+m298_34+m299_34+m300_34+m301_34+m302_34+m303_34+m304_34+m305_34+m306_34+m307_34+m308_34+m309_34+m310_34+m311_34+m312_34+m313_34+m314_34+m315_34+m316_34+m317_34+m318_34+m319_34+m320_34+m321_34+m322_34+m323_34+m324_34+m325_34+m326_34+m327_34+m328_34+m329_34+m330_34+m331_34+m332_34+m333_34+m334_34+m335_34+m336_34+m337_34+m338_34+m339_34+m340_34+m341_34+m342_34+m343_34+m344_34+m345_34+m346_34+m347_34+m348_34+m349_34+m350_34+m351_34+m352_34+m353_34+m354_34+m355_34+m356_34+m357_34+m358_34+m359_34+m360_34+m361_34+m362_34+m363_34+m364_34+m365_34+m366_34+m367_34+m368_34+m369_34+m370_34+m371_34+m372_34+m373_34+m374_34+m375_34+m376_34+m377_34+m378_34+m379_34+m380_34+m381_34+b34;
   always @(posedge clk) out35 <= m1_35+m2_35+m3_35+m4_35+m5_35+m6_35+m7_35+m8_35+m9_35+m10_35+m11_35+m12_35+m13_35+m14_35+m15_35+m16_35+m17_35+m18_35+m19_35+m20_35+m21_35+m22_35+m23_35+m24_35+m25_35+m26_35+m27_35+m28_35+m29_35+m30_35+m31_35+m32_35+m33_35+m34_35+m35_35+m36_35+m37_35+m38_35+m39_35+m40_35+m41_35+m42_35+m43_35+m44_35+m45_35+m46_35+m47_35+m48_35+m49_35+m50_35+m51_35+m52_35+m53_35+m54_35+m55_35+m56_35+m57_35+m58_35+m59_35+m60_35+m61_35+m62_35+m63_35+m64_35+m65_35+m66_35+m67_35+m68_35+m69_35+m70_35+m71_35+m72_35+m73_35+m74_35+m75_35+m76_35+m77_35+m78_35+m79_35+m80_35+m81_35+m82_35+m83_35+m84_35+m85_35+m86_35+m87_35+m88_35+m89_35+m90_35+m91_35+m92_35+m93_35+m94_35+m95_35+m96_35+m97_35+m98_35+m99_35+m100_35+m101_35+m102_35+m103_35+m104_35+m105_35+m106_35+m107_35+m108_35+m109_35+m110_35+m111_35+m112_35+m113_35+m114_35+m115_35+m116_35+m117_35+m118_35+m119_35+m120_35+m121_35+m122_35+m123_35+m124_35+m125_35+m126_35+m127_35+m128_35+m129_35+m130_35+m131_35+m132_35+m133_35+m134_35+m135_35+m136_35+m137_35+m138_35+m139_35+m140_35+m141_35+m142_35+m143_35+m144_35+m145_35+m146_35+m147_35+m148_35+m149_35+m150_35+m151_35+m152_35+m153_35+m154_35+m155_35+m156_35+m157_35+m158_35+m159_35+m160_35+m161_35+m162_35+m163_35+m164_35+m165_35+m166_35+m167_35+m168_35+m169_35+m170_35+m171_35+m172_35+m173_35+m174_35+m175_35+m176_35+m177_35+m178_35+m179_35+m180_35+m181_35+m182_35+m183_35+m184_35+m185_35+m186_35+m187_35+m188_35+m189_35+m190_35+m191_35+m192_35+m193_35+m194_35+m195_35+m196_35+m197_35+m198_35+m199_35+m200_35+m201_35+m202_35+m203_35+m204_35+m205_35+m206_35+m207_35+m208_35+m209_35+m210_35+m211_35+m212_35+m213_35+m214_35+m215_35+m216_35+m217_35+m218_35+m219_35+m220_35+m221_35+m222_35+m223_35+m224_35+m225_35+m226_35+m227_35+m228_35+m229_35+m230_35+m231_35+m232_35+m233_35+m234_35+m235_35+m236_35+m237_35+m238_35+m239_35+m240_35+m241_35+m242_35+m243_35+m244_35+m245_35+m246_35+m247_35+m248_35+m249_35+m250_35+m251_35+m252_35+m253_35+m254_35+m255_35+m256_35+m257_35+m258_35+m259_35+m260_35+m261_35+m262_35+m263_35+m264_35+m265_35+m266_35+m267_35+m268_35+m269_35+m270_35+m271_35+m272_35+m273_35+m274_35+m275_35+m276_35+m277_35+m278_35+m279_35+m280_35+m281_35+m282_35+m283_35+m284_35+m285_35+m286_35+m287_35+m288_35+m289_35+m290_35+m291_35+m292_35+m293_35+m294_35+m295_35+m296_35+m297_35+m298_35+m299_35+m300_35+m301_35+m302_35+m303_35+m304_35+m305_35+m306_35+m307_35+m308_35+m309_35+m310_35+m311_35+m312_35+m313_35+m314_35+m315_35+m316_35+m317_35+m318_35+m319_35+m320_35+m321_35+m322_35+m323_35+m324_35+m325_35+m326_35+m327_35+m328_35+m329_35+m330_35+m331_35+m332_35+m333_35+m334_35+m335_35+m336_35+m337_35+m338_35+m339_35+m340_35+m341_35+m342_35+m343_35+m344_35+m345_35+m346_35+m347_35+m348_35+m349_35+m350_35+m351_35+m352_35+m353_35+m354_35+m355_35+m356_35+m357_35+m358_35+m359_35+m360_35+m361_35+m362_35+m363_35+m364_35+m365_35+m366_35+m367_35+m368_35+m369_35+m370_35+m371_35+m372_35+m373_35+m374_35+m375_35+m376_35+m377_35+m378_35+m379_35+m380_35+m381_35+b35;
   always @(posedge clk) out36 <= m1_36+m2_36+m3_36+m4_36+m5_36+m6_36+m7_36+m8_36+m9_36+m10_36+m11_36+m12_36+m13_36+m14_36+m15_36+m16_36+m17_36+m18_36+m19_36+m20_36+m21_36+m22_36+m23_36+m24_36+m25_36+m26_36+m27_36+m28_36+m29_36+m30_36+m31_36+m32_36+m33_36+m34_36+m35_36+m36_36+m37_36+m38_36+m39_36+m40_36+m41_36+m42_36+m43_36+m44_36+m45_36+m46_36+m47_36+m48_36+m49_36+m50_36+m51_36+m52_36+m53_36+m54_36+m55_36+m56_36+m57_36+m58_36+m59_36+m60_36+m61_36+m62_36+m63_36+m64_36+m65_36+m66_36+m67_36+m68_36+m69_36+m70_36+m71_36+m72_36+m73_36+m74_36+m75_36+m76_36+m77_36+m78_36+m79_36+m80_36+m81_36+m82_36+m83_36+m84_36+m85_36+m86_36+m87_36+m88_36+m89_36+m90_36+m91_36+m92_36+m93_36+m94_36+m95_36+m96_36+m97_36+m98_36+m99_36+m100_36+m101_36+m102_36+m103_36+m104_36+m105_36+m106_36+m107_36+m108_36+m109_36+m110_36+m111_36+m112_36+m113_36+m114_36+m115_36+m116_36+m117_36+m118_36+m119_36+m120_36+m121_36+m122_36+m123_36+m124_36+m125_36+m126_36+m127_36+m128_36+m129_36+m130_36+m131_36+m132_36+m133_36+m134_36+m135_36+m136_36+m137_36+m138_36+m139_36+m140_36+m141_36+m142_36+m143_36+m144_36+m145_36+m146_36+m147_36+m148_36+m149_36+m150_36+m151_36+m152_36+m153_36+m154_36+m155_36+m156_36+m157_36+m158_36+m159_36+m160_36+m161_36+m162_36+m163_36+m164_36+m165_36+m166_36+m167_36+m168_36+m169_36+m170_36+m171_36+m172_36+m173_36+m174_36+m175_36+m176_36+m177_36+m178_36+m179_36+m180_36+m181_36+m182_36+m183_36+m184_36+m185_36+m186_36+m187_36+m188_36+m189_36+m190_36+m191_36+m192_36+m193_36+m194_36+m195_36+m196_36+m197_36+m198_36+m199_36+m200_36+m201_36+m202_36+m203_36+m204_36+m205_36+m206_36+m207_36+m208_36+m209_36+m210_36+m211_36+m212_36+m213_36+m214_36+m215_36+m216_36+m217_36+m218_36+m219_36+m220_36+m221_36+m222_36+m223_36+m224_36+m225_36+m226_36+m227_36+m228_36+m229_36+m230_36+m231_36+m232_36+m233_36+m234_36+m235_36+m236_36+m237_36+m238_36+m239_36+m240_36+m241_36+m242_36+m243_36+m244_36+m245_36+m246_36+m247_36+m248_36+m249_36+m250_36+m251_36+m252_36+m253_36+m254_36+m255_36+m256_36+m257_36+m258_36+m259_36+m260_36+m261_36+m262_36+m263_36+m264_36+m265_36+m266_36+m267_36+m268_36+m269_36+m270_36+m271_36+m272_36+m273_36+m274_36+m275_36+m276_36+m277_36+m278_36+m279_36+m280_36+m281_36+m282_36+m283_36+m284_36+m285_36+m286_36+m287_36+m288_36+m289_36+m290_36+m291_36+m292_36+m293_36+m294_36+m295_36+m296_36+m297_36+m298_36+m299_36+m300_36+m301_36+m302_36+m303_36+m304_36+m305_36+m306_36+m307_36+m308_36+m309_36+m310_36+m311_36+m312_36+m313_36+m314_36+m315_36+m316_36+m317_36+m318_36+m319_36+m320_36+m321_36+m322_36+m323_36+m324_36+m325_36+m326_36+m327_36+m328_36+m329_36+m330_36+m331_36+m332_36+m333_36+m334_36+m335_36+m336_36+m337_36+m338_36+m339_36+m340_36+m341_36+m342_36+m343_36+m344_36+m345_36+m346_36+m347_36+m348_36+m349_36+m350_36+m351_36+m352_36+m353_36+m354_36+m355_36+m356_36+m357_36+m358_36+m359_36+m360_36+m361_36+m362_36+m363_36+m364_36+m365_36+m366_36+m367_36+m368_36+m369_36+m370_36+m371_36+m372_36+m373_36+m374_36+m375_36+m376_36+m377_36+m378_36+m379_36+m380_36+m381_36+b36;
   always @(posedge clk) out37 <= m1_37+m2_37+m3_37+m4_37+m5_37+m6_37+m7_37+m8_37+m9_37+m10_37+m11_37+m12_37+m13_37+m14_37+m15_37+m16_37+m17_37+m18_37+m19_37+m20_37+m21_37+m22_37+m23_37+m24_37+m25_37+m26_37+m27_37+m28_37+m29_37+m30_37+m31_37+m32_37+m33_37+m34_37+m35_37+m36_37+m37_37+m38_37+m39_37+m40_37+m41_37+m42_37+m43_37+m44_37+m45_37+m46_37+m47_37+m48_37+m49_37+m50_37+m51_37+m52_37+m53_37+m54_37+m55_37+m56_37+m57_37+m58_37+m59_37+m60_37+m61_37+m62_37+m63_37+m64_37+m65_37+m66_37+m67_37+m68_37+m69_37+m70_37+m71_37+m72_37+m73_37+m74_37+m75_37+m76_37+m77_37+m78_37+m79_37+m80_37+m81_37+m82_37+m83_37+m84_37+m85_37+m86_37+m87_37+m88_37+m89_37+m90_37+m91_37+m92_37+m93_37+m94_37+m95_37+m96_37+m97_37+m98_37+m99_37+m100_37+m101_37+m102_37+m103_37+m104_37+m105_37+m106_37+m107_37+m108_37+m109_37+m110_37+m111_37+m112_37+m113_37+m114_37+m115_37+m116_37+m117_37+m118_37+m119_37+m120_37+m121_37+m122_37+m123_37+m124_37+m125_37+m126_37+m127_37+m128_37+m129_37+m130_37+m131_37+m132_37+m133_37+m134_37+m135_37+m136_37+m137_37+m138_37+m139_37+m140_37+m141_37+m142_37+m143_37+m144_37+m145_37+m146_37+m147_37+m148_37+m149_37+m150_37+m151_37+m152_37+m153_37+m154_37+m155_37+m156_37+m157_37+m158_37+m159_37+m160_37+m161_37+m162_37+m163_37+m164_37+m165_37+m166_37+m167_37+m168_37+m169_37+m170_37+m171_37+m172_37+m173_37+m174_37+m175_37+m176_37+m177_37+m178_37+m179_37+m180_37+m181_37+m182_37+m183_37+m184_37+m185_37+m186_37+m187_37+m188_37+m189_37+m190_37+m191_37+m192_37+m193_37+m194_37+m195_37+m196_37+m197_37+m198_37+m199_37+m200_37+m201_37+m202_37+m203_37+m204_37+m205_37+m206_37+m207_37+m208_37+m209_37+m210_37+m211_37+m212_37+m213_37+m214_37+m215_37+m216_37+m217_37+m218_37+m219_37+m220_37+m221_37+m222_37+m223_37+m224_37+m225_37+m226_37+m227_37+m228_37+m229_37+m230_37+m231_37+m232_37+m233_37+m234_37+m235_37+m236_37+m237_37+m238_37+m239_37+m240_37+m241_37+m242_37+m243_37+m244_37+m245_37+m246_37+m247_37+m248_37+m249_37+m250_37+m251_37+m252_37+m253_37+m254_37+m255_37+m256_37+m257_37+m258_37+m259_37+m260_37+m261_37+m262_37+m263_37+m264_37+m265_37+m266_37+m267_37+m268_37+m269_37+m270_37+m271_37+m272_37+m273_37+m274_37+m275_37+m276_37+m277_37+m278_37+m279_37+m280_37+m281_37+m282_37+m283_37+m284_37+m285_37+m286_37+m287_37+m288_37+m289_37+m290_37+m291_37+m292_37+m293_37+m294_37+m295_37+m296_37+m297_37+m298_37+m299_37+m300_37+m301_37+m302_37+m303_37+m304_37+m305_37+m306_37+m307_37+m308_37+m309_37+m310_37+m311_37+m312_37+m313_37+m314_37+m315_37+m316_37+m317_37+m318_37+m319_37+m320_37+m321_37+m322_37+m323_37+m324_37+m325_37+m326_37+m327_37+m328_37+m329_37+m330_37+m331_37+m332_37+m333_37+m334_37+m335_37+m336_37+m337_37+m338_37+m339_37+m340_37+m341_37+m342_37+m343_37+m344_37+m345_37+m346_37+m347_37+m348_37+m349_37+m350_37+m351_37+m352_37+m353_37+m354_37+m355_37+m356_37+m357_37+m358_37+m359_37+m360_37+m361_37+m362_37+m363_37+m364_37+m365_37+m366_37+m367_37+m368_37+m369_37+m370_37+m371_37+m372_37+m373_37+m374_37+m375_37+m376_37+m377_37+m378_37+m379_37+m380_37+m381_37+b37;
   always @(posedge clk) out38 <= m1_38+m2_38+m3_38+m4_38+m5_38+m6_38+m7_38+m8_38+m9_38+m10_38+m11_38+m12_38+m13_38+m14_38+m15_38+m16_38+m17_38+m18_38+m19_38+m20_38+m21_38+m22_38+m23_38+m24_38+m25_38+m26_38+m27_38+m28_38+m29_38+m30_38+m31_38+m32_38+m33_38+m34_38+m35_38+m36_38+m37_38+m38_38+m39_38+m40_38+m41_38+m42_38+m43_38+m44_38+m45_38+m46_38+m47_38+m48_38+m49_38+m50_38+m51_38+m52_38+m53_38+m54_38+m55_38+m56_38+m57_38+m58_38+m59_38+m60_38+m61_38+m62_38+m63_38+m64_38+m65_38+m66_38+m67_38+m68_38+m69_38+m70_38+m71_38+m72_38+m73_38+m74_38+m75_38+m76_38+m77_38+m78_38+m79_38+m80_38+m81_38+m82_38+m83_38+m84_38+m85_38+m86_38+m87_38+m88_38+m89_38+m90_38+m91_38+m92_38+m93_38+m94_38+m95_38+m96_38+m97_38+m98_38+m99_38+m100_38+m101_38+m102_38+m103_38+m104_38+m105_38+m106_38+m107_38+m108_38+m109_38+m110_38+m111_38+m112_38+m113_38+m114_38+m115_38+m116_38+m117_38+m118_38+m119_38+m120_38+m121_38+m122_38+m123_38+m124_38+m125_38+m126_38+m127_38+m128_38+m129_38+m130_38+m131_38+m132_38+m133_38+m134_38+m135_38+m136_38+m137_38+m138_38+m139_38+m140_38+m141_38+m142_38+m143_38+m144_38+m145_38+m146_38+m147_38+m148_38+m149_38+m150_38+m151_38+m152_38+m153_38+m154_38+m155_38+m156_38+m157_38+m158_38+m159_38+m160_38+m161_38+m162_38+m163_38+m164_38+m165_38+m166_38+m167_38+m168_38+m169_38+m170_38+m171_38+m172_38+m173_38+m174_38+m175_38+m176_38+m177_38+m178_38+m179_38+m180_38+m181_38+m182_38+m183_38+m184_38+m185_38+m186_38+m187_38+m188_38+m189_38+m190_38+m191_38+m192_38+m193_38+m194_38+m195_38+m196_38+m197_38+m198_38+m199_38+m200_38+m201_38+m202_38+m203_38+m204_38+m205_38+m206_38+m207_38+m208_38+m209_38+m210_38+m211_38+m212_38+m213_38+m214_38+m215_38+m216_38+m217_38+m218_38+m219_38+m220_38+m221_38+m222_38+m223_38+m224_38+m225_38+m226_38+m227_38+m228_38+m229_38+m230_38+m231_38+m232_38+m233_38+m234_38+m235_38+m236_38+m237_38+m238_38+m239_38+m240_38+m241_38+m242_38+m243_38+m244_38+m245_38+m246_38+m247_38+m248_38+m249_38+m250_38+m251_38+m252_38+m253_38+m254_38+m255_38+m256_38+m257_38+m258_38+m259_38+m260_38+m261_38+m262_38+m263_38+m264_38+m265_38+m266_38+m267_38+m268_38+m269_38+m270_38+m271_38+m272_38+m273_38+m274_38+m275_38+m276_38+m277_38+m278_38+m279_38+m280_38+m281_38+m282_38+m283_38+m284_38+m285_38+m286_38+m287_38+m288_38+m289_38+m290_38+m291_38+m292_38+m293_38+m294_38+m295_38+m296_38+m297_38+m298_38+m299_38+m300_38+m301_38+m302_38+m303_38+m304_38+m305_38+m306_38+m307_38+m308_38+m309_38+m310_38+m311_38+m312_38+m313_38+m314_38+m315_38+m316_38+m317_38+m318_38+m319_38+m320_38+m321_38+m322_38+m323_38+m324_38+m325_38+m326_38+m327_38+m328_38+m329_38+m330_38+m331_38+m332_38+m333_38+m334_38+m335_38+m336_38+m337_38+m338_38+m339_38+m340_38+m341_38+m342_38+m343_38+m344_38+m345_38+m346_38+m347_38+m348_38+m349_38+m350_38+m351_38+m352_38+m353_38+m354_38+m355_38+m356_38+m357_38+m358_38+m359_38+m360_38+m361_38+m362_38+m363_38+m364_38+m365_38+m366_38+m367_38+m368_38+m369_38+m370_38+m371_38+m372_38+m373_38+m374_38+m375_38+m376_38+m377_38+m378_38+m379_38+m380_38+m381_38+b38;
   always @(posedge clk) out39 <= m1_39+m2_39+m3_39+m4_39+m5_39+m6_39+m7_39+m8_39+m9_39+m10_39+m11_39+m12_39+m13_39+m14_39+m15_39+m16_39+m17_39+m18_39+m19_39+m20_39+m21_39+m22_39+m23_39+m24_39+m25_39+m26_39+m27_39+m28_39+m29_39+m30_39+m31_39+m32_39+m33_39+m34_39+m35_39+m36_39+m37_39+m38_39+m39_39+m40_39+m41_39+m42_39+m43_39+m44_39+m45_39+m46_39+m47_39+m48_39+m49_39+m50_39+m51_39+m52_39+m53_39+m54_39+m55_39+m56_39+m57_39+m58_39+m59_39+m60_39+m61_39+m62_39+m63_39+m64_39+m65_39+m66_39+m67_39+m68_39+m69_39+m70_39+m71_39+m72_39+m73_39+m74_39+m75_39+m76_39+m77_39+m78_39+m79_39+m80_39+m81_39+m82_39+m83_39+m84_39+m85_39+m86_39+m87_39+m88_39+m89_39+m90_39+m91_39+m92_39+m93_39+m94_39+m95_39+m96_39+m97_39+m98_39+m99_39+m100_39+m101_39+m102_39+m103_39+m104_39+m105_39+m106_39+m107_39+m108_39+m109_39+m110_39+m111_39+m112_39+m113_39+m114_39+m115_39+m116_39+m117_39+m118_39+m119_39+m120_39+m121_39+m122_39+m123_39+m124_39+m125_39+m126_39+m127_39+m128_39+m129_39+m130_39+m131_39+m132_39+m133_39+m134_39+m135_39+m136_39+m137_39+m138_39+m139_39+m140_39+m141_39+m142_39+m143_39+m144_39+m145_39+m146_39+m147_39+m148_39+m149_39+m150_39+m151_39+m152_39+m153_39+m154_39+m155_39+m156_39+m157_39+m158_39+m159_39+m160_39+m161_39+m162_39+m163_39+m164_39+m165_39+m166_39+m167_39+m168_39+m169_39+m170_39+m171_39+m172_39+m173_39+m174_39+m175_39+m176_39+m177_39+m178_39+m179_39+m180_39+m181_39+m182_39+m183_39+m184_39+m185_39+m186_39+m187_39+m188_39+m189_39+m190_39+m191_39+m192_39+m193_39+m194_39+m195_39+m196_39+m197_39+m198_39+m199_39+m200_39+m201_39+m202_39+m203_39+m204_39+m205_39+m206_39+m207_39+m208_39+m209_39+m210_39+m211_39+m212_39+m213_39+m214_39+m215_39+m216_39+m217_39+m218_39+m219_39+m220_39+m221_39+m222_39+m223_39+m224_39+m225_39+m226_39+m227_39+m228_39+m229_39+m230_39+m231_39+m232_39+m233_39+m234_39+m235_39+m236_39+m237_39+m238_39+m239_39+m240_39+m241_39+m242_39+m243_39+m244_39+m245_39+m246_39+m247_39+m248_39+m249_39+m250_39+m251_39+m252_39+m253_39+m254_39+m255_39+m256_39+m257_39+m258_39+m259_39+m260_39+m261_39+m262_39+m263_39+m264_39+m265_39+m266_39+m267_39+m268_39+m269_39+m270_39+m271_39+m272_39+m273_39+m274_39+m275_39+m276_39+m277_39+m278_39+m279_39+m280_39+m281_39+m282_39+m283_39+m284_39+m285_39+m286_39+m287_39+m288_39+m289_39+m290_39+m291_39+m292_39+m293_39+m294_39+m295_39+m296_39+m297_39+m298_39+m299_39+m300_39+m301_39+m302_39+m303_39+m304_39+m305_39+m306_39+m307_39+m308_39+m309_39+m310_39+m311_39+m312_39+m313_39+m314_39+m315_39+m316_39+m317_39+m318_39+m319_39+m320_39+m321_39+m322_39+m323_39+m324_39+m325_39+m326_39+m327_39+m328_39+m329_39+m330_39+m331_39+m332_39+m333_39+m334_39+m335_39+m336_39+m337_39+m338_39+m339_39+m340_39+m341_39+m342_39+m343_39+m344_39+m345_39+m346_39+m347_39+m348_39+m349_39+m350_39+m351_39+m352_39+m353_39+m354_39+m355_39+m356_39+m357_39+m358_39+m359_39+m360_39+m361_39+m362_39+m363_39+m364_39+m365_39+m366_39+m367_39+m368_39+m369_39+m370_39+m371_39+m372_39+m373_39+m374_39+m375_39+m376_39+m377_39+m378_39+m379_39+m380_39+m381_39+b39;
   always @(posedge clk) out40 <= m1_40+m2_40+m3_40+m4_40+m5_40+m6_40+m7_40+m8_40+m9_40+m10_40+m11_40+m12_40+m13_40+m14_40+m15_40+m16_40+m17_40+m18_40+m19_40+m20_40+m21_40+m22_40+m23_40+m24_40+m25_40+m26_40+m27_40+m28_40+m29_40+m30_40+m31_40+m32_40+m33_40+m34_40+m35_40+m36_40+m37_40+m38_40+m39_40+m40_40+m41_40+m42_40+m43_40+m44_40+m45_40+m46_40+m47_40+m48_40+m49_40+m50_40+m51_40+m52_40+m53_40+m54_40+m55_40+m56_40+m57_40+m58_40+m59_40+m60_40+m61_40+m62_40+m63_40+m64_40+m65_40+m66_40+m67_40+m68_40+m69_40+m70_40+m71_40+m72_40+m73_40+m74_40+m75_40+m76_40+m77_40+m78_40+m79_40+m80_40+m81_40+m82_40+m83_40+m84_40+m85_40+m86_40+m87_40+m88_40+m89_40+m90_40+m91_40+m92_40+m93_40+m94_40+m95_40+m96_40+m97_40+m98_40+m99_40+m100_40+m101_40+m102_40+m103_40+m104_40+m105_40+m106_40+m107_40+m108_40+m109_40+m110_40+m111_40+m112_40+m113_40+m114_40+m115_40+m116_40+m117_40+m118_40+m119_40+m120_40+m121_40+m122_40+m123_40+m124_40+m125_40+m126_40+m127_40+m128_40+m129_40+m130_40+m131_40+m132_40+m133_40+m134_40+m135_40+m136_40+m137_40+m138_40+m139_40+m140_40+m141_40+m142_40+m143_40+m144_40+m145_40+m146_40+m147_40+m148_40+m149_40+m150_40+m151_40+m152_40+m153_40+m154_40+m155_40+m156_40+m157_40+m158_40+m159_40+m160_40+m161_40+m162_40+m163_40+m164_40+m165_40+m166_40+m167_40+m168_40+m169_40+m170_40+m171_40+m172_40+m173_40+m174_40+m175_40+m176_40+m177_40+m178_40+m179_40+m180_40+m181_40+m182_40+m183_40+m184_40+m185_40+m186_40+m187_40+m188_40+m189_40+m190_40+m191_40+m192_40+m193_40+m194_40+m195_40+m196_40+m197_40+m198_40+m199_40+m200_40+m201_40+m202_40+m203_40+m204_40+m205_40+m206_40+m207_40+m208_40+m209_40+m210_40+m211_40+m212_40+m213_40+m214_40+m215_40+m216_40+m217_40+m218_40+m219_40+m220_40+m221_40+m222_40+m223_40+m224_40+m225_40+m226_40+m227_40+m228_40+m229_40+m230_40+m231_40+m232_40+m233_40+m234_40+m235_40+m236_40+m237_40+m238_40+m239_40+m240_40+m241_40+m242_40+m243_40+m244_40+m245_40+m246_40+m247_40+m248_40+m249_40+m250_40+m251_40+m252_40+m253_40+m254_40+m255_40+m256_40+m257_40+m258_40+m259_40+m260_40+m261_40+m262_40+m263_40+m264_40+m265_40+m266_40+m267_40+m268_40+m269_40+m270_40+m271_40+m272_40+m273_40+m274_40+m275_40+m276_40+m277_40+m278_40+m279_40+m280_40+m281_40+m282_40+m283_40+m284_40+m285_40+m286_40+m287_40+m288_40+m289_40+m290_40+m291_40+m292_40+m293_40+m294_40+m295_40+m296_40+m297_40+m298_40+m299_40+m300_40+m301_40+m302_40+m303_40+m304_40+m305_40+m306_40+m307_40+m308_40+m309_40+m310_40+m311_40+m312_40+m313_40+m314_40+m315_40+m316_40+m317_40+m318_40+m319_40+m320_40+m321_40+m322_40+m323_40+m324_40+m325_40+m326_40+m327_40+m328_40+m329_40+m330_40+m331_40+m332_40+m333_40+m334_40+m335_40+m336_40+m337_40+m338_40+m339_40+m340_40+m341_40+m342_40+m343_40+m344_40+m345_40+m346_40+m347_40+m348_40+m349_40+m350_40+m351_40+m352_40+m353_40+m354_40+m355_40+m356_40+m357_40+m358_40+m359_40+m360_40+m361_40+m362_40+m363_40+m364_40+m365_40+m366_40+m367_40+m368_40+m369_40+m370_40+m371_40+m372_40+m373_40+m374_40+m375_40+m376_40+m377_40+m378_40+m379_40+m380_40+m381_40+b40;
   always @(posedge clk) out41 <= m1_41+m2_41+m3_41+m4_41+m5_41+m6_41+m7_41+m8_41+m9_41+m10_41+m11_41+m12_41+m13_41+m14_41+m15_41+m16_41+m17_41+m18_41+m19_41+m20_41+m21_41+m22_41+m23_41+m24_41+m25_41+m26_41+m27_41+m28_41+m29_41+m30_41+m31_41+m32_41+m33_41+m34_41+m35_41+m36_41+m37_41+m38_41+m39_41+m40_41+m41_41+m42_41+m43_41+m44_41+m45_41+m46_41+m47_41+m48_41+m49_41+m50_41+m51_41+m52_41+m53_41+m54_41+m55_41+m56_41+m57_41+m58_41+m59_41+m60_41+m61_41+m62_41+m63_41+m64_41+m65_41+m66_41+m67_41+m68_41+m69_41+m70_41+m71_41+m72_41+m73_41+m74_41+m75_41+m76_41+m77_41+m78_41+m79_41+m80_41+m81_41+m82_41+m83_41+m84_41+m85_41+m86_41+m87_41+m88_41+m89_41+m90_41+m91_41+m92_41+m93_41+m94_41+m95_41+m96_41+m97_41+m98_41+m99_41+m100_41+m101_41+m102_41+m103_41+m104_41+m105_41+m106_41+m107_41+m108_41+m109_41+m110_41+m111_41+m112_41+m113_41+m114_41+m115_41+m116_41+m117_41+m118_41+m119_41+m120_41+m121_41+m122_41+m123_41+m124_41+m125_41+m126_41+m127_41+m128_41+m129_41+m130_41+m131_41+m132_41+m133_41+m134_41+m135_41+m136_41+m137_41+m138_41+m139_41+m140_41+m141_41+m142_41+m143_41+m144_41+m145_41+m146_41+m147_41+m148_41+m149_41+m150_41+m151_41+m152_41+m153_41+m154_41+m155_41+m156_41+m157_41+m158_41+m159_41+m160_41+m161_41+m162_41+m163_41+m164_41+m165_41+m166_41+m167_41+m168_41+m169_41+m170_41+m171_41+m172_41+m173_41+m174_41+m175_41+m176_41+m177_41+m178_41+m179_41+m180_41+m181_41+m182_41+m183_41+m184_41+m185_41+m186_41+m187_41+m188_41+m189_41+m190_41+m191_41+m192_41+m193_41+m194_41+m195_41+m196_41+m197_41+m198_41+m199_41+m200_41+m201_41+m202_41+m203_41+m204_41+m205_41+m206_41+m207_41+m208_41+m209_41+m210_41+m211_41+m212_41+m213_41+m214_41+m215_41+m216_41+m217_41+m218_41+m219_41+m220_41+m221_41+m222_41+m223_41+m224_41+m225_41+m226_41+m227_41+m228_41+m229_41+m230_41+m231_41+m232_41+m233_41+m234_41+m235_41+m236_41+m237_41+m238_41+m239_41+m240_41+m241_41+m242_41+m243_41+m244_41+m245_41+m246_41+m247_41+m248_41+m249_41+m250_41+m251_41+m252_41+m253_41+m254_41+m255_41+m256_41+m257_41+m258_41+m259_41+m260_41+m261_41+m262_41+m263_41+m264_41+m265_41+m266_41+m267_41+m268_41+m269_41+m270_41+m271_41+m272_41+m273_41+m274_41+m275_41+m276_41+m277_41+m278_41+m279_41+m280_41+m281_41+m282_41+m283_41+m284_41+m285_41+m286_41+m287_41+m288_41+m289_41+m290_41+m291_41+m292_41+m293_41+m294_41+m295_41+m296_41+m297_41+m298_41+m299_41+m300_41+m301_41+m302_41+m303_41+m304_41+m305_41+m306_41+m307_41+m308_41+m309_41+m310_41+m311_41+m312_41+m313_41+m314_41+m315_41+m316_41+m317_41+m318_41+m319_41+m320_41+m321_41+m322_41+m323_41+m324_41+m325_41+m326_41+m327_41+m328_41+m329_41+m330_41+m331_41+m332_41+m333_41+m334_41+m335_41+m336_41+m337_41+m338_41+m339_41+m340_41+m341_41+m342_41+m343_41+m344_41+m345_41+m346_41+m347_41+m348_41+m349_41+m350_41+m351_41+m352_41+m353_41+m354_41+m355_41+m356_41+m357_41+m358_41+m359_41+m360_41+m361_41+m362_41+m363_41+m364_41+m365_41+m366_41+m367_41+m368_41+m369_41+m370_41+m371_41+m372_41+m373_41+m374_41+m375_41+m376_41+m377_41+m378_41+m379_41+m380_41+m381_41+b41;
   always @(posedge clk) out42 <= m1_42+m2_42+m3_42+m4_42+m5_42+m6_42+m7_42+m8_42+m9_42+m10_42+m11_42+m12_42+m13_42+m14_42+m15_42+m16_42+m17_42+m18_42+m19_42+m20_42+m21_42+m22_42+m23_42+m24_42+m25_42+m26_42+m27_42+m28_42+m29_42+m30_42+m31_42+m32_42+m33_42+m34_42+m35_42+m36_42+m37_42+m38_42+m39_42+m40_42+m41_42+m42_42+m43_42+m44_42+m45_42+m46_42+m47_42+m48_42+m49_42+m50_42+m51_42+m52_42+m53_42+m54_42+m55_42+m56_42+m57_42+m58_42+m59_42+m60_42+m61_42+m62_42+m63_42+m64_42+m65_42+m66_42+m67_42+m68_42+m69_42+m70_42+m71_42+m72_42+m73_42+m74_42+m75_42+m76_42+m77_42+m78_42+m79_42+m80_42+m81_42+m82_42+m83_42+m84_42+m85_42+m86_42+m87_42+m88_42+m89_42+m90_42+m91_42+m92_42+m93_42+m94_42+m95_42+m96_42+m97_42+m98_42+m99_42+m100_42+m101_42+m102_42+m103_42+m104_42+m105_42+m106_42+m107_42+m108_42+m109_42+m110_42+m111_42+m112_42+m113_42+m114_42+m115_42+m116_42+m117_42+m118_42+m119_42+m120_42+m121_42+m122_42+m123_42+m124_42+m125_42+m126_42+m127_42+m128_42+m129_42+m130_42+m131_42+m132_42+m133_42+m134_42+m135_42+m136_42+m137_42+m138_42+m139_42+m140_42+m141_42+m142_42+m143_42+m144_42+m145_42+m146_42+m147_42+m148_42+m149_42+m150_42+m151_42+m152_42+m153_42+m154_42+m155_42+m156_42+m157_42+m158_42+m159_42+m160_42+m161_42+m162_42+m163_42+m164_42+m165_42+m166_42+m167_42+m168_42+m169_42+m170_42+m171_42+m172_42+m173_42+m174_42+m175_42+m176_42+m177_42+m178_42+m179_42+m180_42+m181_42+m182_42+m183_42+m184_42+m185_42+m186_42+m187_42+m188_42+m189_42+m190_42+m191_42+m192_42+m193_42+m194_42+m195_42+m196_42+m197_42+m198_42+m199_42+m200_42+m201_42+m202_42+m203_42+m204_42+m205_42+m206_42+m207_42+m208_42+m209_42+m210_42+m211_42+m212_42+m213_42+m214_42+m215_42+m216_42+m217_42+m218_42+m219_42+m220_42+m221_42+m222_42+m223_42+m224_42+m225_42+m226_42+m227_42+m228_42+m229_42+m230_42+m231_42+m232_42+m233_42+m234_42+m235_42+m236_42+m237_42+m238_42+m239_42+m240_42+m241_42+m242_42+m243_42+m244_42+m245_42+m246_42+m247_42+m248_42+m249_42+m250_42+m251_42+m252_42+m253_42+m254_42+m255_42+m256_42+m257_42+m258_42+m259_42+m260_42+m261_42+m262_42+m263_42+m264_42+m265_42+m266_42+m267_42+m268_42+m269_42+m270_42+m271_42+m272_42+m273_42+m274_42+m275_42+m276_42+m277_42+m278_42+m279_42+m280_42+m281_42+m282_42+m283_42+m284_42+m285_42+m286_42+m287_42+m288_42+m289_42+m290_42+m291_42+m292_42+m293_42+m294_42+m295_42+m296_42+m297_42+m298_42+m299_42+m300_42+m301_42+m302_42+m303_42+m304_42+m305_42+m306_42+m307_42+m308_42+m309_42+m310_42+m311_42+m312_42+m313_42+m314_42+m315_42+m316_42+m317_42+m318_42+m319_42+m320_42+m321_42+m322_42+m323_42+m324_42+m325_42+m326_42+m327_42+m328_42+m329_42+m330_42+m331_42+m332_42+m333_42+m334_42+m335_42+m336_42+m337_42+m338_42+m339_42+m340_42+m341_42+m342_42+m343_42+m344_42+m345_42+m346_42+m347_42+m348_42+m349_42+m350_42+m351_42+m352_42+m353_42+m354_42+m355_42+m356_42+m357_42+m358_42+m359_42+m360_42+m361_42+m362_42+m363_42+m364_42+m365_42+m366_42+m367_42+m368_42+m369_42+m370_42+m371_42+m372_42+m373_42+m374_42+m375_42+m376_42+m377_42+m378_42+m379_42+m380_42+m381_42+b42;
   always @(posedge clk) out43 <= m1_43+m2_43+m3_43+m4_43+m5_43+m6_43+m7_43+m8_43+m9_43+m10_43+m11_43+m12_43+m13_43+m14_43+m15_43+m16_43+m17_43+m18_43+m19_43+m20_43+m21_43+m22_43+m23_43+m24_43+m25_43+m26_43+m27_43+m28_43+m29_43+m30_43+m31_43+m32_43+m33_43+m34_43+m35_43+m36_43+m37_43+m38_43+m39_43+m40_43+m41_43+m42_43+m43_43+m44_43+m45_43+m46_43+m47_43+m48_43+m49_43+m50_43+m51_43+m52_43+m53_43+m54_43+m55_43+m56_43+m57_43+m58_43+m59_43+m60_43+m61_43+m62_43+m63_43+m64_43+m65_43+m66_43+m67_43+m68_43+m69_43+m70_43+m71_43+m72_43+m73_43+m74_43+m75_43+m76_43+m77_43+m78_43+m79_43+m80_43+m81_43+m82_43+m83_43+m84_43+m85_43+m86_43+m87_43+m88_43+m89_43+m90_43+m91_43+m92_43+m93_43+m94_43+m95_43+m96_43+m97_43+m98_43+m99_43+m100_43+m101_43+m102_43+m103_43+m104_43+m105_43+m106_43+m107_43+m108_43+m109_43+m110_43+m111_43+m112_43+m113_43+m114_43+m115_43+m116_43+m117_43+m118_43+m119_43+m120_43+m121_43+m122_43+m123_43+m124_43+m125_43+m126_43+m127_43+m128_43+m129_43+m130_43+m131_43+m132_43+m133_43+m134_43+m135_43+m136_43+m137_43+m138_43+m139_43+m140_43+m141_43+m142_43+m143_43+m144_43+m145_43+m146_43+m147_43+m148_43+m149_43+m150_43+m151_43+m152_43+m153_43+m154_43+m155_43+m156_43+m157_43+m158_43+m159_43+m160_43+m161_43+m162_43+m163_43+m164_43+m165_43+m166_43+m167_43+m168_43+m169_43+m170_43+m171_43+m172_43+m173_43+m174_43+m175_43+m176_43+m177_43+m178_43+m179_43+m180_43+m181_43+m182_43+m183_43+m184_43+m185_43+m186_43+m187_43+m188_43+m189_43+m190_43+m191_43+m192_43+m193_43+m194_43+m195_43+m196_43+m197_43+m198_43+m199_43+m200_43+m201_43+m202_43+m203_43+m204_43+m205_43+m206_43+m207_43+m208_43+m209_43+m210_43+m211_43+m212_43+m213_43+m214_43+m215_43+m216_43+m217_43+m218_43+m219_43+m220_43+m221_43+m222_43+m223_43+m224_43+m225_43+m226_43+m227_43+m228_43+m229_43+m230_43+m231_43+m232_43+m233_43+m234_43+m235_43+m236_43+m237_43+m238_43+m239_43+m240_43+m241_43+m242_43+m243_43+m244_43+m245_43+m246_43+m247_43+m248_43+m249_43+m250_43+m251_43+m252_43+m253_43+m254_43+m255_43+m256_43+m257_43+m258_43+m259_43+m260_43+m261_43+m262_43+m263_43+m264_43+m265_43+m266_43+m267_43+m268_43+m269_43+m270_43+m271_43+m272_43+m273_43+m274_43+m275_43+m276_43+m277_43+m278_43+m279_43+m280_43+m281_43+m282_43+m283_43+m284_43+m285_43+m286_43+m287_43+m288_43+m289_43+m290_43+m291_43+m292_43+m293_43+m294_43+m295_43+m296_43+m297_43+m298_43+m299_43+m300_43+m301_43+m302_43+m303_43+m304_43+m305_43+m306_43+m307_43+m308_43+m309_43+m310_43+m311_43+m312_43+m313_43+m314_43+m315_43+m316_43+m317_43+m318_43+m319_43+m320_43+m321_43+m322_43+m323_43+m324_43+m325_43+m326_43+m327_43+m328_43+m329_43+m330_43+m331_43+m332_43+m333_43+m334_43+m335_43+m336_43+m337_43+m338_43+m339_43+m340_43+m341_43+m342_43+m343_43+m344_43+m345_43+m346_43+m347_43+m348_43+m349_43+m350_43+m351_43+m352_43+m353_43+m354_43+m355_43+m356_43+m357_43+m358_43+m359_43+m360_43+m361_43+m362_43+m363_43+m364_43+m365_43+m366_43+m367_43+m368_43+m369_43+m370_43+m371_43+m372_43+m373_43+m374_43+m375_43+m376_43+m377_43+m378_43+m379_43+m380_43+m381_43+b43;
   always @(posedge clk) out44 <= m1_44+m2_44+m3_44+m4_44+m5_44+m6_44+m7_44+m8_44+m9_44+m10_44+m11_44+m12_44+m13_44+m14_44+m15_44+m16_44+m17_44+m18_44+m19_44+m20_44+m21_44+m22_44+m23_44+m24_44+m25_44+m26_44+m27_44+m28_44+m29_44+m30_44+m31_44+m32_44+m33_44+m34_44+m35_44+m36_44+m37_44+m38_44+m39_44+m40_44+m41_44+m42_44+m43_44+m44_44+m45_44+m46_44+m47_44+m48_44+m49_44+m50_44+m51_44+m52_44+m53_44+m54_44+m55_44+m56_44+m57_44+m58_44+m59_44+m60_44+m61_44+m62_44+m63_44+m64_44+m65_44+m66_44+m67_44+m68_44+m69_44+m70_44+m71_44+m72_44+m73_44+m74_44+m75_44+m76_44+m77_44+m78_44+m79_44+m80_44+m81_44+m82_44+m83_44+m84_44+m85_44+m86_44+m87_44+m88_44+m89_44+m90_44+m91_44+m92_44+m93_44+m94_44+m95_44+m96_44+m97_44+m98_44+m99_44+m100_44+m101_44+m102_44+m103_44+m104_44+m105_44+m106_44+m107_44+m108_44+m109_44+m110_44+m111_44+m112_44+m113_44+m114_44+m115_44+m116_44+m117_44+m118_44+m119_44+m120_44+m121_44+m122_44+m123_44+m124_44+m125_44+m126_44+m127_44+m128_44+m129_44+m130_44+m131_44+m132_44+m133_44+m134_44+m135_44+m136_44+m137_44+m138_44+m139_44+m140_44+m141_44+m142_44+m143_44+m144_44+m145_44+m146_44+m147_44+m148_44+m149_44+m150_44+m151_44+m152_44+m153_44+m154_44+m155_44+m156_44+m157_44+m158_44+m159_44+m160_44+m161_44+m162_44+m163_44+m164_44+m165_44+m166_44+m167_44+m168_44+m169_44+m170_44+m171_44+m172_44+m173_44+m174_44+m175_44+m176_44+m177_44+m178_44+m179_44+m180_44+m181_44+m182_44+m183_44+m184_44+m185_44+m186_44+m187_44+m188_44+m189_44+m190_44+m191_44+m192_44+m193_44+m194_44+m195_44+m196_44+m197_44+m198_44+m199_44+m200_44+m201_44+m202_44+m203_44+m204_44+m205_44+m206_44+m207_44+m208_44+m209_44+m210_44+m211_44+m212_44+m213_44+m214_44+m215_44+m216_44+m217_44+m218_44+m219_44+m220_44+m221_44+m222_44+m223_44+m224_44+m225_44+m226_44+m227_44+m228_44+m229_44+m230_44+m231_44+m232_44+m233_44+m234_44+m235_44+m236_44+m237_44+m238_44+m239_44+m240_44+m241_44+m242_44+m243_44+m244_44+m245_44+m246_44+m247_44+m248_44+m249_44+m250_44+m251_44+m252_44+m253_44+m254_44+m255_44+m256_44+m257_44+m258_44+m259_44+m260_44+m261_44+m262_44+m263_44+m264_44+m265_44+m266_44+m267_44+m268_44+m269_44+m270_44+m271_44+m272_44+m273_44+m274_44+m275_44+m276_44+m277_44+m278_44+m279_44+m280_44+m281_44+m282_44+m283_44+m284_44+m285_44+m286_44+m287_44+m288_44+m289_44+m290_44+m291_44+m292_44+m293_44+m294_44+m295_44+m296_44+m297_44+m298_44+m299_44+m300_44+m301_44+m302_44+m303_44+m304_44+m305_44+m306_44+m307_44+m308_44+m309_44+m310_44+m311_44+m312_44+m313_44+m314_44+m315_44+m316_44+m317_44+m318_44+m319_44+m320_44+m321_44+m322_44+m323_44+m324_44+m325_44+m326_44+m327_44+m328_44+m329_44+m330_44+m331_44+m332_44+m333_44+m334_44+m335_44+m336_44+m337_44+m338_44+m339_44+m340_44+m341_44+m342_44+m343_44+m344_44+m345_44+m346_44+m347_44+m348_44+m349_44+m350_44+m351_44+m352_44+m353_44+m354_44+m355_44+m356_44+m357_44+m358_44+m359_44+m360_44+m361_44+m362_44+m363_44+m364_44+m365_44+m366_44+m367_44+m368_44+m369_44+m370_44+m371_44+m372_44+m373_44+m374_44+m375_44+m376_44+m377_44+m378_44+m379_44+m380_44+m381_44+b44;
   always @(posedge clk) out45 <= m1_45+m2_45+m3_45+m4_45+m5_45+m6_45+m7_45+m8_45+m9_45+m10_45+m11_45+m12_45+m13_45+m14_45+m15_45+m16_45+m17_45+m18_45+m19_45+m20_45+m21_45+m22_45+m23_45+m24_45+m25_45+m26_45+m27_45+m28_45+m29_45+m30_45+m31_45+m32_45+m33_45+m34_45+m35_45+m36_45+m37_45+m38_45+m39_45+m40_45+m41_45+m42_45+m43_45+m44_45+m45_45+m46_45+m47_45+m48_45+m49_45+m50_45+m51_45+m52_45+m53_45+m54_45+m55_45+m56_45+m57_45+m58_45+m59_45+m60_45+m61_45+m62_45+m63_45+m64_45+m65_45+m66_45+m67_45+m68_45+m69_45+m70_45+m71_45+m72_45+m73_45+m74_45+m75_45+m76_45+m77_45+m78_45+m79_45+m80_45+m81_45+m82_45+m83_45+m84_45+m85_45+m86_45+m87_45+m88_45+m89_45+m90_45+m91_45+m92_45+m93_45+m94_45+m95_45+m96_45+m97_45+m98_45+m99_45+m100_45+m101_45+m102_45+m103_45+m104_45+m105_45+m106_45+m107_45+m108_45+m109_45+m110_45+m111_45+m112_45+m113_45+m114_45+m115_45+m116_45+m117_45+m118_45+m119_45+m120_45+m121_45+m122_45+m123_45+m124_45+m125_45+m126_45+m127_45+m128_45+m129_45+m130_45+m131_45+m132_45+m133_45+m134_45+m135_45+m136_45+m137_45+m138_45+m139_45+m140_45+m141_45+m142_45+m143_45+m144_45+m145_45+m146_45+m147_45+m148_45+m149_45+m150_45+m151_45+m152_45+m153_45+m154_45+m155_45+m156_45+m157_45+m158_45+m159_45+m160_45+m161_45+m162_45+m163_45+m164_45+m165_45+m166_45+m167_45+m168_45+m169_45+m170_45+m171_45+m172_45+m173_45+m174_45+m175_45+m176_45+m177_45+m178_45+m179_45+m180_45+m181_45+m182_45+m183_45+m184_45+m185_45+m186_45+m187_45+m188_45+m189_45+m190_45+m191_45+m192_45+m193_45+m194_45+m195_45+m196_45+m197_45+m198_45+m199_45+m200_45+m201_45+m202_45+m203_45+m204_45+m205_45+m206_45+m207_45+m208_45+m209_45+m210_45+m211_45+m212_45+m213_45+m214_45+m215_45+m216_45+m217_45+m218_45+m219_45+m220_45+m221_45+m222_45+m223_45+m224_45+m225_45+m226_45+m227_45+m228_45+m229_45+m230_45+m231_45+m232_45+m233_45+m234_45+m235_45+m236_45+m237_45+m238_45+m239_45+m240_45+m241_45+m242_45+m243_45+m244_45+m245_45+m246_45+m247_45+m248_45+m249_45+m250_45+m251_45+m252_45+m253_45+m254_45+m255_45+m256_45+m257_45+m258_45+m259_45+m260_45+m261_45+m262_45+m263_45+m264_45+m265_45+m266_45+m267_45+m268_45+m269_45+m270_45+m271_45+m272_45+m273_45+m274_45+m275_45+m276_45+m277_45+m278_45+m279_45+m280_45+m281_45+m282_45+m283_45+m284_45+m285_45+m286_45+m287_45+m288_45+m289_45+m290_45+m291_45+m292_45+m293_45+m294_45+m295_45+m296_45+m297_45+m298_45+m299_45+m300_45+m301_45+m302_45+m303_45+m304_45+m305_45+m306_45+m307_45+m308_45+m309_45+m310_45+m311_45+m312_45+m313_45+m314_45+m315_45+m316_45+m317_45+m318_45+m319_45+m320_45+m321_45+m322_45+m323_45+m324_45+m325_45+m326_45+m327_45+m328_45+m329_45+m330_45+m331_45+m332_45+m333_45+m334_45+m335_45+m336_45+m337_45+m338_45+m339_45+m340_45+m341_45+m342_45+m343_45+m344_45+m345_45+m346_45+m347_45+m348_45+m349_45+m350_45+m351_45+m352_45+m353_45+m354_45+m355_45+m356_45+m357_45+m358_45+m359_45+m360_45+m361_45+m362_45+m363_45+m364_45+m365_45+m366_45+m367_45+m368_45+m369_45+m370_45+m371_45+m372_45+m373_45+m374_45+m375_45+m376_45+m377_45+m378_45+m379_45+m380_45+m381_45+b45;
   always @(posedge clk) out46 <= m1_46+m2_46+m3_46+m4_46+m5_46+m6_46+m7_46+m8_46+m9_46+m10_46+m11_46+m12_46+m13_46+m14_46+m15_46+m16_46+m17_46+m18_46+m19_46+m20_46+m21_46+m22_46+m23_46+m24_46+m25_46+m26_46+m27_46+m28_46+m29_46+m30_46+m31_46+m32_46+m33_46+m34_46+m35_46+m36_46+m37_46+m38_46+m39_46+m40_46+m41_46+m42_46+m43_46+m44_46+m45_46+m46_46+m47_46+m48_46+m49_46+m50_46+m51_46+m52_46+m53_46+m54_46+m55_46+m56_46+m57_46+m58_46+m59_46+m60_46+m61_46+m62_46+m63_46+m64_46+m65_46+m66_46+m67_46+m68_46+m69_46+m70_46+m71_46+m72_46+m73_46+m74_46+m75_46+m76_46+m77_46+m78_46+m79_46+m80_46+m81_46+m82_46+m83_46+m84_46+m85_46+m86_46+m87_46+m88_46+m89_46+m90_46+m91_46+m92_46+m93_46+m94_46+m95_46+m96_46+m97_46+m98_46+m99_46+m100_46+m101_46+m102_46+m103_46+m104_46+m105_46+m106_46+m107_46+m108_46+m109_46+m110_46+m111_46+m112_46+m113_46+m114_46+m115_46+m116_46+m117_46+m118_46+m119_46+m120_46+m121_46+m122_46+m123_46+m124_46+m125_46+m126_46+m127_46+m128_46+m129_46+m130_46+m131_46+m132_46+m133_46+m134_46+m135_46+m136_46+m137_46+m138_46+m139_46+m140_46+m141_46+m142_46+m143_46+m144_46+m145_46+m146_46+m147_46+m148_46+m149_46+m150_46+m151_46+m152_46+m153_46+m154_46+m155_46+m156_46+m157_46+m158_46+m159_46+m160_46+m161_46+m162_46+m163_46+m164_46+m165_46+m166_46+m167_46+m168_46+m169_46+m170_46+m171_46+m172_46+m173_46+m174_46+m175_46+m176_46+m177_46+m178_46+m179_46+m180_46+m181_46+m182_46+m183_46+m184_46+m185_46+m186_46+m187_46+m188_46+m189_46+m190_46+m191_46+m192_46+m193_46+m194_46+m195_46+m196_46+m197_46+m198_46+m199_46+m200_46+m201_46+m202_46+m203_46+m204_46+m205_46+m206_46+m207_46+m208_46+m209_46+m210_46+m211_46+m212_46+m213_46+m214_46+m215_46+m216_46+m217_46+m218_46+m219_46+m220_46+m221_46+m222_46+m223_46+m224_46+m225_46+m226_46+m227_46+m228_46+m229_46+m230_46+m231_46+m232_46+m233_46+m234_46+m235_46+m236_46+m237_46+m238_46+m239_46+m240_46+m241_46+m242_46+m243_46+m244_46+m245_46+m246_46+m247_46+m248_46+m249_46+m250_46+m251_46+m252_46+m253_46+m254_46+m255_46+m256_46+m257_46+m258_46+m259_46+m260_46+m261_46+m262_46+m263_46+m264_46+m265_46+m266_46+m267_46+m268_46+m269_46+m270_46+m271_46+m272_46+m273_46+m274_46+m275_46+m276_46+m277_46+m278_46+m279_46+m280_46+m281_46+m282_46+m283_46+m284_46+m285_46+m286_46+m287_46+m288_46+m289_46+m290_46+m291_46+m292_46+m293_46+m294_46+m295_46+m296_46+m297_46+m298_46+m299_46+m300_46+m301_46+m302_46+m303_46+m304_46+m305_46+m306_46+m307_46+m308_46+m309_46+m310_46+m311_46+m312_46+m313_46+m314_46+m315_46+m316_46+m317_46+m318_46+m319_46+m320_46+m321_46+m322_46+m323_46+m324_46+m325_46+m326_46+m327_46+m328_46+m329_46+m330_46+m331_46+m332_46+m333_46+m334_46+m335_46+m336_46+m337_46+m338_46+m339_46+m340_46+m341_46+m342_46+m343_46+m344_46+m345_46+m346_46+m347_46+m348_46+m349_46+m350_46+m351_46+m352_46+m353_46+m354_46+m355_46+m356_46+m357_46+m358_46+m359_46+m360_46+m361_46+m362_46+m363_46+m364_46+m365_46+m366_46+m367_46+m368_46+m369_46+m370_46+m371_46+m372_46+m373_46+m374_46+m375_46+m376_46+m377_46+m378_46+m379_46+m380_46+m381_46+b46;
   always @(posedge clk) out47 <= m1_47+m2_47+m3_47+m4_47+m5_47+m6_47+m7_47+m8_47+m9_47+m10_47+m11_47+m12_47+m13_47+m14_47+m15_47+m16_47+m17_47+m18_47+m19_47+m20_47+m21_47+m22_47+m23_47+m24_47+m25_47+m26_47+m27_47+m28_47+m29_47+m30_47+m31_47+m32_47+m33_47+m34_47+m35_47+m36_47+m37_47+m38_47+m39_47+m40_47+m41_47+m42_47+m43_47+m44_47+m45_47+m46_47+m47_47+m48_47+m49_47+m50_47+m51_47+m52_47+m53_47+m54_47+m55_47+m56_47+m57_47+m58_47+m59_47+m60_47+m61_47+m62_47+m63_47+m64_47+m65_47+m66_47+m67_47+m68_47+m69_47+m70_47+m71_47+m72_47+m73_47+m74_47+m75_47+m76_47+m77_47+m78_47+m79_47+m80_47+m81_47+m82_47+m83_47+m84_47+m85_47+m86_47+m87_47+m88_47+m89_47+m90_47+m91_47+m92_47+m93_47+m94_47+m95_47+m96_47+m97_47+m98_47+m99_47+m100_47+m101_47+m102_47+m103_47+m104_47+m105_47+m106_47+m107_47+m108_47+m109_47+m110_47+m111_47+m112_47+m113_47+m114_47+m115_47+m116_47+m117_47+m118_47+m119_47+m120_47+m121_47+m122_47+m123_47+m124_47+m125_47+m126_47+m127_47+m128_47+m129_47+m130_47+m131_47+m132_47+m133_47+m134_47+m135_47+m136_47+m137_47+m138_47+m139_47+m140_47+m141_47+m142_47+m143_47+m144_47+m145_47+m146_47+m147_47+m148_47+m149_47+m150_47+m151_47+m152_47+m153_47+m154_47+m155_47+m156_47+m157_47+m158_47+m159_47+m160_47+m161_47+m162_47+m163_47+m164_47+m165_47+m166_47+m167_47+m168_47+m169_47+m170_47+m171_47+m172_47+m173_47+m174_47+m175_47+m176_47+m177_47+m178_47+m179_47+m180_47+m181_47+m182_47+m183_47+m184_47+m185_47+m186_47+m187_47+m188_47+m189_47+m190_47+m191_47+m192_47+m193_47+m194_47+m195_47+m196_47+m197_47+m198_47+m199_47+m200_47+m201_47+m202_47+m203_47+m204_47+m205_47+m206_47+m207_47+m208_47+m209_47+m210_47+m211_47+m212_47+m213_47+m214_47+m215_47+m216_47+m217_47+m218_47+m219_47+m220_47+m221_47+m222_47+m223_47+m224_47+m225_47+m226_47+m227_47+m228_47+m229_47+m230_47+m231_47+m232_47+m233_47+m234_47+m235_47+m236_47+m237_47+m238_47+m239_47+m240_47+m241_47+m242_47+m243_47+m244_47+m245_47+m246_47+m247_47+m248_47+m249_47+m250_47+m251_47+m252_47+m253_47+m254_47+m255_47+m256_47+m257_47+m258_47+m259_47+m260_47+m261_47+m262_47+m263_47+m264_47+m265_47+m266_47+m267_47+m268_47+m269_47+m270_47+m271_47+m272_47+m273_47+m274_47+m275_47+m276_47+m277_47+m278_47+m279_47+m280_47+m281_47+m282_47+m283_47+m284_47+m285_47+m286_47+m287_47+m288_47+m289_47+m290_47+m291_47+m292_47+m293_47+m294_47+m295_47+m296_47+m297_47+m298_47+m299_47+m300_47+m301_47+m302_47+m303_47+m304_47+m305_47+m306_47+m307_47+m308_47+m309_47+m310_47+m311_47+m312_47+m313_47+m314_47+m315_47+m316_47+m317_47+m318_47+m319_47+m320_47+m321_47+m322_47+m323_47+m324_47+m325_47+m326_47+m327_47+m328_47+m329_47+m330_47+m331_47+m332_47+m333_47+m334_47+m335_47+m336_47+m337_47+m338_47+m339_47+m340_47+m341_47+m342_47+m343_47+m344_47+m345_47+m346_47+m347_47+m348_47+m349_47+m350_47+m351_47+m352_47+m353_47+m354_47+m355_47+m356_47+m357_47+m358_47+m359_47+m360_47+m361_47+m362_47+m363_47+m364_47+m365_47+m366_47+m367_47+m368_47+m369_47+m370_47+m371_47+m372_47+m373_47+m374_47+m375_47+m376_47+m377_47+m378_47+m379_47+m380_47+m381_47+b47;
   always @(posedge clk) out48 <= m1_48+m2_48+m3_48+m4_48+m5_48+m6_48+m7_48+m8_48+m9_48+m10_48+m11_48+m12_48+m13_48+m14_48+m15_48+m16_48+m17_48+m18_48+m19_48+m20_48+m21_48+m22_48+m23_48+m24_48+m25_48+m26_48+m27_48+m28_48+m29_48+m30_48+m31_48+m32_48+m33_48+m34_48+m35_48+m36_48+m37_48+m38_48+m39_48+m40_48+m41_48+m42_48+m43_48+m44_48+m45_48+m46_48+m47_48+m48_48+m49_48+m50_48+m51_48+m52_48+m53_48+m54_48+m55_48+m56_48+m57_48+m58_48+m59_48+m60_48+m61_48+m62_48+m63_48+m64_48+m65_48+m66_48+m67_48+m68_48+m69_48+m70_48+m71_48+m72_48+m73_48+m74_48+m75_48+m76_48+m77_48+m78_48+m79_48+m80_48+m81_48+m82_48+m83_48+m84_48+m85_48+m86_48+m87_48+m88_48+m89_48+m90_48+m91_48+m92_48+m93_48+m94_48+m95_48+m96_48+m97_48+m98_48+m99_48+m100_48+m101_48+m102_48+m103_48+m104_48+m105_48+m106_48+m107_48+m108_48+m109_48+m110_48+m111_48+m112_48+m113_48+m114_48+m115_48+m116_48+m117_48+m118_48+m119_48+m120_48+m121_48+m122_48+m123_48+m124_48+m125_48+m126_48+m127_48+m128_48+m129_48+m130_48+m131_48+m132_48+m133_48+m134_48+m135_48+m136_48+m137_48+m138_48+m139_48+m140_48+m141_48+m142_48+m143_48+m144_48+m145_48+m146_48+m147_48+m148_48+m149_48+m150_48+m151_48+m152_48+m153_48+m154_48+m155_48+m156_48+m157_48+m158_48+m159_48+m160_48+m161_48+m162_48+m163_48+m164_48+m165_48+m166_48+m167_48+m168_48+m169_48+m170_48+m171_48+m172_48+m173_48+m174_48+m175_48+m176_48+m177_48+m178_48+m179_48+m180_48+m181_48+m182_48+m183_48+m184_48+m185_48+m186_48+m187_48+m188_48+m189_48+m190_48+m191_48+m192_48+m193_48+m194_48+m195_48+m196_48+m197_48+m198_48+m199_48+m200_48+m201_48+m202_48+m203_48+m204_48+m205_48+m206_48+m207_48+m208_48+m209_48+m210_48+m211_48+m212_48+m213_48+m214_48+m215_48+m216_48+m217_48+m218_48+m219_48+m220_48+m221_48+m222_48+m223_48+m224_48+m225_48+m226_48+m227_48+m228_48+m229_48+m230_48+m231_48+m232_48+m233_48+m234_48+m235_48+m236_48+m237_48+m238_48+m239_48+m240_48+m241_48+m242_48+m243_48+m244_48+m245_48+m246_48+m247_48+m248_48+m249_48+m250_48+m251_48+m252_48+m253_48+m254_48+m255_48+m256_48+m257_48+m258_48+m259_48+m260_48+m261_48+m262_48+m263_48+m264_48+m265_48+m266_48+m267_48+m268_48+m269_48+m270_48+m271_48+m272_48+m273_48+m274_48+m275_48+m276_48+m277_48+m278_48+m279_48+m280_48+m281_48+m282_48+m283_48+m284_48+m285_48+m286_48+m287_48+m288_48+m289_48+m290_48+m291_48+m292_48+m293_48+m294_48+m295_48+m296_48+m297_48+m298_48+m299_48+m300_48+m301_48+m302_48+m303_48+m304_48+m305_48+m306_48+m307_48+m308_48+m309_48+m310_48+m311_48+m312_48+m313_48+m314_48+m315_48+m316_48+m317_48+m318_48+m319_48+m320_48+m321_48+m322_48+m323_48+m324_48+m325_48+m326_48+m327_48+m328_48+m329_48+m330_48+m331_48+m332_48+m333_48+m334_48+m335_48+m336_48+m337_48+m338_48+m339_48+m340_48+m341_48+m342_48+m343_48+m344_48+m345_48+m346_48+m347_48+m348_48+m349_48+m350_48+m351_48+m352_48+m353_48+m354_48+m355_48+m356_48+m357_48+m358_48+m359_48+m360_48+m361_48+m362_48+m363_48+m364_48+m365_48+m366_48+m367_48+m368_48+m369_48+m370_48+m371_48+m372_48+m373_48+m374_48+m375_48+m376_48+m377_48+m378_48+m379_48+m380_48+m381_48+b48;
   always @(posedge clk) out49 <= m1_49+m2_49+m3_49+m4_49+m5_49+m6_49+m7_49+m8_49+m9_49+m10_49+m11_49+m12_49+m13_49+m14_49+m15_49+m16_49+m17_49+m18_49+m19_49+m20_49+m21_49+m22_49+m23_49+m24_49+m25_49+m26_49+m27_49+m28_49+m29_49+m30_49+m31_49+m32_49+m33_49+m34_49+m35_49+m36_49+m37_49+m38_49+m39_49+m40_49+m41_49+m42_49+m43_49+m44_49+m45_49+m46_49+m47_49+m48_49+m49_49+m50_49+m51_49+m52_49+m53_49+m54_49+m55_49+m56_49+m57_49+m58_49+m59_49+m60_49+m61_49+m62_49+m63_49+m64_49+m65_49+m66_49+m67_49+m68_49+m69_49+m70_49+m71_49+m72_49+m73_49+m74_49+m75_49+m76_49+m77_49+m78_49+m79_49+m80_49+m81_49+m82_49+m83_49+m84_49+m85_49+m86_49+m87_49+m88_49+m89_49+m90_49+m91_49+m92_49+m93_49+m94_49+m95_49+m96_49+m97_49+m98_49+m99_49+m100_49+m101_49+m102_49+m103_49+m104_49+m105_49+m106_49+m107_49+m108_49+m109_49+m110_49+m111_49+m112_49+m113_49+m114_49+m115_49+m116_49+m117_49+m118_49+m119_49+m120_49+m121_49+m122_49+m123_49+m124_49+m125_49+m126_49+m127_49+m128_49+m129_49+m130_49+m131_49+m132_49+m133_49+m134_49+m135_49+m136_49+m137_49+m138_49+m139_49+m140_49+m141_49+m142_49+m143_49+m144_49+m145_49+m146_49+m147_49+m148_49+m149_49+m150_49+m151_49+m152_49+m153_49+m154_49+m155_49+m156_49+m157_49+m158_49+m159_49+m160_49+m161_49+m162_49+m163_49+m164_49+m165_49+m166_49+m167_49+m168_49+m169_49+m170_49+m171_49+m172_49+m173_49+m174_49+m175_49+m176_49+m177_49+m178_49+m179_49+m180_49+m181_49+m182_49+m183_49+m184_49+m185_49+m186_49+m187_49+m188_49+m189_49+m190_49+m191_49+m192_49+m193_49+m194_49+m195_49+m196_49+m197_49+m198_49+m199_49+m200_49+m201_49+m202_49+m203_49+m204_49+m205_49+m206_49+m207_49+m208_49+m209_49+m210_49+m211_49+m212_49+m213_49+m214_49+m215_49+m216_49+m217_49+m218_49+m219_49+m220_49+m221_49+m222_49+m223_49+m224_49+m225_49+m226_49+m227_49+m228_49+m229_49+m230_49+m231_49+m232_49+m233_49+m234_49+m235_49+m236_49+m237_49+m238_49+m239_49+m240_49+m241_49+m242_49+m243_49+m244_49+m245_49+m246_49+m247_49+m248_49+m249_49+m250_49+m251_49+m252_49+m253_49+m254_49+m255_49+m256_49+m257_49+m258_49+m259_49+m260_49+m261_49+m262_49+m263_49+m264_49+m265_49+m266_49+m267_49+m268_49+m269_49+m270_49+m271_49+m272_49+m273_49+m274_49+m275_49+m276_49+m277_49+m278_49+m279_49+m280_49+m281_49+m282_49+m283_49+m284_49+m285_49+m286_49+m287_49+m288_49+m289_49+m290_49+m291_49+m292_49+m293_49+m294_49+m295_49+m296_49+m297_49+m298_49+m299_49+m300_49+m301_49+m302_49+m303_49+m304_49+m305_49+m306_49+m307_49+m308_49+m309_49+m310_49+m311_49+m312_49+m313_49+m314_49+m315_49+m316_49+m317_49+m318_49+m319_49+m320_49+m321_49+m322_49+m323_49+m324_49+m325_49+m326_49+m327_49+m328_49+m329_49+m330_49+m331_49+m332_49+m333_49+m334_49+m335_49+m336_49+m337_49+m338_49+m339_49+m340_49+m341_49+m342_49+m343_49+m344_49+m345_49+m346_49+m347_49+m348_49+m349_49+m350_49+m351_49+m352_49+m353_49+m354_49+m355_49+m356_49+m357_49+m358_49+m359_49+m360_49+m361_49+m362_49+m363_49+m364_49+m365_49+m366_49+m367_49+m368_49+m369_49+m370_49+m371_49+m372_49+m373_49+m374_49+m375_49+m376_49+m377_49+m378_49+m379_49+m380_49+m381_49+b49;
   always @(posedge clk) out50 <= m1_50+m2_50+m3_50+m4_50+m5_50+m6_50+m7_50+m8_50+m9_50+m10_50+m11_50+m12_50+m13_50+m14_50+m15_50+m16_50+m17_50+m18_50+m19_50+m20_50+m21_50+m22_50+m23_50+m24_50+m25_50+m26_50+m27_50+m28_50+m29_50+m30_50+m31_50+m32_50+m33_50+m34_50+m35_50+m36_50+m37_50+m38_50+m39_50+m40_50+m41_50+m42_50+m43_50+m44_50+m45_50+m46_50+m47_50+m48_50+m49_50+m50_50+m51_50+m52_50+m53_50+m54_50+m55_50+m56_50+m57_50+m58_50+m59_50+m60_50+m61_50+m62_50+m63_50+m64_50+m65_50+m66_50+m67_50+m68_50+m69_50+m70_50+m71_50+m72_50+m73_50+m74_50+m75_50+m76_50+m77_50+m78_50+m79_50+m80_50+m81_50+m82_50+m83_50+m84_50+m85_50+m86_50+m87_50+m88_50+m89_50+m90_50+m91_50+m92_50+m93_50+m94_50+m95_50+m96_50+m97_50+m98_50+m99_50+m100_50+m101_50+m102_50+m103_50+m104_50+m105_50+m106_50+m107_50+m108_50+m109_50+m110_50+m111_50+m112_50+m113_50+m114_50+m115_50+m116_50+m117_50+m118_50+m119_50+m120_50+m121_50+m122_50+m123_50+m124_50+m125_50+m126_50+m127_50+m128_50+m129_50+m130_50+m131_50+m132_50+m133_50+m134_50+m135_50+m136_50+m137_50+m138_50+m139_50+m140_50+m141_50+m142_50+m143_50+m144_50+m145_50+m146_50+m147_50+m148_50+m149_50+m150_50+m151_50+m152_50+m153_50+m154_50+m155_50+m156_50+m157_50+m158_50+m159_50+m160_50+m161_50+m162_50+m163_50+m164_50+m165_50+m166_50+m167_50+m168_50+m169_50+m170_50+m171_50+m172_50+m173_50+m174_50+m175_50+m176_50+m177_50+m178_50+m179_50+m180_50+m181_50+m182_50+m183_50+m184_50+m185_50+m186_50+m187_50+m188_50+m189_50+m190_50+m191_50+m192_50+m193_50+m194_50+m195_50+m196_50+m197_50+m198_50+m199_50+m200_50+m201_50+m202_50+m203_50+m204_50+m205_50+m206_50+m207_50+m208_50+m209_50+m210_50+m211_50+m212_50+m213_50+m214_50+m215_50+m216_50+m217_50+m218_50+m219_50+m220_50+m221_50+m222_50+m223_50+m224_50+m225_50+m226_50+m227_50+m228_50+m229_50+m230_50+m231_50+m232_50+m233_50+m234_50+m235_50+m236_50+m237_50+m238_50+m239_50+m240_50+m241_50+m242_50+m243_50+m244_50+m245_50+m246_50+m247_50+m248_50+m249_50+m250_50+m251_50+m252_50+m253_50+m254_50+m255_50+m256_50+m257_50+m258_50+m259_50+m260_50+m261_50+m262_50+m263_50+m264_50+m265_50+m266_50+m267_50+m268_50+m269_50+m270_50+m271_50+m272_50+m273_50+m274_50+m275_50+m276_50+m277_50+m278_50+m279_50+m280_50+m281_50+m282_50+m283_50+m284_50+m285_50+m286_50+m287_50+m288_50+m289_50+m290_50+m291_50+m292_50+m293_50+m294_50+m295_50+m296_50+m297_50+m298_50+m299_50+m300_50+m301_50+m302_50+m303_50+m304_50+m305_50+m306_50+m307_50+m308_50+m309_50+m310_50+m311_50+m312_50+m313_50+m314_50+m315_50+m316_50+m317_50+m318_50+m319_50+m320_50+m321_50+m322_50+m323_50+m324_50+m325_50+m326_50+m327_50+m328_50+m329_50+m330_50+m331_50+m332_50+m333_50+m334_50+m335_50+m336_50+m337_50+m338_50+m339_50+m340_50+m341_50+m342_50+m343_50+m344_50+m345_50+m346_50+m347_50+m348_50+m349_50+m350_50+m351_50+m352_50+m353_50+m354_50+m355_50+m356_50+m357_50+m358_50+m359_50+m360_50+m361_50+m362_50+m363_50+m364_50+m365_50+m366_50+m367_50+m368_50+m369_50+m370_50+m371_50+m372_50+m373_50+m374_50+m375_50+m376_50+m377_50+m378_50+m379_50+m380_50+m381_50+b50;
   always @(posedge clk) out51 <= m1_51+m2_51+m3_51+m4_51+m5_51+m6_51+m7_51+m8_51+m9_51+m10_51+m11_51+m12_51+m13_51+m14_51+m15_51+m16_51+m17_51+m18_51+m19_51+m20_51+m21_51+m22_51+m23_51+m24_51+m25_51+m26_51+m27_51+m28_51+m29_51+m30_51+m31_51+m32_51+m33_51+m34_51+m35_51+m36_51+m37_51+m38_51+m39_51+m40_51+m41_51+m42_51+m43_51+m44_51+m45_51+m46_51+m47_51+m48_51+m49_51+m50_51+m51_51+m52_51+m53_51+m54_51+m55_51+m56_51+m57_51+m58_51+m59_51+m60_51+m61_51+m62_51+m63_51+m64_51+m65_51+m66_51+m67_51+m68_51+m69_51+m70_51+m71_51+m72_51+m73_51+m74_51+m75_51+m76_51+m77_51+m78_51+m79_51+m80_51+m81_51+m82_51+m83_51+m84_51+m85_51+m86_51+m87_51+m88_51+m89_51+m90_51+m91_51+m92_51+m93_51+m94_51+m95_51+m96_51+m97_51+m98_51+m99_51+m100_51+m101_51+m102_51+m103_51+m104_51+m105_51+m106_51+m107_51+m108_51+m109_51+m110_51+m111_51+m112_51+m113_51+m114_51+m115_51+m116_51+m117_51+m118_51+m119_51+m120_51+m121_51+m122_51+m123_51+m124_51+m125_51+m126_51+m127_51+m128_51+m129_51+m130_51+m131_51+m132_51+m133_51+m134_51+m135_51+m136_51+m137_51+m138_51+m139_51+m140_51+m141_51+m142_51+m143_51+m144_51+m145_51+m146_51+m147_51+m148_51+m149_51+m150_51+m151_51+m152_51+m153_51+m154_51+m155_51+m156_51+m157_51+m158_51+m159_51+m160_51+m161_51+m162_51+m163_51+m164_51+m165_51+m166_51+m167_51+m168_51+m169_51+m170_51+m171_51+m172_51+m173_51+m174_51+m175_51+m176_51+m177_51+m178_51+m179_51+m180_51+m181_51+m182_51+m183_51+m184_51+m185_51+m186_51+m187_51+m188_51+m189_51+m190_51+m191_51+m192_51+m193_51+m194_51+m195_51+m196_51+m197_51+m198_51+m199_51+m200_51+m201_51+m202_51+m203_51+m204_51+m205_51+m206_51+m207_51+m208_51+m209_51+m210_51+m211_51+m212_51+m213_51+m214_51+m215_51+m216_51+m217_51+m218_51+m219_51+m220_51+m221_51+m222_51+m223_51+m224_51+m225_51+m226_51+m227_51+m228_51+m229_51+m230_51+m231_51+m232_51+m233_51+m234_51+m235_51+m236_51+m237_51+m238_51+m239_51+m240_51+m241_51+m242_51+m243_51+m244_51+m245_51+m246_51+m247_51+m248_51+m249_51+m250_51+m251_51+m252_51+m253_51+m254_51+m255_51+m256_51+m257_51+m258_51+m259_51+m260_51+m261_51+m262_51+m263_51+m264_51+m265_51+m266_51+m267_51+m268_51+m269_51+m270_51+m271_51+m272_51+m273_51+m274_51+m275_51+m276_51+m277_51+m278_51+m279_51+m280_51+m281_51+m282_51+m283_51+m284_51+m285_51+m286_51+m287_51+m288_51+m289_51+m290_51+m291_51+m292_51+m293_51+m294_51+m295_51+m296_51+m297_51+m298_51+m299_51+m300_51+m301_51+m302_51+m303_51+m304_51+m305_51+m306_51+m307_51+m308_51+m309_51+m310_51+m311_51+m312_51+m313_51+m314_51+m315_51+m316_51+m317_51+m318_51+m319_51+m320_51+m321_51+m322_51+m323_51+m324_51+m325_51+m326_51+m327_51+m328_51+m329_51+m330_51+m331_51+m332_51+m333_51+m334_51+m335_51+m336_51+m337_51+m338_51+m339_51+m340_51+m341_51+m342_51+m343_51+m344_51+m345_51+m346_51+m347_51+m348_51+m349_51+m350_51+m351_51+m352_51+m353_51+m354_51+m355_51+m356_51+m357_51+m358_51+m359_51+m360_51+m361_51+m362_51+m363_51+m364_51+m365_51+m366_51+m367_51+m368_51+m369_51+m370_51+m371_51+m372_51+m373_51+m374_51+m375_51+m376_51+m377_51+m378_51+m379_51+m380_51+m381_51+b51;
   always @(posedge clk) out52 <= m1_52+m2_52+m3_52+m4_52+m5_52+m6_52+m7_52+m8_52+m9_52+m10_52+m11_52+m12_52+m13_52+m14_52+m15_52+m16_52+m17_52+m18_52+m19_52+m20_52+m21_52+m22_52+m23_52+m24_52+m25_52+m26_52+m27_52+m28_52+m29_52+m30_52+m31_52+m32_52+m33_52+m34_52+m35_52+m36_52+m37_52+m38_52+m39_52+m40_52+m41_52+m42_52+m43_52+m44_52+m45_52+m46_52+m47_52+m48_52+m49_52+m50_52+m51_52+m52_52+m53_52+m54_52+m55_52+m56_52+m57_52+m58_52+m59_52+m60_52+m61_52+m62_52+m63_52+m64_52+m65_52+m66_52+m67_52+m68_52+m69_52+m70_52+m71_52+m72_52+m73_52+m74_52+m75_52+m76_52+m77_52+m78_52+m79_52+m80_52+m81_52+m82_52+m83_52+m84_52+m85_52+m86_52+m87_52+m88_52+m89_52+m90_52+m91_52+m92_52+m93_52+m94_52+m95_52+m96_52+m97_52+m98_52+m99_52+m100_52+m101_52+m102_52+m103_52+m104_52+m105_52+m106_52+m107_52+m108_52+m109_52+m110_52+m111_52+m112_52+m113_52+m114_52+m115_52+m116_52+m117_52+m118_52+m119_52+m120_52+m121_52+m122_52+m123_52+m124_52+m125_52+m126_52+m127_52+m128_52+m129_52+m130_52+m131_52+m132_52+m133_52+m134_52+m135_52+m136_52+m137_52+m138_52+m139_52+m140_52+m141_52+m142_52+m143_52+m144_52+m145_52+m146_52+m147_52+m148_52+m149_52+m150_52+m151_52+m152_52+m153_52+m154_52+m155_52+m156_52+m157_52+m158_52+m159_52+m160_52+m161_52+m162_52+m163_52+m164_52+m165_52+m166_52+m167_52+m168_52+m169_52+m170_52+m171_52+m172_52+m173_52+m174_52+m175_52+m176_52+m177_52+m178_52+m179_52+m180_52+m181_52+m182_52+m183_52+m184_52+m185_52+m186_52+m187_52+m188_52+m189_52+m190_52+m191_52+m192_52+m193_52+m194_52+m195_52+m196_52+m197_52+m198_52+m199_52+m200_52+m201_52+m202_52+m203_52+m204_52+m205_52+m206_52+m207_52+m208_52+m209_52+m210_52+m211_52+m212_52+m213_52+m214_52+m215_52+m216_52+m217_52+m218_52+m219_52+m220_52+m221_52+m222_52+m223_52+m224_52+m225_52+m226_52+m227_52+m228_52+m229_52+m230_52+m231_52+m232_52+m233_52+m234_52+m235_52+m236_52+m237_52+m238_52+m239_52+m240_52+m241_52+m242_52+m243_52+m244_52+m245_52+m246_52+m247_52+m248_52+m249_52+m250_52+m251_52+m252_52+m253_52+m254_52+m255_52+m256_52+m257_52+m258_52+m259_52+m260_52+m261_52+m262_52+m263_52+m264_52+m265_52+m266_52+m267_52+m268_52+m269_52+m270_52+m271_52+m272_52+m273_52+m274_52+m275_52+m276_52+m277_52+m278_52+m279_52+m280_52+m281_52+m282_52+m283_52+m284_52+m285_52+m286_52+m287_52+m288_52+m289_52+m290_52+m291_52+m292_52+m293_52+m294_52+m295_52+m296_52+m297_52+m298_52+m299_52+m300_52+m301_52+m302_52+m303_52+m304_52+m305_52+m306_52+m307_52+m308_52+m309_52+m310_52+m311_52+m312_52+m313_52+m314_52+m315_52+m316_52+m317_52+m318_52+m319_52+m320_52+m321_52+m322_52+m323_52+m324_52+m325_52+m326_52+m327_52+m328_52+m329_52+m330_52+m331_52+m332_52+m333_52+m334_52+m335_52+m336_52+m337_52+m338_52+m339_52+m340_52+m341_52+m342_52+m343_52+m344_52+m345_52+m346_52+m347_52+m348_52+m349_52+m350_52+m351_52+m352_52+m353_52+m354_52+m355_52+m356_52+m357_52+m358_52+m359_52+m360_52+m361_52+m362_52+m363_52+m364_52+m365_52+m366_52+m367_52+m368_52+m369_52+m370_52+m371_52+m372_52+m373_52+m374_52+m375_52+m376_52+m377_52+m378_52+m379_52+m380_52+m381_52+b52;
   always @(posedge clk) out53 <= m1_53+m2_53+m3_53+m4_53+m5_53+m6_53+m7_53+m8_53+m9_53+m10_53+m11_53+m12_53+m13_53+m14_53+m15_53+m16_53+m17_53+m18_53+m19_53+m20_53+m21_53+m22_53+m23_53+m24_53+m25_53+m26_53+m27_53+m28_53+m29_53+m30_53+m31_53+m32_53+m33_53+m34_53+m35_53+m36_53+m37_53+m38_53+m39_53+m40_53+m41_53+m42_53+m43_53+m44_53+m45_53+m46_53+m47_53+m48_53+m49_53+m50_53+m51_53+m52_53+m53_53+m54_53+m55_53+m56_53+m57_53+m58_53+m59_53+m60_53+m61_53+m62_53+m63_53+m64_53+m65_53+m66_53+m67_53+m68_53+m69_53+m70_53+m71_53+m72_53+m73_53+m74_53+m75_53+m76_53+m77_53+m78_53+m79_53+m80_53+m81_53+m82_53+m83_53+m84_53+m85_53+m86_53+m87_53+m88_53+m89_53+m90_53+m91_53+m92_53+m93_53+m94_53+m95_53+m96_53+m97_53+m98_53+m99_53+m100_53+m101_53+m102_53+m103_53+m104_53+m105_53+m106_53+m107_53+m108_53+m109_53+m110_53+m111_53+m112_53+m113_53+m114_53+m115_53+m116_53+m117_53+m118_53+m119_53+m120_53+m121_53+m122_53+m123_53+m124_53+m125_53+m126_53+m127_53+m128_53+m129_53+m130_53+m131_53+m132_53+m133_53+m134_53+m135_53+m136_53+m137_53+m138_53+m139_53+m140_53+m141_53+m142_53+m143_53+m144_53+m145_53+m146_53+m147_53+m148_53+m149_53+m150_53+m151_53+m152_53+m153_53+m154_53+m155_53+m156_53+m157_53+m158_53+m159_53+m160_53+m161_53+m162_53+m163_53+m164_53+m165_53+m166_53+m167_53+m168_53+m169_53+m170_53+m171_53+m172_53+m173_53+m174_53+m175_53+m176_53+m177_53+m178_53+m179_53+m180_53+m181_53+m182_53+m183_53+m184_53+m185_53+m186_53+m187_53+m188_53+m189_53+m190_53+m191_53+m192_53+m193_53+m194_53+m195_53+m196_53+m197_53+m198_53+m199_53+m200_53+m201_53+m202_53+m203_53+m204_53+m205_53+m206_53+m207_53+m208_53+m209_53+m210_53+m211_53+m212_53+m213_53+m214_53+m215_53+m216_53+m217_53+m218_53+m219_53+m220_53+m221_53+m222_53+m223_53+m224_53+m225_53+m226_53+m227_53+m228_53+m229_53+m230_53+m231_53+m232_53+m233_53+m234_53+m235_53+m236_53+m237_53+m238_53+m239_53+m240_53+m241_53+m242_53+m243_53+m244_53+m245_53+m246_53+m247_53+m248_53+m249_53+m250_53+m251_53+m252_53+m253_53+m254_53+m255_53+m256_53+m257_53+m258_53+m259_53+m260_53+m261_53+m262_53+m263_53+m264_53+m265_53+m266_53+m267_53+m268_53+m269_53+m270_53+m271_53+m272_53+m273_53+m274_53+m275_53+m276_53+m277_53+m278_53+m279_53+m280_53+m281_53+m282_53+m283_53+m284_53+m285_53+m286_53+m287_53+m288_53+m289_53+m290_53+m291_53+m292_53+m293_53+m294_53+m295_53+m296_53+m297_53+m298_53+m299_53+m300_53+m301_53+m302_53+m303_53+m304_53+m305_53+m306_53+m307_53+m308_53+m309_53+m310_53+m311_53+m312_53+m313_53+m314_53+m315_53+m316_53+m317_53+m318_53+m319_53+m320_53+m321_53+m322_53+m323_53+m324_53+m325_53+m326_53+m327_53+m328_53+m329_53+m330_53+m331_53+m332_53+m333_53+m334_53+m335_53+m336_53+m337_53+m338_53+m339_53+m340_53+m341_53+m342_53+m343_53+m344_53+m345_53+m346_53+m347_53+m348_53+m349_53+m350_53+m351_53+m352_53+m353_53+m354_53+m355_53+m356_53+m357_53+m358_53+m359_53+m360_53+m361_53+m362_53+m363_53+m364_53+m365_53+m366_53+m367_53+m368_53+m369_53+m370_53+m371_53+m372_53+m373_53+m374_53+m375_53+m376_53+m377_53+m378_53+m379_53+m380_53+m381_53+b53;
   always @(posedge clk) out54 <= m1_54+m2_54+m3_54+m4_54+m5_54+m6_54+m7_54+m8_54+m9_54+m10_54+m11_54+m12_54+m13_54+m14_54+m15_54+m16_54+m17_54+m18_54+m19_54+m20_54+m21_54+m22_54+m23_54+m24_54+m25_54+m26_54+m27_54+m28_54+m29_54+m30_54+m31_54+m32_54+m33_54+m34_54+m35_54+m36_54+m37_54+m38_54+m39_54+m40_54+m41_54+m42_54+m43_54+m44_54+m45_54+m46_54+m47_54+m48_54+m49_54+m50_54+m51_54+m52_54+m53_54+m54_54+m55_54+m56_54+m57_54+m58_54+m59_54+m60_54+m61_54+m62_54+m63_54+m64_54+m65_54+m66_54+m67_54+m68_54+m69_54+m70_54+m71_54+m72_54+m73_54+m74_54+m75_54+m76_54+m77_54+m78_54+m79_54+m80_54+m81_54+m82_54+m83_54+m84_54+m85_54+m86_54+m87_54+m88_54+m89_54+m90_54+m91_54+m92_54+m93_54+m94_54+m95_54+m96_54+m97_54+m98_54+m99_54+m100_54+m101_54+m102_54+m103_54+m104_54+m105_54+m106_54+m107_54+m108_54+m109_54+m110_54+m111_54+m112_54+m113_54+m114_54+m115_54+m116_54+m117_54+m118_54+m119_54+m120_54+m121_54+m122_54+m123_54+m124_54+m125_54+m126_54+m127_54+m128_54+m129_54+m130_54+m131_54+m132_54+m133_54+m134_54+m135_54+m136_54+m137_54+m138_54+m139_54+m140_54+m141_54+m142_54+m143_54+m144_54+m145_54+m146_54+m147_54+m148_54+m149_54+m150_54+m151_54+m152_54+m153_54+m154_54+m155_54+m156_54+m157_54+m158_54+m159_54+m160_54+m161_54+m162_54+m163_54+m164_54+m165_54+m166_54+m167_54+m168_54+m169_54+m170_54+m171_54+m172_54+m173_54+m174_54+m175_54+m176_54+m177_54+m178_54+m179_54+m180_54+m181_54+m182_54+m183_54+m184_54+m185_54+m186_54+m187_54+m188_54+m189_54+m190_54+m191_54+m192_54+m193_54+m194_54+m195_54+m196_54+m197_54+m198_54+m199_54+m200_54+m201_54+m202_54+m203_54+m204_54+m205_54+m206_54+m207_54+m208_54+m209_54+m210_54+m211_54+m212_54+m213_54+m214_54+m215_54+m216_54+m217_54+m218_54+m219_54+m220_54+m221_54+m222_54+m223_54+m224_54+m225_54+m226_54+m227_54+m228_54+m229_54+m230_54+m231_54+m232_54+m233_54+m234_54+m235_54+m236_54+m237_54+m238_54+m239_54+m240_54+m241_54+m242_54+m243_54+m244_54+m245_54+m246_54+m247_54+m248_54+m249_54+m250_54+m251_54+m252_54+m253_54+m254_54+m255_54+m256_54+m257_54+m258_54+m259_54+m260_54+m261_54+m262_54+m263_54+m264_54+m265_54+m266_54+m267_54+m268_54+m269_54+m270_54+m271_54+m272_54+m273_54+m274_54+m275_54+m276_54+m277_54+m278_54+m279_54+m280_54+m281_54+m282_54+m283_54+m284_54+m285_54+m286_54+m287_54+m288_54+m289_54+m290_54+m291_54+m292_54+m293_54+m294_54+m295_54+m296_54+m297_54+m298_54+m299_54+m300_54+m301_54+m302_54+m303_54+m304_54+m305_54+m306_54+m307_54+m308_54+m309_54+m310_54+m311_54+m312_54+m313_54+m314_54+m315_54+m316_54+m317_54+m318_54+m319_54+m320_54+m321_54+m322_54+m323_54+m324_54+m325_54+m326_54+m327_54+m328_54+m329_54+m330_54+m331_54+m332_54+m333_54+m334_54+m335_54+m336_54+m337_54+m338_54+m339_54+m340_54+m341_54+m342_54+m343_54+m344_54+m345_54+m346_54+m347_54+m348_54+m349_54+m350_54+m351_54+m352_54+m353_54+m354_54+m355_54+m356_54+m357_54+m358_54+m359_54+m360_54+m361_54+m362_54+m363_54+m364_54+m365_54+m366_54+m367_54+m368_54+m369_54+m370_54+m371_54+m372_54+m373_54+m374_54+m375_54+m376_54+m377_54+m378_54+m379_54+m380_54+m381_54+b54;
   always @(posedge clk) out55 <= m1_55+m2_55+m3_55+m4_55+m5_55+m6_55+m7_55+m8_55+m9_55+m10_55+m11_55+m12_55+m13_55+m14_55+m15_55+m16_55+m17_55+m18_55+m19_55+m20_55+m21_55+m22_55+m23_55+m24_55+m25_55+m26_55+m27_55+m28_55+m29_55+m30_55+m31_55+m32_55+m33_55+m34_55+m35_55+m36_55+m37_55+m38_55+m39_55+m40_55+m41_55+m42_55+m43_55+m44_55+m45_55+m46_55+m47_55+m48_55+m49_55+m50_55+m51_55+m52_55+m53_55+m54_55+m55_55+m56_55+m57_55+m58_55+m59_55+m60_55+m61_55+m62_55+m63_55+m64_55+m65_55+m66_55+m67_55+m68_55+m69_55+m70_55+m71_55+m72_55+m73_55+m74_55+m75_55+m76_55+m77_55+m78_55+m79_55+m80_55+m81_55+m82_55+m83_55+m84_55+m85_55+m86_55+m87_55+m88_55+m89_55+m90_55+m91_55+m92_55+m93_55+m94_55+m95_55+m96_55+m97_55+m98_55+m99_55+m100_55+m101_55+m102_55+m103_55+m104_55+m105_55+m106_55+m107_55+m108_55+m109_55+m110_55+m111_55+m112_55+m113_55+m114_55+m115_55+m116_55+m117_55+m118_55+m119_55+m120_55+m121_55+m122_55+m123_55+m124_55+m125_55+m126_55+m127_55+m128_55+m129_55+m130_55+m131_55+m132_55+m133_55+m134_55+m135_55+m136_55+m137_55+m138_55+m139_55+m140_55+m141_55+m142_55+m143_55+m144_55+m145_55+m146_55+m147_55+m148_55+m149_55+m150_55+m151_55+m152_55+m153_55+m154_55+m155_55+m156_55+m157_55+m158_55+m159_55+m160_55+m161_55+m162_55+m163_55+m164_55+m165_55+m166_55+m167_55+m168_55+m169_55+m170_55+m171_55+m172_55+m173_55+m174_55+m175_55+m176_55+m177_55+m178_55+m179_55+m180_55+m181_55+m182_55+m183_55+m184_55+m185_55+m186_55+m187_55+m188_55+m189_55+m190_55+m191_55+m192_55+m193_55+m194_55+m195_55+m196_55+m197_55+m198_55+m199_55+m200_55+m201_55+m202_55+m203_55+m204_55+m205_55+m206_55+m207_55+m208_55+m209_55+m210_55+m211_55+m212_55+m213_55+m214_55+m215_55+m216_55+m217_55+m218_55+m219_55+m220_55+m221_55+m222_55+m223_55+m224_55+m225_55+m226_55+m227_55+m228_55+m229_55+m230_55+m231_55+m232_55+m233_55+m234_55+m235_55+m236_55+m237_55+m238_55+m239_55+m240_55+m241_55+m242_55+m243_55+m244_55+m245_55+m246_55+m247_55+m248_55+m249_55+m250_55+m251_55+m252_55+m253_55+m254_55+m255_55+m256_55+m257_55+m258_55+m259_55+m260_55+m261_55+m262_55+m263_55+m264_55+m265_55+m266_55+m267_55+m268_55+m269_55+m270_55+m271_55+m272_55+m273_55+m274_55+m275_55+m276_55+m277_55+m278_55+m279_55+m280_55+m281_55+m282_55+m283_55+m284_55+m285_55+m286_55+m287_55+m288_55+m289_55+m290_55+m291_55+m292_55+m293_55+m294_55+m295_55+m296_55+m297_55+m298_55+m299_55+m300_55+m301_55+m302_55+m303_55+m304_55+m305_55+m306_55+m307_55+m308_55+m309_55+m310_55+m311_55+m312_55+m313_55+m314_55+m315_55+m316_55+m317_55+m318_55+m319_55+m320_55+m321_55+m322_55+m323_55+m324_55+m325_55+m326_55+m327_55+m328_55+m329_55+m330_55+m331_55+m332_55+m333_55+m334_55+m335_55+m336_55+m337_55+m338_55+m339_55+m340_55+m341_55+m342_55+m343_55+m344_55+m345_55+m346_55+m347_55+m348_55+m349_55+m350_55+m351_55+m352_55+m353_55+m354_55+m355_55+m356_55+m357_55+m358_55+m359_55+m360_55+m361_55+m362_55+m363_55+m364_55+m365_55+m366_55+m367_55+m368_55+m369_55+m370_55+m371_55+m372_55+m373_55+m374_55+m375_55+m376_55+m377_55+m378_55+m379_55+m380_55+m381_55+b55;
   always @(posedge clk) out56 <= m1_56+m2_56+m3_56+m4_56+m5_56+m6_56+m7_56+m8_56+m9_56+m10_56+m11_56+m12_56+m13_56+m14_56+m15_56+m16_56+m17_56+m18_56+m19_56+m20_56+m21_56+m22_56+m23_56+m24_56+m25_56+m26_56+m27_56+m28_56+m29_56+m30_56+m31_56+m32_56+m33_56+m34_56+m35_56+m36_56+m37_56+m38_56+m39_56+m40_56+m41_56+m42_56+m43_56+m44_56+m45_56+m46_56+m47_56+m48_56+m49_56+m50_56+m51_56+m52_56+m53_56+m54_56+m55_56+m56_56+m57_56+m58_56+m59_56+m60_56+m61_56+m62_56+m63_56+m64_56+m65_56+m66_56+m67_56+m68_56+m69_56+m70_56+m71_56+m72_56+m73_56+m74_56+m75_56+m76_56+m77_56+m78_56+m79_56+m80_56+m81_56+m82_56+m83_56+m84_56+m85_56+m86_56+m87_56+m88_56+m89_56+m90_56+m91_56+m92_56+m93_56+m94_56+m95_56+m96_56+m97_56+m98_56+m99_56+m100_56+m101_56+m102_56+m103_56+m104_56+m105_56+m106_56+m107_56+m108_56+m109_56+m110_56+m111_56+m112_56+m113_56+m114_56+m115_56+m116_56+m117_56+m118_56+m119_56+m120_56+m121_56+m122_56+m123_56+m124_56+m125_56+m126_56+m127_56+m128_56+m129_56+m130_56+m131_56+m132_56+m133_56+m134_56+m135_56+m136_56+m137_56+m138_56+m139_56+m140_56+m141_56+m142_56+m143_56+m144_56+m145_56+m146_56+m147_56+m148_56+m149_56+m150_56+m151_56+m152_56+m153_56+m154_56+m155_56+m156_56+m157_56+m158_56+m159_56+m160_56+m161_56+m162_56+m163_56+m164_56+m165_56+m166_56+m167_56+m168_56+m169_56+m170_56+m171_56+m172_56+m173_56+m174_56+m175_56+m176_56+m177_56+m178_56+m179_56+m180_56+m181_56+m182_56+m183_56+m184_56+m185_56+m186_56+m187_56+m188_56+m189_56+m190_56+m191_56+m192_56+m193_56+m194_56+m195_56+m196_56+m197_56+m198_56+m199_56+m200_56+m201_56+m202_56+m203_56+m204_56+m205_56+m206_56+m207_56+m208_56+m209_56+m210_56+m211_56+m212_56+m213_56+m214_56+m215_56+m216_56+m217_56+m218_56+m219_56+m220_56+m221_56+m222_56+m223_56+m224_56+m225_56+m226_56+m227_56+m228_56+m229_56+m230_56+m231_56+m232_56+m233_56+m234_56+m235_56+m236_56+m237_56+m238_56+m239_56+m240_56+m241_56+m242_56+m243_56+m244_56+m245_56+m246_56+m247_56+m248_56+m249_56+m250_56+m251_56+m252_56+m253_56+m254_56+m255_56+m256_56+m257_56+m258_56+m259_56+m260_56+m261_56+m262_56+m263_56+m264_56+m265_56+m266_56+m267_56+m268_56+m269_56+m270_56+m271_56+m272_56+m273_56+m274_56+m275_56+m276_56+m277_56+m278_56+m279_56+m280_56+m281_56+m282_56+m283_56+m284_56+m285_56+m286_56+m287_56+m288_56+m289_56+m290_56+m291_56+m292_56+m293_56+m294_56+m295_56+m296_56+m297_56+m298_56+m299_56+m300_56+m301_56+m302_56+m303_56+m304_56+m305_56+m306_56+m307_56+m308_56+m309_56+m310_56+m311_56+m312_56+m313_56+m314_56+m315_56+m316_56+m317_56+m318_56+m319_56+m320_56+m321_56+m322_56+m323_56+m324_56+m325_56+m326_56+m327_56+m328_56+m329_56+m330_56+m331_56+m332_56+m333_56+m334_56+m335_56+m336_56+m337_56+m338_56+m339_56+m340_56+m341_56+m342_56+m343_56+m344_56+m345_56+m346_56+m347_56+m348_56+m349_56+m350_56+m351_56+m352_56+m353_56+m354_56+m355_56+m356_56+m357_56+m358_56+m359_56+m360_56+m361_56+m362_56+m363_56+m364_56+m365_56+m366_56+m367_56+m368_56+m369_56+m370_56+m371_56+m372_56+m373_56+m374_56+m375_56+m376_56+m377_56+m378_56+m379_56+m380_56+m381_56+b56;
   always @(posedge clk) out57 <= m1_57+m2_57+m3_57+m4_57+m5_57+m6_57+m7_57+m8_57+m9_57+m10_57+m11_57+m12_57+m13_57+m14_57+m15_57+m16_57+m17_57+m18_57+m19_57+m20_57+m21_57+m22_57+m23_57+m24_57+m25_57+m26_57+m27_57+m28_57+m29_57+m30_57+m31_57+m32_57+m33_57+m34_57+m35_57+m36_57+m37_57+m38_57+m39_57+m40_57+m41_57+m42_57+m43_57+m44_57+m45_57+m46_57+m47_57+m48_57+m49_57+m50_57+m51_57+m52_57+m53_57+m54_57+m55_57+m56_57+m57_57+m58_57+m59_57+m60_57+m61_57+m62_57+m63_57+m64_57+m65_57+m66_57+m67_57+m68_57+m69_57+m70_57+m71_57+m72_57+m73_57+m74_57+m75_57+m76_57+m77_57+m78_57+m79_57+m80_57+m81_57+m82_57+m83_57+m84_57+m85_57+m86_57+m87_57+m88_57+m89_57+m90_57+m91_57+m92_57+m93_57+m94_57+m95_57+m96_57+m97_57+m98_57+m99_57+m100_57+m101_57+m102_57+m103_57+m104_57+m105_57+m106_57+m107_57+m108_57+m109_57+m110_57+m111_57+m112_57+m113_57+m114_57+m115_57+m116_57+m117_57+m118_57+m119_57+m120_57+m121_57+m122_57+m123_57+m124_57+m125_57+m126_57+m127_57+m128_57+m129_57+m130_57+m131_57+m132_57+m133_57+m134_57+m135_57+m136_57+m137_57+m138_57+m139_57+m140_57+m141_57+m142_57+m143_57+m144_57+m145_57+m146_57+m147_57+m148_57+m149_57+m150_57+m151_57+m152_57+m153_57+m154_57+m155_57+m156_57+m157_57+m158_57+m159_57+m160_57+m161_57+m162_57+m163_57+m164_57+m165_57+m166_57+m167_57+m168_57+m169_57+m170_57+m171_57+m172_57+m173_57+m174_57+m175_57+m176_57+m177_57+m178_57+m179_57+m180_57+m181_57+m182_57+m183_57+m184_57+m185_57+m186_57+m187_57+m188_57+m189_57+m190_57+m191_57+m192_57+m193_57+m194_57+m195_57+m196_57+m197_57+m198_57+m199_57+m200_57+m201_57+m202_57+m203_57+m204_57+m205_57+m206_57+m207_57+m208_57+m209_57+m210_57+m211_57+m212_57+m213_57+m214_57+m215_57+m216_57+m217_57+m218_57+m219_57+m220_57+m221_57+m222_57+m223_57+m224_57+m225_57+m226_57+m227_57+m228_57+m229_57+m230_57+m231_57+m232_57+m233_57+m234_57+m235_57+m236_57+m237_57+m238_57+m239_57+m240_57+m241_57+m242_57+m243_57+m244_57+m245_57+m246_57+m247_57+m248_57+m249_57+m250_57+m251_57+m252_57+m253_57+m254_57+m255_57+m256_57+m257_57+m258_57+m259_57+m260_57+m261_57+m262_57+m263_57+m264_57+m265_57+m266_57+m267_57+m268_57+m269_57+m270_57+m271_57+m272_57+m273_57+m274_57+m275_57+m276_57+m277_57+m278_57+m279_57+m280_57+m281_57+m282_57+m283_57+m284_57+m285_57+m286_57+m287_57+m288_57+m289_57+m290_57+m291_57+m292_57+m293_57+m294_57+m295_57+m296_57+m297_57+m298_57+m299_57+m300_57+m301_57+m302_57+m303_57+m304_57+m305_57+m306_57+m307_57+m308_57+m309_57+m310_57+m311_57+m312_57+m313_57+m314_57+m315_57+m316_57+m317_57+m318_57+m319_57+m320_57+m321_57+m322_57+m323_57+m324_57+m325_57+m326_57+m327_57+m328_57+m329_57+m330_57+m331_57+m332_57+m333_57+m334_57+m335_57+m336_57+m337_57+m338_57+m339_57+m340_57+m341_57+m342_57+m343_57+m344_57+m345_57+m346_57+m347_57+m348_57+m349_57+m350_57+m351_57+m352_57+m353_57+m354_57+m355_57+m356_57+m357_57+m358_57+m359_57+m360_57+m361_57+m362_57+m363_57+m364_57+m365_57+m366_57+m367_57+m368_57+m369_57+m370_57+m371_57+m372_57+m373_57+m374_57+m375_57+m376_57+m377_57+m378_57+m379_57+m380_57+m381_57+b57;
   always @(posedge clk) out58 <= m1_58+m2_58+m3_58+m4_58+m5_58+m6_58+m7_58+m8_58+m9_58+m10_58+m11_58+m12_58+m13_58+m14_58+m15_58+m16_58+m17_58+m18_58+m19_58+m20_58+m21_58+m22_58+m23_58+m24_58+m25_58+m26_58+m27_58+m28_58+m29_58+m30_58+m31_58+m32_58+m33_58+m34_58+m35_58+m36_58+m37_58+m38_58+m39_58+m40_58+m41_58+m42_58+m43_58+m44_58+m45_58+m46_58+m47_58+m48_58+m49_58+m50_58+m51_58+m52_58+m53_58+m54_58+m55_58+m56_58+m57_58+m58_58+m59_58+m60_58+m61_58+m62_58+m63_58+m64_58+m65_58+m66_58+m67_58+m68_58+m69_58+m70_58+m71_58+m72_58+m73_58+m74_58+m75_58+m76_58+m77_58+m78_58+m79_58+m80_58+m81_58+m82_58+m83_58+m84_58+m85_58+m86_58+m87_58+m88_58+m89_58+m90_58+m91_58+m92_58+m93_58+m94_58+m95_58+m96_58+m97_58+m98_58+m99_58+m100_58+m101_58+m102_58+m103_58+m104_58+m105_58+m106_58+m107_58+m108_58+m109_58+m110_58+m111_58+m112_58+m113_58+m114_58+m115_58+m116_58+m117_58+m118_58+m119_58+m120_58+m121_58+m122_58+m123_58+m124_58+m125_58+m126_58+m127_58+m128_58+m129_58+m130_58+m131_58+m132_58+m133_58+m134_58+m135_58+m136_58+m137_58+m138_58+m139_58+m140_58+m141_58+m142_58+m143_58+m144_58+m145_58+m146_58+m147_58+m148_58+m149_58+m150_58+m151_58+m152_58+m153_58+m154_58+m155_58+m156_58+m157_58+m158_58+m159_58+m160_58+m161_58+m162_58+m163_58+m164_58+m165_58+m166_58+m167_58+m168_58+m169_58+m170_58+m171_58+m172_58+m173_58+m174_58+m175_58+m176_58+m177_58+m178_58+m179_58+m180_58+m181_58+m182_58+m183_58+m184_58+m185_58+m186_58+m187_58+m188_58+m189_58+m190_58+m191_58+m192_58+m193_58+m194_58+m195_58+m196_58+m197_58+m198_58+m199_58+m200_58+m201_58+m202_58+m203_58+m204_58+m205_58+m206_58+m207_58+m208_58+m209_58+m210_58+m211_58+m212_58+m213_58+m214_58+m215_58+m216_58+m217_58+m218_58+m219_58+m220_58+m221_58+m222_58+m223_58+m224_58+m225_58+m226_58+m227_58+m228_58+m229_58+m230_58+m231_58+m232_58+m233_58+m234_58+m235_58+m236_58+m237_58+m238_58+m239_58+m240_58+m241_58+m242_58+m243_58+m244_58+m245_58+m246_58+m247_58+m248_58+m249_58+m250_58+m251_58+m252_58+m253_58+m254_58+m255_58+m256_58+m257_58+m258_58+m259_58+m260_58+m261_58+m262_58+m263_58+m264_58+m265_58+m266_58+m267_58+m268_58+m269_58+m270_58+m271_58+m272_58+m273_58+m274_58+m275_58+m276_58+m277_58+m278_58+m279_58+m280_58+m281_58+m282_58+m283_58+m284_58+m285_58+m286_58+m287_58+m288_58+m289_58+m290_58+m291_58+m292_58+m293_58+m294_58+m295_58+m296_58+m297_58+m298_58+m299_58+m300_58+m301_58+m302_58+m303_58+m304_58+m305_58+m306_58+m307_58+m308_58+m309_58+m310_58+m311_58+m312_58+m313_58+m314_58+m315_58+m316_58+m317_58+m318_58+m319_58+m320_58+m321_58+m322_58+m323_58+m324_58+m325_58+m326_58+m327_58+m328_58+m329_58+m330_58+m331_58+m332_58+m333_58+m334_58+m335_58+m336_58+m337_58+m338_58+m339_58+m340_58+m341_58+m342_58+m343_58+m344_58+m345_58+m346_58+m347_58+m348_58+m349_58+m350_58+m351_58+m352_58+m353_58+m354_58+m355_58+m356_58+m357_58+m358_58+m359_58+m360_58+m361_58+m362_58+m363_58+m364_58+m365_58+m366_58+m367_58+m368_58+m369_58+m370_58+m371_58+m372_58+m373_58+m374_58+m375_58+m376_58+m377_58+m378_58+m379_58+m380_58+m381_58+b58;
   always @(posedge clk) out59 <= m1_59+m2_59+m3_59+m4_59+m5_59+m6_59+m7_59+m8_59+m9_59+m10_59+m11_59+m12_59+m13_59+m14_59+m15_59+m16_59+m17_59+m18_59+m19_59+m20_59+m21_59+m22_59+m23_59+m24_59+m25_59+m26_59+m27_59+m28_59+m29_59+m30_59+m31_59+m32_59+m33_59+m34_59+m35_59+m36_59+m37_59+m38_59+m39_59+m40_59+m41_59+m42_59+m43_59+m44_59+m45_59+m46_59+m47_59+m48_59+m49_59+m50_59+m51_59+m52_59+m53_59+m54_59+m55_59+m56_59+m57_59+m58_59+m59_59+m60_59+m61_59+m62_59+m63_59+m64_59+m65_59+m66_59+m67_59+m68_59+m69_59+m70_59+m71_59+m72_59+m73_59+m74_59+m75_59+m76_59+m77_59+m78_59+m79_59+m80_59+m81_59+m82_59+m83_59+m84_59+m85_59+m86_59+m87_59+m88_59+m89_59+m90_59+m91_59+m92_59+m93_59+m94_59+m95_59+m96_59+m97_59+m98_59+m99_59+m100_59+m101_59+m102_59+m103_59+m104_59+m105_59+m106_59+m107_59+m108_59+m109_59+m110_59+m111_59+m112_59+m113_59+m114_59+m115_59+m116_59+m117_59+m118_59+m119_59+m120_59+m121_59+m122_59+m123_59+m124_59+m125_59+m126_59+m127_59+m128_59+m129_59+m130_59+m131_59+m132_59+m133_59+m134_59+m135_59+m136_59+m137_59+m138_59+m139_59+m140_59+m141_59+m142_59+m143_59+m144_59+m145_59+m146_59+m147_59+m148_59+m149_59+m150_59+m151_59+m152_59+m153_59+m154_59+m155_59+m156_59+m157_59+m158_59+m159_59+m160_59+m161_59+m162_59+m163_59+m164_59+m165_59+m166_59+m167_59+m168_59+m169_59+m170_59+m171_59+m172_59+m173_59+m174_59+m175_59+m176_59+m177_59+m178_59+m179_59+m180_59+m181_59+m182_59+m183_59+m184_59+m185_59+m186_59+m187_59+m188_59+m189_59+m190_59+m191_59+m192_59+m193_59+m194_59+m195_59+m196_59+m197_59+m198_59+m199_59+m200_59+m201_59+m202_59+m203_59+m204_59+m205_59+m206_59+m207_59+m208_59+m209_59+m210_59+m211_59+m212_59+m213_59+m214_59+m215_59+m216_59+m217_59+m218_59+m219_59+m220_59+m221_59+m222_59+m223_59+m224_59+m225_59+m226_59+m227_59+m228_59+m229_59+m230_59+m231_59+m232_59+m233_59+m234_59+m235_59+m236_59+m237_59+m238_59+m239_59+m240_59+m241_59+m242_59+m243_59+m244_59+m245_59+m246_59+m247_59+m248_59+m249_59+m250_59+m251_59+m252_59+m253_59+m254_59+m255_59+m256_59+m257_59+m258_59+m259_59+m260_59+m261_59+m262_59+m263_59+m264_59+m265_59+m266_59+m267_59+m268_59+m269_59+m270_59+m271_59+m272_59+m273_59+m274_59+m275_59+m276_59+m277_59+m278_59+m279_59+m280_59+m281_59+m282_59+m283_59+m284_59+m285_59+m286_59+m287_59+m288_59+m289_59+m290_59+m291_59+m292_59+m293_59+m294_59+m295_59+m296_59+m297_59+m298_59+m299_59+m300_59+m301_59+m302_59+m303_59+m304_59+m305_59+m306_59+m307_59+m308_59+m309_59+m310_59+m311_59+m312_59+m313_59+m314_59+m315_59+m316_59+m317_59+m318_59+m319_59+m320_59+m321_59+m322_59+m323_59+m324_59+m325_59+m326_59+m327_59+m328_59+m329_59+m330_59+m331_59+m332_59+m333_59+m334_59+m335_59+m336_59+m337_59+m338_59+m339_59+m340_59+m341_59+m342_59+m343_59+m344_59+m345_59+m346_59+m347_59+m348_59+m349_59+m350_59+m351_59+m352_59+m353_59+m354_59+m355_59+m356_59+m357_59+m358_59+m359_59+m360_59+m361_59+m362_59+m363_59+m364_59+m365_59+m366_59+m367_59+m368_59+m369_59+m370_59+m371_59+m372_59+m373_59+m374_59+m375_59+m376_59+m377_59+m378_59+m379_59+m380_59+m381_59+b59;
   always @(posedge clk) out60 <= m1_60+m2_60+m3_60+m4_60+m5_60+m6_60+m7_60+m8_60+m9_60+m10_60+m11_60+m12_60+m13_60+m14_60+m15_60+m16_60+m17_60+m18_60+m19_60+m20_60+m21_60+m22_60+m23_60+m24_60+m25_60+m26_60+m27_60+m28_60+m29_60+m30_60+m31_60+m32_60+m33_60+m34_60+m35_60+m36_60+m37_60+m38_60+m39_60+m40_60+m41_60+m42_60+m43_60+m44_60+m45_60+m46_60+m47_60+m48_60+m49_60+m50_60+m51_60+m52_60+m53_60+m54_60+m55_60+m56_60+m57_60+m58_60+m59_60+m60_60+m61_60+m62_60+m63_60+m64_60+m65_60+m66_60+m67_60+m68_60+m69_60+m70_60+m71_60+m72_60+m73_60+m74_60+m75_60+m76_60+m77_60+m78_60+m79_60+m80_60+m81_60+m82_60+m83_60+m84_60+m85_60+m86_60+m87_60+m88_60+m89_60+m90_60+m91_60+m92_60+m93_60+m94_60+m95_60+m96_60+m97_60+m98_60+m99_60+m100_60+m101_60+m102_60+m103_60+m104_60+m105_60+m106_60+m107_60+m108_60+m109_60+m110_60+m111_60+m112_60+m113_60+m114_60+m115_60+m116_60+m117_60+m118_60+m119_60+m120_60+m121_60+m122_60+m123_60+m124_60+m125_60+m126_60+m127_60+m128_60+m129_60+m130_60+m131_60+m132_60+m133_60+m134_60+m135_60+m136_60+m137_60+m138_60+m139_60+m140_60+m141_60+m142_60+m143_60+m144_60+m145_60+m146_60+m147_60+m148_60+m149_60+m150_60+m151_60+m152_60+m153_60+m154_60+m155_60+m156_60+m157_60+m158_60+m159_60+m160_60+m161_60+m162_60+m163_60+m164_60+m165_60+m166_60+m167_60+m168_60+m169_60+m170_60+m171_60+m172_60+m173_60+m174_60+m175_60+m176_60+m177_60+m178_60+m179_60+m180_60+m181_60+m182_60+m183_60+m184_60+m185_60+m186_60+m187_60+m188_60+m189_60+m190_60+m191_60+m192_60+m193_60+m194_60+m195_60+m196_60+m197_60+m198_60+m199_60+m200_60+m201_60+m202_60+m203_60+m204_60+m205_60+m206_60+m207_60+m208_60+m209_60+m210_60+m211_60+m212_60+m213_60+m214_60+m215_60+m216_60+m217_60+m218_60+m219_60+m220_60+m221_60+m222_60+m223_60+m224_60+m225_60+m226_60+m227_60+m228_60+m229_60+m230_60+m231_60+m232_60+m233_60+m234_60+m235_60+m236_60+m237_60+m238_60+m239_60+m240_60+m241_60+m242_60+m243_60+m244_60+m245_60+m246_60+m247_60+m248_60+m249_60+m250_60+m251_60+m252_60+m253_60+m254_60+m255_60+m256_60+m257_60+m258_60+m259_60+m260_60+m261_60+m262_60+m263_60+m264_60+m265_60+m266_60+m267_60+m268_60+m269_60+m270_60+m271_60+m272_60+m273_60+m274_60+m275_60+m276_60+m277_60+m278_60+m279_60+m280_60+m281_60+m282_60+m283_60+m284_60+m285_60+m286_60+m287_60+m288_60+m289_60+m290_60+m291_60+m292_60+m293_60+m294_60+m295_60+m296_60+m297_60+m298_60+m299_60+m300_60+m301_60+m302_60+m303_60+m304_60+m305_60+m306_60+m307_60+m308_60+m309_60+m310_60+m311_60+m312_60+m313_60+m314_60+m315_60+m316_60+m317_60+m318_60+m319_60+m320_60+m321_60+m322_60+m323_60+m324_60+m325_60+m326_60+m327_60+m328_60+m329_60+m330_60+m331_60+m332_60+m333_60+m334_60+m335_60+m336_60+m337_60+m338_60+m339_60+m340_60+m341_60+m342_60+m343_60+m344_60+m345_60+m346_60+m347_60+m348_60+m349_60+m350_60+m351_60+m352_60+m353_60+m354_60+m355_60+m356_60+m357_60+m358_60+m359_60+m360_60+m361_60+m362_60+m363_60+m364_60+m365_60+m366_60+m367_60+m368_60+m369_60+m370_60+m371_60+m372_60+m373_60+m374_60+m375_60+m376_60+m377_60+m378_60+m379_60+m380_60+m381_60+b60;
   always @(posedge clk) out61 <= m1_61+m2_61+m3_61+m4_61+m5_61+m6_61+m7_61+m8_61+m9_61+m10_61+m11_61+m12_61+m13_61+m14_61+m15_61+m16_61+m17_61+m18_61+m19_61+m20_61+m21_61+m22_61+m23_61+m24_61+m25_61+m26_61+m27_61+m28_61+m29_61+m30_61+m31_61+m32_61+m33_61+m34_61+m35_61+m36_61+m37_61+m38_61+m39_61+m40_61+m41_61+m42_61+m43_61+m44_61+m45_61+m46_61+m47_61+m48_61+m49_61+m50_61+m51_61+m52_61+m53_61+m54_61+m55_61+m56_61+m57_61+m58_61+m59_61+m60_61+m61_61+m62_61+m63_61+m64_61+m65_61+m66_61+m67_61+m68_61+m69_61+m70_61+m71_61+m72_61+m73_61+m74_61+m75_61+m76_61+m77_61+m78_61+m79_61+m80_61+m81_61+m82_61+m83_61+m84_61+m85_61+m86_61+m87_61+m88_61+m89_61+m90_61+m91_61+m92_61+m93_61+m94_61+m95_61+m96_61+m97_61+m98_61+m99_61+m100_61+m101_61+m102_61+m103_61+m104_61+m105_61+m106_61+m107_61+m108_61+m109_61+m110_61+m111_61+m112_61+m113_61+m114_61+m115_61+m116_61+m117_61+m118_61+m119_61+m120_61+m121_61+m122_61+m123_61+m124_61+m125_61+m126_61+m127_61+m128_61+m129_61+m130_61+m131_61+m132_61+m133_61+m134_61+m135_61+m136_61+m137_61+m138_61+m139_61+m140_61+m141_61+m142_61+m143_61+m144_61+m145_61+m146_61+m147_61+m148_61+m149_61+m150_61+m151_61+m152_61+m153_61+m154_61+m155_61+m156_61+m157_61+m158_61+m159_61+m160_61+m161_61+m162_61+m163_61+m164_61+m165_61+m166_61+m167_61+m168_61+m169_61+m170_61+m171_61+m172_61+m173_61+m174_61+m175_61+m176_61+m177_61+m178_61+m179_61+m180_61+m181_61+m182_61+m183_61+m184_61+m185_61+m186_61+m187_61+m188_61+m189_61+m190_61+m191_61+m192_61+m193_61+m194_61+m195_61+m196_61+m197_61+m198_61+m199_61+m200_61+m201_61+m202_61+m203_61+m204_61+m205_61+m206_61+m207_61+m208_61+m209_61+m210_61+m211_61+m212_61+m213_61+m214_61+m215_61+m216_61+m217_61+m218_61+m219_61+m220_61+m221_61+m222_61+m223_61+m224_61+m225_61+m226_61+m227_61+m228_61+m229_61+m230_61+m231_61+m232_61+m233_61+m234_61+m235_61+m236_61+m237_61+m238_61+m239_61+m240_61+m241_61+m242_61+m243_61+m244_61+m245_61+m246_61+m247_61+m248_61+m249_61+m250_61+m251_61+m252_61+m253_61+m254_61+m255_61+m256_61+m257_61+m258_61+m259_61+m260_61+m261_61+m262_61+m263_61+m264_61+m265_61+m266_61+m267_61+m268_61+m269_61+m270_61+m271_61+m272_61+m273_61+m274_61+m275_61+m276_61+m277_61+m278_61+m279_61+m280_61+m281_61+m282_61+m283_61+m284_61+m285_61+m286_61+m287_61+m288_61+m289_61+m290_61+m291_61+m292_61+m293_61+m294_61+m295_61+m296_61+m297_61+m298_61+m299_61+m300_61+m301_61+m302_61+m303_61+m304_61+m305_61+m306_61+m307_61+m308_61+m309_61+m310_61+m311_61+m312_61+m313_61+m314_61+m315_61+m316_61+m317_61+m318_61+m319_61+m320_61+m321_61+m322_61+m323_61+m324_61+m325_61+m326_61+m327_61+m328_61+m329_61+m330_61+m331_61+m332_61+m333_61+m334_61+m335_61+m336_61+m337_61+m338_61+m339_61+m340_61+m341_61+m342_61+m343_61+m344_61+m345_61+m346_61+m347_61+m348_61+m349_61+m350_61+m351_61+m352_61+m353_61+m354_61+m355_61+m356_61+m357_61+m358_61+m359_61+m360_61+m361_61+m362_61+m363_61+m364_61+m365_61+m366_61+m367_61+m368_61+m369_61+m370_61+m371_61+m372_61+m373_61+m374_61+m375_61+m376_61+m377_61+m378_61+m379_61+m380_61+m381_61+b61;
   always @(posedge clk) out62 <= m1_62+m2_62+m3_62+m4_62+m5_62+m6_62+m7_62+m8_62+m9_62+m10_62+m11_62+m12_62+m13_62+m14_62+m15_62+m16_62+m17_62+m18_62+m19_62+m20_62+m21_62+m22_62+m23_62+m24_62+m25_62+m26_62+m27_62+m28_62+m29_62+m30_62+m31_62+m32_62+m33_62+m34_62+m35_62+m36_62+m37_62+m38_62+m39_62+m40_62+m41_62+m42_62+m43_62+m44_62+m45_62+m46_62+m47_62+m48_62+m49_62+m50_62+m51_62+m52_62+m53_62+m54_62+m55_62+m56_62+m57_62+m58_62+m59_62+m60_62+m61_62+m62_62+m63_62+m64_62+m65_62+m66_62+m67_62+m68_62+m69_62+m70_62+m71_62+m72_62+m73_62+m74_62+m75_62+m76_62+m77_62+m78_62+m79_62+m80_62+m81_62+m82_62+m83_62+m84_62+m85_62+m86_62+m87_62+m88_62+m89_62+m90_62+m91_62+m92_62+m93_62+m94_62+m95_62+m96_62+m97_62+m98_62+m99_62+m100_62+m101_62+m102_62+m103_62+m104_62+m105_62+m106_62+m107_62+m108_62+m109_62+m110_62+m111_62+m112_62+m113_62+m114_62+m115_62+m116_62+m117_62+m118_62+m119_62+m120_62+m121_62+m122_62+m123_62+m124_62+m125_62+m126_62+m127_62+m128_62+m129_62+m130_62+m131_62+m132_62+m133_62+m134_62+m135_62+m136_62+m137_62+m138_62+m139_62+m140_62+m141_62+m142_62+m143_62+m144_62+m145_62+m146_62+m147_62+m148_62+m149_62+m150_62+m151_62+m152_62+m153_62+m154_62+m155_62+m156_62+m157_62+m158_62+m159_62+m160_62+m161_62+m162_62+m163_62+m164_62+m165_62+m166_62+m167_62+m168_62+m169_62+m170_62+m171_62+m172_62+m173_62+m174_62+m175_62+m176_62+m177_62+m178_62+m179_62+m180_62+m181_62+m182_62+m183_62+m184_62+m185_62+m186_62+m187_62+m188_62+m189_62+m190_62+m191_62+m192_62+m193_62+m194_62+m195_62+m196_62+m197_62+m198_62+m199_62+m200_62+m201_62+m202_62+m203_62+m204_62+m205_62+m206_62+m207_62+m208_62+m209_62+m210_62+m211_62+m212_62+m213_62+m214_62+m215_62+m216_62+m217_62+m218_62+m219_62+m220_62+m221_62+m222_62+m223_62+m224_62+m225_62+m226_62+m227_62+m228_62+m229_62+m230_62+m231_62+m232_62+m233_62+m234_62+m235_62+m236_62+m237_62+m238_62+m239_62+m240_62+m241_62+m242_62+m243_62+m244_62+m245_62+m246_62+m247_62+m248_62+m249_62+m250_62+m251_62+m252_62+m253_62+m254_62+m255_62+m256_62+m257_62+m258_62+m259_62+m260_62+m261_62+m262_62+m263_62+m264_62+m265_62+m266_62+m267_62+m268_62+m269_62+m270_62+m271_62+m272_62+m273_62+m274_62+m275_62+m276_62+m277_62+m278_62+m279_62+m280_62+m281_62+m282_62+m283_62+m284_62+m285_62+m286_62+m287_62+m288_62+m289_62+m290_62+m291_62+m292_62+m293_62+m294_62+m295_62+m296_62+m297_62+m298_62+m299_62+m300_62+m301_62+m302_62+m303_62+m304_62+m305_62+m306_62+m307_62+m308_62+m309_62+m310_62+m311_62+m312_62+m313_62+m314_62+m315_62+m316_62+m317_62+m318_62+m319_62+m320_62+m321_62+m322_62+m323_62+m324_62+m325_62+m326_62+m327_62+m328_62+m329_62+m330_62+m331_62+m332_62+m333_62+m334_62+m335_62+m336_62+m337_62+m338_62+m339_62+m340_62+m341_62+m342_62+m343_62+m344_62+m345_62+m346_62+m347_62+m348_62+m349_62+m350_62+m351_62+m352_62+m353_62+m354_62+m355_62+m356_62+m357_62+m358_62+m359_62+m360_62+m361_62+m362_62+m363_62+m364_62+m365_62+m366_62+m367_62+m368_62+m369_62+m370_62+m371_62+m372_62+m373_62+m374_62+m375_62+m376_62+m377_62+m378_62+m379_62+m380_62+m381_62+b62;
   always @(posedge clk) out63 <= m1_63+m2_63+m3_63+m4_63+m5_63+m6_63+m7_63+m8_63+m9_63+m10_63+m11_63+m12_63+m13_63+m14_63+m15_63+m16_63+m17_63+m18_63+m19_63+m20_63+m21_63+m22_63+m23_63+m24_63+m25_63+m26_63+m27_63+m28_63+m29_63+m30_63+m31_63+m32_63+m33_63+m34_63+m35_63+m36_63+m37_63+m38_63+m39_63+m40_63+m41_63+m42_63+m43_63+m44_63+m45_63+m46_63+m47_63+m48_63+m49_63+m50_63+m51_63+m52_63+m53_63+m54_63+m55_63+m56_63+m57_63+m58_63+m59_63+m60_63+m61_63+m62_63+m63_63+m64_63+m65_63+m66_63+m67_63+m68_63+m69_63+m70_63+m71_63+m72_63+m73_63+m74_63+m75_63+m76_63+m77_63+m78_63+m79_63+m80_63+m81_63+m82_63+m83_63+m84_63+m85_63+m86_63+m87_63+m88_63+m89_63+m90_63+m91_63+m92_63+m93_63+m94_63+m95_63+m96_63+m97_63+m98_63+m99_63+m100_63+m101_63+m102_63+m103_63+m104_63+m105_63+m106_63+m107_63+m108_63+m109_63+m110_63+m111_63+m112_63+m113_63+m114_63+m115_63+m116_63+m117_63+m118_63+m119_63+m120_63+m121_63+m122_63+m123_63+m124_63+m125_63+m126_63+m127_63+m128_63+m129_63+m130_63+m131_63+m132_63+m133_63+m134_63+m135_63+m136_63+m137_63+m138_63+m139_63+m140_63+m141_63+m142_63+m143_63+m144_63+m145_63+m146_63+m147_63+m148_63+m149_63+m150_63+m151_63+m152_63+m153_63+m154_63+m155_63+m156_63+m157_63+m158_63+m159_63+m160_63+m161_63+m162_63+m163_63+m164_63+m165_63+m166_63+m167_63+m168_63+m169_63+m170_63+m171_63+m172_63+m173_63+m174_63+m175_63+m176_63+m177_63+m178_63+m179_63+m180_63+m181_63+m182_63+m183_63+m184_63+m185_63+m186_63+m187_63+m188_63+m189_63+m190_63+m191_63+m192_63+m193_63+m194_63+m195_63+m196_63+m197_63+m198_63+m199_63+m200_63+m201_63+m202_63+m203_63+m204_63+m205_63+m206_63+m207_63+m208_63+m209_63+m210_63+m211_63+m212_63+m213_63+m214_63+m215_63+m216_63+m217_63+m218_63+m219_63+m220_63+m221_63+m222_63+m223_63+m224_63+m225_63+m226_63+m227_63+m228_63+m229_63+m230_63+m231_63+m232_63+m233_63+m234_63+m235_63+m236_63+m237_63+m238_63+m239_63+m240_63+m241_63+m242_63+m243_63+m244_63+m245_63+m246_63+m247_63+m248_63+m249_63+m250_63+m251_63+m252_63+m253_63+m254_63+m255_63+m256_63+m257_63+m258_63+m259_63+m260_63+m261_63+m262_63+m263_63+m264_63+m265_63+m266_63+m267_63+m268_63+m269_63+m270_63+m271_63+m272_63+m273_63+m274_63+m275_63+m276_63+m277_63+m278_63+m279_63+m280_63+m281_63+m282_63+m283_63+m284_63+m285_63+m286_63+m287_63+m288_63+m289_63+m290_63+m291_63+m292_63+m293_63+m294_63+m295_63+m296_63+m297_63+m298_63+m299_63+m300_63+m301_63+m302_63+m303_63+m304_63+m305_63+m306_63+m307_63+m308_63+m309_63+m310_63+m311_63+m312_63+m313_63+m314_63+m315_63+m316_63+m317_63+m318_63+m319_63+m320_63+m321_63+m322_63+m323_63+m324_63+m325_63+m326_63+m327_63+m328_63+m329_63+m330_63+m331_63+m332_63+m333_63+m334_63+m335_63+m336_63+m337_63+m338_63+m339_63+m340_63+m341_63+m342_63+m343_63+m344_63+m345_63+m346_63+m347_63+m348_63+m349_63+m350_63+m351_63+m352_63+m353_63+m354_63+m355_63+m356_63+m357_63+m358_63+m359_63+m360_63+m361_63+m362_63+m363_63+m364_63+m365_63+m366_63+m367_63+m368_63+m369_63+m370_63+m371_63+m372_63+m373_63+m374_63+m375_63+m376_63+m377_63+m378_63+m379_63+m380_63+m381_63+b63;
   always @(posedge clk) out64 <= m1_64+m2_64+m3_64+m4_64+m5_64+m6_64+m7_64+m8_64+m9_64+m10_64+m11_64+m12_64+m13_64+m14_64+m15_64+m16_64+m17_64+m18_64+m19_64+m20_64+m21_64+m22_64+m23_64+m24_64+m25_64+m26_64+m27_64+m28_64+m29_64+m30_64+m31_64+m32_64+m33_64+m34_64+m35_64+m36_64+m37_64+m38_64+m39_64+m40_64+m41_64+m42_64+m43_64+m44_64+m45_64+m46_64+m47_64+m48_64+m49_64+m50_64+m51_64+m52_64+m53_64+m54_64+m55_64+m56_64+m57_64+m58_64+m59_64+m60_64+m61_64+m62_64+m63_64+m64_64+m65_64+m66_64+m67_64+m68_64+m69_64+m70_64+m71_64+m72_64+m73_64+m74_64+m75_64+m76_64+m77_64+m78_64+m79_64+m80_64+m81_64+m82_64+m83_64+m84_64+m85_64+m86_64+m87_64+m88_64+m89_64+m90_64+m91_64+m92_64+m93_64+m94_64+m95_64+m96_64+m97_64+m98_64+m99_64+m100_64+m101_64+m102_64+m103_64+m104_64+m105_64+m106_64+m107_64+m108_64+m109_64+m110_64+m111_64+m112_64+m113_64+m114_64+m115_64+m116_64+m117_64+m118_64+m119_64+m120_64+m121_64+m122_64+m123_64+m124_64+m125_64+m126_64+m127_64+m128_64+m129_64+m130_64+m131_64+m132_64+m133_64+m134_64+m135_64+m136_64+m137_64+m138_64+m139_64+m140_64+m141_64+m142_64+m143_64+m144_64+m145_64+m146_64+m147_64+m148_64+m149_64+m150_64+m151_64+m152_64+m153_64+m154_64+m155_64+m156_64+m157_64+m158_64+m159_64+m160_64+m161_64+m162_64+m163_64+m164_64+m165_64+m166_64+m167_64+m168_64+m169_64+m170_64+m171_64+m172_64+m173_64+m174_64+m175_64+m176_64+m177_64+m178_64+m179_64+m180_64+m181_64+m182_64+m183_64+m184_64+m185_64+m186_64+m187_64+m188_64+m189_64+m190_64+m191_64+m192_64+m193_64+m194_64+m195_64+m196_64+m197_64+m198_64+m199_64+m200_64+m201_64+m202_64+m203_64+m204_64+m205_64+m206_64+m207_64+m208_64+m209_64+m210_64+m211_64+m212_64+m213_64+m214_64+m215_64+m216_64+m217_64+m218_64+m219_64+m220_64+m221_64+m222_64+m223_64+m224_64+m225_64+m226_64+m227_64+m228_64+m229_64+m230_64+m231_64+m232_64+m233_64+m234_64+m235_64+m236_64+m237_64+m238_64+m239_64+m240_64+m241_64+m242_64+m243_64+m244_64+m245_64+m246_64+m247_64+m248_64+m249_64+m250_64+m251_64+m252_64+m253_64+m254_64+m255_64+m256_64+m257_64+m258_64+m259_64+m260_64+m261_64+m262_64+m263_64+m264_64+m265_64+m266_64+m267_64+m268_64+m269_64+m270_64+m271_64+m272_64+m273_64+m274_64+m275_64+m276_64+m277_64+m278_64+m279_64+m280_64+m281_64+m282_64+m283_64+m284_64+m285_64+m286_64+m287_64+m288_64+m289_64+m290_64+m291_64+m292_64+m293_64+m294_64+m295_64+m296_64+m297_64+m298_64+m299_64+m300_64+m301_64+m302_64+m303_64+m304_64+m305_64+m306_64+m307_64+m308_64+m309_64+m310_64+m311_64+m312_64+m313_64+m314_64+m315_64+m316_64+m317_64+m318_64+m319_64+m320_64+m321_64+m322_64+m323_64+m324_64+m325_64+m326_64+m327_64+m328_64+m329_64+m330_64+m331_64+m332_64+m333_64+m334_64+m335_64+m336_64+m337_64+m338_64+m339_64+m340_64+m341_64+m342_64+m343_64+m344_64+m345_64+m346_64+m347_64+m348_64+m349_64+m350_64+m351_64+m352_64+m353_64+m354_64+m355_64+m356_64+m357_64+m358_64+m359_64+m360_64+m361_64+m362_64+m363_64+m364_64+m365_64+m366_64+m367_64+m368_64+m369_64+m370_64+m371_64+m372_64+m373_64+m374_64+m375_64+m376_64+m377_64+m378_64+m379_64+m380_64+m381_64+b64;
   always @(posedge clk) out65 <= m1_65+m2_65+m3_65+m4_65+m5_65+m6_65+m7_65+m8_65+m9_65+m10_65+m11_65+m12_65+m13_65+m14_65+m15_65+m16_65+m17_65+m18_65+m19_65+m20_65+m21_65+m22_65+m23_65+m24_65+m25_65+m26_65+m27_65+m28_65+m29_65+m30_65+m31_65+m32_65+m33_65+m34_65+m35_65+m36_65+m37_65+m38_65+m39_65+m40_65+m41_65+m42_65+m43_65+m44_65+m45_65+m46_65+m47_65+m48_65+m49_65+m50_65+m51_65+m52_65+m53_65+m54_65+m55_65+m56_65+m57_65+m58_65+m59_65+m60_65+m61_65+m62_65+m63_65+m64_65+m65_65+m66_65+m67_65+m68_65+m69_65+m70_65+m71_65+m72_65+m73_65+m74_65+m75_65+m76_65+m77_65+m78_65+m79_65+m80_65+m81_65+m82_65+m83_65+m84_65+m85_65+m86_65+m87_65+m88_65+m89_65+m90_65+m91_65+m92_65+m93_65+m94_65+m95_65+m96_65+m97_65+m98_65+m99_65+m100_65+m101_65+m102_65+m103_65+m104_65+m105_65+m106_65+m107_65+m108_65+m109_65+m110_65+m111_65+m112_65+m113_65+m114_65+m115_65+m116_65+m117_65+m118_65+m119_65+m120_65+m121_65+m122_65+m123_65+m124_65+m125_65+m126_65+m127_65+m128_65+m129_65+m130_65+m131_65+m132_65+m133_65+m134_65+m135_65+m136_65+m137_65+m138_65+m139_65+m140_65+m141_65+m142_65+m143_65+m144_65+m145_65+m146_65+m147_65+m148_65+m149_65+m150_65+m151_65+m152_65+m153_65+m154_65+m155_65+m156_65+m157_65+m158_65+m159_65+m160_65+m161_65+m162_65+m163_65+m164_65+m165_65+m166_65+m167_65+m168_65+m169_65+m170_65+m171_65+m172_65+m173_65+m174_65+m175_65+m176_65+m177_65+m178_65+m179_65+m180_65+m181_65+m182_65+m183_65+m184_65+m185_65+m186_65+m187_65+m188_65+m189_65+m190_65+m191_65+m192_65+m193_65+m194_65+m195_65+m196_65+m197_65+m198_65+m199_65+m200_65+m201_65+m202_65+m203_65+m204_65+m205_65+m206_65+m207_65+m208_65+m209_65+m210_65+m211_65+m212_65+m213_65+m214_65+m215_65+m216_65+m217_65+m218_65+m219_65+m220_65+m221_65+m222_65+m223_65+m224_65+m225_65+m226_65+m227_65+m228_65+m229_65+m230_65+m231_65+m232_65+m233_65+m234_65+m235_65+m236_65+m237_65+m238_65+m239_65+m240_65+m241_65+m242_65+m243_65+m244_65+m245_65+m246_65+m247_65+m248_65+m249_65+m250_65+m251_65+m252_65+m253_65+m254_65+m255_65+m256_65+m257_65+m258_65+m259_65+m260_65+m261_65+m262_65+m263_65+m264_65+m265_65+m266_65+m267_65+m268_65+m269_65+m270_65+m271_65+m272_65+m273_65+m274_65+m275_65+m276_65+m277_65+m278_65+m279_65+m280_65+m281_65+m282_65+m283_65+m284_65+m285_65+m286_65+m287_65+m288_65+m289_65+m290_65+m291_65+m292_65+m293_65+m294_65+m295_65+m296_65+m297_65+m298_65+m299_65+m300_65+m301_65+m302_65+m303_65+m304_65+m305_65+m306_65+m307_65+m308_65+m309_65+m310_65+m311_65+m312_65+m313_65+m314_65+m315_65+m316_65+m317_65+m318_65+m319_65+m320_65+m321_65+m322_65+m323_65+m324_65+m325_65+m326_65+m327_65+m328_65+m329_65+m330_65+m331_65+m332_65+m333_65+m334_65+m335_65+m336_65+m337_65+m338_65+m339_65+m340_65+m341_65+m342_65+m343_65+m344_65+m345_65+m346_65+m347_65+m348_65+m349_65+m350_65+m351_65+m352_65+m353_65+m354_65+m355_65+m356_65+m357_65+m358_65+m359_65+m360_65+m361_65+m362_65+m363_65+m364_65+m365_65+m366_65+m367_65+m368_65+m369_65+m370_65+m371_65+m372_65+m373_65+m374_65+m375_65+m376_65+m377_65+m378_65+m379_65+m380_65+m381_65+b65;
   always @(posedge clk) out66 <= m1_66+m2_66+m3_66+m4_66+m5_66+m6_66+m7_66+m8_66+m9_66+m10_66+m11_66+m12_66+m13_66+m14_66+m15_66+m16_66+m17_66+m18_66+m19_66+m20_66+m21_66+m22_66+m23_66+m24_66+m25_66+m26_66+m27_66+m28_66+m29_66+m30_66+m31_66+m32_66+m33_66+m34_66+m35_66+m36_66+m37_66+m38_66+m39_66+m40_66+m41_66+m42_66+m43_66+m44_66+m45_66+m46_66+m47_66+m48_66+m49_66+m50_66+m51_66+m52_66+m53_66+m54_66+m55_66+m56_66+m57_66+m58_66+m59_66+m60_66+m61_66+m62_66+m63_66+m64_66+m65_66+m66_66+m67_66+m68_66+m69_66+m70_66+m71_66+m72_66+m73_66+m74_66+m75_66+m76_66+m77_66+m78_66+m79_66+m80_66+m81_66+m82_66+m83_66+m84_66+m85_66+m86_66+m87_66+m88_66+m89_66+m90_66+m91_66+m92_66+m93_66+m94_66+m95_66+m96_66+m97_66+m98_66+m99_66+m100_66+m101_66+m102_66+m103_66+m104_66+m105_66+m106_66+m107_66+m108_66+m109_66+m110_66+m111_66+m112_66+m113_66+m114_66+m115_66+m116_66+m117_66+m118_66+m119_66+m120_66+m121_66+m122_66+m123_66+m124_66+m125_66+m126_66+m127_66+m128_66+m129_66+m130_66+m131_66+m132_66+m133_66+m134_66+m135_66+m136_66+m137_66+m138_66+m139_66+m140_66+m141_66+m142_66+m143_66+m144_66+m145_66+m146_66+m147_66+m148_66+m149_66+m150_66+m151_66+m152_66+m153_66+m154_66+m155_66+m156_66+m157_66+m158_66+m159_66+m160_66+m161_66+m162_66+m163_66+m164_66+m165_66+m166_66+m167_66+m168_66+m169_66+m170_66+m171_66+m172_66+m173_66+m174_66+m175_66+m176_66+m177_66+m178_66+m179_66+m180_66+m181_66+m182_66+m183_66+m184_66+m185_66+m186_66+m187_66+m188_66+m189_66+m190_66+m191_66+m192_66+m193_66+m194_66+m195_66+m196_66+m197_66+m198_66+m199_66+m200_66+m201_66+m202_66+m203_66+m204_66+m205_66+m206_66+m207_66+m208_66+m209_66+m210_66+m211_66+m212_66+m213_66+m214_66+m215_66+m216_66+m217_66+m218_66+m219_66+m220_66+m221_66+m222_66+m223_66+m224_66+m225_66+m226_66+m227_66+m228_66+m229_66+m230_66+m231_66+m232_66+m233_66+m234_66+m235_66+m236_66+m237_66+m238_66+m239_66+m240_66+m241_66+m242_66+m243_66+m244_66+m245_66+m246_66+m247_66+m248_66+m249_66+m250_66+m251_66+m252_66+m253_66+m254_66+m255_66+m256_66+m257_66+m258_66+m259_66+m260_66+m261_66+m262_66+m263_66+m264_66+m265_66+m266_66+m267_66+m268_66+m269_66+m270_66+m271_66+m272_66+m273_66+m274_66+m275_66+m276_66+m277_66+m278_66+m279_66+m280_66+m281_66+m282_66+m283_66+m284_66+m285_66+m286_66+m287_66+m288_66+m289_66+m290_66+m291_66+m292_66+m293_66+m294_66+m295_66+m296_66+m297_66+m298_66+m299_66+m300_66+m301_66+m302_66+m303_66+m304_66+m305_66+m306_66+m307_66+m308_66+m309_66+m310_66+m311_66+m312_66+m313_66+m314_66+m315_66+m316_66+m317_66+m318_66+m319_66+m320_66+m321_66+m322_66+m323_66+m324_66+m325_66+m326_66+m327_66+m328_66+m329_66+m330_66+m331_66+m332_66+m333_66+m334_66+m335_66+m336_66+m337_66+m338_66+m339_66+m340_66+m341_66+m342_66+m343_66+m344_66+m345_66+m346_66+m347_66+m348_66+m349_66+m350_66+m351_66+m352_66+m353_66+m354_66+m355_66+m356_66+m357_66+m358_66+m359_66+m360_66+m361_66+m362_66+m363_66+m364_66+m365_66+m366_66+m367_66+m368_66+m369_66+m370_66+m371_66+m372_66+m373_66+m374_66+m375_66+m376_66+m377_66+m378_66+m379_66+m380_66+m381_66+b66;
   always @(posedge clk) out67 <= m1_67+m2_67+m3_67+m4_67+m5_67+m6_67+m7_67+m8_67+m9_67+m10_67+m11_67+m12_67+m13_67+m14_67+m15_67+m16_67+m17_67+m18_67+m19_67+m20_67+m21_67+m22_67+m23_67+m24_67+m25_67+m26_67+m27_67+m28_67+m29_67+m30_67+m31_67+m32_67+m33_67+m34_67+m35_67+m36_67+m37_67+m38_67+m39_67+m40_67+m41_67+m42_67+m43_67+m44_67+m45_67+m46_67+m47_67+m48_67+m49_67+m50_67+m51_67+m52_67+m53_67+m54_67+m55_67+m56_67+m57_67+m58_67+m59_67+m60_67+m61_67+m62_67+m63_67+m64_67+m65_67+m66_67+m67_67+m68_67+m69_67+m70_67+m71_67+m72_67+m73_67+m74_67+m75_67+m76_67+m77_67+m78_67+m79_67+m80_67+m81_67+m82_67+m83_67+m84_67+m85_67+m86_67+m87_67+m88_67+m89_67+m90_67+m91_67+m92_67+m93_67+m94_67+m95_67+m96_67+m97_67+m98_67+m99_67+m100_67+m101_67+m102_67+m103_67+m104_67+m105_67+m106_67+m107_67+m108_67+m109_67+m110_67+m111_67+m112_67+m113_67+m114_67+m115_67+m116_67+m117_67+m118_67+m119_67+m120_67+m121_67+m122_67+m123_67+m124_67+m125_67+m126_67+m127_67+m128_67+m129_67+m130_67+m131_67+m132_67+m133_67+m134_67+m135_67+m136_67+m137_67+m138_67+m139_67+m140_67+m141_67+m142_67+m143_67+m144_67+m145_67+m146_67+m147_67+m148_67+m149_67+m150_67+m151_67+m152_67+m153_67+m154_67+m155_67+m156_67+m157_67+m158_67+m159_67+m160_67+m161_67+m162_67+m163_67+m164_67+m165_67+m166_67+m167_67+m168_67+m169_67+m170_67+m171_67+m172_67+m173_67+m174_67+m175_67+m176_67+m177_67+m178_67+m179_67+m180_67+m181_67+m182_67+m183_67+m184_67+m185_67+m186_67+m187_67+m188_67+m189_67+m190_67+m191_67+m192_67+m193_67+m194_67+m195_67+m196_67+m197_67+m198_67+m199_67+m200_67+m201_67+m202_67+m203_67+m204_67+m205_67+m206_67+m207_67+m208_67+m209_67+m210_67+m211_67+m212_67+m213_67+m214_67+m215_67+m216_67+m217_67+m218_67+m219_67+m220_67+m221_67+m222_67+m223_67+m224_67+m225_67+m226_67+m227_67+m228_67+m229_67+m230_67+m231_67+m232_67+m233_67+m234_67+m235_67+m236_67+m237_67+m238_67+m239_67+m240_67+m241_67+m242_67+m243_67+m244_67+m245_67+m246_67+m247_67+m248_67+m249_67+m250_67+m251_67+m252_67+m253_67+m254_67+m255_67+m256_67+m257_67+m258_67+m259_67+m260_67+m261_67+m262_67+m263_67+m264_67+m265_67+m266_67+m267_67+m268_67+m269_67+m270_67+m271_67+m272_67+m273_67+m274_67+m275_67+m276_67+m277_67+m278_67+m279_67+m280_67+m281_67+m282_67+m283_67+m284_67+m285_67+m286_67+m287_67+m288_67+m289_67+m290_67+m291_67+m292_67+m293_67+m294_67+m295_67+m296_67+m297_67+m298_67+m299_67+m300_67+m301_67+m302_67+m303_67+m304_67+m305_67+m306_67+m307_67+m308_67+m309_67+m310_67+m311_67+m312_67+m313_67+m314_67+m315_67+m316_67+m317_67+m318_67+m319_67+m320_67+m321_67+m322_67+m323_67+m324_67+m325_67+m326_67+m327_67+m328_67+m329_67+m330_67+m331_67+m332_67+m333_67+m334_67+m335_67+m336_67+m337_67+m338_67+m339_67+m340_67+m341_67+m342_67+m343_67+m344_67+m345_67+m346_67+m347_67+m348_67+m349_67+m350_67+m351_67+m352_67+m353_67+m354_67+m355_67+m356_67+m357_67+m358_67+m359_67+m360_67+m361_67+m362_67+m363_67+m364_67+m365_67+m366_67+m367_67+m368_67+m369_67+m370_67+m371_67+m372_67+m373_67+m374_67+m375_67+m376_67+m377_67+m378_67+m379_67+m380_67+m381_67+b67;
   always @(posedge clk) out68 <= m1_68+m2_68+m3_68+m4_68+m5_68+m6_68+m7_68+m8_68+m9_68+m10_68+m11_68+m12_68+m13_68+m14_68+m15_68+m16_68+m17_68+m18_68+m19_68+m20_68+m21_68+m22_68+m23_68+m24_68+m25_68+m26_68+m27_68+m28_68+m29_68+m30_68+m31_68+m32_68+m33_68+m34_68+m35_68+m36_68+m37_68+m38_68+m39_68+m40_68+m41_68+m42_68+m43_68+m44_68+m45_68+m46_68+m47_68+m48_68+m49_68+m50_68+m51_68+m52_68+m53_68+m54_68+m55_68+m56_68+m57_68+m58_68+m59_68+m60_68+m61_68+m62_68+m63_68+m64_68+m65_68+m66_68+m67_68+m68_68+m69_68+m70_68+m71_68+m72_68+m73_68+m74_68+m75_68+m76_68+m77_68+m78_68+m79_68+m80_68+m81_68+m82_68+m83_68+m84_68+m85_68+m86_68+m87_68+m88_68+m89_68+m90_68+m91_68+m92_68+m93_68+m94_68+m95_68+m96_68+m97_68+m98_68+m99_68+m100_68+m101_68+m102_68+m103_68+m104_68+m105_68+m106_68+m107_68+m108_68+m109_68+m110_68+m111_68+m112_68+m113_68+m114_68+m115_68+m116_68+m117_68+m118_68+m119_68+m120_68+m121_68+m122_68+m123_68+m124_68+m125_68+m126_68+m127_68+m128_68+m129_68+m130_68+m131_68+m132_68+m133_68+m134_68+m135_68+m136_68+m137_68+m138_68+m139_68+m140_68+m141_68+m142_68+m143_68+m144_68+m145_68+m146_68+m147_68+m148_68+m149_68+m150_68+m151_68+m152_68+m153_68+m154_68+m155_68+m156_68+m157_68+m158_68+m159_68+m160_68+m161_68+m162_68+m163_68+m164_68+m165_68+m166_68+m167_68+m168_68+m169_68+m170_68+m171_68+m172_68+m173_68+m174_68+m175_68+m176_68+m177_68+m178_68+m179_68+m180_68+m181_68+m182_68+m183_68+m184_68+m185_68+m186_68+m187_68+m188_68+m189_68+m190_68+m191_68+m192_68+m193_68+m194_68+m195_68+m196_68+m197_68+m198_68+m199_68+m200_68+m201_68+m202_68+m203_68+m204_68+m205_68+m206_68+m207_68+m208_68+m209_68+m210_68+m211_68+m212_68+m213_68+m214_68+m215_68+m216_68+m217_68+m218_68+m219_68+m220_68+m221_68+m222_68+m223_68+m224_68+m225_68+m226_68+m227_68+m228_68+m229_68+m230_68+m231_68+m232_68+m233_68+m234_68+m235_68+m236_68+m237_68+m238_68+m239_68+m240_68+m241_68+m242_68+m243_68+m244_68+m245_68+m246_68+m247_68+m248_68+m249_68+m250_68+m251_68+m252_68+m253_68+m254_68+m255_68+m256_68+m257_68+m258_68+m259_68+m260_68+m261_68+m262_68+m263_68+m264_68+m265_68+m266_68+m267_68+m268_68+m269_68+m270_68+m271_68+m272_68+m273_68+m274_68+m275_68+m276_68+m277_68+m278_68+m279_68+m280_68+m281_68+m282_68+m283_68+m284_68+m285_68+m286_68+m287_68+m288_68+m289_68+m290_68+m291_68+m292_68+m293_68+m294_68+m295_68+m296_68+m297_68+m298_68+m299_68+m300_68+m301_68+m302_68+m303_68+m304_68+m305_68+m306_68+m307_68+m308_68+m309_68+m310_68+m311_68+m312_68+m313_68+m314_68+m315_68+m316_68+m317_68+m318_68+m319_68+m320_68+m321_68+m322_68+m323_68+m324_68+m325_68+m326_68+m327_68+m328_68+m329_68+m330_68+m331_68+m332_68+m333_68+m334_68+m335_68+m336_68+m337_68+m338_68+m339_68+m340_68+m341_68+m342_68+m343_68+m344_68+m345_68+m346_68+m347_68+m348_68+m349_68+m350_68+m351_68+m352_68+m353_68+m354_68+m355_68+m356_68+m357_68+m358_68+m359_68+m360_68+m361_68+m362_68+m363_68+m364_68+m365_68+m366_68+m367_68+m368_68+m369_68+m370_68+m371_68+m372_68+m373_68+m374_68+m375_68+m376_68+m377_68+m378_68+m379_68+m380_68+m381_68+b68;
   always @(posedge clk) out69 <= m1_69+m2_69+m3_69+m4_69+m5_69+m6_69+m7_69+m8_69+m9_69+m10_69+m11_69+m12_69+m13_69+m14_69+m15_69+m16_69+m17_69+m18_69+m19_69+m20_69+m21_69+m22_69+m23_69+m24_69+m25_69+m26_69+m27_69+m28_69+m29_69+m30_69+m31_69+m32_69+m33_69+m34_69+m35_69+m36_69+m37_69+m38_69+m39_69+m40_69+m41_69+m42_69+m43_69+m44_69+m45_69+m46_69+m47_69+m48_69+m49_69+m50_69+m51_69+m52_69+m53_69+m54_69+m55_69+m56_69+m57_69+m58_69+m59_69+m60_69+m61_69+m62_69+m63_69+m64_69+m65_69+m66_69+m67_69+m68_69+m69_69+m70_69+m71_69+m72_69+m73_69+m74_69+m75_69+m76_69+m77_69+m78_69+m79_69+m80_69+m81_69+m82_69+m83_69+m84_69+m85_69+m86_69+m87_69+m88_69+m89_69+m90_69+m91_69+m92_69+m93_69+m94_69+m95_69+m96_69+m97_69+m98_69+m99_69+m100_69+m101_69+m102_69+m103_69+m104_69+m105_69+m106_69+m107_69+m108_69+m109_69+m110_69+m111_69+m112_69+m113_69+m114_69+m115_69+m116_69+m117_69+m118_69+m119_69+m120_69+m121_69+m122_69+m123_69+m124_69+m125_69+m126_69+m127_69+m128_69+m129_69+m130_69+m131_69+m132_69+m133_69+m134_69+m135_69+m136_69+m137_69+m138_69+m139_69+m140_69+m141_69+m142_69+m143_69+m144_69+m145_69+m146_69+m147_69+m148_69+m149_69+m150_69+m151_69+m152_69+m153_69+m154_69+m155_69+m156_69+m157_69+m158_69+m159_69+m160_69+m161_69+m162_69+m163_69+m164_69+m165_69+m166_69+m167_69+m168_69+m169_69+m170_69+m171_69+m172_69+m173_69+m174_69+m175_69+m176_69+m177_69+m178_69+m179_69+m180_69+m181_69+m182_69+m183_69+m184_69+m185_69+m186_69+m187_69+m188_69+m189_69+m190_69+m191_69+m192_69+m193_69+m194_69+m195_69+m196_69+m197_69+m198_69+m199_69+m200_69+m201_69+m202_69+m203_69+m204_69+m205_69+m206_69+m207_69+m208_69+m209_69+m210_69+m211_69+m212_69+m213_69+m214_69+m215_69+m216_69+m217_69+m218_69+m219_69+m220_69+m221_69+m222_69+m223_69+m224_69+m225_69+m226_69+m227_69+m228_69+m229_69+m230_69+m231_69+m232_69+m233_69+m234_69+m235_69+m236_69+m237_69+m238_69+m239_69+m240_69+m241_69+m242_69+m243_69+m244_69+m245_69+m246_69+m247_69+m248_69+m249_69+m250_69+m251_69+m252_69+m253_69+m254_69+m255_69+m256_69+m257_69+m258_69+m259_69+m260_69+m261_69+m262_69+m263_69+m264_69+m265_69+m266_69+m267_69+m268_69+m269_69+m270_69+m271_69+m272_69+m273_69+m274_69+m275_69+m276_69+m277_69+m278_69+m279_69+m280_69+m281_69+m282_69+m283_69+m284_69+m285_69+m286_69+m287_69+m288_69+m289_69+m290_69+m291_69+m292_69+m293_69+m294_69+m295_69+m296_69+m297_69+m298_69+m299_69+m300_69+m301_69+m302_69+m303_69+m304_69+m305_69+m306_69+m307_69+m308_69+m309_69+m310_69+m311_69+m312_69+m313_69+m314_69+m315_69+m316_69+m317_69+m318_69+m319_69+m320_69+m321_69+m322_69+m323_69+m324_69+m325_69+m326_69+m327_69+m328_69+m329_69+m330_69+m331_69+m332_69+m333_69+m334_69+m335_69+m336_69+m337_69+m338_69+m339_69+m340_69+m341_69+m342_69+m343_69+m344_69+m345_69+m346_69+m347_69+m348_69+m349_69+m350_69+m351_69+m352_69+m353_69+m354_69+m355_69+m356_69+m357_69+m358_69+m359_69+m360_69+m361_69+m362_69+m363_69+m364_69+m365_69+m366_69+m367_69+m368_69+m369_69+m370_69+m371_69+m372_69+m373_69+m374_69+m375_69+m376_69+m377_69+m378_69+m379_69+m380_69+m381_69+b69;
   always @(posedge clk) out70 <= m1_70+m2_70+m3_70+m4_70+m5_70+m6_70+m7_70+m8_70+m9_70+m10_70+m11_70+m12_70+m13_70+m14_70+m15_70+m16_70+m17_70+m18_70+m19_70+m20_70+m21_70+m22_70+m23_70+m24_70+m25_70+m26_70+m27_70+m28_70+m29_70+m30_70+m31_70+m32_70+m33_70+m34_70+m35_70+m36_70+m37_70+m38_70+m39_70+m40_70+m41_70+m42_70+m43_70+m44_70+m45_70+m46_70+m47_70+m48_70+m49_70+m50_70+m51_70+m52_70+m53_70+m54_70+m55_70+m56_70+m57_70+m58_70+m59_70+m60_70+m61_70+m62_70+m63_70+m64_70+m65_70+m66_70+m67_70+m68_70+m69_70+m70_70+m71_70+m72_70+m73_70+m74_70+m75_70+m76_70+m77_70+m78_70+m79_70+m80_70+m81_70+m82_70+m83_70+m84_70+m85_70+m86_70+m87_70+m88_70+m89_70+m90_70+m91_70+m92_70+m93_70+m94_70+m95_70+m96_70+m97_70+m98_70+m99_70+m100_70+m101_70+m102_70+m103_70+m104_70+m105_70+m106_70+m107_70+m108_70+m109_70+m110_70+m111_70+m112_70+m113_70+m114_70+m115_70+m116_70+m117_70+m118_70+m119_70+m120_70+m121_70+m122_70+m123_70+m124_70+m125_70+m126_70+m127_70+m128_70+m129_70+m130_70+m131_70+m132_70+m133_70+m134_70+m135_70+m136_70+m137_70+m138_70+m139_70+m140_70+m141_70+m142_70+m143_70+m144_70+m145_70+m146_70+m147_70+m148_70+m149_70+m150_70+m151_70+m152_70+m153_70+m154_70+m155_70+m156_70+m157_70+m158_70+m159_70+m160_70+m161_70+m162_70+m163_70+m164_70+m165_70+m166_70+m167_70+m168_70+m169_70+m170_70+m171_70+m172_70+m173_70+m174_70+m175_70+m176_70+m177_70+m178_70+m179_70+m180_70+m181_70+m182_70+m183_70+m184_70+m185_70+m186_70+m187_70+m188_70+m189_70+m190_70+m191_70+m192_70+m193_70+m194_70+m195_70+m196_70+m197_70+m198_70+m199_70+m200_70+m201_70+m202_70+m203_70+m204_70+m205_70+m206_70+m207_70+m208_70+m209_70+m210_70+m211_70+m212_70+m213_70+m214_70+m215_70+m216_70+m217_70+m218_70+m219_70+m220_70+m221_70+m222_70+m223_70+m224_70+m225_70+m226_70+m227_70+m228_70+m229_70+m230_70+m231_70+m232_70+m233_70+m234_70+m235_70+m236_70+m237_70+m238_70+m239_70+m240_70+m241_70+m242_70+m243_70+m244_70+m245_70+m246_70+m247_70+m248_70+m249_70+m250_70+m251_70+m252_70+m253_70+m254_70+m255_70+m256_70+m257_70+m258_70+m259_70+m260_70+m261_70+m262_70+m263_70+m264_70+m265_70+m266_70+m267_70+m268_70+m269_70+m270_70+m271_70+m272_70+m273_70+m274_70+m275_70+m276_70+m277_70+m278_70+m279_70+m280_70+m281_70+m282_70+m283_70+m284_70+m285_70+m286_70+m287_70+m288_70+m289_70+m290_70+m291_70+m292_70+m293_70+m294_70+m295_70+m296_70+m297_70+m298_70+m299_70+m300_70+m301_70+m302_70+m303_70+m304_70+m305_70+m306_70+m307_70+m308_70+m309_70+m310_70+m311_70+m312_70+m313_70+m314_70+m315_70+m316_70+m317_70+m318_70+m319_70+m320_70+m321_70+m322_70+m323_70+m324_70+m325_70+m326_70+m327_70+m328_70+m329_70+m330_70+m331_70+m332_70+m333_70+m334_70+m335_70+m336_70+m337_70+m338_70+m339_70+m340_70+m341_70+m342_70+m343_70+m344_70+m345_70+m346_70+m347_70+m348_70+m349_70+m350_70+m351_70+m352_70+m353_70+m354_70+m355_70+m356_70+m357_70+m358_70+m359_70+m360_70+m361_70+m362_70+m363_70+m364_70+m365_70+m366_70+m367_70+m368_70+m369_70+m370_70+m371_70+m372_70+m373_70+m374_70+m375_70+m376_70+m377_70+m378_70+m379_70+m380_70+m381_70+b70;
   always @(posedge clk) out71 <= m1_71+m2_71+m3_71+m4_71+m5_71+m6_71+m7_71+m8_71+m9_71+m10_71+m11_71+m12_71+m13_71+m14_71+m15_71+m16_71+m17_71+m18_71+m19_71+m20_71+m21_71+m22_71+m23_71+m24_71+m25_71+m26_71+m27_71+m28_71+m29_71+m30_71+m31_71+m32_71+m33_71+m34_71+m35_71+m36_71+m37_71+m38_71+m39_71+m40_71+m41_71+m42_71+m43_71+m44_71+m45_71+m46_71+m47_71+m48_71+m49_71+m50_71+m51_71+m52_71+m53_71+m54_71+m55_71+m56_71+m57_71+m58_71+m59_71+m60_71+m61_71+m62_71+m63_71+m64_71+m65_71+m66_71+m67_71+m68_71+m69_71+m70_71+m71_71+m72_71+m73_71+m74_71+m75_71+m76_71+m77_71+m78_71+m79_71+m80_71+m81_71+m82_71+m83_71+m84_71+m85_71+m86_71+m87_71+m88_71+m89_71+m90_71+m91_71+m92_71+m93_71+m94_71+m95_71+m96_71+m97_71+m98_71+m99_71+m100_71+m101_71+m102_71+m103_71+m104_71+m105_71+m106_71+m107_71+m108_71+m109_71+m110_71+m111_71+m112_71+m113_71+m114_71+m115_71+m116_71+m117_71+m118_71+m119_71+m120_71+m121_71+m122_71+m123_71+m124_71+m125_71+m126_71+m127_71+m128_71+m129_71+m130_71+m131_71+m132_71+m133_71+m134_71+m135_71+m136_71+m137_71+m138_71+m139_71+m140_71+m141_71+m142_71+m143_71+m144_71+m145_71+m146_71+m147_71+m148_71+m149_71+m150_71+m151_71+m152_71+m153_71+m154_71+m155_71+m156_71+m157_71+m158_71+m159_71+m160_71+m161_71+m162_71+m163_71+m164_71+m165_71+m166_71+m167_71+m168_71+m169_71+m170_71+m171_71+m172_71+m173_71+m174_71+m175_71+m176_71+m177_71+m178_71+m179_71+m180_71+m181_71+m182_71+m183_71+m184_71+m185_71+m186_71+m187_71+m188_71+m189_71+m190_71+m191_71+m192_71+m193_71+m194_71+m195_71+m196_71+m197_71+m198_71+m199_71+m200_71+m201_71+m202_71+m203_71+m204_71+m205_71+m206_71+m207_71+m208_71+m209_71+m210_71+m211_71+m212_71+m213_71+m214_71+m215_71+m216_71+m217_71+m218_71+m219_71+m220_71+m221_71+m222_71+m223_71+m224_71+m225_71+m226_71+m227_71+m228_71+m229_71+m230_71+m231_71+m232_71+m233_71+m234_71+m235_71+m236_71+m237_71+m238_71+m239_71+m240_71+m241_71+m242_71+m243_71+m244_71+m245_71+m246_71+m247_71+m248_71+m249_71+m250_71+m251_71+m252_71+m253_71+m254_71+m255_71+m256_71+m257_71+m258_71+m259_71+m260_71+m261_71+m262_71+m263_71+m264_71+m265_71+m266_71+m267_71+m268_71+m269_71+m270_71+m271_71+m272_71+m273_71+m274_71+m275_71+m276_71+m277_71+m278_71+m279_71+m280_71+m281_71+m282_71+m283_71+m284_71+m285_71+m286_71+m287_71+m288_71+m289_71+m290_71+m291_71+m292_71+m293_71+m294_71+m295_71+m296_71+m297_71+m298_71+m299_71+m300_71+m301_71+m302_71+m303_71+m304_71+m305_71+m306_71+m307_71+m308_71+m309_71+m310_71+m311_71+m312_71+m313_71+m314_71+m315_71+m316_71+m317_71+m318_71+m319_71+m320_71+m321_71+m322_71+m323_71+m324_71+m325_71+m326_71+m327_71+m328_71+m329_71+m330_71+m331_71+m332_71+m333_71+m334_71+m335_71+m336_71+m337_71+m338_71+m339_71+m340_71+m341_71+m342_71+m343_71+m344_71+m345_71+m346_71+m347_71+m348_71+m349_71+m350_71+m351_71+m352_71+m353_71+m354_71+m355_71+m356_71+m357_71+m358_71+m359_71+m360_71+m361_71+m362_71+m363_71+m364_71+m365_71+m366_71+m367_71+m368_71+m369_71+m370_71+m371_71+m372_71+m373_71+m374_71+m375_71+m376_71+m377_71+m378_71+m379_71+m380_71+m381_71+b71;
   always @(posedge clk) out72 <= m1_72+m2_72+m3_72+m4_72+m5_72+m6_72+m7_72+m8_72+m9_72+m10_72+m11_72+m12_72+m13_72+m14_72+m15_72+m16_72+m17_72+m18_72+m19_72+m20_72+m21_72+m22_72+m23_72+m24_72+m25_72+m26_72+m27_72+m28_72+m29_72+m30_72+m31_72+m32_72+m33_72+m34_72+m35_72+m36_72+m37_72+m38_72+m39_72+m40_72+m41_72+m42_72+m43_72+m44_72+m45_72+m46_72+m47_72+m48_72+m49_72+m50_72+m51_72+m52_72+m53_72+m54_72+m55_72+m56_72+m57_72+m58_72+m59_72+m60_72+m61_72+m62_72+m63_72+m64_72+m65_72+m66_72+m67_72+m68_72+m69_72+m70_72+m71_72+m72_72+m73_72+m74_72+m75_72+m76_72+m77_72+m78_72+m79_72+m80_72+m81_72+m82_72+m83_72+m84_72+m85_72+m86_72+m87_72+m88_72+m89_72+m90_72+m91_72+m92_72+m93_72+m94_72+m95_72+m96_72+m97_72+m98_72+m99_72+m100_72+m101_72+m102_72+m103_72+m104_72+m105_72+m106_72+m107_72+m108_72+m109_72+m110_72+m111_72+m112_72+m113_72+m114_72+m115_72+m116_72+m117_72+m118_72+m119_72+m120_72+m121_72+m122_72+m123_72+m124_72+m125_72+m126_72+m127_72+m128_72+m129_72+m130_72+m131_72+m132_72+m133_72+m134_72+m135_72+m136_72+m137_72+m138_72+m139_72+m140_72+m141_72+m142_72+m143_72+m144_72+m145_72+m146_72+m147_72+m148_72+m149_72+m150_72+m151_72+m152_72+m153_72+m154_72+m155_72+m156_72+m157_72+m158_72+m159_72+m160_72+m161_72+m162_72+m163_72+m164_72+m165_72+m166_72+m167_72+m168_72+m169_72+m170_72+m171_72+m172_72+m173_72+m174_72+m175_72+m176_72+m177_72+m178_72+m179_72+m180_72+m181_72+m182_72+m183_72+m184_72+m185_72+m186_72+m187_72+m188_72+m189_72+m190_72+m191_72+m192_72+m193_72+m194_72+m195_72+m196_72+m197_72+m198_72+m199_72+m200_72+m201_72+m202_72+m203_72+m204_72+m205_72+m206_72+m207_72+m208_72+m209_72+m210_72+m211_72+m212_72+m213_72+m214_72+m215_72+m216_72+m217_72+m218_72+m219_72+m220_72+m221_72+m222_72+m223_72+m224_72+m225_72+m226_72+m227_72+m228_72+m229_72+m230_72+m231_72+m232_72+m233_72+m234_72+m235_72+m236_72+m237_72+m238_72+m239_72+m240_72+m241_72+m242_72+m243_72+m244_72+m245_72+m246_72+m247_72+m248_72+m249_72+m250_72+m251_72+m252_72+m253_72+m254_72+m255_72+m256_72+m257_72+m258_72+m259_72+m260_72+m261_72+m262_72+m263_72+m264_72+m265_72+m266_72+m267_72+m268_72+m269_72+m270_72+m271_72+m272_72+m273_72+m274_72+m275_72+m276_72+m277_72+m278_72+m279_72+m280_72+m281_72+m282_72+m283_72+m284_72+m285_72+m286_72+m287_72+m288_72+m289_72+m290_72+m291_72+m292_72+m293_72+m294_72+m295_72+m296_72+m297_72+m298_72+m299_72+m300_72+m301_72+m302_72+m303_72+m304_72+m305_72+m306_72+m307_72+m308_72+m309_72+m310_72+m311_72+m312_72+m313_72+m314_72+m315_72+m316_72+m317_72+m318_72+m319_72+m320_72+m321_72+m322_72+m323_72+m324_72+m325_72+m326_72+m327_72+m328_72+m329_72+m330_72+m331_72+m332_72+m333_72+m334_72+m335_72+m336_72+m337_72+m338_72+m339_72+m340_72+m341_72+m342_72+m343_72+m344_72+m345_72+m346_72+m347_72+m348_72+m349_72+m350_72+m351_72+m352_72+m353_72+m354_72+m355_72+m356_72+m357_72+m358_72+m359_72+m360_72+m361_72+m362_72+m363_72+m364_72+m365_72+m366_72+m367_72+m368_72+m369_72+m370_72+m371_72+m372_72+m373_72+m374_72+m375_72+m376_72+m377_72+m378_72+m379_72+m380_72+m381_72+b72;
   always @(posedge clk) out73 <= m1_73+m2_73+m3_73+m4_73+m5_73+m6_73+m7_73+m8_73+m9_73+m10_73+m11_73+m12_73+m13_73+m14_73+m15_73+m16_73+m17_73+m18_73+m19_73+m20_73+m21_73+m22_73+m23_73+m24_73+m25_73+m26_73+m27_73+m28_73+m29_73+m30_73+m31_73+m32_73+m33_73+m34_73+m35_73+m36_73+m37_73+m38_73+m39_73+m40_73+m41_73+m42_73+m43_73+m44_73+m45_73+m46_73+m47_73+m48_73+m49_73+m50_73+m51_73+m52_73+m53_73+m54_73+m55_73+m56_73+m57_73+m58_73+m59_73+m60_73+m61_73+m62_73+m63_73+m64_73+m65_73+m66_73+m67_73+m68_73+m69_73+m70_73+m71_73+m72_73+m73_73+m74_73+m75_73+m76_73+m77_73+m78_73+m79_73+m80_73+m81_73+m82_73+m83_73+m84_73+m85_73+m86_73+m87_73+m88_73+m89_73+m90_73+m91_73+m92_73+m93_73+m94_73+m95_73+m96_73+m97_73+m98_73+m99_73+m100_73+m101_73+m102_73+m103_73+m104_73+m105_73+m106_73+m107_73+m108_73+m109_73+m110_73+m111_73+m112_73+m113_73+m114_73+m115_73+m116_73+m117_73+m118_73+m119_73+m120_73+m121_73+m122_73+m123_73+m124_73+m125_73+m126_73+m127_73+m128_73+m129_73+m130_73+m131_73+m132_73+m133_73+m134_73+m135_73+m136_73+m137_73+m138_73+m139_73+m140_73+m141_73+m142_73+m143_73+m144_73+m145_73+m146_73+m147_73+m148_73+m149_73+m150_73+m151_73+m152_73+m153_73+m154_73+m155_73+m156_73+m157_73+m158_73+m159_73+m160_73+m161_73+m162_73+m163_73+m164_73+m165_73+m166_73+m167_73+m168_73+m169_73+m170_73+m171_73+m172_73+m173_73+m174_73+m175_73+m176_73+m177_73+m178_73+m179_73+m180_73+m181_73+m182_73+m183_73+m184_73+m185_73+m186_73+m187_73+m188_73+m189_73+m190_73+m191_73+m192_73+m193_73+m194_73+m195_73+m196_73+m197_73+m198_73+m199_73+m200_73+m201_73+m202_73+m203_73+m204_73+m205_73+m206_73+m207_73+m208_73+m209_73+m210_73+m211_73+m212_73+m213_73+m214_73+m215_73+m216_73+m217_73+m218_73+m219_73+m220_73+m221_73+m222_73+m223_73+m224_73+m225_73+m226_73+m227_73+m228_73+m229_73+m230_73+m231_73+m232_73+m233_73+m234_73+m235_73+m236_73+m237_73+m238_73+m239_73+m240_73+m241_73+m242_73+m243_73+m244_73+m245_73+m246_73+m247_73+m248_73+m249_73+m250_73+m251_73+m252_73+m253_73+m254_73+m255_73+m256_73+m257_73+m258_73+m259_73+m260_73+m261_73+m262_73+m263_73+m264_73+m265_73+m266_73+m267_73+m268_73+m269_73+m270_73+m271_73+m272_73+m273_73+m274_73+m275_73+m276_73+m277_73+m278_73+m279_73+m280_73+m281_73+m282_73+m283_73+m284_73+m285_73+m286_73+m287_73+m288_73+m289_73+m290_73+m291_73+m292_73+m293_73+m294_73+m295_73+m296_73+m297_73+m298_73+m299_73+m300_73+m301_73+m302_73+m303_73+m304_73+m305_73+m306_73+m307_73+m308_73+m309_73+m310_73+m311_73+m312_73+m313_73+m314_73+m315_73+m316_73+m317_73+m318_73+m319_73+m320_73+m321_73+m322_73+m323_73+m324_73+m325_73+m326_73+m327_73+m328_73+m329_73+m330_73+m331_73+m332_73+m333_73+m334_73+m335_73+m336_73+m337_73+m338_73+m339_73+m340_73+m341_73+m342_73+m343_73+m344_73+m345_73+m346_73+m347_73+m348_73+m349_73+m350_73+m351_73+m352_73+m353_73+m354_73+m355_73+m356_73+m357_73+m358_73+m359_73+m360_73+m361_73+m362_73+m363_73+m364_73+m365_73+m366_73+m367_73+m368_73+m369_73+m370_73+m371_73+m372_73+m373_73+m374_73+m375_73+m376_73+m377_73+m378_73+m379_73+m380_73+m381_73+b73;
   always @(posedge clk) out74 <= m1_74+m2_74+m3_74+m4_74+m5_74+m6_74+m7_74+m8_74+m9_74+m10_74+m11_74+m12_74+m13_74+m14_74+m15_74+m16_74+m17_74+m18_74+m19_74+m20_74+m21_74+m22_74+m23_74+m24_74+m25_74+m26_74+m27_74+m28_74+m29_74+m30_74+m31_74+m32_74+m33_74+m34_74+m35_74+m36_74+m37_74+m38_74+m39_74+m40_74+m41_74+m42_74+m43_74+m44_74+m45_74+m46_74+m47_74+m48_74+m49_74+m50_74+m51_74+m52_74+m53_74+m54_74+m55_74+m56_74+m57_74+m58_74+m59_74+m60_74+m61_74+m62_74+m63_74+m64_74+m65_74+m66_74+m67_74+m68_74+m69_74+m70_74+m71_74+m72_74+m73_74+m74_74+m75_74+m76_74+m77_74+m78_74+m79_74+m80_74+m81_74+m82_74+m83_74+m84_74+m85_74+m86_74+m87_74+m88_74+m89_74+m90_74+m91_74+m92_74+m93_74+m94_74+m95_74+m96_74+m97_74+m98_74+m99_74+m100_74+m101_74+m102_74+m103_74+m104_74+m105_74+m106_74+m107_74+m108_74+m109_74+m110_74+m111_74+m112_74+m113_74+m114_74+m115_74+m116_74+m117_74+m118_74+m119_74+m120_74+m121_74+m122_74+m123_74+m124_74+m125_74+m126_74+m127_74+m128_74+m129_74+m130_74+m131_74+m132_74+m133_74+m134_74+m135_74+m136_74+m137_74+m138_74+m139_74+m140_74+m141_74+m142_74+m143_74+m144_74+m145_74+m146_74+m147_74+m148_74+m149_74+m150_74+m151_74+m152_74+m153_74+m154_74+m155_74+m156_74+m157_74+m158_74+m159_74+m160_74+m161_74+m162_74+m163_74+m164_74+m165_74+m166_74+m167_74+m168_74+m169_74+m170_74+m171_74+m172_74+m173_74+m174_74+m175_74+m176_74+m177_74+m178_74+m179_74+m180_74+m181_74+m182_74+m183_74+m184_74+m185_74+m186_74+m187_74+m188_74+m189_74+m190_74+m191_74+m192_74+m193_74+m194_74+m195_74+m196_74+m197_74+m198_74+m199_74+m200_74+m201_74+m202_74+m203_74+m204_74+m205_74+m206_74+m207_74+m208_74+m209_74+m210_74+m211_74+m212_74+m213_74+m214_74+m215_74+m216_74+m217_74+m218_74+m219_74+m220_74+m221_74+m222_74+m223_74+m224_74+m225_74+m226_74+m227_74+m228_74+m229_74+m230_74+m231_74+m232_74+m233_74+m234_74+m235_74+m236_74+m237_74+m238_74+m239_74+m240_74+m241_74+m242_74+m243_74+m244_74+m245_74+m246_74+m247_74+m248_74+m249_74+m250_74+m251_74+m252_74+m253_74+m254_74+m255_74+m256_74+m257_74+m258_74+m259_74+m260_74+m261_74+m262_74+m263_74+m264_74+m265_74+m266_74+m267_74+m268_74+m269_74+m270_74+m271_74+m272_74+m273_74+m274_74+m275_74+m276_74+m277_74+m278_74+m279_74+m280_74+m281_74+m282_74+m283_74+m284_74+m285_74+m286_74+m287_74+m288_74+m289_74+m290_74+m291_74+m292_74+m293_74+m294_74+m295_74+m296_74+m297_74+m298_74+m299_74+m300_74+m301_74+m302_74+m303_74+m304_74+m305_74+m306_74+m307_74+m308_74+m309_74+m310_74+m311_74+m312_74+m313_74+m314_74+m315_74+m316_74+m317_74+m318_74+m319_74+m320_74+m321_74+m322_74+m323_74+m324_74+m325_74+m326_74+m327_74+m328_74+m329_74+m330_74+m331_74+m332_74+m333_74+m334_74+m335_74+m336_74+m337_74+m338_74+m339_74+m340_74+m341_74+m342_74+m343_74+m344_74+m345_74+m346_74+m347_74+m348_74+m349_74+m350_74+m351_74+m352_74+m353_74+m354_74+m355_74+m356_74+m357_74+m358_74+m359_74+m360_74+m361_74+m362_74+m363_74+m364_74+m365_74+m366_74+m367_74+m368_74+m369_74+m370_74+m371_74+m372_74+m373_74+m374_74+m375_74+m376_74+m377_74+m378_74+m379_74+m380_74+m381_74+b74;
   always @(posedge clk) out75 <= m1_75+m2_75+m3_75+m4_75+m5_75+m6_75+m7_75+m8_75+m9_75+m10_75+m11_75+m12_75+m13_75+m14_75+m15_75+m16_75+m17_75+m18_75+m19_75+m20_75+m21_75+m22_75+m23_75+m24_75+m25_75+m26_75+m27_75+m28_75+m29_75+m30_75+m31_75+m32_75+m33_75+m34_75+m35_75+m36_75+m37_75+m38_75+m39_75+m40_75+m41_75+m42_75+m43_75+m44_75+m45_75+m46_75+m47_75+m48_75+m49_75+m50_75+m51_75+m52_75+m53_75+m54_75+m55_75+m56_75+m57_75+m58_75+m59_75+m60_75+m61_75+m62_75+m63_75+m64_75+m65_75+m66_75+m67_75+m68_75+m69_75+m70_75+m71_75+m72_75+m73_75+m74_75+m75_75+m76_75+m77_75+m78_75+m79_75+m80_75+m81_75+m82_75+m83_75+m84_75+m85_75+m86_75+m87_75+m88_75+m89_75+m90_75+m91_75+m92_75+m93_75+m94_75+m95_75+m96_75+m97_75+m98_75+m99_75+m100_75+m101_75+m102_75+m103_75+m104_75+m105_75+m106_75+m107_75+m108_75+m109_75+m110_75+m111_75+m112_75+m113_75+m114_75+m115_75+m116_75+m117_75+m118_75+m119_75+m120_75+m121_75+m122_75+m123_75+m124_75+m125_75+m126_75+m127_75+m128_75+m129_75+m130_75+m131_75+m132_75+m133_75+m134_75+m135_75+m136_75+m137_75+m138_75+m139_75+m140_75+m141_75+m142_75+m143_75+m144_75+m145_75+m146_75+m147_75+m148_75+m149_75+m150_75+m151_75+m152_75+m153_75+m154_75+m155_75+m156_75+m157_75+m158_75+m159_75+m160_75+m161_75+m162_75+m163_75+m164_75+m165_75+m166_75+m167_75+m168_75+m169_75+m170_75+m171_75+m172_75+m173_75+m174_75+m175_75+m176_75+m177_75+m178_75+m179_75+m180_75+m181_75+m182_75+m183_75+m184_75+m185_75+m186_75+m187_75+m188_75+m189_75+m190_75+m191_75+m192_75+m193_75+m194_75+m195_75+m196_75+m197_75+m198_75+m199_75+m200_75+m201_75+m202_75+m203_75+m204_75+m205_75+m206_75+m207_75+m208_75+m209_75+m210_75+m211_75+m212_75+m213_75+m214_75+m215_75+m216_75+m217_75+m218_75+m219_75+m220_75+m221_75+m222_75+m223_75+m224_75+m225_75+m226_75+m227_75+m228_75+m229_75+m230_75+m231_75+m232_75+m233_75+m234_75+m235_75+m236_75+m237_75+m238_75+m239_75+m240_75+m241_75+m242_75+m243_75+m244_75+m245_75+m246_75+m247_75+m248_75+m249_75+m250_75+m251_75+m252_75+m253_75+m254_75+m255_75+m256_75+m257_75+m258_75+m259_75+m260_75+m261_75+m262_75+m263_75+m264_75+m265_75+m266_75+m267_75+m268_75+m269_75+m270_75+m271_75+m272_75+m273_75+m274_75+m275_75+m276_75+m277_75+m278_75+m279_75+m280_75+m281_75+m282_75+m283_75+m284_75+m285_75+m286_75+m287_75+m288_75+m289_75+m290_75+m291_75+m292_75+m293_75+m294_75+m295_75+m296_75+m297_75+m298_75+m299_75+m300_75+m301_75+m302_75+m303_75+m304_75+m305_75+m306_75+m307_75+m308_75+m309_75+m310_75+m311_75+m312_75+m313_75+m314_75+m315_75+m316_75+m317_75+m318_75+m319_75+m320_75+m321_75+m322_75+m323_75+m324_75+m325_75+m326_75+m327_75+m328_75+m329_75+m330_75+m331_75+m332_75+m333_75+m334_75+m335_75+m336_75+m337_75+m338_75+m339_75+m340_75+m341_75+m342_75+m343_75+m344_75+m345_75+m346_75+m347_75+m348_75+m349_75+m350_75+m351_75+m352_75+m353_75+m354_75+m355_75+m356_75+m357_75+m358_75+m359_75+m360_75+m361_75+m362_75+m363_75+m364_75+m365_75+m366_75+m367_75+m368_75+m369_75+m370_75+m371_75+m372_75+m373_75+m374_75+m375_75+m376_75+m377_75+m378_75+m379_75+m380_75+m381_75+b75;
   always @(posedge clk) out76 <= m1_76+m2_76+m3_76+m4_76+m5_76+m6_76+m7_76+m8_76+m9_76+m10_76+m11_76+m12_76+m13_76+m14_76+m15_76+m16_76+m17_76+m18_76+m19_76+m20_76+m21_76+m22_76+m23_76+m24_76+m25_76+m26_76+m27_76+m28_76+m29_76+m30_76+m31_76+m32_76+m33_76+m34_76+m35_76+m36_76+m37_76+m38_76+m39_76+m40_76+m41_76+m42_76+m43_76+m44_76+m45_76+m46_76+m47_76+m48_76+m49_76+m50_76+m51_76+m52_76+m53_76+m54_76+m55_76+m56_76+m57_76+m58_76+m59_76+m60_76+m61_76+m62_76+m63_76+m64_76+m65_76+m66_76+m67_76+m68_76+m69_76+m70_76+m71_76+m72_76+m73_76+m74_76+m75_76+m76_76+m77_76+m78_76+m79_76+m80_76+m81_76+m82_76+m83_76+m84_76+m85_76+m86_76+m87_76+m88_76+m89_76+m90_76+m91_76+m92_76+m93_76+m94_76+m95_76+m96_76+m97_76+m98_76+m99_76+m100_76+m101_76+m102_76+m103_76+m104_76+m105_76+m106_76+m107_76+m108_76+m109_76+m110_76+m111_76+m112_76+m113_76+m114_76+m115_76+m116_76+m117_76+m118_76+m119_76+m120_76+m121_76+m122_76+m123_76+m124_76+m125_76+m126_76+m127_76+m128_76+m129_76+m130_76+m131_76+m132_76+m133_76+m134_76+m135_76+m136_76+m137_76+m138_76+m139_76+m140_76+m141_76+m142_76+m143_76+m144_76+m145_76+m146_76+m147_76+m148_76+m149_76+m150_76+m151_76+m152_76+m153_76+m154_76+m155_76+m156_76+m157_76+m158_76+m159_76+m160_76+m161_76+m162_76+m163_76+m164_76+m165_76+m166_76+m167_76+m168_76+m169_76+m170_76+m171_76+m172_76+m173_76+m174_76+m175_76+m176_76+m177_76+m178_76+m179_76+m180_76+m181_76+m182_76+m183_76+m184_76+m185_76+m186_76+m187_76+m188_76+m189_76+m190_76+m191_76+m192_76+m193_76+m194_76+m195_76+m196_76+m197_76+m198_76+m199_76+m200_76+m201_76+m202_76+m203_76+m204_76+m205_76+m206_76+m207_76+m208_76+m209_76+m210_76+m211_76+m212_76+m213_76+m214_76+m215_76+m216_76+m217_76+m218_76+m219_76+m220_76+m221_76+m222_76+m223_76+m224_76+m225_76+m226_76+m227_76+m228_76+m229_76+m230_76+m231_76+m232_76+m233_76+m234_76+m235_76+m236_76+m237_76+m238_76+m239_76+m240_76+m241_76+m242_76+m243_76+m244_76+m245_76+m246_76+m247_76+m248_76+m249_76+m250_76+m251_76+m252_76+m253_76+m254_76+m255_76+m256_76+m257_76+m258_76+m259_76+m260_76+m261_76+m262_76+m263_76+m264_76+m265_76+m266_76+m267_76+m268_76+m269_76+m270_76+m271_76+m272_76+m273_76+m274_76+m275_76+m276_76+m277_76+m278_76+m279_76+m280_76+m281_76+m282_76+m283_76+m284_76+m285_76+m286_76+m287_76+m288_76+m289_76+m290_76+m291_76+m292_76+m293_76+m294_76+m295_76+m296_76+m297_76+m298_76+m299_76+m300_76+m301_76+m302_76+m303_76+m304_76+m305_76+m306_76+m307_76+m308_76+m309_76+m310_76+m311_76+m312_76+m313_76+m314_76+m315_76+m316_76+m317_76+m318_76+m319_76+m320_76+m321_76+m322_76+m323_76+m324_76+m325_76+m326_76+m327_76+m328_76+m329_76+m330_76+m331_76+m332_76+m333_76+m334_76+m335_76+m336_76+m337_76+m338_76+m339_76+m340_76+m341_76+m342_76+m343_76+m344_76+m345_76+m346_76+m347_76+m348_76+m349_76+m350_76+m351_76+m352_76+m353_76+m354_76+m355_76+m356_76+m357_76+m358_76+m359_76+m360_76+m361_76+m362_76+m363_76+m364_76+m365_76+m366_76+m367_76+m368_76+m369_76+m370_76+m371_76+m372_76+m373_76+m374_76+m375_76+m376_76+m377_76+m378_76+m379_76+m380_76+m381_76+b76;
   always @(posedge clk) out77 <= m1_77+m2_77+m3_77+m4_77+m5_77+m6_77+m7_77+m8_77+m9_77+m10_77+m11_77+m12_77+m13_77+m14_77+m15_77+m16_77+m17_77+m18_77+m19_77+m20_77+m21_77+m22_77+m23_77+m24_77+m25_77+m26_77+m27_77+m28_77+m29_77+m30_77+m31_77+m32_77+m33_77+m34_77+m35_77+m36_77+m37_77+m38_77+m39_77+m40_77+m41_77+m42_77+m43_77+m44_77+m45_77+m46_77+m47_77+m48_77+m49_77+m50_77+m51_77+m52_77+m53_77+m54_77+m55_77+m56_77+m57_77+m58_77+m59_77+m60_77+m61_77+m62_77+m63_77+m64_77+m65_77+m66_77+m67_77+m68_77+m69_77+m70_77+m71_77+m72_77+m73_77+m74_77+m75_77+m76_77+m77_77+m78_77+m79_77+m80_77+m81_77+m82_77+m83_77+m84_77+m85_77+m86_77+m87_77+m88_77+m89_77+m90_77+m91_77+m92_77+m93_77+m94_77+m95_77+m96_77+m97_77+m98_77+m99_77+m100_77+m101_77+m102_77+m103_77+m104_77+m105_77+m106_77+m107_77+m108_77+m109_77+m110_77+m111_77+m112_77+m113_77+m114_77+m115_77+m116_77+m117_77+m118_77+m119_77+m120_77+m121_77+m122_77+m123_77+m124_77+m125_77+m126_77+m127_77+m128_77+m129_77+m130_77+m131_77+m132_77+m133_77+m134_77+m135_77+m136_77+m137_77+m138_77+m139_77+m140_77+m141_77+m142_77+m143_77+m144_77+m145_77+m146_77+m147_77+m148_77+m149_77+m150_77+m151_77+m152_77+m153_77+m154_77+m155_77+m156_77+m157_77+m158_77+m159_77+m160_77+m161_77+m162_77+m163_77+m164_77+m165_77+m166_77+m167_77+m168_77+m169_77+m170_77+m171_77+m172_77+m173_77+m174_77+m175_77+m176_77+m177_77+m178_77+m179_77+m180_77+m181_77+m182_77+m183_77+m184_77+m185_77+m186_77+m187_77+m188_77+m189_77+m190_77+m191_77+m192_77+m193_77+m194_77+m195_77+m196_77+m197_77+m198_77+m199_77+m200_77+m201_77+m202_77+m203_77+m204_77+m205_77+m206_77+m207_77+m208_77+m209_77+m210_77+m211_77+m212_77+m213_77+m214_77+m215_77+m216_77+m217_77+m218_77+m219_77+m220_77+m221_77+m222_77+m223_77+m224_77+m225_77+m226_77+m227_77+m228_77+m229_77+m230_77+m231_77+m232_77+m233_77+m234_77+m235_77+m236_77+m237_77+m238_77+m239_77+m240_77+m241_77+m242_77+m243_77+m244_77+m245_77+m246_77+m247_77+m248_77+m249_77+m250_77+m251_77+m252_77+m253_77+m254_77+m255_77+m256_77+m257_77+m258_77+m259_77+m260_77+m261_77+m262_77+m263_77+m264_77+m265_77+m266_77+m267_77+m268_77+m269_77+m270_77+m271_77+m272_77+m273_77+m274_77+m275_77+m276_77+m277_77+m278_77+m279_77+m280_77+m281_77+m282_77+m283_77+m284_77+m285_77+m286_77+m287_77+m288_77+m289_77+m290_77+m291_77+m292_77+m293_77+m294_77+m295_77+m296_77+m297_77+m298_77+m299_77+m300_77+m301_77+m302_77+m303_77+m304_77+m305_77+m306_77+m307_77+m308_77+m309_77+m310_77+m311_77+m312_77+m313_77+m314_77+m315_77+m316_77+m317_77+m318_77+m319_77+m320_77+m321_77+m322_77+m323_77+m324_77+m325_77+m326_77+m327_77+m328_77+m329_77+m330_77+m331_77+m332_77+m333_77+m334_77+m335_77+m336_77+m337_77+m338_77+m339_77+m340_77+m341_77+m342_77+m343_77+m344_77+m345_77+m346_77+m347_77+m348_77+m349_77+m350_77+m351_77+m352_77+m353_77+m354_77+m355_77+m356_77+m357_77+m358_77+m359_77+m360_77+m361_77+m362_77+m363_77+m364_77+m365_77+m366_77+m367_77+m368_77+m369_77+m370_77+m371_77+m372_77+m373_77+m374_77+m375_77+m376_77+m377_77+m378_77+m379_77+m380_77+m381_77+b77;
   always @(posedge clk) out78 <= m1_78+m2_78+m3_78+m4_78+m5_78+m6_78+m7_78+m8_78+m9_78+m10_78+m11_78+m12_78+m13_78+m14_78+m15_78+m16_78+m17_78+m18_78+m19_78+m20_78+m21_78+m22_78+m23_78+m24_78+m25_78+m26_78+m27_78+m28_78+m29_78+m30_78+m31_78+m32_78+m33_78+m34_78+m35_78+m36_78+m37_78+m38_78+m39_78+m40_78+m41_78+m42_78+m43_78+m44_78+m45_78+m46_78+m47_78+m48_78+m49_78+m50_78+m51_78+m52_78+m53_78+m54_78+m55_78+m56_78+m57_78+m58_78+m59_78+m60_78+m61_78+m62_78+m63_78+m64_78+m65_78+m66_78+m67_78+m68_78+m69_78+m70_78+m71_78+m72_78+m73_78+m74_78+m75_78+m76_78+m77_78+m78_78+m79_78+m80_78+m81_78+m82_78+m83_78+m84_78+m85_78+m86_78+m87_78+m88_78+m89_78+m90_78+m91_78+m92_78+m93_78+m94_78+m95_78+m96_78+m97_78+m98_78+m99_78+m100_78+m101_78+m102_78+m103_78+m104_78+m105_78+m106_78+m107_78+m108_78+m109_78+m110_78+m111_78+m112_78+m113_78+m114_78+m115_78+m116_78+m117_78+m118_78+m119_78+m120_78+m121_78+m122_78+m123_78+m124_78+m125_78+m126_78+m127_78+m128_78+m129_78+m130_78+m131_78+m132_78+m133_78+m134_78+m135_78+m136_78+m137_78+m138_78+m139_78+m140_78+m141_78+m142_78+m143_78+m144_78+m145_78+m146_78+m147_78+m148_78+m149_78+m150_78+m151_78+m152_78+m153_78+m154_78+m155_78+m156_78+m157_78+m158_78+m159_78+m160_78+m161_78+m162_78+m163_78+m164_78+m165_78+m166_78+m167_78+m168_78+m169_78+m170_78+m171_78+m172_78+m173_78+m174_78+m175_78+m176_78+m177_78+m178_78+m179_78+m180_78+m181_78+m182_78+m183_78+m184_78+m185_78+m186_78+m187_78+m188_78+m189_78+m190_78+m191_78+m192_78+m193_78+m194_78+m195_78+m196_78+m197_78+m198_78+m199_78+m200_78+m201_78+m202_78+m203_78+m204_78+m205_78+m206_78+m207_78+m208_78+m209_78+m210_78+m211_78+m212_78+m213_78+m214_78+m215_78+m216_78+m217_78+m218_78+m219_78+m220_78+m221_78+m222_78+m223_78+m224_78+m225_78+m226_78+m227_78+m228_78+m229_78+m230_78+m231_78+m232_78+m233_78+m234_78+m235_78+m236_78+m237_78+m238_78+m239_78+m240_78+m241_78+m242_78+m243_78+m244_78+m245_78+m246_78+m247_78+m248_78+m249_78+m250_78+m251_78+m252_78+m253_78+m254_78+m255_78+m256_78+m257_78+m258_78+m259_78+m260_78+m261_78+m262_78+m263_78+m264_78+m265_78+m266_78+m267_78+m268_78+m269_78+m270_78+m271_78+m272_78+m273_78+m274_78+m275_78+m276_78+m277_78+m278_78+m279_78+m280_78+m281_78+m282_78+m283_78+m284_78+m285_78+m286_78+m287_78+m288_78+m289_78+m290_78+m291_78+m292_78+m293_78+m294_78+m295_78+m296_78+m297_78+m298_78+m299_78+m300_78+m301_78+m302_78+m303_78+m304_78+m305_78+m306_78+m307_78+m308_78+m309_78+m310_78+m311_78+m312_78+m313_78+m314_78+m315_78+m316_78+m317_78+m318_78+m319_78+m320_78+m321_78+m322_78+m323_78+m324_78+m325_78+m326_78+m327_78+m328_78+m329_78+m330_78+m331_78+m332_78+m333_78+m334_78+m335_78+m336_78+m337_78+m338_78+m339_78+m340_78+m341_78+m342_78+m343_78+m344_78+m345_78+m346_78+m347_78+m348_78+m349_78+m350_78+m351_78+m352_78+m353_78+m354_78+m355_78+m356_78+m357_78+m358_78+m359_78+m360_78+m361_78+m362_78+m363_78+m364_78+m365_78+m366_78+m367_78+m368_78+m369_78+m370_78+m371_78+m372_78+m373_78+m374_78+m375_78+m376_78+m377_78+m378_78+m379_78+m380_78+m381_78+b78;
   always @(posedge clk) out79 <= m1_79+m2_79+m3_79+m4_79+m5_79+m6_79+m7_79+m8_79+m9_79+m10_79+m11_79+m12_79+m13_79+m14_79+m15_79+m16_79+m17_79+m18_79+m19_79+m20_79+m21_79+m22_79+m23_79+m24_79+m25_79+m26_79+m27_79+m28_79+m29_79+m30_79+m31_79+m32_79+m33_79+m34_79+m35_79+m36_79+m37_79+m38_79+m39_79+m40_79+m41_79+m42_79+m43_79+m44_79+m45_79+m46_79+m47_79+m48_79+m49_79+m50_79+m51_79+m52_79+m53_79+m54_79+m55_79+m56_79+m57_79+m58_79+m59_79+m60_79+m61_79+m62_79+m63_79+m64_79+m65_79+m66_79+m67_79+m68_79+m69_79+m70_79+m71_79+m72_79+m73_79+m74_79+m75_79+m76_79+m77_79+m78_79+m79_79+m80_79+m81_79+m82_79+m83_79+m84_79+m85_79+m86_79+m87_79+m88_79+m89_79+m90_79+m91_79+m92_79+m93_79+m94_79+m95_79+m96_79+m97_79+m98_79+m99_79+m100_79+m101_79+m102_79+m103_79+m104_79+m105_79+m106_79+m107_79+m108_79+m109_79+m110_79+m111_79+m112_79+m113_79+m114_79+m115_79+m116_79+m117_79+m118_79+m119_79+m120_79+m121_79+m122_79+m123_79+m124_79+m125_79+m126_79+m127_79+m128_79+m129_79+m130_79+m131_79+m132_79+m133_79+m134_79+m135_79+m136_79+m137_79+m138_79+m139_79+m140_79+m141_79+m142_79+m143_79+m144_79+m145_79+m146_79+m147_79+m148_79+m149_79+m150_79+m151_79+m152_79+m153_79+m154_79+m155_79+m156_79+m157_79+m158_79+m159_79+m160_79+m161_79+m162_79+m163_79+m164_79+m165_79+m166_79+m167_79+m168_79+m169_79+m170_79+m171_79+m172_79+m173_79+m174_79+m175_79+m176_79+m177_79+m178_79+m179_79+m180_79+m181_79+m182_79+m183_79+m184_79+m185_79+m186_79+m187_79+m188_79+m189_79+m190_79+m191_79+m192_79+m193_79+m194_79+m195_79+m196_79+m197_79+m198_79+m199_79+m200_79+m201_79+m202_79+m203_79+m204_79+m205_79+m206_79+m207_79+m208_79+m209_79+m210_79+m211_79+m212_79+m213_79+m214_79+m215_79+m216_79+m217_79+m218_79+m219_79+m220_79+m221_79+m222_79+m223_79+m224_79+m225_79+m226_79+m227_79+m228_79+m229_79+m230_79+m231_79+m232_79+m233_79+m234_79+m235_79+m236_79+m237_79+m238_79+m239_79+m240_79+m241_79+m242_79+m243_79+m244_79+m245_79+m246_79+m247_79+m248_79+m249_79+m250_79+m251_79+m252_79+m253_79+m254_79+m255_79+m256_79+m257_79+m258_79+m259_79+m260_79+m261_79+m262_79+m263_79+m264_79+m265_79+m266_79+m267_79+m268_79+m269_79+m270_79+m271_79+m272_79+m273_79+m274_79+m275_79+m276_79+m277_79+m278_79+m279_79+m280_79+m281_79+m282_79+m283_79+m284_79+m285_79+m286_79+m287_79+m288_79+m289_79+m290_79+m291_79+m292_79+m293_79+m294_79+m295_79+m296_79+m297_79+m298_79+m299_79+m300_79+m301_79+m302_79+m303_79+m304_79+m305_79+m306_79+m307_79+m308_79+m309_79+m310_79+m311_79+m312_79+m313_79+m314_79+m315_79+m316_79+m317_79+m318_79+m319_79+m320_79+m321_79+m322_79+m323_79+m324_79+m325_79+m326_79+m327_79+m328_79+m329_79+m330_79+m331_79+m332_79+m333_79+m334_79+m335_79+m336_79+m337_79+m338_79+m339_79+m340_79+m341_79+m342_79+m343_79+m344_79+m345_79+m346_79+m347_79+m348_79+m349_79+m350_79+m351_79+m352_79+m353_79+m354_79+m355_79+m356_79+m357_79+m358_79+m359_79+m360_79+m361_79+m362_79+m363_79+m364_79+m365_79+m366_79+m367_79+m368_79+m369_79+m370_79+m371_79+m372_79+m373_79+m374_79+m375_79+m376_79+m377_79+m378_79+m379_79+m380_79+m381_79+b79;
   always @(posedge clk) out80 <= m1_80+m2_80+m3_80+m4_80+m5_80+m6_80+m7_80+m8_80+m9_80+m10_80+m11_80+m12_80+m13_80+m14_80+m15_80+m16_80+m17_80+m18_80+m19_80+m20_80+m21_80+m22_80+m23_80+m24_80+m25_80+m26_80+m27_80+m28_80+m29_80+m30_80+m31_80+m32_80+m33_80+m34_80+m35_80+m36_80+m37_80+m38_80+m39_80+m40_80+m41_80+m42_80+m43_80+m44_80+m45_80+m46_80+m47_80+m48_80+m49_80+m50_80+m51_80+m52_80+m53_80+m54_80+m55_80+m56_80+m57_80+m58_80+m59_80+m60_80+m61_80+m62_80+m63_80+m64_80+m65_80+m66_80+m67_80+m68_80+m69_80+m70_80+m71_80+m72_80+m73_80+m74_80+m75_80+m76_80+m77_80+m78_80+m79_80+m80_80+m81_80+m82_80+m83_80+m84_80+m85_80+m86_80+m87_80+m88_80+m89_80+m90_80+m91_80+m92_80+m93_80+m94_80+m95_80+m96_80+m97_80+m98_80+m99_80+m100_80+m101_80+m102_80+m103_80+m104_80+m105_80+m106_80+m107_80+m108_80+m109_80+m110_80+m111_80+m112_80+m113_80+m114_80+m115_80+m116_80+m117_80+m118_80+m119_80+m120_80+m121_80+m122_80+m123_80+m124_80+m125_80+m126_80+m127_80+m128_80+m129_80+m130_80+m131_80+m132_80+m133_80+m134_80+m135_80+m136_80+m137_80+m138_80+m139_80+m140_80+m141_80+m142_80+m143_80+m144_80+m145_80+m146_80+m147_80+m148_80+m149_80+m150_80+m151_80+m152_80+m153_80+m154_80+m155_80+m156_80+m157_80+m158_80+m159_80+m160_80+m161_80+m162_80+m163_80+m164_80+m165_80+m166_80+m167_80+m168_80+m169_80+m170_80+m171_80+m172_80+m173_80+m174_80+m175_80+m176_80+m177_80+m178_80+m179_80+m180_80+m181_80+m182_80+m183_80+m184_80+m185_80+m186_80+m187_80+m188_80+m189_80+m190_80+m191_80+m192_80+m193_80+m194_80+m195_80+m196_80+m197_80+m198_80+m199_80+m200_80+m201_80+m202_80+m203_80+m204_80+m205_80+m206_80+m207_80+m208_80+m209_80+m210_80+m211_80+m212_80+m213_80+m214_80+m215_80+m216_80+m217_80+m218_80+m219_80+m220_80+m221_80+m222_80+m223_80+m224_80+m225_80+m226_80+m227_80+m228_80+m229_80+m230_80+m231_80+m232_80+m233_80+m234_80+m235_80+m236_80+m237_80+m238_80+m239_80+m240_80+m241_80+m242_80+m243_80+m244_80+m245_80+m246_80+m247_80+m248_80+m249_80+m250_80+m251_80+m252_80+m253_80+m254_80+m255_80+m256_80+m257_80+m258_80+m259_80+m260_80+m261_80+m262_80+m263_80+m264_80+m265_80+m266_80+m267_80+m268_80+m269_80+m270_80+m271_80+m272_80+m273_80+m274_80+m275_80+m276_80+m277_80+m278_80+m279_80+m280_80+m281_80+m282_80+m283_80+m284_80+m285_80+m286_80+m287_80+m288_80+m289_80+m290_80+m291_80+m292_80+m293_80+m294_80+m295_80+m296_80+m297_80+m298_80+m299_80+m300_80+m301_80+m302_80+m303_80+m304_80+m305_80+m306_80+m307_80+m308_80+m309_80+m310_80+m311_80+m312_80+m313_80+m314_80+m315_80+m316_80+m317_80+m318_80+m319_80+m320_80+m321_80+m322_80+m323_80+m324_80+m325_80+m326_80+m327_80+m328_80+m329_80+m330_80+m331_80+m332_80+m333_80+m334_80+m335_80+m336_80+m337_80+m338_80+m339_80+m340_80+m341_80+m342_80+m343_80+m344_80+m345_80+m346_80+m347_80+m348_80+m349_80+m350_80+m351_80+m352_80+m353_80+m354_80+m355_80+m356_80+m357_80+m358_80+m359_80+m360_80+m361_80+m362_80+m363_80+m364_80+m365_80+m366_80+m367_80+m368_80+m369_80+m370_80+m371_80+m372_80+m373_80+m374_80+m375_80+m376_80+m377_80+m378_80+m379_80+m380_80+m381_80+b80;
   always @(posedge clk) out81 <= m1_81+m2_81+m3_81+m4_81+m5_81+m6_81+m7_81+m8_81+m9_81+m10_81+m11_81+m12_81+m13_81+m14_81+m15_81+m16_81+m17_81+m18_81+m19_81+m20_81+m21_81+m22_81+m23_81+m24_81+m25_81+m26_81+m27_81+m28_81+m29_81+m30_81+m31_81+m32_81+m33_81+m34_81+m35_81+m36_81+m37_81+m38_81+m39_81+m40_81+m41_81+m42_81+m43_81+m44_81+m45_81+m46_81+m47_81+m48_81+m49_81+m50_81+m51_81+m52_81+m53_81+m54_81+m55_81+m56_81+m57_81+m58_81+m59_81+m60_81+m61_81+m62_81+m63_81+m64_81+m65_81+m66_81+m67_81+m68_81+m69_81+m70_81+m71_81+m72_81+m73_81+m74_81+m75_81+m76_81+m77_81+m78_81+m79_81+m80_81+m81_81+m82_81+m83_81+m84_81+m85_81+m86_81+m87_81+m88_81+m89_81+m90_81+m91_81+m92_81+m93_81+m94_81+m95_81+m96_81+m97_81+m98_81+m99_81+m100_81+m101_81+m102_81+m103_81+m104_81+m105_81+m106_81+m107_81+m108_81+m109_81+m110_81+m111_81+m112_81+m113_81+m114_81+m115_81+m116_81+m117_81+m118_81+m119_81+m120_81+m121_81+m122_81+m123_81+m124_81+m125_81+m126_81+m127_81+m128_81+m129_81+m130_81+m131_81+m132_81+m133_81+m134_81+m135_81+m136_81+m137_81+m138_81+m139_81+m140_81+m141_81+m142_81+m143_81+m144_81+m145_81+m146_81+m147_81+m148_81+m149_81+m150_81+m151_81+m152_81+m153_81+m154_81+m155_81+m156_81+m157_81+m158_81+m159_81+m160_81+m161_81+m162_81+m163_81+m164_81+m165_81+m166_81+m167_81+m168_81+m169_81+m170_81+m171_81+m172_81+m173_81+m174_81+m175_81+m176_81+m177_81+m178_81+m179_81+m180_81+m181_81+m182_81+m183_81+m184_81+m185_81+m186_81+m187_81+m188_81+m189_81+m190_81+m191_81+m192_81+m193_81+m194_81+m195_81+m196_81+m197_81+m198_81+m199_81+m200_81+m201_81+m202_81+m203_81+m204_81+m205_81+m206_81+m207_81+m208_81+m209_81+m210_81+m211_81+m212_81+m213_81+m214_81+m215_81+m216_81+m217_81+m218_81+m219_81+m220_81+m221_81+m222_81+m223_81+m224_81+m225_81+m226_81+m227_81+m228_81+m229_81+m230_81+m231_81+m232_81+m233_81+m234_81+m235_81+m236_81+m237_81+m238_81+m239_81+m240_81+m241_81+m242_81+m243_81+m244_81+m245_81+m246_81+m247_81+m248_81+m249_81+m250_81+m251_81+m252_81+m253_81+m254_81+m255_81+m256_81+m257_81+m258_81+m259_81+m260_81+m261_81+m262_81+m263_81+m264_81+m265_81+m266_81+m267_81+m268_81+m269_81+m270_81+m271_81+m272_81+m273_81+m274_81+m275_81+m276_81+m277_81+m278_81+m279_81+m280_81+m281_81+m282_81+m283_81+m284_81+m285_81+m286_81+m287_81+m288_81+m289_81+m290_81+m291_81+m292_81+m293_81+m294_81+m295_81+m296_81+m297_81+m298_81+m299_81+m300_81+m301_81+m302_81+m303_81+m304_81+m305_81+m306_81+m307_81+m308_81+m309_81+m310_81+m311_81+m312_81+m313_81+m314_81+m315_81+m316_81+m317_81+m318_81+m319_81+m320_81+m321_81+m322_81+m323_81+m324_81+m325_81+m326_81+m327_81+m328_81+m329_81+m330_81+m331_81+m332_81+m333_81+m334_81+m335_81+m336_81+m337_81+m338_81+m339_81+m340_81+m341_81+m342_81+m343_81+m344_81+m345_81+m346_81+m347_81+m348_81+m349_81+m350_81+m351_81+m352_81+m353_81+m354_81+m355_81+m356_81+m357_81+m358_81+m359_81+m360_81+m361_81+m362_81+m363_81+m364_81+m365_81+m366_81+m367_81+m368_81+m369_81+m370_81+m371_81+m372_81+m373_81+m374_81+m375_81+m376_81+m377_81+m378_81+m379_81+m380_81+m381_81+b81;
   always @(posedge clk) out82 <= m1_82+m2_82+m3_82+m4_82+m5_82+m6_82+m7_82+m8_82+m9_82+m10_82+m11_82+m12_82+m13_82+m14_82+m15_82+m16_82+m17_82+m18_82+m19_82+m20_82+m21_82+m22_82+m23_82+m24_82+m25_82+m26_82+m27_82+m28_82+m29_82+m30_82+m31_82+m32_82+m33_82+m34_82+m35_82+m36_82+m37_82+m38_82+m39_82+m40_82+m41_82+m42_82+m43_82+m44_82+m45_82+m46_82+m47_82+m48_82+m49_82+m50_82+m51_82+m52_82+m53_82+m54_82+m55_82+m56_82+m57_82+m58_82+m59_82+m60_82+m61_82+m62_82+m63_82+m64_82+m65_82+m66_82+m67_82+m68_82+m69_82+m70_82+m71_82+m72_82+m73_82+m74_82+m75_82+m76_82+m77_82+m78_82+m79_82+m80_82+m81_82+m82_82+m83_82+m84_82+m85_82+m86_82+m87_82+m88_82+m89_82+m90_82+m91_82+m92_82+m93_82+m94_82+m95_82+m96_82+m97_82+m98_82+m99_82+m100_82+m101_82+m102_82+m103_82+m104_82+m105_82+m106_82+m107_82+m108_82+m109_82+m110_82+m111_82+m112_82+m113_82+m114_82+m115_82+m116_82+m117_82+m118_82+m119_82+m120_82+m121_82+m122_82+m123_82+m124_82+m125_82+m126_82+m127_82+m128_82+m129_82+m130_82+m131_82+m132_82+m133_82+m134_82+m135_82+m136_82+m137_82+m138_82+m139_82+m140_82+m141_82+m142_82+m143_82+m144_82+m145_82+m146_82+m147_82+m148_82+m149_82+m150_82+m151_82+m152_82+m153_82+m154_82+m155_82+m156_82+m157_82+m158_82+m159_82+m160_82+m161_82+m162_82+m163_82+m164_82+m165_82+m166_82+m167_82+m168_82+m169_82+m170_82+m171_82+m172_82+m173_82+m174_82+m175_82+m176_82+m177_82+m178_82+m179_82+m180_82+m181_82+m182_82+m183_82+m184_82+m185_82+m186_82+m187_82+m188_82+m189_82+m190_82+m191_82+m192_82+m193_82+m194_82+m195_82+m196_82+m197_82+m198_82+m199_82+m200_82+m201_82+m202_82+m203_82+m204_82+m205_82+m206_82+m207_82+m208_82+m209_82+m210_82+m211_82+m212_82+m213_82+m214_82+m215_82+m216_82+m217_82+m218_82+m219_82+m220_82+m221_82+m222_82+m223_82+m224_82+m225_82+m226_82+m227_82+m228_82+m229_82+m230_82+m231_82+m232_82+m233_82+m234_82+m235_82+m236_82+m237_82+m238_82+m239_82+m240_82+m241_82+m242_82+m243_82+m244_82+m245_82+m246_82+m247_82+m248_82+m249_82+m250_82+m251_82+m252_82+m253_82+m254_82+m255_82+m256_82+m257_82+m258_82+m259_82+m260_82+m261_82+m262_82+m263_82+m264_82+m265_82+m266_82+m267_82+m268_82+m269_82+m270_82+m271_82+m272_82+m273_82+m274_82+m275_82+m276_82+m277_82+m278_82+m279_82+m280_82+m281_82+m282_82+m283_82+m284_82+m285_82+m286_82+m287_82+m288_82+m289_82+m290_82+m291_82+m292_82+m293_82+m294_82+m295_82+m296_82+m297_82+m298_82+m299_82+m300_82+m301_82+m302_82+m303_82+m304_82+m305_82+m306_82+m307_82+m308_82+m309_82+m310_82+m311_82+m312_82+m313_82+m314_82+m315_82+m316_82+m317_82+m318_82+m319_82+m320_82+m321_82+m322_82+m323_82+m324_82+m325_82+m326_82+m327_82+m328_82+m329_82+m330_82+m331_82+m332_82+m333_82+m334_82+m335_82+m336_82+m337_82+m338_82+m339_82+m340_82+m341_82+m342_82+m343_82+m344_82+m345_82+m346_82+m347_82+m348_82+m349_82+m350_82+m351_82+m352_82+m353_82+m354_82+m355_82+m356_82+m357_82+m358_82+m359_82+m360_82+m361_82+m362_82+m363_82+m364_82+m365_82+m366_82+m367_82+m368_82+m369_82+m370_82+m371_82+m372_82+m373_82+m374_82+m375_82+m376_82+m377_82+m378_82+m379_82+m380_82+m381_82+b82;
   always @(posedge clk) out83 <= m1_83+m2_83+m3_83+m4_83+m5_83+m6_83+m7_83+m8_83+m9_83+m10_83+m11_83+m12_83+m13_83+m14_83+m15_83+m16_83+m17_83+m18_83+m19_83+m20_83+m21_83+m22_83+m23_83+m24_83+m25_83+m26_83+m27_83+m28_83+m29_83+m30_83+m31_83+m32_83+m33_83+m34_83+m35_83+m36_83+m37_83+m38_83+m39_83+m40_83+m41_83+m42_83+m43_83+m44_83+m45_83+m46_83+m47_83+m48_83+m49_83+m50_83+m51_83+m52_83+m53_83+m54_83+m55_83+m56_83+m57_83+m58_83+m59_83+m60_83+m61_83+m62_83+m63_83+m64_83+m65_83+m66_83+m67_83+m68_83+m69_83+m70_83+m71_83+m72_83+m73_83+m74_83+m75_83+m76_83+m77_83+m78_83+m79_83+m80_83+m81_83+m82_83+m83_83+m84_83+m85_83+m86_83+m87_83+m88_83+m89_83+m90_83+m91_83+m92_83+m93_83+m94_83+m95_83+m96_83+m97_83+m98_83+m99_83+m100_83+m101_83+m102_83+m103_83+m104_83+m105_83+m106_83+m107_83+m108_83+m109_83+m110_83+m111_83+m112_83+m113_83+m114_83+m115_83+m116_83+m117_83+m118_83+m119_83+m120_83+m121_83+m122_83+m123_83+m124_83+m125_83+m126_83+m127_83+m128_83+m129_83+m130_83+m131_83+m132_83+m133_83+m134_83+m135_83+m136_83+m137_83+m138_83+m139_83+m140_83+m141_83+m142_83+m143_83+m144_83+m145_83+m146_83+m147_83+m148_83+m149_83+m150_83+m151_83+m152_83+m153_83+m154_83+m155_83+m156_83+m157_83+m158_83+m159_83+m160_83+m161_83+m162_83+m163_83+m164_83+m165_83+m166_83+m167_83+m168_83+m169_83+m170_83+m171_83+m172_83+m173_83+m174_83+m175_83+m176_83+m177_83+m178_83+m179_83+m180_83+m181_83+m182_83+m183_83+m184_83+m185_83+m186_83+m187_83+m188_83+m189_83+m190_83+m191_83+m192_83+m193_83+m194_83+m195_83+m196_83+m197_83+m198_83+m199_83+m200_83+m201_83+m202_83+m203_83+m204_83+m205_83+m206_83+m207_83+m208_83+m209_83+m210_83+m211_83+m212_83+m213_83+m214_83+m215_83+m216_83+m217_83+m218_83+m219_83+m220_83+m221_83+m222_83+m223_83+m224_83+m225_83+m226_83+m227_83+m228_83+m229_83+m230_83+m231_83+m232_83+m233_83+m234_83+m235_83+m236_83+m237_83+m238_83+m239_83+m240_83+m241_83+m242_83+m243_83+m244_83+m245_83+m246_83+m247_83+m248_83+m249_83+m250_83+m251_83+m252_83+m253_83+m254_83+m255_83+m256_83+m257_83+m258_83+m259_83+m260_83+m261_83+m262_83+m263_83+m264_83+m265_83+m266_83+m267_83+m268_83+m269_83+m270_83+m271_83+m272_83+m273_83+m274_83+m275_83+m276_83+m277_83+m278_83+m279_83+m280_83+m281_83+m282_83+m283_83+m284_83+m285_83+m286_83+m287_83+m288_83+m289_83+m290_83+m291_83+m292_83+m293_83+m294_83+m295_83+m296_83+m297_83+m298_83+m299_83+m300_83+m301_83+m302_83+m303_83+m304_83+m305_83+m306_83+m307_83+m308_83+m309_83+m310_83+m311_83+m312_83+m313_83+m314_83+m315_83+m316_83+m317_83+m318_83+m319_83+m320_83+m321_83+m322_83+m323_83+m324_83+m325_83+m326_83+m327_83+m328_83+m329_83+m330_83+m331_83+m332_83+m333_83+m334_83+m335_83+m336_83+m337_83+m338_83+m339_83+m340_83+m341_83+m342_83+m343_83+m344_83+m345_83+m346_83+m347_83+m348_83+m349_83+m350_83+m351_83+m352_83+m353_83+m354_83+m355_83+m356_83+m357_83+m358_83+m359_83+m360_83+m361_83+m362_83+m363_83+m364_83+m365_83+m366_83+m367_83+m368_83+m369_83+m370_83+m371_83+m372_83+m373_83+m374_83+m375_83+m376_83+m377_83+m378_83+m379_83+m380_83+m381_83+b83;
   always @(posedge clk) out84 <= m1_84+m2_84+m3_84+m4_84+m5_84+m6_84+m7_84+m8_84+m9_84+m10_84+m11_84+m12_84+m13_84+m14_84+m15_84+m16_84+m17_84+m18_84+m19_84+m20_84+m21_84+m22_84+m23_84+m24_84+m25_84+m26_84+m27_84+m28_84+m29_84+m30_84+m31_84+m32_84+m33_84+m34_84+m35_84+m36_84+m37_84+m38_84+m39_84+m40_84+m41_84+m42_84+m43_84+m44_84+m45_84+m46_84+m47_84+m48_84+m49_84+m50_84+m51_84+m52_84+m53_84+m54_84+m55_84+m56_84+m57_84+m58_84+m59_84+m60_84+m61_84+m62_84+m63_84+m64_84+m65_84+m66_84+m67_84+m68_84+m69_84+m70_84+m71_84+m72_84+m73_84+m74_84+m75_84+m76_84+m77_84+m78_84+m79_84+m80_84+m81_84+m82_84+m83_84+m84_84+m85_84+m86_84+m87_84+m88_84+m89_84+m90_84+m91_84+m92_84+m93_84+m94_84+m95_84+m96_84+m97_84+m98_84+m99_84+m100_84+m101_84+m102_84+m103_84+m104_84+m105_84+m106_84+m107_84+m108_84+m109_84+m110_84+m111_84+m112_84+m113_84+m114_84+m115_84+m116_84+m117_84+m118_84+m119_84+m120_84+m121_84+m122_84+m123_84+m124_84+m125_84+m126_84+m127_84+m128_84+m129_84+m130_84+m131_84+m132_84+m133_84+m134_84+m135_84+m136_84+m137_84+m138_84+m139_84+m140_84+m141_84+m142_84+m143_84+m144_84+m145_84+m146_84+m147_84+m148_84+m149_84+m150_84+m151_84+m152_84+m153_84+m154_84+m155_84+m156_84+m157_84+m158_84+m159_84+m160_84+m161_84+m162_84+m163_84+m164_84+m165_84+m166_84+m167_84+m168_84+m169_84+m170_84+m171_84+m172_84+m173_84+m174_84+m175_84+m176_84+m177_84+m178_84+m179_84+m180_84+m181_84+m182_84+m183_84+m184_84+m185_84+m186_84+m187_84+m188_84+m189_84+m190_84+m191_84+m192_84+m193_84+m194_84+m195_84+m196_84+m197_84+m198_84+m199_84+m200_84+m201_84+m202_84+m203_84+m204_84+m205_84+m206_84+m207_84+m208_84+m209_84+m210_84+m211_84+m212_84+m213_84+m214_84+m215_84+m216_84+m217_84+m218_84+m219_84+m220_84+m221_84+m222_84+m223_84+m224_84+m225_84+m226_84+m227_84+m228_84+m229_84+m230_84+m231_84+m232_84+m233_84+m234_84+m235_84+m236_84+m237_84+m238_84+m239_84+m240_84+m241_84+m242_84+m243_84+m244_84+m245_84+m246_84+m247_84+m248_84+m249_84+m250_84+m251_84+m252_84+m253_84+m254_84+m255_84+m256_84+m257_84+m258_84+m259_84+m260_84+m261_84+m262_84+m263_84+m264_84+m265_84+m266_84+m267_84+m268_84+m269_84+m270_84+m271_84+m272_84+m273_84+m274_84+m275_84+m276_84+m277_84+m278_84+m279_84+m280_84+m281_84+m282_84+m283_84+m284_84+m285_84+m286_84+m287_84+m288_84+m289_84+m290_84+m291_84+m292_84+m293_84+m294_84+m295_84+m296_84+m297_84+m298_84+m299_84+m300_84+m301_84+m302_84+m303_84+m304_84+m305_84+m306_84+m307_84+m308_84+m309_84+m310_84+m311_84+m312_84+m313_84+m314_84+m315_84+m316_84+m317_84+m318_84+m319_84+m320_84+m321_84+m322_84+m323_84+m324_84+m325_84+m326_84+m327_84+m328_84+m329_84+m330_84+m331_84+m332_84+m333_84+m334_84+m335_84+m336_84+m337_84+m338_84+m339_84+m340_84+m341_84+m342_84+m343_84+m344_84+m345_84+m346_84+m347_84+m348_84+m349_84+m350_84+m351_84+m352_84+m353_84+m354_84+m355_84+m356_84+m357_84+m358_84+m359_84+m360_84+m361_84+m362_84+m363_84+m364_84+m365_84+m366_84+m367_84+m368_84+m369_84+m370_84+m371_84+m372_84+m373_84+m374_84+m375_84+m376_84+m377_84+m378_84+m379_84+m380_84+m381_84+b84;
   always @(posedge clk) out85 <= m1_85+m2_85+m3_85+m4_85+m5_85+m6_85+m7_85+m8_85+m9_85+m10_85+m11_85+m12_85+m13_85+m14_85+m15_85+m16_85+m17_85+m18_85+m19_85+m20_85+m21_85+m22_85+m23_85+m24_85+m25_85+m26_85+m27_85+m28_85+m29_85+m30_85+m31_85+m32_85+m33_85+m34_85+m35_85+m36_85+m37_85+m38_85+m39_85+m40_85+m41_85+m42_85+m43_85+m44_85+m45_85+m46_85+m47_85+m48_85+m49_85+m50_85+m51_85+m52_85+m53_85+m54_85+m55_85+m56_85+m57_85+m58_85+m59_85+m60_85+m61_85+m62_85+m63_85+m64_85+m65_85+m66_85+m67_85+m68_85+m69_85+m70_85+m71_85+m72_85+m73_85+m74_85+m75_85+m76_85+m77_85+m78_85+m79_85+m80_85+m81_85+m82_85+m83_85+m84_85+m85_85+m86_85+m87_85+m88_85+m89_85+m90_85+m91_85+m92_85+m93_85+m94_85+m95_85+m96_85+m97_85+m98_85+m99_85+m100_85+m101_85+m102_85+m103_85+m104_85+m105_85+m106_85+m107_85+m108_85+m109_85+m110_85+m111_85+m112_85+m113_85+m114_85+m115_85+m116_85+m117_85+m118_85+m119_85+m120_85+m121_85+m122_85+m123_85+m124_85+m125_85+m126_85+m127_85+m128_85+m129_85+m130_85+m131_85+m132_85+m133_85+m134_85+m135_85+m136_85+m137_85+m138_85+m139_85+m140_85+m141_85+m142_85+m143_85+m144_85+m145_85+m146_85+m147_85+m148_85+m149_85+m150_85+m151_85+m152_85+m153_85+m154_85+m155_85+m156_85+m157_85+m158_85+m159_85+m160_85+m161_85+m162_85+m163_85+m164_85+m165_85+m166_85+m167_85+m168_85+m169_85+m170_85+m171_85+m172_85+m173_85+m174_85+m175_85+m176_85+m177_85+m178_85+m179_85+m180_85+m181_85+m182_85+m183_85+m184_85+m185_85+m186_85+m187_85+m188_85+m189_85+m190_85+m191_85+m192_85+m193_85+m194_85+m195_85+m196_85+m197_85+m198_85+m199_85+m200_85+m201_85+m202_85+m203_85+m204_85+m205_85+m206_85+m207_85+m208_85+m209_85+m210_85+m211_85+m212_85+m213_85+m214_85+m215_85+m216_85+m217_85+m218_85+m219_85+m220_85+m221_85+m222_85+m223_85+m224_85+m225_85+m226_85+m227_85+m228_85+m229_85+m230_85+m231_85+m232_85+m233_85+m234_85+m235_85+m236_85+m237_85+m238_85+m239_85+m240_85+m241_85+m242_85+m243_85+m244_85+m245_85+m246_85+m247_85+m248_85+m249_85+m250_85+m251_85+m252_85+m253_85+m254_85+m255_85+m256_85+m257_85+m258_85+m259_85+m260_85+m261_85+m262_85+m263_85+m264_85+m265_85+m266_85+m267_85+m268_85+m269_85+m270_85+m271_85+m272_85+m273_85+m274_85+m275_85+m276_85+m277_85+m278_85+m279_85+m280_85+m281_85+m282_85+m283_85+m284_85+m285_85+m286_85+m287_85+m288_85+m289_85+m290_85+m291_85+m292_85+m293_85+m294_85+m295_85+m296_85+m297_85+m298_85+m299_85+m300_85+m301_85+m302_85+m303_85+m304_85+m305_85+m306_85+m307_85+m308_85+m309_85+m310_85+m311_85+m312_85+m313_85+m314_85+m315_85+m316_85+m317_85+m318_85+m319_85+m320_85+m321_85+m322_85+m323_85+m324_85+m325_85+m326_85+m327_85+m328_85+m329_85+m330_85+m331_85+m332_85+m333_85+m334_85+m335_85+m336_85+m337_85+m338_85+m339_85+m340_85+m341_85+m342_85+m343_85+m344_85+m345_85+m346_85+m347_85+m348_85+m349_85+m350_85+m351_85+m352_85+m353_85+m354_85+m355_85+m356_85+m357_85+m358_85+m359_85+m360_85+m361_85+m362_85+m363_85+m364_85+m365_85+m366_85+m367_85+m368_85+m369_85+m370_85+m371_85+m372_85+m373_85+m374_85+m375_85+m376_85+m377_85+m378_85+m379_85+m380_85+m381_85+b85;
   always @(posedge clk) out86 <= m1_86+m2_86+m3_86+m4_86+m5_86+m6_86+m7_86+m8_86+m9_86+m10_86+m11_86+m12_86+m13_86+m14_86+m15_86+m16_86+m17_86+m18_86+m19_86+m20_86+m21_86+m22_86+m23_86+m24_86+m25_86+m26_86+m27_86+m28_86+m29_86+m30_86+m31_86+m32_86+m33_86+m34_86+m35_86+m36_86+m37_86+m38_86+m39_86+m40_86+m41_86+m42_86+m43_86+m44_86+m45_86+m46_86+m47_86+m48_86+m49_86+m50_86+m51_86+m52_86+m53_86+m54_86+m55_86+m56_86+m57_86+m58_86+m59_86+m60_86+m61_86+m62_86+m63_86+m64_86+m65_86+m66_86+m67_86+m68_86+m69_86+m70_86+m71_86+m72_86+m73_86+m74_86+m75_86+m76_86+m77_86+m78_86+m79_86+m80_86+m81_86+m82_86+m83_86+m84_86+m85_86+m86_86+m87_86+m88_86+m89_86+m90_86+m91_86+m92_86+m93_86+m94_86+m95_86+m96_86+m97_86+m98_86+m99_86+m100_86+m101_86+m102_86+m103_86+m104_86+m105_86+m106_86+m107_86+m108_86+m109_86+m110_86+m111_86+m112_86+m113_86+m114_86+m115_86+m116_86+m117_86+m118_86+m119_86+m120_86+m121_86+m122_86+m123_86+m124_86+m125_86+m126_86+m127_86+m128_86+m129_86+m130_86+m131_86+m132_86+m133_86+m134_86+m135_86+m136_86+m137_86+m138_86+m139_86+m140_86+m141_86+m142_86+m143_86+m144_86+m145_86+m146_86+m147_86+m148_86+m149_86+m150_86+m151_86+m152_86+m153_86+m154_86+m155_86+m156_86+m157_86+m158_86+m159_86+m160_86+m161_86+m162_86+m163_86+m164_86+m165_86+m166_86+m167_86+m168_86+m169_86+m170_86+m171_86+m172_86+m173_86+m174_86+m175_86+m176_86+m177_86+m178_86+m179_86+m180_86+m181_86+m182_86+m183_86+m184_86+m185_86+m186_86+m187_86+m188_86+m189_86+m190_86+m191_86+m192_86+m193_86+m194_86+m195_86+m196_86+m197_86+m198_86+m199_86+m200_86+m201_86+m202_86+m203_86+m204_86+m205_86+m206_86+m207_86+m208_86+m209_86+m210_86+m211_86+m212_86+m213_86+m214_86+m215_86+m216_86+m217_86+m218_86+m219_86+m220_86+m221_86+m222_86+m223_86+m224_86+m225_86+m226_86+m227_86+m228_86+m229_86+m230_86+m231_86+m232_86+m233_86+m234_86+m235_86+m236_86+m237_86+m238_86+m239_86+m240_86+m241_86+m242_86+m243_86+m244_86+m245_86+m246_86+m247_86+m248_86+m249_86+m250_86+m251_86+m252_86+m253_86+m254_86+m255_86+m256_86+m257_86+m258_86+m259_86+m260_86+m261_86+m262_86+m263_86+m264_86+m265_86+m266_86+m267_86+m268_86+m269_86+m270_86+m271_86+m272_86+m273_86+m274_86+m275_86+m276_86+m277_86+m278_86+m279_86+m280_86+m281_86+m282_86+m283_86+m284_86+m285_86+m286_86+m287_86+m288_86+m289_86+m290_86+m291_86+m292_86+m293_86+m294_86+m295_86+m296_86+m297_86+m298_86+m299_86+m300_86+m301_86+m302_86+m303_86+m304_86+m305_86+m306_86+m307_86+m308_86+m309_86+m310_86+m311_86+m312_86+m313_86+m314_86+m315_86+m316_86+m317_86+m318_86+m319_86+m320_86+m321_86+m322_86+m323_86+m324_86+m325_86+m326_86+m327_86+m328_86+m329_86+m330_86+m331_86+m332_86+m333_86+m334_86+m335_86+m336_86+m337_86+m338_86+m339_86+m340_86+m341_86+m342_86+m343_86+m344_86+m345_86+m346_86+m347_86+m348_86+m349_86+m350_86+m351_86+m352_86+m353_86+m354_86+m355_86+m356_86+m357_86+m358_86+m359_86+m360_86+m361_86+m362_86+m363_86+m364_86+m365_86+m366_86+m367_86+m368_86+m369_86+m370_86+m371_86+m372_86+m373_86+m374_86+m375_86+m376_86+m377_86+m378_86+m379_86+m380_86+m381_86+b86;
   always @(posedge clk) out87 <= m1_87+m2_87+m3_87+m4_87+m5_87+m6_87+m7_87+m8_87+m9_87+m10_87+m11_87+m12_87+m13_87+m14_87+m15_87+m16_87+m17_87+m18_87+m19_87+m20_87+m21_87+m22_87+m23_87+m24_87+m25_87+m26_87+m27_87+m28_87+m29_87+m30_87+m31_87+m32_87+m33_87+m34_87+m35_87+m36_87+m37_87+m38_87+m39_87+m40_87+m41_87+m42_87+m43_87+m44_87+m45_87+m46_87+m47_87+m48_87+m49_87+m50_87+m51_87+m52_87+m53_87+m54_87+m55_87+m56_87+m57_87+m58_87+m59_87+m60_87+m61_87+m62_87+m63_87+m64_87+m65_87+m66_87+m67_87+m68_87+m69_87+m70_87+m71_87+m72_87+m73_87+m74_87+m75_87+m76_87+m77_87+m78_87+m79_87+m80_87+m81_87+m82_87+m83_87+m84_87+m85_87+m86_87+m87_87+m88_87+m89_87+m90_87+m91_87+m92_87+m93_87+m94_87+m95_87+m96_87+m97_87+m98_87+m99_87+m100_87+m101_87+m102_87+m103_87+m104_87+m105_87+m106_87+m107_87+m108_87+m109_87+m110_87+m111_87+m112_87+m113_87+m114_87+m115_87+m116_87+m117_87+m118_87+m119_87+m120_87+m121_87+m122_87+m123_87+m124_87+m125_87+m126_87+m127_87+m128_87+m129_87+m130_87+m131_87+m132_87+m133_87+m134_87+m135_87+m136_87+m137_87+m138_87+m139_87+m140_87+m141_87+m142_87+m143_87+m144_87+m145_87+m146_87+m147_87+m148_87+m149_87+m150_87+m151_87+m152_87+m153_87+m154_87+m155_87+m156_87+m157_87+m158_87+m159_87+m160_87+m161_87+m162_87+m163_87+m164_87+m165_87+m166_87+m167_87+m168_87+m169_87+m170_87+m171_87+m172_87+m173_87+m174_87+m175_87+m176_87+m177_87+m178_87+m179_87+m180_87+m181_87+m182_87+m183_87+m184_87+m185_87+m186_87+m187_87+m188_87+m189_87+m190_87+m191_87+m192_87+m193_87+m194_87+m195_87+m196_87+m197_87+m198_87+m199_87+m200_87+m201_87+m202_87+m203_87+m204_87+m205_87+m206_87+m207_87+m208_87+m209_87+m210_87+m211_87+m212_87+m213_87+m214_87+m215_87+m216_87+m217_87+m218_87+m219_87+m220_87+m221_87+m222_87+m223_87+m224_87+m225_87+m226_87+m227_87+m228_87+m229_87+m230_87+m231_87+m232_87+m233_87+m234_87+m235_87+m236_87+m237_87+m238_87+m239_87+m240_87+m241_87+m242_87+m243_87+m244_87+m245_87+m246_87+m247_87+m248_87+m249_87+m250_87+m251_87+m252_87+m253_87+m254_87+m255_87+m256_87+m257_87+m258_87+m259_87+m260_87+m261_87+m262_87+m263_87+m264_87+m265_87+m266_87+m267_87+m268_87+m269_87+m270_87+m271_87+m272_87+m273_87+m274_87+m275_87+m276_87+m277_87+m278_87+m279_87+m280_87+m281_87+m282_87+m283_87+m284_87+m285_87+m286_87+m287_87+m288_87+m289_87+m290_87+m291_87+m292_87+m293_87+m294_87+m295_87+m296_87+m297_87+m298_87+m299_87+m300_87+m301_87+m302_87+m303_87+m304_87+m305_87+m306_87+m307_87+m308_87+m309_87+m310_87+m311_87+m312_87+m313_87+m314_87+m315_87+m316_87+m317_87+m318_87+m319_87+m320_87+m321_87+m322_87+m323_87+m324_87+m325_87+m326_87+m327_87+m328_87+m329_87+m330_87+m331_87+m332_87+m333_87+m334_87+m335_87+m336_87+m337_87+m338_87+m339_87+m340_87+m341_87+m342_87+m343_87+m344_87+m345_87+m346_87+m347_87+m348_87+m349_87+m350_87+m351_87+m352_87+m353_87+m354_87+m355_87+m356_87+m357_87+m358_87+m359_87+m360_87+m361_87+m362_87+m363_87+m364_87+m365_87+m366_87+m367_87+m368_87+m369_87+m370_87+m371_87+m372_87+m373_87+m374_87+m375_87+m376_87+m377_87+m378_87+m379_87+m380_87+m381_87+b87;
   always @(posedge clk) out88 <= m1_88+m2_88+m3_88+m4_88+m5_88+m6_88+m7_88+m8_88+m9_88+m10_88+m11_88+m12_88+m13_88+m14_88+m15_88+m16_88+m17_88+m18_88+m19_88+m20_88+m21_88+m22_88+m23_88+m24_88+m25_88+m26_88+m27_88+m28_88+m29_88+m30_88+m31_88+m32_88+m33_88+m34_88+m35_88+m36_88+m37_88+m38_88+m39_88+m40_88+m41_88+m42_88+m43_88+m44_88+m45_88+m46_88+m47_88+m48_88+m49_88+m50_88+m51_88+m52_88+m53_88+m54_88+m55_88+m56_88+m57_88+m58_88+m59_88+m60_88+m61_88+m62_88+m63_88+m64_88+m65_88+m66_88+m67_88+m68_88+m69_88+m70_88+m71_88+m72_88+m73_88+m74_88+m75_88+m76_88+m77_88+m78_88+m79_88+m80_88+m81_88+m82_88+m83_88+m84_88+m85_88+m86_88+m87_88+m88_88+m89_88+m90_88+m91_88+m92_88+m93_88+m94_88+m95_88+m96_88+m97_88+m98_88+m99_88+m100_88+m101_88+m102_88+m103_88+m104_88+m105_88+m106_88+m107_88+m108_88+m109_88+m110_88+m111_88+m112_88+m113_88+m114_88+m115_88+m116_88+m117_88+m118_88+m119_88+m120_88+m121_88+m122_88+m123_88+m124_88+m125_88+m126_88+m127_88+m128_88+m129_88+m130_88+m131_88+m132_88+m133_88+m134_88+m135_88+m136_88+m137_88+m138_88+m139_88+m140_88+m141_88+m142_88+m143_88+m144_88+m145_88+m146_88+m147_88+m148_88+m149_88+m150_88+m151_88+m152_88+m153_88+m154_88+m155_88+m156_88+m157_88+m158_88+m159_88+m160_88+m161_88+m162_88+m163_88+m164_88+m165_88+m166_88+m167_88+m168_88+m169_88+m170_88+m171_88+m172_88+m173_88+m174_88+m175_88+m176_88+m177_88+m178_88+m179_88+m180_88+m181_88+m182_88+m183_88+m184_88+m185_88+m186_88+m187_88+m188_88+m189_88+m190_88+m191_88+m192_88+m193_88+m194_88+m195_88+m196_88+m197_88+m198_88+m199_88+m200_88+m201_88+m202_88+m203_88+m204_88+m205_88+m206_88+m207_88+m208_88+m209_88+m210_88+m211_88+m212_88+m213_88+m214_88+m215_88+m216_88+m217_88+m218_88+m219_88+m220_88+m221_88+m222_88+m223_88+m224_88+m225_88+m226_88+m227_88+m228_88+m229_88+m230_88+m231_88+m232_88+m233_88+m234_88+m235_88+m236_88+m237_88+m238_88+m239_88+m240_88+m241_88+m242_88+m243_88+m244_88+m245_88+m246_88+m247_88+m248_88+m249_88+m250_88+m251_88+m252_88+m253_88+m254_88+m255_88+m256_88+m257_88+m258_88+m259_88+m260_88+m261_88+m262_88+m263_88+m264_88+m265_88+m266_88+m267_88+m268_88+m269_88+m270_88+m271_88+m272_88+m273_88+m274_88+m275_88+m276_88+m277_88+m278_88+m279_88+m280_88+m281_88+m282_88+m283_88+m284_88+m285_88+m286_88+m287_88+m288_88+m289_88+m290_88+m291_88+m292_88+m293_88+m294_88+m295_88+m296_88+m297_88+m298_88+m299_88+m300_88+m301_88+m302_88+m303_88+m304_88+m305_88+m306_88+m307_88+m308_88+m309_88+m310_88+m311_88+m312_88+m313_88+m314_88+m315_88+m316_88+m317_88+m318_88+m319_88+m320_88+m321_88+m322_88+m323_88+m324_88+m325_88+m326_88+m327_88+m328_88+m329_88+m330_88+m331_88+m332_88+m333_88+m334_88+m335_88+m336_88+m337_88+m338_88+m339_88+m340_88+m341_88+m342_88+m343_88+m344_88+m345_88+m346_88+m347_88+m348_88+m349_88+m350_88+m351_88+m352_88+m353_88+m354_88+m355_88+m356_88+m357_88+m358_88+m359_88+m360_88+m361_88+m362_88+m363_88+m364_88+m365_88+m366_88+m367_88+m368_88+m369_88+m370_88+m371_88+m372_88+m373_88+m374_88+m375_88+m376_88+m377_88+m378_88+m379_88+m380_88+m381_88+b88;
   always @(posedge clk) out89 <= m1_89+m2_89+m3_89+m4_89+m5_89+m6_89+m7_89+m8_89+m9_89+m10_89+m11_89+m12_89+m13_89+m14_89+m15_89+m16_89+m17_89+m18_89+m19_89+m20_89+m21_89+m22_89+m23_89+m24_89+m25_89+m26_89+m27_89+m28_89+m29_89+m30_89+m31_89+m32_89+m33_89+m34_89+m35_89+m36_89+m37_89+m38_89+m39_89+m40_89+m41_89+m42_89+m43_89+m44_89+m45_89+m46_89+m47_89+m48_89+m49_89+m50_89+m51_89+m52_89+m53_89+m54_89+m55_89+m56_89+m57_89+m58_89+m59_89+m60_89+m61_89+m62_89+m63_89+m64_89+m65_89+m66_89+m67_89+m68_89+m69_89+m70_89+m71_89+m72_89+m73_89+m74_89+m75_89+m76_89+m77_89+m78_89+m79_89+m80_89+m81_89+m82_89+m83_89+m84_89+m85_89+m86_89+m87_89+m88_89+m89_89+m90_89+m91_89+m92_89+m93_89+m94_89+m95_89+m96_89+m97_89+m98_89+m99_89+m100_89+m101_89+m102_89+m103_89+m104_89+m105_89+m106_89+m107_89+m108_89+m109_89+m110_89+m111_89+m112_89+m113_89+m114_89+m115_89+m116_89+m117_89+m118_89+m119_89+m120_89+m121_89+m122_89+m123_89+m124_89+m125_89+m126_89+m127_89+m128_89+m129_89+m130_89+m131_89+m132_89+m133_89+m134_89+m135_89+m136_89+m137_89+m138_89+m139_89+m140_89+m141_89+m142_89+m143_89+m144_89+m145_89+m146_89+m147_89+m148_89+m149_89+m150_89+m151_89+m152_89+m153_89+m154_89+m155_89+m156_89+m157_89+m158_89+m159_89+m160_89+m161_89+m162_89+m163_89+m164_89+m165_89+m166_89+m167_89+m168_89+m169_89+m170_89+m171_89+m172_89+m173_89+m174_89+m175_89+m176_89+m177_89+m178_89+m179_89+m180_89+m181_89+m182_89+m183_89+m184_89+m185_89+m186_89+m187_89+m188_89+m189_89+m190_89+m191_89+m192_89+m193_89+m194_89+m195_89+m196_89+m197_89+m198_89+m199_89+m200_89+m201_89+m202_89+m203_89+m204_89+m205_89+m206_89+m207_89+m208_89+m209_89+m210_89+m211_89+m212_89+m213_89+m214_89+m215_89+m216_89+m217_89+m218_89+m219_89+m220_89+m221_89+m222_89+m223_89+m224_89+m225_89+m226_89+m227_89+m228_89+m229_89+m230_89+m231_89+m232_89+m233_89+m234_89+m235_89+m236_89+m237_89+m238_89+m239_89+m240_89+m241_89+m242_89+m243_89+m244_89+m245_89+m246_89+m247_89+m248_89+m249_89+m250_89+m251_89+m252_89+m253_89+m254_89+m255_89+m256_89+m257_89+m258_89+m259_89+m260_89+m261_89+m262_89+m263_89+m264_89+m265_89+m266_89+m267_89+m268_89+m269_89+m270_89+m271_89+m272_89+m273_89+m274_89+m275_89+m276_89+m277_89+m278_89+m279_89+m280_89+m281_89+m282_89+m283_89+m284_89+m285_89+m286_89+m287_89+m288_89+m289_89+m290_89+m291_89+m292_89+m293_89+m294_89+m295_89+m296_89+m297_89+m298_89+m299_89+m300_89+m301_89+m302_89+m303_89+m304_89+m305_89+m306_89+m307_89+m308_89+m309_89+m310_89+m311_89+m312_89+m313_89+m314_89+m315_89+m316_89+m317_89+m318_89+m319_89+m320_89+m321_89+m322_89+m323_89+m324_89+m325_89+m326_89+m327_89+m328_89+m329_89+m330_89+m331_89+m332_89+m333_89+m334_89+m335_89+m336_89+m337_89+m338_89+m339_89+m340_89+m341_89+m342_89+m343_89+m344_89+m345_89+m346_89+m347_89+m348_89+m349_89+m350_89+m351_89+m352_89+m353_89+m354_89+m355_89+m356_89+m357_89+m358_89+m359_89+m360_89+m361_89+m362_89+m363_89+m364_89+m365_89+m366_89+m367_89+m368_89+m369_89+m370_89+m371_89+m372_89+m373_89+m374_89+m375_89+m376_89+m377_89+m378_89+m379_89+m380_89+m381_89+b89;
   always @(posedge clk) out90 <= m1_90+m2_90+m3_90+m4_90+m5_90+m6_90+m7_90+m8_90+m9_90+m10_90+m11_90+m12_90+m13_90+m14_90+m15_90+m16_90+m17_90+m18_90+m19_90+m20_90+m21_90+m22_90+m23_90+m24_90+m25_90+m26_90+m27_90+m28_90+m29_90+m30_90+m31_90+m32_90+m33_90+m34_90+m35_90+m36_90+m37_90+m38_90+m39_90+m40_90+m41_90+m42_90+m43_90+m44_90+m45_90+m46_90+m47_90+m48_90+m49_90+m50_90+m51_90+m52_90+m53_90+m54_90+m55_90+m56_90+m57_90+m58_90+m59_90+m60_90+m61_90+m62_90+m63_90+m64_90+m65_90+m66_90+m67_90+m68_90+m69_90+m70_90+m71_90+m72_90+m73_90+m74_90+m75_90+m76_90+m77_90+m78_90+m79_90+m80_90+m81_90+m82_90+m83_90+m84_90+m85_90+m86_90+m87_90+m88_90+m89_90+m90_90+m91_90+m92_90+m93_90+m94_90+m95_90+m96_90+m97_90+m98_90+m99_90+m100_90+m101_90+m102_90+m103_90+m104_90+m105_90+m106_90+m107_90+m108_90+m109_90+m110_90+m111_90+m112_90+m113_90+m114_90+m115_90+m116_90+m117_90+m118_90+m119_90+m120_90+m121_90+m122_90+m123_90+m124_90+m125_90+m126_90+m127_90+m128_90+m129_90+m130_90+m131_90+m132_90+m133_90+m134_90+m135_90+m136_90+m137_90+m138_90+m139_90+m140_90+m141_90+m142_90+m143_90+m144_90+m145_90+m146_90+m147_90+m148_90+m149_90+m150_90+m151_90+m152_90+m153_90+m154_90+m155_90+m156_90+m157_90+m158_90+m159_90+m160_90+m161_90+m162_90+m163_90+m164_90+m165_90+m166_90+m167_90+m168_90+m169_90+m170_90+m171_90+m172_90+m173_90+m174_90+m175_90+m176_90+m177_90+m178_90+m179_90+m180_90+m181_90+m182_90+m183_90+m184_90+m185_90+m186_90+m187_90+m188_90+m189_90+m190_90+m191_90+m192_90+m193_90+m194_90+m195_90+m196_90+m197_90+m198_90+m199_90+m200_90+m201_90+m202_90+m203_90+m204_90+m205_90+m206_90+m207_90+m208_90+m209_90+m210_90+m211_90+m212_90+m213_90+m214_90+m215_90+m216_90+m217_90+m218_90+m219_90+m220_90+m221_90+m222_90+m223_90+m224_90+m225_90+m226_90+m227_90+m228_90+m229_90+m230_90+m231_90+m232_90+m233_90+m234_90+m235_90+m236_90+m237_90+m238_90+m239_90+m240_90+m241_90+m242_90+m243_90+m244_90+m245_90+m246_90+m247_90+m248_90+m249_90+m250_90+m251_90+m252_90+m253_90+m254_90+m255_90+m256_90+m257_90+m258_90+m259_90+m260_90+m261_90+m262_90+m263_90+m264_90+m265_90+m266_90+m267_90+m268_90+m269_90+m270_90+m271_90+m272_90+m273_90+m274_90+m275_90+m276_90+m277_90+m278_90+m279_90+m280_90+m281_90+m282_90+m283_90+m284_90+m285_90+m286_90+m287_90+m288_90+m289_90+m290_90+m291_90+m292_90+m293_90+m294_90+m295_90+m296_90+m297_90+m298_90+m299_90+m300_90+m301_90+m302_90+m303_90+m304_90+m305_90+m306_90+m307_90+m308_90+m309_90+m310_90+m311_90+m312_90+m313_90+m314_90+m315_90+m316_90+m317_90+m318_90+m319_90+m320_90+m321_90+m322_90+m323_90+m324_90+m325_90+m326_90+m327_90+m328_90+m329_90+m330_90+m331_90+m332_90+m333_90+m334_90+m335_90+m336_90+m337_90+m338_90+m339_90+m340_90+m341_90+m342_90+m343_90+m344_90+m345_90+m346_90+m347_90+m348_90+m349_90+m350_90+m351_90+m352_90+m353_90+m354_90+m355_90+m356_90+m357_90+m358_90+m359_90+m360_90+m361_90+m362_90+m363_90+m364_90+m365_90+m366_90+m367_90+m368_90+m369_90+m370_90+m371_90+m372_90+m373_90+m374_90+m375_90+m376_90+m377_90+m378_90+m379_90+m380_90+m381_90+b90;
   always @(posedge clk) out91 <= m1_91+m2_91+m3_91+m4_91+m5_91+m6_91+m7_91+m8_91+m9_91+m10_91+m11_91+m12_91+m13_91+m14_91+m15_91+m16_91+m17_91+m18_91+m19_91+m20_91+m21_91+m22_91+m23_91+m24_91+m25_91+m26_91+m27_91+m28_91+m29_91+m30_91+m31_91+m32_91+m33_91+m34_91+m35_91+m36_91+m37_91+m38_91+m39_91+m40_91+m41_91+m42_91+m43_91+m44_91+m45_91+m46_91+m47_91+m48_91+m49_91+m50_91+m51_91+m52_91+m53_91+m54_91+m55_91+m56_91+m57_91+m58_91+m59_91+m60_91+m61_91+m62_91+m63_91+m64_91+m65_91+m66_91+m67_91+m68_91+m69_91+m70_91+m71_91+m72_91+m73_91+m74_91+m75_91+m76_91+m77_91+m78_91+m79_91+m80_91+m81_91+m82_91+m83_91+m84_91+m85_91+m86_91+m87_91+m88_91+m89_91+m90_91+m91_91+m92_91+m93_91+m94_91+m95_91+m96_91+m97_91+m98_91+m99_91+m100_91+m101_91+m102_91+m103_91+m104_91+m105_91+m106_91+m107_91+m108_91+m109_91+m110_91+m111_91+m112_91+m113_91+m114_91+m115_91+m116_91+m117_91+m118_91+m119_91+m120_91+m121_91+m122_91+m123_91+m124_91+m125_91+m126_91+m127_91+m128_91+m129_91+m130_91+m131_91+m132_91+m133_91+m134_91+m135_91+m136_91+m137_91+m138_91+m139_91+m140_91+m141_91+m142_91+m143_91+m144_91+m145_91+m146_91+m147_91+m148_91+m149_91+m150_91+m151_91+m152_91+m153_91+m154_91+m155_91+m156_91+m157_91+m158_91+m159_91+m160_91+m161_91+m162_91+m163_91+m164_91+m165_91+m166_91+m167_91+m168_91+m169_91+m170_91+m171_91+m172_91+m173_91+m174_91+m175_91+m176_91+m177_91+m178_91+m179_91+m180_91+m181_91+m182_91+m183_91+m184_91+m185_91+m186_91+m187_91+m188_91+m189_91+m190_91+m191_91+m192_91+m193_91+m194_91+m195_91+m196_91+m197_91+m198_91+m199_91+m200_91+m201_91+m202_91+m203_91+m204_91+m205_91+m206_91+m207_91+m208_91+m209_91+m210_91+m211_91+m212_91+m213_91+m214_91+m215_91+m216_91+m217_91+m218_91+m219_91+m220_91+m221_91+m222_91+m223_91+m224_91+m225_91+m226_91+m227_91+m228_91+m229_91+m230_91+m231_91+m232_91+m233_91+m234_91+m235_91+m236_91+m237_91+m238_91+m239_91+m240_91+m241_91+m242_91+m243_91+m244_91+m245_91+m246_91+m247_91+m248_91+m249_91+m250_91+m251_91+m252_91+m253_91+m254_91+m255_91+m256_91+m257_91+m258_91+m259_91+m260_91+m261_91+m262_91+m263_91+m264_91+m265_91+m266_91+m267_91+m268_91+m269_91+m270_91+m271_91+m272_91+m273_91+m274_91+m275_91+m276_91+m277_91+m278_91+m279_91+m280_91+m281_91+m282_91+m283_91+m284_91+m285_91+m286_91+m287_91+m288_91+m289_91+m290_91+m291_91+m292_91+m293_91+m294_91+m295_91+m296_91+m297_91+m298_91+m299_91+m300_91+m301_91+m302_91+m303_91+m304_91+m305_91+m306_91+m307_91+m308_91+m309_91+m310_91+m311_91+m312_91+m313_91+m314_91+m315_91+m316_91+m317_91+m318_91+m319_91+m320_91+m321_91+m322_91+m323_91+m324_91+m325_91+m326_91+m327_91+m328_91+m329_91+m330_91+m331_91+m332_91+m333_91+m334_91+m335_91+m336_91+m337_91+m338_91+m339_91+m340_91+m341_91+m342_91+m343_91+m344_91+m345_91+m346_91+m347_91+m348_91+m349_91+m350_91+m351_91+m352_91+m353_91+m354_91+m355_91+m356_91+m357_91+m358_91+m359_91+m360_91+m361_91+m362_91+m363_91+m364_91+m365_91+m366_91+m367_91+m368_91+m369_91+m370_91+m371_91+m372_91+m373_91+m374_91+m375_91+m376_91+m377_91+m378_91+m379_91+m380_91+m381_91+b91;
   always @(posedge clk) out92 <= m1_92+m2_92+m3_92+m4_92+m5_92+m6_92+m7_92+m8_92+m9_92+m10_92+m11_92+m12_92+m13_92+m14_92+m15_92+m16_92+m17_92+m18_92+m19_92+m20_92+m21_92+m22_92+m23_92+m24_92+m25_92+m26_92+m27_92+m28_92+m29_92+m30_92+m31_92+m32_92+m33_92+m34_92+m35_92+m36_92+m37_92+m38_92+m39_92+m40_92+m41_92+m42_92+m43_92+m44_92+m45_92+m46_92+m47_92+m48_92+m49_92+m50_92+m51_92+m52_92+m53_92+m54_92+m55_92+m56_92+m57_92+m58_92+m59_92+m60_92+m61_92+m62_92+m63_92+m64_92+m65_92+m66_92+m67_92+m68_92+m69_92+m70_92+m71_92+m72_92+m73_92+m74_92+m75_92+m76_92+m77_92+m78_92+m79_92+m80_92+m81_92+m82_92+m83_92+m84_92+m85_92+m86_92+m87_92+m88_92+m89_92+m90_92+m91_92+m92_92+m93_92+m94_92+m95_92+m96_92+m97_92+m98_92+m99_92+m100_92+m101_92+m102_92+m103_92+m104_92+m105_92+m106_92+m107_92+m108_92+m109_92+m110_92+m111_92+m112_92+m113_92+m114_92+m115_92+m116_92+m117_92+m118_92+m119_92+m120_92+m121_92+m122_92+m123_92+m124_92+m125_92+m126_92+m127_92+m128_92+m129_92+m130_92+m131_92+m132_92+m133_92+m134_92+m135_92+m136_92+m137_92+m138_92+m139_92+m140_92+m141_92+m142_92+m143_92+m144_92+m145_92+m146_92+m147_92+m148_92+m149_92+m150_92+m151_92+m152_92+m153_92+m154_92+m155_92+m156_92+m157_92+m158_92+m159_92+m160_92+m161_92+m162_92+m163_92+m164_92+m165_92+m166_92+m167_92+m168_92+m169_92+m170_92+m171_92+m172_92+m173_92+m174_92+m175_92+m176_92+m177_92+m178_92+m179_92+m180_92+m181_92+m182_92+m183_92+m184_92+m185_92+m186_92+m187_92+m188_92+m189_92+m190_92+m191_92+m192_92+m193_92+m194_92+m195_92+m196_92+m197_92+m198_92+m199_92+m200_92+m201_92+m202_92+m203_92+m204_92+m205_92+m206_92+m207_92+m208_92+m209_92+m210_92+m211_92+m212_92+m213_92+m214_92+m215_92+m216_92+m217_92+m218_92+m219_92+m220_92+m221_92+m222_92+m223_92+m224_92+m225_92+m226_92+m227_92+m228_92+m229_92+m230_92+m231_92+m232_92+m233_92+m234_92+m235_92+m236_92+m237_92+m238_92+m239_92+m240_92+m241_92+m242_92+m243_92+m244_92+m245_92+m246_92+m247_92+m248_92+m249_92+m250_92+m251_92+m252_92+m253_92+m254_92+m255_92+m256_92+m257_92+m258_92+m259_92+m260_92+m261_92+m262_92+m263_92+m264_92+m265_92+m266_92+m267_92+m268_92+m269_92+m270_92+m271_92+m272_92+m273_92+m274_92+m275_92+m276_92+m277_92+m278_92+m279_92+m280_92+m281_92+m282_92+m283_92+m284_92+m285_92+m286_92+m287_92+m288_92+m289_92+m290_92+m291_92+m292_92+m293_92+m294_92+m295_92+m296_92+m297_92+m298_92+m299_92+m300_92+m301_92+m302_92+m303_92+m304_92+m305_92+m306_92+m307_92+m308_92+m309_92+m310_92+m311_92+m312_92+m313_92+m314_92+m315_92+m316_92+m317_92+m318_92+m319_92+m320_92+m321_92+m322_92+m323_92+m324_92+m325_92+m326_92+m327_92+m328_92+m329_92+m330_92+m331_92+m332_92+m333_92+m334_92+m335_92+m336_92+m337_92+m338_92+m339_92+m340_92+m341_92+m342_92+m343_92+m344_92+m345_92+m346_92+m347_92+m348_92+m349_92+m350_92+m351_92+m352_92+m353_92+m354_92+m355_92+m356_92+m357_92+m358_92+m359_92+m360_92+m361_92+m362_92+m363_92+m364_92+m365_92+m366_92+m367_92+m368_92+m369_92+m370_92+m371_92+m372_92+m373_92+m374_92+m375_92+m376_92+m377_92+m378_92+m379_92+m380_92+m381_92+b92;
   always @(posedge clk) out93 <= m1_93+m2_93+m3_93+m4_93+m5_93+m6_93+m7_93+m8_93+m9_93+m10_93+m11_93+m12_93+m13_93+m14_93+m15_93+m16_93+m17_93+m18_93+m19_93+m20_93+m21_93+m22_93+m23_93+m24_93+m25_93+m26_93+m27_93+m28_93+m29_93+m30_93+m31_93+m32_93+m33_93+m34_93+m35_93+m36_93+m37_93+m38_93+m39_93+m40_93+m41_93+m42_93+m43_93+m44_93+m45_93+m46_93+m47_93+m48_93+m49_93+m50_93+m51_93+m52_93+m53_93+m54_93+m55_93+m56_93+m57_93+m58_93+m59_93+m60_93+m61_93+m62_93+m63_93+m64_93+m65_93+m66_93+m67_93+m68_93+m69_93+m70_93+m71_93+m72_93+m73_93+m74_93+m75_93+m76_93+m77_93+m78_93+m79_93+m80_93+m81_93+m82_93+m83_93+m84_93+m85_93+m86_93+m87_93+m88_93+m89_93+m90_93+m91_93+m92_93+m93_93+m94_93+m95_93+m96_93+m97_93+m98_93+m99_93+m100_93+m101_93+m102_93+m103_93+m104_93+m105_93+m106_93+m107_93+m108_93+m109_93+m110_93+m111_93+m112_93+m113_93+m114_93+m115_93+m116_93+m117_93+m118_93+m119_93+m120_93+m121_93+m122_93+m123_93+m124_93+m125_93+m126_93+m127_93+m128_93+m129_93+m130_93+m131_93+m132_93+m133_93+m134_93+m135_93+m136_93+m137_93+m138_93+m139_93+m140_93+m141_93+m142_93+m143_93+m144_93+m145_93+m146_93+m147_93+m148_93+m149_93+m150_93+m151_93+m152_93+m153_93+m154_93+m155_93+m156_93+m157_93+m158_93+m159_93+m160_93+m161_93+m162_93+m163_93+m164_93+m165_93+m166_93+m167_93+m168_93+m169_93+m170_93+m171_93+m172_93+m173_93+m174_93+m175_93+m176_93+m177_93+m178_93+m179_93+m180_93+m181_93+m182_93+m183_93+m184_93+m185_93+m186_93+m187_93+m188_93+m189_93+m190_93+m191_93+m192_93+m193_93+m194_93+m195_93+m196_93+m197_93+m198_93+m199_93+m200_93+m201_93+m202_93+m203_93+m204_93+m205_93+m206_93+m207_93+m208_93+m209_93+m210_93+m211_93+m212_93+m213_93+m214_93+m215_93+m216_93+m217_93+m218_93+m219_93+m220_93+m221_93+m222_93+m223_93+m224_93+m225_93+m226_93+m227_93+m228_93+m229_93+m230_93+m231_93+m232_93+m233_93+m234_93+m235_93+m236_93+m237_93+m238_93+m239_93+m240_93+m241_93+m242_93+m243_93+m244_93+m245_93+m246_93+m247_93+m248_93+m249_93+m250_93+m251_93+m252_93+m253_93+m254_93+m255_93+m256_93+m257_93+m258_93+m259_93+m260_93+m261_93+m262_93+m263_93+m264_93+m265_93+m266_93+m267_93+m268_93+m269_93+m270_93+m271_93+m272_93+m273_93+m274_93+m275_93+m276_93+m277_93+m278_93+m279_93+m280_93+m281_93+m282_93+m283_93+m284_93+m285_93+m286_93+m287_93+m288_93+m289_93+m290_93+m291_93+m292_93+m293_93+m294_93+m295_93+m296_93+m297_93+m298_93+m299_93+m300_93+m301_93+m302_93+m303_93+m304_93+m305_93+m306_93+m307_93+m308_93+m309_93+m310_93+m311_93+m312_93+m313_93+m314_93+m315_93+m316_93+m317_93+m318_93+m319_93+m320_93+m321_93+m322_93+m323_93+m324_93+m325_93+m326_93+m327_93+m328_93+m329_93+m330_93+m331_93+m332_93+m333_93+m334_93+m335_93+m336_93+m337_93+m338_93+m339_93+m340_93+m341_93+m342_93+m343_93+m344_93+m345_93+m346_93+m347_93+m348_93+m349_93+m350_93+m351_93+m352_93+m353_93+m354_93+m355_93+m356_93+m357_93+m358_93+m359_93+m360_93+m361_93+m362_93+m363_93+m364_93+m365_93+m366_93+m367_93+m368_93+m369_93+m370_93+m371_93+m372_93+m373_93+m374_93+m375_93+m376_93+m377_93+m378_93+m379_93+m380_93+m381_93+b93;
   always @(posedge clk) out94 <= m1_94+m2_94+m3_94+m4_94+m5_94+m6_94+m7_94+m8_94+m9_94+m10_94+m11_94+m12_94+m13_94+m14_94+m15_94+m16_94+m17_94+m18_94+m19_94+m20_94+m21_94+m22_94+m23_94+m24_94+m25_94+m26_94+m27_94+m28_94+m29_94+m30_94+m31_94+m32_94+m33_94+m34_94+m35_94+m36_94+m37_94+m38_94+m39_94+m40_94+m41_94+m42_94+m43_94+m44_94+m45_94+m46_94+m47_94+m48_94+m49_94+m50_94+m51_94+m52_94+m53_94+m54_94+m55_94+m56_94+m57_94+m58_94+m59_94+m60_94+m61_94+m62_94+m63_94+m64_94+m65_94+m66_94+m67_94+m68_94+m69_94+m70_94+m71_94+m72_94+m73_94+m74_94+m75_94+m76_94+m77_94+m78_94+m79_94+m80_94+m81_94+m82_94+m83_94+m84_94+m85_94+m86_94+m87_94+m88_94+m89_94+m90_94+m91_94+m92_94+m93_94+m94_94+m95_94+m96_94+m97_94+m98_94+m99_94+m100_94+m101_94+m102_94+m103_94+m104_94+m105_94+m106_94+m107_94+m108_94+m109_94+m110_94+m111_94+m112_94+m113_94+m114_94+m115_94+m116_94+m117_94+m118_94+m119_94+m120_94+m121_94+m122_94+m123_94+m124_94+m125_94+m126_94+m127_94+m128_94+m129_94+m130_94+m131_94+m132_94+m133_94+m134_94+m135_94+m136_94+m137_94+m138_94+m139_94+m140_94+m141_94+m142_94+m143_94+m144_94+m145_94+m146_94+m147_94+m148_94+m149_94+m150_94+m151_94+m152_94+m153_94+m154_94+m155_94+m156_94+m157_94+m158_94+m159_94+m160_94+m161_94+m162_94+m163_94+m164_94+m165_94+m166_94+m167_94+m168_94+m169_94+m170_94+m171_94+m172_94+m173_94+m174_94+m175_94+m176_94+m177_94+m178_94+m179_94+m180_94+m181_94+m182_94+m183_94+m184_94+m185_94+m186_94+m187_94+m188_94+m189_94+m190_94+m191_94+m192_94+m193_94+m194_94+m195_94+m196_94+m197_94+m198_94+m199_94+m200_94+m201_94+m202_94+m203_94+m204_94+m205_94+m206_94+m207_94+m208_94+m209_94+m210_94+m211_94+m212_94+m213_94+m214_94+m215_94+m216_94+m217_94+m218_94+m219_94+m220_94+m221_94+m222_94+m223_94+m224_94+m225_94+m226_94+m227_94+m228_94+m229_94+m230_94+m231_94+m232_94+m233_94+m234_94+m235_94+m236_94+m237_94+m238_94+m239_94+m240_94+m241_94+m242_94+m243_94+m244_94+m245_94+m246_94+m247_94+m248_94+m249_94+m250_94+m251_94+m252_94+m253_94+m254_94+m255_94+m256_94+m257_94+m258_94+m259_94+m260_94+m261_94+m262_94+m263_94+m264_94+m265_94+m266_94+m267_94+m268_94+m269_94+m270_94+m271_94+m272_94+m273_94+m274_94+m275_94+m276_94+m277_94+m278_94+m279_94+m280_94+m281_94+m282_94+m283_94+m284_94+m285_94+m286_94+m287_94+m288_94+m289_94+m290_94+m291_94+m292_94+m293_94+m294_94+m295_94+m296_94+m297_94+m298_94+m299_94+m300_94+m301_94+m302_94+m303_94+m304_94+m305_94+m306_94+m307_94+m308_94+m309_94+m310_94+m311_94+m312_94+m313_94+m314_94+m315_94+m316_94+m317_94+m318_94+m319_94+m320_94+m321_94+m322_94+m323_94+m324_94+m325_94+m326_94+m327_94+m328_94+m329_94+m330_94+m331_94+m332_94+m333_94+m334_94+m335_94+m336_94+m337_94+m338_94+m339_94+m340_94+m341_94+m342_94+m343_94+m344_94+m345_94+m346_94+m347_94+m348_94+m349_94+m350_94+m351_94+m352_94+m353_94+m354_94+m355_94+m356_94+m357_94+m358_94+m359_94+m360_94+m361_94+m362_94+m363_94+m364_94+m365_94+m366_94+m367_94+m368_94+m369_94+m370_94+m371_94+m372_94+m373_94+m374_94+m375_94+m376_94+m377_94+m378_94+m379_94+m380_94+m381_94+b94;
   always @(posedge clk) out95 <= m1_95+m2_95+m3_95+m4_95+m5_95+m6_95+m7_95+m8_95+m9_95+m10_95+m11_95+m12_95+m13_95+m14_95+m15_95+m16_95+m17_95+m18_95+m19_95+m20_95+m21_95+m22_95+m23_95+m24_95+m25_95+m26_95+m27_95+m28_95+m29_95+m30_95+m31_95+m32_95+m33_95+m34_95+m35_95+m36_95+m37_95+m38_95+m39_95+m40_95+m41_95+m42_95+m43_95+m44_95+m45_95+m46_95+m47_95+m48_95+m49_95+m50_95+m51_95+m52_95+m53_95+m54_95+m55_95+m56_95+m57_95+m58_95+m59_95+m60_95+m61_95+m62_95+m63_95+m64_95+m65_95+m66_95+m67_95+m68_95+m69_95+m70_95+m71_95+m72_95+m73_95+m74_95+m75_95+m76_95+m77_95+m78_95+m79_95+m80_95+m81_95+m82_95+m83_95+m84_95+m85_95+m86_95+m87_95+m88_95+m89_95+m90_95+m91_95+m92_95+m93_95+m94_95+m95_95+m96_95+m97_95+m98_95+m99_95+m100_95+m101_95+m102_95+m103_95+m104_95+m105_95+m106_95+m107_95+m108_95+m109_95+m110_95+m111_95+m112_95+m113_95+m114_95+m115_95+m116_95+m117_95+m118_95+m119_95+m120_95+m121_95+m122_95+m123_95+m124_95+m125_95+m126_95+m127_95+m128_95+m129_95+m130_95+m131_95+m132_95+m133_95+m134_95+m135_95+m136_95+m137_95+m138_95+m139_95+m140_95+m141_95+m142_95+m143_95+m144_95+m145_95+m146_95+m147_95+m148_95+m149_95+m150_95+m151_95+m152_95+m153_95+m154_95+m155_95+m156_95+m157_95+m158_95+m159_95+m160_95+m161_95+m162_95+m163_95+m164_95+m165_95+m166_95+m167_95+m168_95+m169_95+m170_95+m171_95+m172_95+m173_95+m174_95+m175_95+m176_95+m177_95+m178_95+m179_95+m180_95+m181_95+m182_95+m183_95+m184_95+m185_95+m186_95+m187_95+m188_95+m189_95+m190_95+m191_95+m192_95+m193_95+m194_95+m195_95+m196_95+m197_95+m198_95+m199_95+m200_95+m201_95+m202_95+m203_95+m204_95+m205_95+m206_95+m207_95+m208_95+m209_95+m210_95+m211_95+m212_95+m213_95+m214_95+m215_95+m216_95+m217_95+m218_95+m219_95+m220_95+m221_95+m222_95+m223_95+m224_95+m225_95+m226_95+m227_95+m228_95+m229_95+m230_95+m231_95+m232_95+m233_95+m234_95+m235_95+m236_95+m237_95+m238_95+m239_95+m240_95+m241_95+m242_95+m243_95+m244_95+m245_95+m246_95+m247_95+m248_95+m249_95+m250_95+m251_95+m252_95+m253_95+m254_95+m255_95+m256_95+m257_95+m258_95+m259_95+m260_95+m261_95+m262_95+m263_95+m264_95+m265_95+m266_95+m267_95+m268_95+m269_95+m270_95+m271_95+m272_95+m273_95+m274_95+m275_95+m276_95+m277_95+m278_95+m279_95+m280_95+m281_95+m282_95+m283_95+m284_95+m285_95+m286_95+m287_95+m288_95+m289_95+m290_95+m291_95+m292_95+m293_95+m294_95+m295_95+m296_95+m297_95+m298_95+m299_95+m300_95+m301_95+m302_95+m303_95+m304_95+m305_95+m306_95+m307_95+m308_95+m309_95+m310_95+m311_95+m312_95+m313_95+m314_95+m315_95+m316_95+m317_95+m318_95+m319_95+m320_95+m321_95+m322_95+m323_95+m324_95+m325_95+m326_95+m327_95+m328_95+m329_95+m330_95+m331_95+m332_95+m333_95+m334_95+m335_95+m336_95+m337_95+m338_95+m339_95+m340_95+m341_95+m342_95+m343_95+m344_95+m345_95+m346_95+m347_95+m348_95+m349_95+m350_95+m351_95+m352_95+m353_95+m354_95+m355_95+m356_95+m357_95+m358_95+m359_95+m360_95+m361_95+m362_95+m363_95+m364_95+m365_95+m366_95+m367_95+m368_95+m369_95+m370_95+m371_95+m372_95+m373_95+m374_95+m375_95+m376_95+m377_95+m378_95+m379_95+m380_95+m381_95+b95;
   always @(posedge clk) out96 <= m1_96+m2_96+m3_96+m4_96+m5_96+m6_96+m7_96+m8_96+m9_96+m10_96+m11_96+m12_96+m13_96+m14_96+m15_96+m16_96+m17_96+m18_96+m19_96+m20_96+m21_96+m22_96+m23_96+m24_96+m25_96+m26_96+m27_96+m28_96+m29_96+m30_96+m31_96+m32_96+m33_96+m34_96+m35_96+m36_96+m37_96+m38_96+m39_96+m40_96+m41_96+m42_96+m43_96+m44_96+m45_96+m46_96+m47_96+m48_96+m49_96+m50_96+m51_96+m52_96+m53_96+m54_96+m55_96+m56_96+m57_96+m58_96+m59_96+m60_96+m61_96+m62_96+m63_96+m64_96+m65_96+m66_96+m67_96+m68_96+m69_96+m70_96+m71_96+m72_96+m73_96+m74_96+m75_96+m76_96+m77_96+m78_96+m79_96+m80_96+m81_96+m82_96+m83_96+m84_96+m85_96+m86_96+m87_96+m88_96+m89_96+m90_96+m91_96+m92_96+m93_96+m94_96+m95_96+m96_96+m97_96+m98_96+m99_96+m100_96+m101_96+m102_96+m103_96+m104_96+m105_96+m106_96+m107_96+m108_96+m109_96+m110_96+m111_96+m112_96+m113_96+m114_96+m115_96+m116_96+m117_96+m118_96+m119_96+m120_96+m121_96+m122_96+m123_96+m124_96+m125_96+m126_96+m127_96+m128_96+m129_96+m130_96+m131_96+m132_96+m133_96+m134_96+m135_96+m136_96+m137_96+m138_96+m139_96+m140_96+m141_96+m142_96+m143_96+m144_96+m145_96+m146_96+m147_96+m148_96+m149_96+m150_96+m151_96+m152_96+m153_96+m154_96+m155_96+m156_96+m157_96+m158_96+m159_96+m160_96+m161_96+m162_96+m163_96+m164_96+m165_96+m166_96+m167_96+m168_96+m169_96+m170_96+m171_96+m172_96+m173_96+m174_96+m175_96+m176_96+m177_96+m178_96+m179_96+m180_96+m181_96+m182_96+m183_96+m184_96+m185_96+m186_96+m187_96+m188_96+m189_96+m190_96+m191_96+m192_96+m193_96+m194_96+m195_96+m196_96+m197_96+m198_96+m199_96+m200_96+m201_96+m202_96+m203_96+m204_96+m205_96+m206_96+m207_96+m208_96+m209_96+m210_96+m211_96+m212_96+m213_96+m214_96+m215_96+m216_96+m217_96+m218_96+m219_96+m220_96+m221_96+m222_96+m223_96+m224_96+m225_96+m226_96+m227_96+m228_96+m229_96+m230_96+m231_96+m232_96+m233_96+m234_96+m235_96+m236_96+m237_96+m238_96+m239_96+m240_96+m241_96+m242_96+m243_96+m244_96+m245_96+m246_96+m247_96+m248_96+m249_96+m250_96+m251_96+m252_96+m253_96+m254_96+m255_96+m256_96+m257_96+m258_96+m259_96+m260_96+m261_96+m262_96+m263_96+m264_96+m265_96+m266_96+m267_96+m268_96+m269_96+m270_96+m271_96+m272_96+m273_96+m274_96+m275_96+m276_96+m277_96+m278_96+m279_96+m280_96+m281_96+m282_96+m283_96+m284_96+m285_96+m286_96+m287_96+m288_96+m289_96+m290_96+m291_96+m292_96+m293_96+m294_96+m295_96+m296_96+m297_96+m298_96+m299_96+m300_96+m301_96+m302_96+m303_96+m304_96+m305_96+m306_96+m307_96+m308_96+m309_96+m310_96+m311_96+m312_96+m313_96+m314_96+m315_96+m316_96+m317_96+m318_96+m319_96+m320_96+m321_96+m322_96+m323_96+m324_96+m325_96+m326_96+m327_96+m328_96+m329_96+m330_96+m331_96+m332_96+m333_96+m334_96+m335_96+m336_96+m337_96+m338_96+m339_96+m340_96+m341_96+m342_96+m343_96+m344_96+m345_96+m346_96+m347_96+m348_96+m349_96+m350_96+m351_96+m352_96+m353_96+m354_96+m355_96+m356_96+m357_96+m358_96+m359_96+m360_96+m361_96+m362_96+m363_96+m364_96+m365_96+m366_96+m367_96+m368_96+m369_96+m370_96+m371_96+m372_96+m373_96+m374_96+m375_96+m376_96+m377_96+m378_96+m379_96+m380_96+m381_96+b96;
   always @(posedge clk) out97 <= m1_97+m2_97+m3_97+m4_97+m5_97+m6_97+m7_97+m8_97+m9_97+m10_97+m11_97+m12_97+m13_97+m14_97+m15_97+m16_97+m17_97+m18_97+m19_97+m20_97+m21_97+m22_97+m23_97+m24_97+m25_97+m26_97+m27_97+m28_97+m29_97+m30_97+m31_97+m32_97+m33_97+m34_97+m35_97+m36_97+m37_97+m38_97+m39_97+m40_97+m41_97+m42_97+m43_97+m44_97+m45_97+m46_97+m47_97+m48_97+m49_97+m50_97+m51_97+m52_97+m53_97+m54_97+m55_97+m56_97+m57_97+m58_97+m59_97+m60_97+m61_97+m62_97+m63_97+m64_97+m65_97+m66_97+m67_97+m68_97+m69_97+m70_97+m71_97+m72_97+m73_97+m74_97+m75_97+m76_97+m77_97+m78_97+m79_97+m80_97+m81_97+m82_97+m83_97+m84_97+m85_97+m86_97+m87_97+m88_97+m89_97+m90_97+m91_97+m92_97+m93_97+m94_97+m95_97+m96_97+m97_97+m98_97+m99_97+m100_97+m101_97+m102_97+m103_97+m104_97+m105_97+m106_97+m107_97+m108_97+m109_97+m110_97+m111_97+m112_97+m113_97+m114_97+m115_97+m116_97+m117_97+m118_97+m119_97+m120_97+m121_97+m122_97+m123_97+m124_97+m125_97+m126_97+m127_97+m128_97+m129_97+m130_97+m131_97+m132_97+m133_97+m134_97+m135_97+m136_97+m137_97+m138_97+m139_97+m140_97+m141_97+m142_97+m143_97+m144_97+m145_97+m146_97+m147_97+m148_97+m149_97+m150_97+m151_97+m152_97+m153_97+m154_97+m155_97+m156_97+m157_97+m158_97+m159_97+m160_97+m161_97+m162_97+m163_97+m164_97+m165_97+m166_97+m167_97+m168_97+m169_97+m170_97+m171_97+m172_97+m173_97+m174_97+m175_97+m176_97+m177_97+m178_97+m179_97+m180_97+m181_97+m182_97+m183_97+m184_97+m185_97+m186_97+m187_97+m188_97+m189_97+m190_97+m191_97+m192_97+m193_97+m194_97+m195_97+m196_97+m197_97+m198_97+m199_97+m200_97+m201_97+m202_97+m203_97+m204_97+m205_97+m206_97+m207_97+m208_97+m209_97+m210_97+m211_97+m212_97+m213_97+m214_97+m215_97+m216_97+m217_97+m218_97+m219_97+m220_97+m221_97+m222_97+m223_97+m224_97+m225_97+m226_97+m227_97+m228_97+m229_97+m230_97+m231_97+m232_97+m233_97+m234_97+m235_97+m236_97+m237_97+m238_97+m239_97+m240_97+m241_97+m242_97+m243_97+m244_97+m245_97+m246_97+m247_97+m248_97+m249_97+m250_97+m251_97+m252_97+m253_97+m254_97+m255_97+m256_97+m257_97+m258_97+m259_97+m260_97+m261_97+m262_97+m263_97+m264_97+m265_97+m266_97+m267_97+m268_97+m269_97+m270_97+m271_97+m272_97+m273_97+m274_97+m275_97+m276_97+m277_97+m278_97+m279_97+m280_97+m281_97+m282_97+m283_97+m284_97+m285_97+m286_97+m287_97+m288_97+m289_97+m290_97+m291_97+m292_97+m293_97+m294_97+m295_97+m296_97+m297_97+m298_97+m299_97+m300_97+m301_97+m302_97+m303_97+m304_97+m305_97+m306_97+m307_97+m308_97+m309_97+m310_97+m311_97+m312_97+m313_97+m314_97+m315_97+m316_97+m317_97+m318_97+m319_97+m320_97+m321_97+m322_97+m323_97+m324_97+m325_97+m326_97+m327_97+m328_97+m329_97+m330_97+m331_97+m332_97+m333_97+m334_97+m335_97+m336_97+m337_97+m338_97+m339_97+m340_97+m341_97+m342_97+m343_97+m344_97+m345_97+m346_97+m347_97+m348_97+m349_97+m350_97+m351_97+m352_97+m353_97+m354_97+m355_97+m356_97+m357_97+m358_97+m359_97+m360_97+m361_97+m362_97+m363_97+m364_97+m365_97+m366_97+m367_97+m368_97+m369_97+m370_97+m371_97+m372_97+m373_97+m374_97+m375_97+m376_97+m377_97+m378_97+m379_97+m380_97+m381_97+b97;
   always @(posedge clk) out98 <= m1_98+m2_98+m3_98+m4_98+m5_98+m6_98+m7_98+m8_98+m9_98+m10_98+m11_98+m12_98+m13_98+m14_98+m15_98+m16_98+m17_98+m18_98+m19_98+m20_98+m21_98+m22_98+m23_98+m24_98+m25_98+m26_98+m27_98+m28_98+m29_98+m30_98+m31_98+m32_98+m33_98+m34_98+m35_98+m36_98+m37_98+m38_98+m39_98+m40_98+m41_98+m42_98+m43_98+m44_98+m45_98+m46_98+m47_98+m48_98+m49_98+m50_98+m51_98+m52_98+m53_98+m54_98+m55_98+m56_98+m57_98+m58_98+m59_98+m60_98+m61_98+m62_98+m63_98+m64_98+m65_98+m66_98+m67_98+m68_98+m69_98+m70_98+m71_98+m72_98+m73_98+m74_98+m75_98+m76_98+m77_98+m78_98+m79_98+m80_98+m81_98+m82_98+m83_98+m84_98+m85_98+m86_98+m87_98+m88_98+m89_98+m90_98+m91_98+m92_98+m93_98+m94_98+m95_98+m96_98+m97_98+m98_98+m99_98+m100_98+m101_98+m102_98+m103_98+m104_98+m105_98+m106_98+m107_98+m108_98+m109_98+m110_98+m111_98+m112_98+m113_98+m114_98+m115_98+m116_98+m117_98+m118_98+m119_98+m120_98+m121_98+m122_98+m123_98+m124_98+m125_98+m126_98+m127_98+m128_98+m129_98+m130_98+m131_98+m132_98+m133_98+m134_98+m135_98+m136_98+m137_98+m138_98+m139_98+m140_98+m141_98+m142_98+m143_98+m144_98+m145_98+m146_98+m147_98+m148_98+m149_98+m150_98+m151_98+m152_98+m153_98+m154_98+m155_98+m156_98+m157_98+m158_98+m159_98+m160_98+m161_98+m162_98+m163_98+m164_98+m165_98+m166_98+m167_98+m168_98+m169_98+m170_98+m171_98+m172_98+m173_98+m174_98+m175_98+m176_98+m177_98+m178_98+m179_98+m180_98+m181_98+m182_98+m183_98+m184_98+m185_98+m186_98+m187_98+m188_98+m189_98+m190_98+m191_98+m192_98+m193_98+m194_98+m195_98+m196_98+m197_98+m198_98+m199_98+m200_98+m201_98+m202_98+m203_98+m204_98+m205_98+m206_98+m207_98+m208_98+m209_98+m210_98+m211_98+m212_98+m213_98+m214_98+m215_98+m216_98+m217_98+m218_98+m219_98+m220_98+m221_98+m222_98+m223_98+m224_98+m225_98+m226_98+m227_98+m228_98+m229_98+m230_98+m231_98+m232_98+m233_98+m234_98+m235_98+m236_98+m237_98+m238_98+m239_98+m240_98+m241_98+m242_98+m243_98+m244_98+m245_98+m246_98+m247_98+m248_98+m249_98+m250_98+m251_98+m252_98+m253_98+m254_98+m255_98+m256_98+m257_98+m258_98+m259_98+m260_98+m261_98+m262_98+m263_98+m264_98+m265_98+m266_98+m267_98+m268_98+m269_98+m270_98+m271_98+m272_98+m273_98+m274_98+m275_98+m276_98+m277_98+m278_98+m279_98+m280_98+m281_98+m282_98+m283_98+m284_98+m285_98+m286_98+m287_98+m288_98+m289_98+m290_98+m291_98+m292_98+m293_98+m294_98+m295_98+m296_98+m297_98+m298_98+m299_98+m300_98+m301_98+m302_98+m303_98+m304_98+m305_98+m306_98+m307_98+m308_98+m309_98+m310_98+m311_98+m312_98+m313_98+m314_98+m315_98+m316_98+m317_98+m318_98+m319_98+m320_98+m321_98+m322_98+m323_98+m324_98+m325_98+m326_98+m327_98+m328_98+m329_98+m330_98+m331_98+m332_98+m333_98+m334_98+m335_98+m336_98+m337_98+m338_98+m339_98+m340_98+m341_98+m342_98+m343_98+m344_98+m345_98+m346_98+m347_98+m348_98+m349_98+m350_98+m351_98+m352_98+m353_98+m354_98+m355_98+m356_98+m357_98+m358_98+m359_98+m360_98+m361_98+m362_98+m363_98+m364_98+m365_98+m366_98+m367_98+m368_98+m369_98+m370_98+m371_98+m372_98+m373_98+m374_98+m375_98+m376_98+m377_98+m378_98+m379_98+m380_98+m381_98+b98;
   always @(posedge clk) out99 <= m1_99+m2_99+m3_99+m4_99+m5_99+m6_99+m7_99+m8_99+m9_99+m10_99+m11_99+m12_99+m13_99+m14_99+m15_99+m16_99+m17_99+m18_99+m19_99+m20_99+m21_99+m22_99+m23_99+m24_99+m25_99+m26_99+m27_99+m28_99+m29_99+m30_99+m31_99+m32_99+m33_99+m34_99+m35_99+m36_99+m37_99+m38_99+m39_99+m40_99+m41_99+m42_99+m43_99+m44_99+m45_99+m46_99+m47_99+m48_99+m49_99+m50_99+m51_99+m52_99+m53_99+m54_99+m55_99+m56_99+m57_99+m58_99+m59_99+m60_99+m61_99+m62_99+m63_99+m64_99+m65_99+m66_99+m67_99+m68_99+m69_99+m70_99+m71_99+m72_99+m73_99+m74_99+m75_99+m76_99+m77_99+m78_99+m79_99+m80_99+m81_99+m82_99+m83_99+m84_99+m85_99+m86_99+m87_99+m88_99+m89_99+m90_99+m91_99+m92_99+m93_99+m94_99+m95_99+m96_99+m97_99+m98_99+m99_99+m100_99+m101_99+m102_99+m103_99+m104_99+m105_99+m106_99+m107_99+m108_99+m109_99+m110_99+m111_99+m112_99+m113_99+m114_99+m115_99+m116_99+m117_99+m118_99+m119_99+m120_99+m121_99+m122_99+m123_99+m124_99+m125_99+m126_99+m127_99+m128_99+m129_99+m130_99+m131_99+m132_99+m133_99+m134_99+m135_99+m136_99+m137_99+m138_99+m139_99+m140_99+m141_99+m142_99+m143_99+m144_99+m145_99+m146_99+m147_99+m148_99+m149_99+m150_99+m151_99+m152_99+m153_99+m154_99+m155_99+m156_99+m157_99+m158_99+m159_99+m160_99+m161_99+m162_99+m163_99+m164_99+m165_99+m166_99+m167_99+m168_99+m169_99+m170_99+m171_99+m172_99+m173_99+m174_99+m175_99+m176_99+m177_99+m178_99+m179_99+m180_99+m181_99+m182_99+m183_99+m184_99+m185_99+m186_99+m187_99+m188_99+m189_99+m190_99+m191_99+m192_99+m193_99+m194_99+m195_99+m196_99+m197_99+m198_99+m199_99+m200_99+m201_99+m202_99+m203_99+m204_99+m205_99+m206_99+m207_99+m208_99+m209_99+m210_99+m211_99+m212_99+m213_99+m214_99+m215_99+m216_99+m217_99+m218_99+m219_99+m220_99+m221_99+m222_99+m223_99+m224_99+m225_99+m226_99+m227_99+m228_99+m229_99+m230_99+m231_99+m232_99+m233_99+m234_99+m235_99+m236_99+m237_99+m238_99+m239_99+m240_99+m241_99+m242_99+m243_99+m244_99+m245_99+m246_99+m247_99+m248_99+m249_99+m250_99+m251_99+m252_99+m253_99+m254_99+m255_99+m256_99+m257_99+m258_99+m259_99+m260_99+m261_99+m262_99+m263_99+m264_99+m265_99+m266_99+m267_99+m268_99+m269_99+m270_99+m271_99+m272_99+m273_99+m274_99+m275_99+m276_99+m277_99+m278_99+m279_99+m280_99+m281_99+m282_99+m283_99+m284_99+m285_99+m286_99+m287_99+m288_99+m289_99+m290_99+m291_99+m292_99+m293_99+m294_99+m295_99+m296_99+m297_99+m298_99+m299_99+m300_99+m301_99+m302_99+m303_99+m304_99+m305_99+m306_99+m307_99+m308_99+m309_99+m310_99+m311_99+m312_99+m313_99+m314_99+m315_99+m316_99+m317_99+m318_99+m319_99+m320_99+m321_99+m322_99+m323_99+m324_99+m325_99+m326_99+m327_99+m328_99+m329_99+m330_99+m331_99+m332_99+m333_99+m334_99+m335_99+m336_99+m337_99+m338_99+m339_99+m340_99+m341_99+m342_99+m343_99+m344_99+m345_99+m346_99+m347_99+m348_99+m349_99+m350_99+m351_99+m352_99+m353_99+m354_99+m355_99+m356_99+m357_99+m358_99+m359_99+m360_99+m361_99+m362_99+m363_99+m364_99+m365_99+m366_99+m367_99+m368_99+m369_99+m370_99+m371_99+m372_99+m373_99+m374_99+m375_99+m376_99+m377_99+m378_99+m379_99+m380_99+m381_99+b99;
   always @(posedge clk) out100 <= m1_100+m2_100+m3_100+m4_100+m5_100+m6_100+m7_100+m8_100+m9_100+m10_100+m11_100+m12_100+m13_100+m14_100+m15_100+m16_100+m17_100+m18_100+m19_100+m20_100+m21_100+m22_100+m23_100+m24_100+m25_100+m26_100+m27_100+m28_100+m29_100+m30_100+m31_100+m32_100+m33_100+m34_100+m35_100+m36_100+m37_100+m38_100+m39_100+m40_100+m41_100+m42_100+m43_100+m44_100+m45_100+m46_100+m47_100+m48_100+m49_100+m50_100+m51_100+m52_100+m53_100+m54_100+m55_100+m56_100+m57_100+m58_100+m59_100+m60_100+m61_100+m62_100+m63_100+m64_100+m65_100+m66_100+m67_100+m68_100+m69_100+m70_100+m71_100+m72_100+m73_100+m74_100+m75_100+m76_100+m77_100+m78_100+m79_100+m80_100+m81_100+m82_100+m83_100+m84_100+m85_100+m86_100+m87_100+m88_100+m89_100+m90_100+m91_100+m92_100+m93_100+m94_100+m95_100+m96_100+m97_100+m98_100+m99_100+m100_100+m101_100+m102_100+m103_100+m104_100+m105_100+m106_100+m107_100+m108_100+m109_100+m110_100+m111_100+m112_100+m113_100+m114_100+m115_100+m116_100+m117_100+m118_100+m119_100+m120_100+m121_100+m122_100+m123_100+m124_100+m125_100+m126_100+m127_100+m128_100+m129_100+m130_100+m131_100+m132_100+m133_100+m134_100+m135_100+m136_100+m137_100+m138_100+m139_100+m140_100+m141_100+m142_100+m143_100+m144_100+m145_100+m146_100+m147_100+m148_100+m149_100+m150_100+m151_100+m152_100+m153_100+m154_100+m155_100+m156_100+m157_100+m158_100+m159_100+m160_100+m161_100+m162_100+m163_100+m164_100+m165_100+m166_100+m167_100+m168_100+m169_100+m170_100+m171_100+m172_100+m173_100+m174_100+m175_100+m176_100+m177_100+m178_100+m179_100+m180_100+m181_100+m182_100+m183_100+m184_100+m185_100+m186_100+m187_100+m188_100+m189_100+m190_100+m191_100+m192_100+m193_100+m194_100+m195_100+m196_100+m197_100+m198_100+m199_100+m200_100+m201_100+m202_100+m203_100+m204_100+m205_100+m206_100+m207_100+m208_100+m209_100+m210_100+m211_100+m212_100+m213_100+m214_100+m215_100+m216_100+m217_100+m218_100+m219_100+m220_100+m221_100+m222_100+m223_100+m224_100+m225_100+m226_100+m227_100+m228_100+m229_100+m230_100+m231_100+m232_100+m233_100+m234_100+m235_100+m236_100+m237_100+m238_100+m239_100+m240_100+m241_100+m242_100+m243_100+m244_100+m245_100+m246_100+m247_100+m248_100+m249_100+m250_100+m251_100+m252_100+m253_100+m254_100+m255_100+m256_100+m257_100+m258_100+m259_100+m260_100+m261_100+m262_100+m263_100+m264_100+m265_100+m266_100+m267_100+m268_100+m269_100+m270_100+m271_100+m272_100+m273_100+m274_100+m275_100+m276_100+m277_100+m278_100+m279_100+m280_100+m281_100+m282_100+m283_100+m284_100+m285_100+m286_100+m287_100+m288_100+m289_100+m290_100+m291_100+m292_100+m293_100+m294_100+m295_100+m296_100+m297_100+m298_100+m299_100+m300_100+m301_100+m302_100+m303_100+m304_100+m305_100+m306_100+m307_100+m308_100+m309_100+m310_100+m311_100+m312_100+m313_100+m314_100+m315_100+m316_100+m317_100+m318_100+m319_100+m320_100+m321_100+m322_100+m323_100+m324_100+m325_100+m326_100+m327_100+m328_100+m329_100+m330_100+m331_100+m332_100+m333_100+m334_100+m335_100+m336_100+m337_100+m338_100+m339_100+m340_100+m341_100+m342_100+m343_100+m344_100+m345_100+m346_100+m347_100+m348_100+m349_100+m350_100+m351_100+m352_100+m353_100+m354_100+m355_100+m356_100+m357_100+m358_100+m359_100+m360_100+m361_100+m362_100+m363_100+m364_100+m365_100+m366_100+m367_100+m368_100+m369_100+m370_100+m371_100+m372_100+m373_100+m374_100+m375_100+m376_100+m377_100+m378_100+m379_100+m380_100+m381_100+b100;
   always @(posedge clk) out101 <= m1_101+m2_101+m3_101+m4_101+m5_101+m6_101+m7_101+m8_101+m9_101+m10_101+m11_101+m12_101+m13_101+m14_101+m15_101+m16_101+m17_101+m18_101+m19_101+m20_101+m21_101+m22_101+m23_101+m24_101+m25_101+m26_101+m27_101+m28_101+m29_101+m30_101+m31_101+m32_101+m33_101+m34_101+m35_101+m36_101+m37_101+m38_101+m39_101+m40_101+m41_101+m42_101+m43_101+m44_101+m45_101+m46_101+m47_101+m48_101+m49_101+m50_101+m51_101+m52_101+m53_101+m54_101+m55_101+m56_101+m57_101+m58_101+m59_101+m60_101+m61_101+m62_101+m63_101+m64_101+m65_101+m66_101+m67_101+m68_101+m69_101+m70_101+m71_101+m72_101+m73_101+m74_101+m75_101+m76_101+m77_101+m78_101+m79_101+m80_101+m81_101+m82_101+m83_101+m84_101+m85_101+m86_101+m87_101+m88_101+m89_101+m90_101+m91_101+m92_101+m93_101+m94_101+m95_101+m96_101+m97_101+m98_101+m99_101+m100_101+m101_101+m102_101+m103_101+m104_101+m105_101+m106_101+m107_101+m108_101+m109_101+m110_101+m111_101+m112_101+m113_101+m114_101+m115_101+m116_101+m117_101+m118_101+m119_101+m120_101+m121_101+m122_101+m123_101+m124_101+m125_101+m126_101+m127_101+m128_101+m129_101+m130_101+m131_101+m132_101+m133_101+m134_101+m135_101+m136_101+m137_101+m138_101+m139_101+m140_101+m141_101+m142_101+m143_101+m144_101+m145_101+m146_101+m147_101+m148_101+m149_101+m150_101+m151_101+m152_101+m153_101+m154_101+m155_101+m156_101+m157_101+m158_101+m159_101+m160_101+m161_101+m162_101+m163_101+m164_101+m165_101+m166_101+m167_101+m168_101+m169_101+m170_101+m171_101+m172_101+m173_101+m174_101+m175_101+m176_101+m177_101+m178_101+m179_101+m180_101+m181_101+m182_101+m183_101+m184_101+m185_101+m186_101+m187_101+m188_101+m189_101+m190_101+m191_101+m192_101+m193_101+m194_101+m195_101+m196_101+m197_101+m198_101+m199_101+m200_101+m201_101+m202_101+m203_101+m204_101+m205_101+m206_101+m207_101+m208_101+m209_101+m210_101+m211_101+m212_101+m213_101+m214_101+m215_101+m216_101+m217_101+m218_101+m219_101+m220_101+m221_101+m222_101+m223_101+m224_101+m225_101+m226_101+m227_101+m228_101+m229_101+m230_101+m231_101+m232_101+m233_101+m234_101+m235_101+m236_101+m237_101+m238_101+m239_101+m240_101+m241_101+m242_101+m243_101+m244_101+m245_101+m246_101+m247_101+m248_101+m249_101+m250_101+m251_101+m252_101+m253_101+m254_101+m255_101+m256_101+m257_101+m258_101+m259_101+m260_101+m261_101+m262_101+m263_101+m264_101+m265_101+m266_101+m267_101+m268_101+m269_101+m270_101+m271_101+m272_101+m273_101+m274_101+m275_101+m276_101+m277_101+m278_101+m279_101+m280_101+m281_101+m282_101+m283_101+m284_101+m285_101+m286_101+m287_101+m288_101+m289_101+m290_101+m291_101+m292_101+m293_101+m294_101+m295_101+m296_101+m297_101+m298_101+m299_101+m300_101+m301_101+m302_101+m303_101+m304_101+m305_101+m306_101+m307_101+m308_101+m309_101+m310_101+m311_101+m312_101+m313_101+m314_101+m315_101+m316_101+m317_101+m318_101+m319_101+m320_101+m321_101+m322_101+m323_101+m324_101+m325_101+m326_101+m327_101+m328_101+m329_101+m330_101+m331_101+m332_101+m333_101+m334_101+m335_101+m336_101+m337_101+m338_101+m339_101+m340_101+m341_101+m342_101+m343_101+m344_101+m345_101+m346_101+m347_101+m348_101+m349_101+m350_101+m351_101+m352_101+m353_101+m354_101+m355_101+m356_101+m357_101+m358_101+m359_101+m360_101+m361_101+m362_101+m363_101+m364_101+m365_101+m366_101+m367_101+m368_101+m369_101+m370_101+m371_101+m372_101+m373_101+m374_101+m375_101+m376_101+m377_101+m378_101+m379_101+m380_101+m381_101+b101;
   always @(posedge clk) out102 <= m1_102+m2_102+m3_102+m4_102+m5_102+m6_102+m7_102+m8_102+m9_102+m10_102+m11_102+m12_102+m13_102+m14_102+m15_102+m16_102+m17_102+m18_102+m19_102+m20_102+m21_102+m22_102+m23_102+m24_102+m25_102+m26_102+m27_102+m28_102+m29_102+m30_102+m31_102+m32_102+m33_102+m34_102+m35_102+m36_102+m37_102+m38_102+m39_102+m40_102+m41_102+m42_102+m43_102+m44_102+m45_102+m46_102+m47_102+m48_102+m49_102+m50_102+m51_102+m52_102+m53_102+m54_102+m55_102+m56_102+m57_102+m58_102+m59_102+m60_102+m61_102+m62_102+m63_102+m64_102+m65_102+m66_102+m67_102+m68_102+m69_102+m70_102+m71_102+m72_102+m73_102+m74_102+m75_102+m76_102+m77_102+m78_102+m79_102+m80_102+m81_102+m82_102+m83_102+m84_102+m85_102+m86_102+m87_102+m88_102+m89_102+m90_102+m91_102+m92_102+m93_102+m94_102+m95_102+m96_102+m97_102+m98_102+m99_102+m100_102+m101_102+m102_102+m103_102+m104_102+m105_102+m106_102+m107_102+m108_102+m109_102+m110_102+m111_102+m112_102+m113_102+m114_102+m115_102+m116_102+m117_102+m118_102+m119_102+m120_102+m121_102+m122_102+m123_102+m124_102+m125_102+m126_102+m127_102+m128_102+m129_102+m130_102+m131_102+m132_102+m133_102+m134_102+m135_102+m136_102+m137_102+m138_102+m139_102+m140_102+m141_102+m142_102+m143_102+m144_102+m145_102+m146_102+m147_102+m148_102+m149_102+m150_102+m151_102+m152_102+m153_102+m154_102+m155_102+m156_102+m157_102+m158_102+m159_102+m160_102+m161_102+m162_102+m163_102+m164_102+m165_102+m166_102+m167_102+m168_102+m169_102+m170_102+m171_102+m172_102+m173_102+m174_102+m175_102+m176_102+m177_102+m178_102+m179_102+m180_102+m181_102+m182_102+m183_102+m184_102+m185_102+m186_102+m187_102+m188_102+m189_102+m190_102+m191_102+m192_102+m193_102+m194_102+m195_102+m196_102+m197_102+m198_102+m199_102+m200_102+m201_102+m202_102+m203_102+m204_102+m205_102+m206_102+m207_102+m208_102+m209_102+m210_102+m211_102+m212_102+m213_102+m214_102+m215_102+m216_102+m217_102+m218_102+m219_102+m220_102+m221_102+m222_102+m223_102+m224_102+m225_102+m226_102+m227_102+m228_102+m229_102+m230_102+m231_102+m232_102+m233_102+m234_102+m235_102+m236_102+m237_102+m238_102+m239_102+m240_102+m241_102+m242_102+m243_102+m244_102+m245_102+m246_102+m247_102+m248_102+m249_102+m250_102+m251_102+m252_102+m253_102+m254_102+m255_102+m256_102+m257_102+m258_102+m259_102+m260_102+m261_102+m262_102+m263_102+m264_102+m265_102+m266_102+m267_102+m268_102+m269_102+m270_102+m271_102+m272_102+m273_102+m274_102+m275_102+m276_102+m277_102+m278_102+m279_102+m280_102+m281_102+m282_102+m283_102+m284_102+m285_102+m286_102+m287_102+m288_102+m289_102+m290_102+m291_102+m292_102+m293_102+m294_102+m295_102+m296_102+m297_102+m298_102+m299_102+m300_102+m301_102+m302_102+m303_102+m304_102+m305_102+m306_102+m307_102+m308_102+m309_102+m310_102+m311_102+m312_102+m313_102+m314_102+m315_102+m316_102+m317_102+m318_102+m319_102+m320_102+m321_102+m322_102+m323_102+m324_102+m325_102+m326_102+m327_102+m328_102+m329_102+m330_102+m331_102+m332_102+m333_102+m334_102+m335_102+m336_102+m337_102+m338_102+m339_102+m340_102+m341_102+m342_102+m343_102+m344_102+m345_102+m346_102+m347_102+m348_102+m349_102+m350_102+m351_102+m352_102+m353_102+m354_102+m355_102+m356_102+m357_102+m358_102+m359_102+m360_102+m361_102+m362_102+m363_102+m364_102+m365_102+m366_102+m367_102+m368_102+m369_102+m370_102+m371_102+m372_102+m373_102+m374_102+m375_102+m376_102+m377_102+m378_102+m379_102+m380_102+m381_102+b102;
   always @(posedge clk) out103 <= m1_103+m2_103+m3_103+m4_103+m5_103+m6_103+m7_103+m8_103+m9_103+m10_103+m11_103+m12_103+m13_103+m14_103+m15_103+m16_103+m17_103+m18_103+m19_103+m20_103+m21_103+m22_103+m23_103+m24_103+m25_103+m26_103+m27_103+m28_103+m29_103+m30_103+m31_103+m32_103+m33_103+m34_103+m35_103+m36_103+m37_103+m38_103+m39_103+m40_103+m41_103+m42_103+m43_103+m44_103+m45_103+m46_103+m47_103+m48_103+m49_103+m50_103+m51_103+m52_103+m53_103+m54_103+m55_103+m56_103+m57_103+m58_103+m59_103+m60_103+m61_103+m62_103+m63_103+m64_103+m65_103+m66_103+m67_103+m68_103+m69_103+m70_103+m71_103+m72_103+m73_103+m74_103+m75_103+m76_103+m77_103+m78_103+m79_103+m80_103+m81_103+m82_103+m83_103+m84_103+m85_103+m86_103+m87_103+m88_103+m89_103+m90_103+m91_103+m92_103+m93_103+m94_103+m95_103+m96_103+m97_103+m98_103+m99_103+m100_103+m101_103+m102_103+m103_103+m104_103+m105_103+m106_103+m107_103+m108_103+m109_103+m110_103+m111_103+m112_103+m113_103+m114_103+m115_103+m116_103+m117_103+m118_103+m119_103+m120_103+m121_103+m122_103+m123_103+m124_103+m125_103+m126_103+m127_103+m128_103+m129_103+m130_103+m131_103+m132_103+m133_103+m134_103+m135_103+m136_103+m137_103+m138_103+m139_103+m140_103+m141_103+m142_103+m143_103+m144_103+m145_103+m146_103+m147_103+m148_103+m149_103+m150_103+m151_103+m152_103+m153_103+m154_103+m155_103+m156_103+m157_103+m158_103+m159_103+m160_103+m161_103+m162_103+m163_103+m164_103+m165_103+m166_103+m167_103+m168_103+m169_103+m170_103+m171_103+m172_103+m173_103+m174_103+m175_103+m176_103+m177_103+m178_103+m179_103+m180_103+m181_103+m182_103+m183_103+m184_103+m185_103+m186_103+m187_103+m188_103+m189_103+m190_103+m191_103+m192_103+m193_103+m194_103+m195_103+m196_103+m197_103+m198_103+m199_103+m200_103+m201_103+m202_103+m203_103+m204_103+m205_103+m206_103+m207_103+m208_103+m209_103+m210_103+m211_103+m212_103+m213_103+m214_103+m215_103+m216_103+m217_103+m218_103+m219_103+m220_103+m221_103+m222_103+m223_103+m224_103+m225_103+m226_103+m227_103+m228_103+m229_103+m230_103+m231_103+m232_103+m233_103+m234_103+m235_103+m236_103+m237_103+m238_103+m239_103+m240_103+m241_103+m242_103+m243_103+m244_103+m245_103+m246_103+m247_103+m248_103+m249_103+m250_103+m251_103+m252_103+m253_103+m254_103+m255_103+m256_103+m257_103+m258_103+m259_103+m260_103+m261_103+m262_103+m263_103+m264_103+m265_103+m266_103+m267_103+m268_103+m269_103+m270_103+m271_103+m272_103+m273_103+m274_103+m275_103+m276_103+m277_103+m278_103+m279_103+m280_103+m281_103+m282_103+m283_103+m284_103+m285_103+m286_103+m287_103+m288_103+m289_103+m290_103+m291_103+m292_103+m293_103+m294_103+m295_103+m296_103+m297_103+m298_103+m299_103+m300_103+m301_103+m302_103+m303_103+m304_103+m305_103+m306_103+m307_103+m308_103+m309_103+m310_103+m311_103+m312_103+m313_103+m314_103+m315_103+m316_103+m317_103+m318_103+m319_103+m320_103+m321_103+m322_103+m323_103+m324_103+m325_103+m326_103+m327_103+m328_103+m329_103+m330_103+m331_103+m332_103+m333_103+m334_103+m335_103+m336_103+m337_103+m338_103+m339_103+m340_103+m341_103+m342_103+m343_103+m344_103+m345_103+m346_103+m347_103+m348_103+m349_103+m350_103+m351_103+m352_103+m353_103+m354_103+m355_103+m356_103+m357_103+m358_103+m359_103+m360_103+m361_103+m362_103+m363_103+m364_103+m365_103+m366_103+m367_103+m368_103+m369_103+m370_103+m371_103+m372_103+m373_103+m374_103+m375_103+m376_103+m377_103+m378_103+m379_103+m380_103+m381_103+b103;
   always @(posedge clk) out104 <= m1_104+m2_104+m3_104+m4_104+m5_104+m6_104+m7_104+m8_104+m9_104+m10_104+m11_104+m12_104+m13_104+m14_104+m15_104+m16_104+m17_104+m18_104+m19_104+m20_104+m21_104+m22_104+m23_104+m24_104+m25_104+m26_104+m27_104+m28_104+m29_104+m30_104+m31_104+m32_104+m33_104+m34_104+m35_104+m36_104+m37_104+m38_104+m39_104+m40_104+m41_104+m42_104+m43_104+m44_104+m45_104+m46_104+m47_104+m48_104+m49_104+m50_104+m51_104+m52_104+m53_104+m54_104+m55_104+m56_104+m57_104+m58_104+m59_104+m60_104+m61_104+m62_104+m63_104+m64_104+m65_104+m66_104+m67_104+m68_104+m69_104+m70_104+m71_104+m72_104+m73_104+m74_104+m75_104+m76_104+m77_104+m78_104+m79_104+m80_104+m81_104+m82_104+m83_104+m84_104+m85_104+m86_104+m87_104+m88_104+m89_104+m90_104+m91_104+m92_104+m93_104+m94_104+m95_104+m96_104+m97_104+m98_104+m99_104+m100_104+m101_104+m102_104+m103_104+m104_104+m105_104+m106_104+m107_104+m108_104+m109_104+m110_104+m111_104+m112_104+m113_104+m114_104+m115_104+m116_104+m117_104+m118_104+m119_104+m120_104+m121_104+m122_104+m123_104+m124_104+m125_104+m126_104+m127_104+m128_104+m129_104+m130_104+m131_104+m132_104+m133_104+m134_104+m135_104+m136_104+m137_104+m138_104+m139_104+m140_104+m141_104+m142_104+m143_104+m144_104+m145_104+m146_104+m147_104+m148_104+m149_104+m150_104+m151_104+m152_104+m153_104+m154_104+m155_104+m156_104+m157_104+m158_104+m159_104+m160_104+m161_104+m162_104+m163_104+m164_104+m165_104+m166_104+m167_104+m168_104+m169_104+m170_104+m171_104+m172_104+m173_104+m174_104+m175_104+m176_104+m177_104+m178_104+m179_104+m180_104+m181_104+m182_104+m183_104+m184_104+m185_104+m186_104+m187_104+m188_104+m189_104+m190_104+m191_104+m192_104+m193_104+m194_104+m195_104+m196_104+m197_104+m198_104+m199_104+m200_104+m201_104+m202_104+m203_104+m204_104+m205_104+m206_104+m207_104+m208_104+m209_104+m210_104+m211_104+m212_104+m213_104+m214_104+m215_104+m216_104+m217_104+m218_104+m219_104+m220_104+m221_104+m222_104+m223_104+m224_104+m225_104+m226_104+m227_104+m228_104+m229_104+m230_104+m231_104+m232_104+m233_104+m234_104+m235_104+m236_104+m237_104+m238_104+m239_104+m240_104+m241_104+m242_104+m243_104+m244_104+m245_104+m246_104+m247_104+m248_104+m249_104+m250_104+m251_104+m252_104+m253_104+m254_104+m255_104+m256_104+m257_104+m258_104+m259_104+m260_104+m261_104+m262_104+m263_104+m264_104+m265_104+m266_104+m267_104+m268_104+m269_104+m270_104+m271_104+m272_104+m273_104+m274_104+m275_104+m276_104+m277_104+m278_104+m279_104+m280_104+m281_104+m282_104+m283_104+m284_104+m285_104+m286_104+m287_104+m288_104+m289_104+m290_104+m291_104+m292_104+m293_104+m294_104+m295_104+m296_104+m297_104+m298_104+m299_104+m300_104+m301_104+m302_104+m303_104+m304_104+m305_104+m306_104+m307_104+m308_104+m309_104+m310_104+m311_104+m312_104+m313_104+m314_104+m315_104+m316_104+m317_104+m318_104+m319_104+m320_104+m321_104+m322_104+m323_104+m324_104+m325_104+m326_104+m327_104+m328_104+m329_104+m330_104+m331_104+m332_104+m333_104+m334_104+m335_104+m336_104+m337_104+m338_104+m339_104+m340_104+m341_104+m342_104+m343_104+m344_104+m345_104+m346_104+m347_104+m348_104+m349_104+m350_104+m351_104+m352_104+m353_104+m354_104+m355_104+m356_104+m357_104+m358_104+m359_104+m360_104+m361_104+m362_104+m363_104+m364_104+m365_104+m366_104+m367_104+m368_104+m369_104+m370_104+m371_104+m372_104+m373_104+m374_104+m375_104+m376_104+m377_104+m378_104+m379_104+m380_104+m381_104+b104;
   always @(posedge clk) out105 <= m1_105+m2_105+m3_105+m4_105+m5_105+m6_105+m7_105+m8_105+m9_105+m10_105+m11_105+m12_105+m13_105+m14_105+m15_105+m16_105+m17_105+m18_105+m19_105+m20_105+m21_105+m22_105+m23_105+m24_105+m25_105+m26_105+m27_105+m28_105+m29_105+m30_105+m31_105+m32_105+m33_105+m34_105+m35_105+m36_105+m37_105+m38_105+m39_105+m40_105+m41_105+m42_105+m43_105+m44_105+m45_105+m46_105+m47_105+m48_105+m49_105+m50_105+m51_105+m52_105+m53_105+m54_105+m55_105+m56_105+m57_105+m58_105+m59_105+m60_105+m61_105+m62_105+m63_105+m64_105+m65_105+m66_105+m67_105+m68_105+m69_105+m70_105+m71_105+m72_105+m73_105+m74_105+m75_105+m76_105+m77_105+m78_105+m79_105+m80_105+m81_105+m82_105+m83_105+m84_105+m85_105+m86_105+m87_105+m88_105+m89_105+m90_105+m91_105+m92_105+m93_105+m94_105+m95_105+m96_105+m97_105+m98_105+m99_105+m100_105+m101_105+m102_105+m103_105+m104_105+m105_105+m106_105+m107_105+m108_105+m109_105+m110_105+m111_105+m112_105+m113_105+m114_105+m115_105+m116_105+m117_105+m118_105+m119_105+m120_105+m121_105+m122_105+m123_105+m124_105+m125_105+m126_105+m127_105+m128_105+m129_105+m130_105+m131_105+m132_105+m133_105+m134_105+m135_105+m136_105+m137_105+m138_105+m139_105+m140_105+m141_105+m142_105+m143_105+m144_105+m145_105+m146_105+m147_105+m148_105+m149_105+m150_105+m151_105+m152_105+m153_105+m154_105+m155_105+m156_105+m157_105+m158_105+m159_105+m160_105+m161_105+m162_105+m163_105+m164_105+m165_105+m166_105+m167_105+m168_105+m169_105+m170_105+m171_105+m172_105+m173_105+m174_105+m175_105+m176_105+m177_105+m178_105+m179_105+m180_105+m181_105+m182_105+m183_105+m184_105+m185_105+m186_105+m187_105+m188_105+m189_105+m190_105+m191_105+m192_105+m193_105+m194_105+m195_105+m196_105+m197_105+m198_105+m199_105+m200_105+m201_105+m202_105+m203_105+m204_105+m205_105+m206_105+m207_105+m208_105+m209_105+m210_105+m211_105+m212_105+m213_105+m214_105+m215_105+m216_105+m217_105+m218_105+m219_105+m220_105+m221_105+m222_105+m223_105+m224_105+m225_105+m226_105+m227_105+m228_105+m229_105+m230_105+m231_105+m232_105+m233_105+m234_105+m235_105+m236_105+m237_105+m238_105+m239_105+m240_105+m241_105+m242_105+m243_105+m244_105+m245_105+m246_105+m247_105+m248_105+m249_105+m250_105+m251_105+m252_105+m253_105+m254_105+m255_105+m256_105+m257_105+m258_105+m259_105+m260_105+m261_105+m262_105+m263_105+m264_105+m265_105+m266_105+m267_105+m268_105+m269_105+m270_105+m271_105+m272_105+m273_105+m274_105+m275_105+m276_105+m277_105+m278_105+m279_105+m280_105+m281_105+m282_105+m283_105+m284_105+m285_105+m286_105+m287_105+m288_105+m289_105+m290_105+m291_105+m292_105+m293_105+m294_105+m295_105+m296_105+m297_105+m298_105+m299_105+m300_105+m301_105+m302_105+m303_105+m304_105+m305_105+m306_105+m307_105+m308_105+m309_105+m310_105+m311_105+m312_105+m313_105+m314_105+m315_105+m316_105+m317_105+m318_105+m319_105+m320_105+m321_105+m322_105+m323_105+m324_105+m325_105+m326_105+m327_105+m328_105+m329_105+m330_105+m331_105+m332_105+m333_105+m334_105+m335_105+m336_105+m337_105+m338_105+m339_105+m340_105+m341_105+m342_105+m343_105+m344_105+m345_105+m346_105+m347_105+m348_105+m349_105+m350_105+m351_105+m352_105+m353_105+m354_105+m355_105+m356_105+m357_105+m358_105+m359_105+m360_105+m361_105+m362_105+m363_105+m364_105+m365_105+m366_105+m367_105+m368_105+m369_105+m370_105+m371_105+m372_105+m373_105+m374_105+m375_105+m376_105+m377_105+m378_105+m379_105+m380_105+m381_105+b105;
   always @(posedge clk) out106 <= m1_106+m2_106+m3_106+m4_106+m5_106+m6_106+m7_106+m8_106+m9_106+m10_106+m11_106+m12_106+m13_106+m14_106+m15_106+m16_106+m17_106+m18_106+m19_106+m20_106+m21_106+m22_106+m23_106+m24_106+m25_106+m26_106+m27_106+m28_106+m29_106+m30_106+m31_106+m32_106+m33_106+m34_106+m35_106+m36_106+m37_106+m38_106+m39_106+m40_106+m41_106+m42_106+m43_106+m44_106+m45_106+m46_106+m47_106+m48_106+m49_106+m50_106+m51_106+m52_106+m53_106+m54_106+m55_106+m56_106+m57_106+m58_106+m59_106+m60_106+m61_106+m62_106+m63_106+m64_106+m65_106+m66_106+m67_106+m68_106+m69_106+m70_106+m71_106+m72_106+m73_106+m74_106+m75_106+m76_106+m77_106+m78_106+m79_106+m80_106+m81_106+m82_106+m83_106+m84_106+m85_106+m86_106+m87_106+m88_106+m89_106+m90_106+m91_106+m92_106+m93_106+m94_106+m95_106+m96_106+m97_106+m98_106+m99_106+m100_106+m101_106+m102_106+m103_106+m104_106+m105_106+m106_106+m107_106+m108_106+m109_106+m110_106+m111_106+m112_106+m113_106+m114_106+m115_106+m116_106+m117_106+m118_106+m119_106+m120_106+m121_106+m122_106+m123_106+m124_106+m125_106+m126_106+m127_106+m128_106+m129_106+m130_106+m131_106+m132_106+m133_106+m134_106+m135_106+m136_106+m137_106+m138_106+m139_106+m140_106+m141_106+m142_106+m143_106+m144_106+m145_106+m146_106+m147_106+m148_106+m149_106+m150_106+m151_106+m152_106+m153_106+m154_106+m155_106+m156_106+m157_106+m158_106+m159_106+m160_106+m161_106+m162_106+m163_106+m164_106+m165_106+m166_106+m167_106+m168_106+m169_106+m170_106+m171_106+m172_106+m173_106+m174_106+m175_106+m176_106+m177_106+m178_106+m179_106+m180_106+m181_106+m182_106+m183_106+m184_106+m185_106+m186_106+m187_106+m188_106+m189_106+m190_106+m191_106+m192_106+m193_106+m194_106+m195_106+m196_106+m197_106+m198_106+m199_106+m200_106+m201_106+m202_106+m203_106+m204_106+m205_106+m206_106+m207_106+m208_106+m209_106+m210_106+m211_106+m212_106+m213_106+m214_106+m215_106+m216_106+m217_106+m218_106+m219_106+m220_106+m221_106+m222_106+m223_106+m224_106+m225_106+m226_106+m227_106+m228_106+m229_106+m230_106+m231_106+m232_106+m233_106+m234_106+m235_106+m236_106+m237_106+m238_106+m239_106+m240_106+m241_106+m242_106+m243_106+m244_106+m245_106+m246_106+m247_106+m248_106+m249_106+m250_106+m251_106+m252_106+m253_106+m254_106+m255_106+m256_106+m257_106+m258_106+m259_106+m260_106+m261_106+m262_106+m263_106+m264_106+m265_106+m266_106+m267_106+m268_106+m269_106+m270_106+m271_106+m272_106+m273_106+m274_106+m275_106+m276_106+m277_106+m278_106+m279_106+m280_106+m281_106+m282_106+m283_106+m284_106+m285_106+m286_106+m287_106+m288_106+m289_106+m290_106+m291_106+m292_106+m293_106+m294_106+m295_106+m296_106+m297_106+m298_106+m299_106+m300_106+m301_106+m302_106+m303_106+m304_106+m305_106+m306_106+m307_106+m308_106+m309_106+m310_106+m311_106+m312_106+m313_106+m314_106+m315_106+m316_106+m317_106+m318_106+m319_106+m320_106+m321_106+m322_106+m323_106+m324_106+m325_106+m326_106+m327_106+m328_106+m329_106+m330_106+m331_106+m332_106+m333_106+m334_106+m335_106+m336_106+m337_106+m338_106+m339_106+m340_106+m341_106+m342_106+m343_106+m344_106+m345_106+m346_106+m347_106+m348_106+m349_106+m350_106+m351_106+m352_106+m353_106+m354_106+m355_106+m356_106+m357_106+m358_106+m359_106+m360_106+m361_106+m362_106+m363_106+m364_106+m365_106+m366_106+m367_106+m368_106+m369_106+m370_106+m371_106+m372_106+m373_106+m374_106+m375_106+m376_106+m377_106+m378_106+m379_106+m380_106+m381_106+b106;
   always @(posedge clk) out107 <= m1_107+m2_107+m3_107+m4_107+m5_107+m6_107+m7_107+m8_107+m9_107+m10_107+m11_107+m12_107+m13_107+m14_107+m15_107+m16_107+m17_107+m18_107+m19_107+m20_107+m21_107+m22_107+m23_107+m24_107+m25_107+m26_107+m27_107+m28_107+m29_107+m30_107+m31_107+m32_107+m33_107+m34_107+m35_107+m36_107+m37_107+m38_107+m39_107+m40_107+m41_107+m42_107+m43_107+m44_107+m45_107+m46_107+m47_107+m48_107+m49_107+m50_107+m51_107+m52_107+m53_107+m54_107+m55_107+m56_107+m57_107+m58_107+m59_107+m60_107+m61_107+m62_107+m63_107+m64_107+m65_107+m66_107+m67_107+m68_107+m69_107+m70_107+m71_107+m72_107+m73_107+m74_107+m75_107+m76_107+m77_107+m78_107+m79_107+m80_107+m81_107+m82_107+m83_107+m84_107+m85_107+m86_107+m87_107+m88_107+m89_107+m90_107+m91_107+m92_107+m93_107+m94_107+m95_107+m96_107+m97_107+m98_107+m99_107+m100_107+m101_107+m102_107+m103_107+m104_107+m105_107+m106_107+m107_107+m108_107+m109_107+m110_107+m111_107+m112_107+m113_107+m114_107+m115_107+m116_107+m117_107+m118_107+m119_107+m120_107+m121_107+m122_107+m123_107+m124_107+m125_107+m126_107+m127_107+m128_107+m129_107+m130_107+m131_107+m132_107+m133_107+m134_107+m135_107+m136_107+m137_107+m138_107+m139_107+m140_107+m141_107+m142_107+m143_107+m144_107+m145_107+m146_107+m147_107+m148_107+m149_107+m150_107+m151_107+m152_107+m153_107+m154_107+m155_107+m156_107+m157_107+m158_107+m159_107+m160_107+m161_107+m162_107+m163_107+m164_107+m165_107+m166_107+m167_107+m168_107+m169_107+m170_107+m171_107+m172_107+m173_107+m174_107+m175_107+m176_107+m177_107+m178_107+m179_107+m180_107+m181_107+m182_107+m183_107+m184_107+m185_107+m186_107+m187_107+m188_107+m189_107+m190_107+m191_107+m192_107+m193_107+m194_107+m195_107+m196_107+m197_107+m198_107+m199_107+m200_107+m201_107+m202_107+m203_107+m204_107+m205_107+m206_107+m207_107+m208_107+m209_107+m210_107+m211_107+m212_107+m213_107+m214_107+m215_107+m216_107+m217_107+m218_107+m219_107+m220_107+m221_107+m222_107+m223_107+m224_107+m225_107+m226_107+m227_107+m228_107+m229_107+m230_107+m231_107+m232_107+m233_107+m234_107+m235_107+m236_107+m237_107+m238_107+m239_107+m240_107+m241_107+m242_107+m243_107+m244_107+m245_107+m246_107+m247_107+m248_107+m249_107+m250_107+m251_107+m252_107+m253_107+m254_107+m255_107+m256_107+m257_107+m258_107+m259_107+m260_107+m261_107+m262_107+m263_107+m264_107+m265_107+m266_107+m267_107+m268_107+m269_107+m270_107+m271_107+m272_107+m273_107+m274_107+m275_107+m276_107+m277_107+m278_107+m279_107+m280_107+m281_107+m282_107+m283_107+m284_107+m285_107+m286_107+m287_107+m288_107+m289_107+m290_107+m291_107+m292_107+m293_107+m294_107+m295_107+m296_107+m297_107+m298_107+m299_107+m300_107+m301_107+m302_107+m303_107+m304_107+m305_107+m306_107+m307_107+m308_107+m309_107+m310_107+m311_107+m312_107+m313_107+m314_107+m315_107+m316_107+m317_107+m318_107+m319_107+m320_107+m321_107+m322_107+m323_107+m324_107+m325_107+m326_107+m327_107+m328_107+m329_107+m330_107+m331_107+m332_107+m333_107+m334_107+m335_107+m336_107+m337_107+m338_107+m339_107+m340_107+m341_107+m342_107+m343_107+m344_107+m345_107+m346_107+m347_107+m348_107+m349_107+m350_107+m351_107+m352_107+m353_107+m354_107+m355_107+m356_107+m357_107+m358_107+m359_107+m360_107+m361_107+m362_107+m363_107+m364_107+m365_107+m366_107+m367_107+m368_107+m369_107+m370_107+m371_107+m372_107+m373_107+m374_107+m375_107+m376_107+m377_107+m378_107+m379_107+m380_107+m381_107+b107;
   always @(posedge clk) out108 <= m1_108+m2_108+m3_108+m4_108+m5_108+m6_108+m7_108+m8_108+m9_108+m10_108+m11_108+m12_108+m13_108+m14_108+m15_108+m16_108+m17_108+m18_108+m19_108+m20_108+m21_108+m22_108+m23_108+m24_108+m25_108+m26_108+m27_108+m28_108+m29_108+m30_108+m31_108+m32_108+m33_108+m34_108+m35_108+m36_108+m37_108+m38_108+m39_108+m40_108+m41_108+m42_108+m43_108+m44_108+m45_108+m46_108+m47_108+m48_108+m49_108+m50_108+m51_108+m52_108+m53_108+m54_108+m55_108+m56_108+m57_108+m58_108+m59_108+m60_108+m61_108+m62_108+m63_108+m64_108+m65_108+m66_108+m67_108+m68_108+m69_108+m70_108+m71_108+m72_108+m73_108+m74_108+m75_108+m76_108+m77_108+m78_108+m79_108+m80_108+m81_108+m82_108+m83_108+m84_108+m85_108+m86_108+m87_108+m88_108+m89_108+m90_108+m91_108+m92_108+m93_108+m94_108+m95_108+m96_108+m97_108+m98_108+m99_108+m100_108+m101_108+m102_108+m103_108+m104_108+m105_108+m106_108+m107_108+m108_108+m109_108+m110_108+m111_108+m112_108+m113_108+m114_108+m115_108+m116_108+m117_108+m118_108+m119_108+m120_108+m121_108+m122_108+m123_108+m124_108+m125_108+m126_108+m127_108+m128_108+m129_108+m130_108+m131_108+m132_108+m133_108+m134_108+m135_108+m136_108+m137_108+m138_108+m139_108+m140_108+m141_108+m142_108+m143_108+m144_108+m145_108+m146_108+m147_108+m148_108+m149_108+m150_108+m151_108+m152_108+m153_108+m154_108+m155_108+m156_108+m157_108+m158_108+m159_108+m160_108+m161_108+m162_108+m163_108+m164_108+m165_108+m166_108+m167_108+m168_108+m169_108+m170_108+m171_108+m172_108+m173_108+m174_108+m175_108+m176_108+m177_108+m178_108+m179_108+m180_108+m181_108+m182_108+m183_108+m184_108+m185_108+m186_108+m187_108+m188_108+m189_108+m190_108+m191_108+m192_108+m193_108+m194_108+m195_108+m196_108+m197_108+m198_108+m199_108+m200_108+m201_108+m202_108+m203_108+m204_108+m205_108+m206_108+m207_108+m208_108+m209_108+m210_108+m211_108+m212_108+m213_108+m214_108+m215_108+m216_108+m217_108+m218_108+m219_108+m220_108+m221_108+m222_108+m223_108+m224_108+m225_108+m226_108+m227_108+m228_108+m229_108+m230_108+m231_108+m232_108+m233_108+m234_108+m235_108+m236_108+m237_108+m238_108+m239_108+m240_108+m241_108+m242_108+m243_108+m244_108+m245_108+m246_108+m247_108+m248_108+m249_108+m250_108+m251_108+m252_108+m253_108+m254_108+m255_108+m256_108+m257_108+m258_108+m259_108+m260_108+m261_108+m262_108+m263_108+m264_108+m265_108+m266_108+m267_108+m268_108+m269_108+m270_108+m271_108+m272_108+m273_108+m274_108+m275_108+m276_108+m277_108+m278_108+m279_108+m280_108+m281_108+m282_108+m283_108+m284_108+m285_108+m286_108+m287_108+m288_108+m289_108+m290_108+m291_108+m292_108+m293_108+m294_108+m295_108+m296_108+m297_108+m298_108+m299_108+m300_108+m301_108+m302_108+m303_108+m304_108+m305_108+m306_108+m307_108+m308_108+m309_108+m310_108+m311_108+m312_108+m313_108+m314_108+m315_108+m316_108+m317_108+m318_108+m319_108+m320_108+m321_108+m322_108+m323_108+m324_108+m325_108+m326_108+m327_108+m328_108+m329_108+m330_108+m331_108+m332_108+m333_108+m334_108+m335_108+m336_108+m337_108+m338_108+m339_108+m340_108+m341_108+m342_108+m343_108+m344_108+m345_108+m346_108+m347_108+m348_108+m349_108+m350_108+m351_108+m352_108+m353_108+m354_108+m355_108+m356_108+m357_108+m358_108+m359_108+m360_108+m361_108+m362_108+m363_108+m364_108+m365_108+m366_108+m367_108+m368_108+m369_108+m370_108+m371_108+m372_108+m373_108+m374_108+m375_108+m376_108+m377_108+m378_108+m379_108+m380_108+m381_108+b108;
   always @(posedge clk) out109 <= m1_109+m2_109+m3_109+m4_109+m5_109+m6_109+m7_109+m8_109+m9_109+m10_109+m11_109+m12_109+m13_109+m14_109+m15_109+m16_109+m17_109+m18_109+m19_109+m20_109+m21_109+m22_109+m23_109+m24_109+m25_109+m26_109+m27_109+m28_109+m29_109+m30_109+m31_109+m32_109+m33_109+m34_109+m35_109+m36_109+m37_109+m38_109+m39_109+m40_109+m41_109+m42_109+m43_109+m44_109+m45_109+m46_109+m47_109+m48_109+m49_109+m50_109+m51_109+m52_109+m53_109+m54_109+m55_109+m56_109+m57_109+m58_109+m59_109+m60_109+m61_109+m62_109+m63_109+m64_109+m65_109+m66_109+m67_109+m68_109+m69_109+m70_109+m71_109+m72_109+m73_109+m74_109+m75_109+m76_109+m77_109+m78_109+m79_109+m80_109+m81_109+m82_109+m83_109+m84_109+m85_109+m86_109+m87_109+m88_109+m89_109+m90_109+m91_109+m92_109+m93_109+m94_109+m95_109+m96_109+m97_109+m98_109+m99_109+m100_109+m101_109+m102_109+m103_109+m104_109+m105_109+m106_109+m107_109+m108_109+m109_109+m110_109+m111_109+m112_109+m113_109+m114_109+m115_109+m116_109+m117_109+m118_109+m119_109+m120_109+m121_109+m122_109+m123_109+m124_109+m125_109+m126_109+m127_109+m128_109+m129_109+m130_109+m131_109+m132_109+m133_109+m134_109+m135_109+m136_109+m137_109+m138_109+m139_109+m140_109+m141_109+m142_109+m143_109+m144_109+m145_109+m146_109+m147_109+m148_109+m149_109+m150_109+m151_109+m152_109+m153_109+m154_109+m155_109+m156_109+m157_109+m158_109+m159_109+m160_109+m161_109+m162_109+m163_109+m164_109+m165_109+m166_109+m167_109+m168_109+m169_109+m170_109+m171_109+m172_109+m173_109+m174_109+m175_109+m176_109+m177_109+m178_109+m179_109+m180_109+m181_109+m182_109+m183_109+m184_109+m185_109+m186_109+m187_109+m188_109+m189_109+m190_109+m191_109+m192_109+m193_109+m194_109+m195_109+m196_109+m197_109+m198_109+m199_109+m200_109+m201_109+m202_109+m203_109+m204_109+m205_109+m206_109+m207_109+m208_109+m209_109+m210_109+m211_109+m212_109+m213_109+m214_109+m215_109+m216_109+m217_109+m218_109+m219_109+m220_109+m221_109+m222_109+m223_109+m224_109+m225_109+m226_109+m227_109+m228_109+m229_109+m230_109+m231_109+m232_109+m233_109+m234_109+m235_109+m236_109+m237_109+m238_109+m239_109+m240_109+m241_109+m242_109+m243_109+m244_109+m245_109+m246_109+m247_109+m248_109+m249_109+m250_109+m251_109+m252_109+m253_109+m254_109+m255_109+m256_109+m257_109+m258_109+m259_109+m260_109+m261_109+m262_109+m263_109+m264_109+m265_109+m266_109+m267_109+m268_109+m269_109+m270_109+m271_109+m272_109+m273_109+m274_109+m275_109+m276_109+m277_109+m278_109+m279_109+m280_109+m281_109+m282_109+m283_109+m284_109+m285_109+m286_109+m287_109+m288_109+m289_109+m290_109+m291_109+m292_109+m293_109+m294_109+m295_109+m296_109+m297_109+m298_109+m299_109+m300_109+m301_109+m302_109+m303_109+m304_109+m305_109+m306_109+m307_109+m308_109+m309_109+m310_109+m311_109+m312_109+m313_109+m314_109+m315_109+m316_109+m317_109+m318_109+m319_109+m320_109+m321_109+m322_109+m323_109+m324_109+m325_109+m326_109+m327_109+m328_109+m329_109+m330_109+m331_109+m332_109+m333_109+m334_109+m335_109+m336_109+m337_109+m338_109+m339_109+m340_109+m341_109+m342_109+m343_109+m344_109+m345_109+m346_109+m347_109+m348_109+m349_109+m350_109+m351_109+m352_109+m353_109+m354_109+m355_109+m356_109+m357_109+m358_109+m359_109+m360_109+m361_109+m362_109+m363_109+m364_109+m365_109+m366_109+m367_109+m368_109+m369_109+m370_109+m371_109+m372_109+m373_109+m374_109+m375_109+m376_109+m377_109+m378_109+m379_109+m380_109+m381_109+b109;
   always @(posedge clk) out110 <= m1_110+m2_110+m3_110+m4_110+m5_110+m6_110+m7_110+m8_110+m9_110+m10_110+m11_110+m12_110+m13_110+m14_110+m15_110+m16_110+m17_110+m18_110+m19_110+m20_110+m21_110+m22_110+m23_110+m24_110+m25_110+m26_110+m27_110+m28_110+m29_110+m30_110+m31_110+m32_110+m33_110+m34_110+m35_110+m36_110+m37_110+m38_110+m39_110+m40_110+m41_110+m42_110+m43_110+m44_110+m45_110+m46_110+m47_110+m48_110+m49_110+m50_110+m51_110+m52_110+m53_110+m54_110+m55_110+m56_110+m57_110+m58_110+m59_110+m60_110+m61_110+m62_110+m63_110+m64_110+m65_110+m66_110+m67_110+m68_110+m69_110+m70_110+m71_110+m72_110+m73_110+m74_110+m75_110+m76_110+m77_110+m78_110+m79_110+m80_110+m81_110+m82_110+m83_110+m84_110+m85_110+m86_110+m87_110+m88_110+m89_110+m90_110+m91_110+m92_110+m93_110+m94_110+m95_110+m96_110+m97_110+m98_110+m99_110+m100_110+m101_110+m102_110+m103_110+m104_110+m105_110+m106_110+m107_110+m108_110+m109_110+m110_110+m111_110+m112_110+m113_110+m114_110+m115_110+m116_110+m117_110+m118_110+m119_110+m120_110+m121_110+m122_110+m123_110+m124_110+m125_110+m126_110+m127_110+m128_110+m129_110+m130_110+m131_110+m132_110+m133_110+m134_110+m135_110+m136_110+m137_110+m138_110+m139_110+m140_110+m141_110+m142_110+m143_110+m144_110+m145_110+m146_110+m147_110+m148_110+m149_110+m150_110+m151_110+m152_110+m153_110+m154_110+m155_110+m156_110+m157_110+m158_110+m159_110+m160_110+m161_110+m162_110+m163_110+m164_110+m165_110+m166_110+m167_110+m168_110+m169_110+m170_110+m171_110+m172_110+m173_110+m174_110+m175_110+m176_110+m177_110+m178_110+m179_110+m180_110+m181_110+m182_110+m183_110+m184_110+m185_110+m186_110+m187_110+m188_110+m189_110+m190_110+m191_110+m192_110+m193_110+m194_110+m195_110+m196_110+m197_110+m198_110+m199_110+m200_110+m201_110+m202_110+m203_110+m204_110+m205_110+m206_110+m207_110+m208_110+m209_110+m210_110+m211_110+m212_110+m213_110+m214_110+m215_110+m216_110+m217_110+m218_110+m219_110+m220_110+m221_110+m222_110+m223_110+m224_110+m225_110+m226_110+m227_110+m228_110+m229_110+m230_110+m231_110+m232_110+m233_110+m234_110+m235_110+m236_110+m237_110+m238_110+m239_110+m240_110+m241_110+m242_110+m243_110+m244_110+m245_110+m246_110+m247_110+m248_110+m249_110+m250_110+m251_110+m252_110+m253_110+m254_110+m255_110+m256_110+m257_110+m258_110+m259_110+m260_110+m261_110+m262_110+m263_110+m264_110+m265_110+m266_110+m267_110+m268_110+m269_110+m270_110+m271_110+m272_110+m273_110+m274_110+m275_110+m276_110+m277_110+m278_110+m279_110+m280_110+m281_110+m282_110+m283_110+m284_110+m285_110+m286_110+m287_110+m288_110+m289_110+m290_110+m291_110+m292_110+m293_110+m294_110+m295_110+m296_110+m297_110+m298_110+m299_110+m300_110+m301_110+m302_110+m303_110+m304_110+m305_110+m306_110+m307_110+m308_110+m309_110+m310_110+m311_110+m312_110+m313_110+m314_110+m315_110+m316_110+m317_110+m318_110+m319_110+m320_110+m321_110+m322_110+m323_110+m324_110+m325_110+m326_110+m327_110+m328_110+m329_110+m330_110+m331_110+m332_110+m333_110+m334_110+m335_110+m336_110+m337_110+m338_110+m339_110+m340_110+m341_110+m342_110+m343_110+m344_110+m345_110+m346_110+m347_110+m348_110+m349_110+m350_110+m351_110+m352_110+m353_110+m354_110+m355_110+m356_110+m357_110+m358_110+m359_110+m360_110+m361_110+m362_110+m363_110+m364_110+m365_110+m366_110+m367_110+m368_110+m369_110+m370_110+m371_110+m372_110+m373_110+m374_110+m375_110+m376_110+m377_110+m378_110+m379_110+m380_110+m381_110+b110;
   always @(posedge clk) out111 <= m1_111+m2_111+m3_111+m4_111+m5_111+m6_111+m7_111+m8_111+m9_111+m10_111+m11_111+m12_111+m13_111+m14_111+m15_111+m16_111+m17_111+m18_111+m19_111+m20_111+m21_111+m22_111+m23_111+m24_111+m25_111+m26_111+m27_111+m28_111+m29_111+m30_111+m31_111+m32_111+m33_111+m34_111+m35_111+m36_111+m37_111+m38_111+m39_111+m40_111+m41_111+m42_111+m43_111+m44_111+m45_111+m46_111+m47_111+m48_111+m49_111+m50_111+m51_111+m52_111+m53_111+m54_111+m55_111+m56_111+m57_111+m58_111+m59_111+m60_111+m61_111+m62_111+m63_111+m64_111+m65_111+m66_111+m67_111+m68_111+m69_111+m70_111+m71_111+m72_111+m73_111+m74_111+m75_111+m76_111+m77_111+m78_111+m79_111+m80_111+m81_111+m82_111+m83_111+m84_111+m85_111+m86_111+m87_111+m88_111+m89_111+m90_111+m91_111+m92_111+m93_111+m94_111+m95_111+m96_111+m97_111+m98_111+m99_111+m100_111+m101_111+m102_111+m103_111+m104_111+m105_111+m106_111+m107_111+m108_111+m109_111+m110_111+m111_111+m112_111+m113_111+m114_111+m115_111+m116_111+m117_111+m118_111+m119_111+m120_111+m121_111+m122_111+m123_111+m124_111+m125_111+m126_111+m127_111+m128_111+m129_111+m130_111+m131_111+m132_111+m133_111+m134_111+m135_111+m136_111+m137_111+m138_111+m139_111+m140_111+m141_111+m142_111+m143_111+m144_111+m145_111+m146_111+m147_111+m148_111+m149_111+m150_111+m151_111+m152_111+m153_111+m154_111+m155_111+m156_111+m157_111+m158_111+m159_111+m160_111+m161_111+m162_111+m163_111+m164_111+m165_111+m166_111+m167_111+m168_111+m169_111+m170_111+m171_111+m172_111+m173_111+m174_111+m175_111+m176_111+m177_111+m178_111+m179_111+m180_111+m181_111+m182_111+m183_111+m184_111+m185_111+m186_111+m187_111+m188_111+m189_111+m190_111+m191_111+m192_111+m193_111+m194_111+m195_111+m196_111+m197_111+m198_111+m199_111+m200_111+m201_111+m202_111+m203_111+m204_111+m205_111+m206_111+m207_111+m208_111+m209_111+m210_111+m211_111+m212_111+m213_111+m214_111+m215_111+m216_111+m217_111+m218_111+m219_111+m220_111+m221_111+m222_111+m223_111+m224_111+m225_111+m226_111+m227_111+m228_111+m229_111+m230_111+m231_111+m232_111+m233_111+m234_111+m235_111+m236_111+m237_111+m238_111+m239_111+m240_111+m241_111+m242_111+m243_111+m244_111+m245_111+m246_111+m247_111+m248_111+m249_111+m250_111+m251_111+m252_111+m253_111+m254_111+m255_111+m256_111+m257_111+m258_111+m259_111+m260_111+m261_111+m262_111+m263_111+m264_111+m265_111+m266_111+m267_111+m268_111+m269_111+m270_111+m271_111+m272_111+m273_111+m274_111+m275_111+m276_111+m277_111+m278_111+m279_111+m280_111+m281_111+m282_111+m283_111+m284_111+m285_111+m286_111+m287_111+m288_111+m289_111+m290_111+m291_111+m292_111+m293_111+m294_111+m295_111+m296_111+m297_111+m298_111+m299_111+m300_111+m301_111+m302_111+m303_111+m304_111+m305_111+m306_111+m307_111+m308_111+m309_111+m310_111+m311_111+m312_111+m313_111+m314_111+m315_111+m316_111+m317_111+m318_111+m319_111+m320_111+m321_111+m322_111+m323_111+m324_111+m325_111+m326_111+m327_111+m328_111+m329_111+m330_111+m331_111+m332_111+m333_111+m334_111+m335_111+m336_111+m337_111+m338_111+m339_111+m340_111+m341_111+m342_111+m343_111+m344_111+m345_111+m346_111+m347_111+m348_111+m349_111+m350_111+m351_111+m352_111+m353_111+m354_111+m355_111+m356_111+m357_111+m358_111+m359_111+m360_111+m361_111+m362_111+m363_111+m364_111+m365_111+m366_111+m367_111+m368_111+m369_111+m370_111+m371_111+m372_111+m373_111+m374_111+m375_111+m376_111+m377_111+m378_111+m379_111+m380_111+m381_111+b111;
   always @(posedge clk) out112 <= m1_112+m2_112+m3_112+m4_112+m5_112+m6_112+m7_112+m8_112+m9_112+m10_112+m11_112+m12_112+m13_112+m14_112+m15_112+m16_112+m17_112+m18_112+m19_112+m20_112+m21_112+m22_112+m23_112+m24_112+m25_112+m26_112+m27_112+m28_112+m29_112+m30_112+m31_112+m32_112+m33_112+m34_112+m35_112+m36_112+m37_112+m38_112+m39_112+m40_112+m41_112+m42_112+m43_112+m44_112+m45_112+m46_112+m47_112+m48_112+m49_112+m50_112+m51_112+m52_112+m53_112+m54_112+m55_112+m56_112+m57_112+m58_112+m59_112+m60_112+m61_112+m62_112+m63_112+m64_112+m65_112+m66_112+m67_112+m68_112+m69_112+m70_112+m71_112+m72_112+m73_112+m74_112+m75_112+m76_112+m77_112+m78_112+m79_112+m80_112+m81_112+m82_112+m83_112+m84_112+m85_112+m86_112+m87_112+m88_112+m89_112+m90_112+m91_112+m92_112+m93_112+m94_112+m95_112+m96_112+m97_112+m98_112+m99_112+m100_112+m101_112+m102_112+m103_112+m104_112+m105_112+m106_112+m107_112+m108_112+m109_112+m110_112+m111_112+m112_112+m113_112+m114_112+m115_112+m116_112+m117_112+m118_112+m119_112+m120_112+m121_112+m122_112+m123_112+m124_112+m125_112+m126_112+m127_112+m128_112+m129_112+m130_112+m131_112+m132_112+m133_112+m134_112+m135_112+m136_112+m137_112+m138_112+m139_112+m140_112+m141_112+m142_112+m143_112+m144_112+m145_112+m146_112+m147_112+m148_112+m149_112+m150_112+m151_112+m152_112+m153_112+m154_112+m155_112+m156_112+m157_112+m158_112+m159_112+m160_112+m161_112+m162_112+m163_112+m164_112+m165_112+m166_112+m167_112+m168_112+m169_112+m170_112+m171_112+m172_112+m173_112+m174_112+m175_112+m176_112+m177_112+m178_112+m179_112+m180_112+m181_112+m182_112+m183_112+m184_112+m185_112+m186_112+m187_112+m188_112+m189_112+m190_112+m191_112+m192_112+m193_112+m194_112+m195_112+m196_112+m197_112+m198_112+m199_112+m200_112+m201_112+m202_112+m203_112+m204_112+m205_112+m206_112+m207_112+m208_112+m209_112+m210_112+m211_112+m212_112+m213_112+m214_112+m215_112+m216_112+m217_112+m218_112+m219_112+m220_112+m221_112+m222_112+m223_112+m224_112+m225_112+m226_112+m227_112+m228_112+m229_112+m230_112+m231_112+m232_112+m233_112+m234_112+m235_112+m236_112+m237_112+m238_112+m239_112+m240_112+m241_112+m242_112+m243_112+m244_112+m245_112+m246_112+m247_112+m248_112+m249_112+m250_112+m251_112+m252_112+m253_112+m254_112+m255_112+m256_112+m257_112+m258_112+m259_112+m260_112+m261_112+m262_112+m263_112+m264_112+m265_112+m266_112+m267_112+m268_112+m269_112+m270_112+m271_112+m272_112+m273_112+m274_112+m275_112+m276_112+m277_112+m278_112+m279_112+m280_112+m281_112+m282_112+m283_112+m284_112+m285_112+m286_112+m287_112+m288_112+m289_112+m290_112+m291_112+m292_112+m293_112+m294_112+m295_112+m296_112+m297_112+m298_112+m299_112+m300_112+m301_112+m302_112+m303_112+m304_112+m305_112+m306_112+m307_112+m308_112+m309_112+m310_112+m311_112+m312_112+m313_112+m314_112+m315_112+m316_112+m317_112+m318_112+m319_112+m320_112+m321_112+m322_112+m323_112+m324_112+m325_112+m326_112+m327_112+m328_112+m329_112+m330_112+m331_112+m332_112+m333_112+m334_112+m335_112+m336_112+m337_112+m338_112+m339_112+m340_112+m341_112+m342_112+m343_112+m344_112+m345_112+m346_112+m347_112+m348_112+m349_112+m350_112+m351_112+m352_112+m353_112+m354_112+m355_112+m356_112+m357_112+m358_112+m359_112+m360_112+m361_112+m362_112+m363_112+m364_112+m365_112+m366_112+m367_112+m368_112+m369_112+m370_112+m371_112+m372_112+m373_112+m374_112+m375_112+m376_112+m377_112+m378_112+m379_112+m380_112+m381_112+b112;
   always @(posedge clk) out113 <= m1_113+m2_113+m3_113+m4_113+m5_113+m6_113+m7_113+m8_113+m9_113+m10_113+m11_113+m12_113+m13_113+m14_113+m15_113+m16_113+m17_113+m18_113+m19_113+m20_113+m21_113+m22_113+m23_113+m24_113+m25_113+m26_113+m27_113+m28_113+m29_113+m30_113+m31_113+m32_113+m33_113+m34_113+m35_113+m36_113+m37_113+m38_113+m39_113+m40_113+m41_113+m42_113+m43_113+m44_113+m45_113+m46_113+m47_113+m48_113+m49_113+m50_113+m51_113+m52_113+m53_113+m54_113+m55_113+m56_113+m57_113+m58_113+m59_113+m60_113+m61_113+m62_113+m63_113+m64_113+m65_113+m66_113+m67_113+m68_113+m69_113+m70_113+m71_113+m72_113+m73_113+m74_113+m75_113+m76_113+m77_113+m78_113+m79_113+m80_113+m81_113+m82_113+m83_113+m84_113+m85_113+m86_113+m87_113+m88_113+m89_113+m90_113+m91_113+m92_113+m93_113+m94_113+m95_113+m96_113+m97_113+m98_113+m99_113+m100_113+m101_113+m102_113+m103_113+m104_113+m105_113+m106_113+m107_113+m108_113+m109_113+m110_113+m111_113+m112_113+m113_113+m114_113+m115_113+m116_113+m117_113+m118_113+m119_113+m120_113+m121_113+m122_113+m123_113+m124_113+m125_113+m126_113+m127_113+m128_113+m129_113+m130_113+m131_113+m132_113+m133_113+m134_113+m135_113+m136_113+m137_113+m138_113+m139_113+m140_113+m141_113+m142_113+m143_113+m144_113+m145_113+m146_113+m147_113+m148_113+m149_113+m150_113+m151_113+m152_113+m153_113+m154_113+m155_113+m156_113+m157_113+m158_113+m159_113+m160_113+m161_113+m162_113+m163_113+m164_113+m165_113+m166_113+m167_113+m168_113+m169_113+m170_113+m171_113+m172_113+m173_113+m174_113+m175_113+m176_113+m177_113+m178_113+m179_113+m180_113+m181_113+m182_113+m183_113+m184_113+m185_113+m186_113+m187_113+m188_113+m189_113+m190_113+m191_113+m192_113+m193_113+m194_113+m195_113+m196_113+m197_113+m198_113+m199_113+m200_113+m201_113+m202_113+m203_113+m204_113+m205_113+m206_113+m207_113+m208_113+m209_113+m210_113+m211_113+m212_113+m213_113+m214_113+m215_113+m216_113+m217_113+m218_113+m219_113+m220_113+m221_113+m222_113+m223_113+m224_113+m225_113+m226_113+m227_113+m228_113+m229_113+m230_113+m231_113+m232_113+m233_113+m234_113+m235_113+m236_113+m237_113+m238_113+m239_113+m240_113+m241_113+m242_113+m243_113+m244_113+m245_113+m246_113+m247_113+m248_113+m249_113+m250_113+m251_113+m252_113+m253_113+m254_113+m255_113+m256_113+m257_113+m258_113+m259_113+m260_113+m261_113+m262_113+m263_113+m264_113+m265_113+m266_113+m267_113+m268_113+m269_113+m270_113+m271_113+m272_113+m273_113+m274_113+m275_113+m276_113+m277_113+m278_113+m279_113+m280_113+m281_113+m282_113+m283_113+m284_113+m285_113+m286_113+m287_113+m288_113+m289_113+m290_113+m291_113+m292_113+m293_113+m294_113+m295_113+m296_113+m297_113+m298_113+m299_113+m300_113+m301_113+m302_113+m303_113+m304_113+m305_113+m306_113+m307_113+m308_113+m309_113+m310_113+m311_113+m312_113+m313_113+m314_113+m315_113+m316_113+m317_113+m318_113+m319_113+m320_113+m321_113+m322_113+m323_113+m324_113+m325_113+m326_113+m327_113+m328_113+m329_113+m330_113+m331_113+m332_113+m333_113+m334_113+m335_113+m336_113+m337_113+m338_113+m339_113+m340_113+m341_113+m342_113+m343_113+m344_113+m345_113+m346_113+m347_113+m348_113+m349_113+m350_113+m351_113+m352_113+m353_113+m354_113+m355_113+m356_113+m357_113+m358_113+m359_113+m360_113+m361_113+m362_113+m363_113+m364_113+m365_113+m366_113+m367_113+m368_113+m369_113+m370_113+m371_113+m372_113+m373_113+m374_113+m375_113+m376_113+m377_113+m378_113+m379_113+m380_113+m381_113+b113;
   always @(posedge clk) out114 <= m1_114+m2_114+m3_114+m4_114+m5_114+m6_114+m7_114+m8_114+m9_114+m10_114+m11_114+m12_114+m13_114+m14_114+m15_114+m16_114+m17_114+m18_114+m19_114+m20_114+m21_114+m22_114+m23_114+m24_114+m25_114+m26_114+m27_114+m28_114+m29_114+m30_114+m31_114+m32_114+m33_114+m34_114+m35_114+m36_114+m37_114+m38_114+m39_114+m40_114+m41_114+m42_114+m43_114+m44_114+m45_114+m46_114+m47_114+m48_114+m49_114+m50_114+m51_114+m52_114+m53_114+m54_114+m55_114+m56_114+m57_114+m58_114+m59_114+m60_114+m61_114+m62_114+m63_114+m64_114+m65_114+m66_114+m67_114+m68_114+m69_114+m70_114+m71_114+m72_114+m73_114+m74_114+m75_114+m76_114+m77_114+m78_114+m79_114+m80_114+m81_114+m82_114+m83_114+m84_114+m85_114+m86_114+m87_114+m88_114+m89_114+m90_114+m91_114+m92_114+m93_114+m94_114+m95_114+m96_114+m97_114+m98_114+m99_114+m100_114+m101_114+m102_114+m103_114+m104_114+m105_114+m106_114+m107_114+m108_114+m109_114+m110_114+m111_114+m112_114+m113_114+m114_114+m115_114+m116_114+m117_114+m118_114+m119_114+m120_114+m121_114+m122_114+m123_114+m124_114+m125_114+m126_114+m127_114+m128_114+m129_114+m130_114+m131_114+m132_114+m133_114+m134_114+m135_114+m136_114+m137_114+m138_114+m139_114+m140_114+m141_114+m142_114+m143_114+m144_114+m145_114+m146_114+m147_114+m148_114+m149_114+m150_114+m151_114+m152_114+m153_114+m154_114+m155_114+m156_114+m157_114+m158_114+m159_114+m160_114+m161_114+m162_114+m163_114+m164_114+m165_114+m166_114+m167_114+m168_114+m169_114+m170_114+m171_114+m172_114+m173_114+m174_114+m175_114+m176_114+m177_114+m178_114+m179_114+m180_114+m181_114+m182_114+m183_114+m184_114+m185_114+m186_114+m187_114+m188_114+m189_114+m190_114+m191_114+m192_114+m193_114+m194_114+m195_114+m196_114+m197_114+m198_114+m199_114+m200_114+m201_114+m202_114+m203_114+m204_114+m205_114+m206_114+m207_114+m208_114+m209_114+m210_114+m211_114+m212_114+m213_114+m214_114+m215_114+m216_114+m217_114+m218_114+m219_114+m220_114+m221_114+m222_114+m223_114+m224_114+m225_114+m226_114+m227_114+m228_114+m229_114+m230_114+m231_114+m232_114+m233_114+m234_114+m235_114+m236_114+m237_114+m238_114+m239_114+m240_114+m241_114+m242_114+m243_114+m244_114+m245_114+m246_114+m247_114+m248_114+m249_114+m250_114+m251_114+m252_114+m253_114+m254_114+m255_114+m256_114+m257_114+m258_114+m259_114+m260_114+m261_114+m262_114+m263_114+m264_114+m265_114+m266_114+m267_114+m268_114+m269_114+m270_114+m271_114+m272_114+m273_114+m274_114+m275_114+m276_114+m277_114+m278_114+m279_114+m280_114+m281_114+m282_114+m283_114+m284_114+m285_114+m286_114+m287_114+m288_114+m289_114+m290_114+m291_114+m292_114+m293_114+m294_114+m295_114+m296_114+m297_114+m298_114+m299_114+m300_114+m301_114+m302_114+m303_114+m304_114+m305_114+m306_114+m307_114+m308_114+m309_114+m310_114+m311_114+m312_114+m313_114+m314_114+m315_114+m316_114+m317_114+m318_114+m319_114+m320_114+m321_114+m322_114+m323_114+m324_114+m325_114+m326_114+m327_114+m328_114+m329_114+m330_114+m331_114+m332_114+m333_114+m334_114+m335_114+m336_114+m337_114+m338_114+m339_114+m340_114+m341_114+m342_114+m343_114+m344_114+m345_114+m346_114+m347_114+m348_114+m349_114+m350_114+m351_114+m352_114+m353_114+m354_114+m355_114+m356_114+m357_114+m358_114+m359_114+m360_114+m361_114+m362_114+m363_114+m364_114+m365_114+m366_114+m367_114+m368_114+m369_114+m370_114+m371_114+m372_114+m373_114+m374_114+m375_114+m376_114+m377_114+m378_114+m379_114+m380_114+m381_114+b114;
   always @(posedge clk) out115 <= m1_115+m2_115+m3_115+m4_115+m5_115+m6_115+m7_115+m8_115+m9_115+m10_115+m11_115+m12_115+m13_115+m14_115+m15_115+m16_115+m17_115+m18_115+m19_115+m20_115+m21_115+m22_115+m23_115+m24_115+m25_115+m26_115+m27_115+m28_115+m29_115+m30_115+m31_115+m32_115+m33_115+m34_115+m35_115+m36_115+m37_115+m38_115+m39_115+m40_115+m41_115+m42_115+m43_115+m44_115+m45_115+m46_115+m47_115+m48_115+m49_115+m50_115+m51_115+m52_115+m53_115+m54_115+m55_115+m56_115+m57_115+m58_115+m59_115+m60_115+m61_115+m62_115+m63_115+m64_115+m65_115+m66_115+m67_115+m68_115+m69_115+m70_115+m71_115+m72_115+m73_115+m74_115+m75_115+m76_115+m77_115+m78_115+m79_115+m80_115+m81_115+m82_115+m83_115+m84_115+m85_115+m86_115+m87_115+m88_115+m89_115+m90_115+m91_115+m92_115+m93_115+m94_115+m95_115+m96_115+m97_115+m98_115+m99_115+m100_115+m101_115+m102_115+m103_115+m104_115+m105_115+m106_115+m107_115+m108_115+m109_115+m110_115+m111_115+m112_115+m113_115+m114_115+m115_115+m116_115+m117_115+m118_115+m119_115+m120_115+m121_115+m122_115+m123_115+m124_115+m125_115+m126_115+m127_115+m128_115+m129_115+m130_115+m131_115+m132_115+m133_115+m134_115+m135_115+m136_115+m137_115+m138_115+m139_115+m140_115+m141_115+m142_115+m143_115+m144_115+m145_115+m146_115+m147_115+m148_115+m149_115+m150_115+m151_115+m152_115+m153_115+m154_115+m155_115+m156_115+m157_115+m158_115+m159_115+m160_115+m161_115+m162_115+m163_115+m164_115+m165_115+m166_115+m167_115+m168_115+m169_115+m170_115+m171_115+m172_115+m173_115+m174_115+m175_115+m176_115+m177_115+m178_115+m179_115+m180_115+m181_115+m182_115+m183_115+m184_115+m185_115+m186_115+m187_115+m188_115+m189_115+m190_115+m191_115+m192_115+m193_115+m194_115+m195_115+m196_115+m197_115+m198_115+m199_115+m200_115+m201_115+m202_115+m203_115+m204_115+m205_115+m206_115+m207_115+m208_115+m209_115+m210_115+m211_115+m212_115+m213_115+m214_115+m215_115+m216_115+m217_115+m218_115+m219_115+m220_115+m221_115+m222_115+m223_115+m224_115+m225_115+m226_115+m227_115+m228_115+m229_115+m230_115+m231_115+m232_115+m233_115+m234_115+m235_115+m236_115+m237_115+m238_115+m239_115+m240_115+m241_115+m242_115+m243_115+m244_115+m245_115+m246_115+m247_115+m248_115+m249_115+m250_115+m251_115+m252_115+m253_115+m254_115+m255_115+m256_115+m257_115+m258_115+m259_115+m260_115+m261_115+m262_115+m263_115+m264_115+m265_115+m266_115+m267_115+m268_115+m269_115+m270_115+m271_115+m272_115+m273_115+m274_115+m275_115+m276_115+m277_115+m278_115+m279_115+m280_115+m281_115+m282_115+m283_115+m284_115+m285_115+m286_115+m287_115+m288_115+m289_115+m290_115+m291_115+m292_115+m293_115+m294_115+m295_115+m296_115+m297_115+m298_115+m299_115+m300_115+m301_115+m302_115+m303_115+m304_115+m305_115+m306_115+m307_115+m308_115+m309_115+m310_115+m311_115+m312_115+m313_115+m314_115+m315_115+m316_115+m317_115+m318_115+m319_115+m320_115+m321_115+m322_115+m323_115+m324_115+m325_115+m326_115+m327_115+m328_115+m329_115+m330_115+m331_115+m332_115+m333_115+m334_115+m335_115+m336_115+m337_115+m338_115+m339_115+m340_115+m341_115+m342_115+m343_115+m344_115+m345_115+m346_115+m347_115+m348_115+m349_115+m350_115+m351_115+m352_115+m353_115+m354_115+m355_115+m356_115+m357_115+m358_115+m359_115+m360_115+m361_115+m362_115+m363_115+m364_115+m365_115+m366_115+m367_115+m368_115+m369_115+m370_115+m371_115+m372_115+m373_115+m374_115+m375_115+m376_115+m377_115+m378_115+m379_115+m380_115+m381_115+b115;
   always @(posedge clk) out116 <= m1_116+m2_116+m3_116+m4_116+m5_116+m6_116+m7_116+m8_116+m9_116+m10_116+m11_116+m12_116+m13_116+m14_116+m15_116+m16_116+m17_116+m18_116+m19_116+m20_116+m21_116+m22_116+m23_116+m24_116+m25_116+m26_116+m27_116+m28_116+m29_116+m30_116+m31_116+m32_116+m33_116+m34_116+m35_116+m36_116+m37_116+m38_116+m39_116+m40_116+m41_116+m42_116+m43_116+m44_116+m45_116+m46_116+m47_116+m48_116+m49_116+m50_116+m51_116+m52_116+m53_116+m54_116+m55_116+m56_116+m57_116+m58_116+m59_116+m60_116+m61_116+m62_116+m63_116+m64_116+m65_116+m66_116+m67_116+m68_116+m69_116+m70_116+m71_116+m72_116+m73_116+m74_116+m75_116+m76_116+m77_116+m78_116+m79_116+m80_116+m81_116+m82_116+m83_116+m84_116+m85_116+m86_116+m87_116+m88_116+m89_116+m90_116+m91_116+m92_116+m93_116+m94_116+m95_116+m96_116+m97_116+m98_116+m99_116+m100_116+m101_116+m102_116+m103_116+m104_116+m105_116+m106_116+m107_116+m108_116+m109_116+m110_116+m111_116+m112_116+m113_116+m114_116+m115_116+m116_116+m117_116+m118_116+m119_116+m120_116+m121_116+m122_116+m123_116+m124_116+m125_116+m126_116+m127_116+m128_116+m129_116+m130_116+m131_116+m132_116+m133_116+m134_116+m135_116+m136_116+m137_116+m138_116+m139_116+m140_116+m141_116+m142_116+m143_116+m144_116+m145_116+m146_116+m147_116+m148_116+m149_116+m150_116+m151_116+m152_116+m153_116+m154_116+m155_116+m156_116+m157_116+m158_116+m159_116+m160_116+m161_116+m162_116+m163_116+m164_116+m165_116+m166_116+m167_116+m168_116+m169_116+m170_116+m171_116+m172_116+m173_116+m174_116+m175_116+m176_116+m177_116+m178_116+m179_116+m180_116+m181_116+m182_116+m183_116+m184_116+m185_116+m186_116+m187_116+m188_116+m189_116+m190_116+m191_116+m192_116+m193_116+m194_116+m195_116+m196_116+m197_116+m198_116+m199_116+m200_116+m201_116+m202_116+m203_116+m204_116+m205_116+m206_116+m207_116+m208_116+m209_116+m210_116+m211_116+m212_116+m213_116+m214_116+m215_116+m216_116+m217_116+m218_116+m219_116+m220_116+m221_116+m222_116+m223_116+m224_116+m225_116+m226_116+m227_116+m228_116+m229_116+m230_116+m231_116+m232_116+m233_116+m234_116+m235_116+m236_116+m237_116+m238_116+m239_116+m240_116+m241_116+m242_116+m243_116+m244_116+m245_116+m246_116+m247_116+m248_116+m249_116+m250_116+m251_116+m252_116+m253_116+m254_116+m255_116+m256_116+m257_116+m258_116+m259_116+m260_116+m261_116+m262_116+m263_116+m264_116+m265_116+m266_116+m267_116+m268_116+m269_116+m270_116+m271_116+m272_116+m273_116+m274_116+m275_116+m276_116+m277_116+m278_116+m279_116+m280_116+m281_116+m282_116+m283_116+m284_116+m285_116+m286_116+m287_116+m288_116+m289_116+m290_116+m291_116+m292_116+m293_116+m294_116+m295_116+m296_116+m297_116+m298_116+m299_116+m300_116+m301_116+m302_116+m303_116+m304_116+m305_116+m306_116+m307_116+m308_116+m309_116+m310_116+m311_116+m312_116+m313_116+m314_116+m315_116+m316_116+m317_116+m318_116+m319_116+m320_116+m321_116+m322_116+m323_116+m324_116+m325_116+m326_116+m327_116+m328_116+m329_116+m330_116+m331_116+m332_116+m333_116+m334_116+m335_116+m336_116+m337_116+m338_116+m339_116+m340_116+m341_116+m342_116+m343_116+m344_116+m345_116+m346_116+m347_116+m348_116+m349_116+m350_116+m351_116+m352_116+m353_116+m354_116+m355_116+m356_116+m357_116+m358_116+m359_116+m360_116+m361_116+m362_116+m363_116+m364_116+m365_116+m366_116+m367_116+m368_116+m369_116+m370_116+m371_116+m372_116+m373_116+m374_116+m375_116+m376_116+m377_116+m378_116+m379_116+m380_116+m381_116+b116;
   always @(posedge clk) out117 <= m1_117+m2_117+m3_117+m4_117+m5_117+m6_117+m7_117+m8_117+m9_117+m10_117+m11_117+m12_117+m13_117+m14_117+m15_117+m16_117+m17_117+m18_117+m19_117+m20_117+m21_117+m22_117+m23_117+m24_117+m25_117+m26_117+m27_117+m28_117+m29_117+m30_117+m31_117+m32_117+m33_117+m34_117+m35_117+m36_117+m37_117+m38_117+m39_117+m40_117+m41_117+m42_117+m43_117+m44_117+m45_117+m46_117+m47_117+m48_117+m49_117+m50_117+m51_117+m52_117+m53_117+m54_117+m55_117+m56_117+m57_117+m58_117+m59_117+m60_117+m61_117+m62_117+m63_117+m64_117+m65_117+m66_117+m67_117+m68_117+m69_117+m70_117+m71_117+m72_117+m73_117+m74_117+m75_117+m76_117+m77_117+m78_117+m79_117+m80_117+m81_117+m82_117+m83_117+m84_117+m85_117+m86_117+m87_117+m88_117+m89_117+m90_117+m91_117+m92_117+m93_117+m94_117+m95_117+m96_117+m97_117+m98_117+m99_117+m100_117+m101_117+m102_117+m103_117+m104_117+m105_117+m106_117+m107_117+m108_117+m109_117+m110_117+m111_117+m112_117+m113_117+m114_117+m115_117+m116_117+m117_117+m118_117+m119_117+m120_117+m121_117+m122_117+m123_117+m124_117+m125_117+m126_117+m127_117+m128_117+m129_117+m130_117+m131_117+m132_117+m133_117+m134_117+m135_117+m136_117+m137_117+m138_117+m139_117+m140_117+m141_117+m142_117+m143_117+m144_117+m145_117+m146_117+m147_117+m148_117+m149_117+m150_117+m151_117+m152_117+m153_117+m154_117+m155_117+m156_117+m157_117+m158_117+m159_117+m160_117+m161_117+m162_117+m163_117+m164_117+m165_117+m166_117+m167_117+m168_117+m169_117+m170_117+m171_117+m172_117+m173_117+m174_117+m175_117+m176_117+m177_117+m178_117+m179_117+m180_117+m181_117+m182_117+m183_117+m184_117+m185_117+m186_117+m187_117+m188_117+m189_117+m190_117+m191_117+m192_117+m193_117+m194_117+m195_117+m196_117+m197_117+m198_117+m199_117+m200_117+m201_117+m202_117+m203_117+m204_117+m205_117+m206_117+m207_117+m208_117+m209_117+m210_117+m211_117+m212_117+m213_117+m214_117+m215_117+m216_117+m217_117+m218_117+m219_117+m220_117+m221_117+m222_117+m223_117+m224_117+m225_117+m226_117+m227_117+m228_117+m229_117+m230_117+m231_117+m232_117+m233_117+m234_117+m235_117+m236_117+m237_117+m238_117+m239_117+m240_117+m241_117+m242_117+m243_117+m244_117+m245_117+m246_117+m247_117+m248_117+m249_117+m250_117+m251_117+m252_117+m253_117+m254_117+m255_117+m256_117+m257_117+m258_117+m259_117+m260_117+m261_117+m262_117+m263_117+m264_117+m265_117+m266_117+m267_117+m268_117+m269_117+m270_117+m271_117+m272_117+m273_117+m274_117+m275_117+m276_117+m277_117+m278_117+m279_117+m280_117+m281_117+m282_117+m283_117+m284_117+m285_117+m286_117+m287_117+m288_117+m289_117+m290_117+m291_117+m292_117+m293_117+m294_117+m295_117+m296_117+m297_117+m298_117+m299_117+m300_117+m301_117+m302_117+m303_117+m304_117+m305_117+m306_117+m307_117+m308_117+m309_117+m310_117+m311_117+m312_117+m313_117+m314_117+m315_117+m316_117+m317_117+m318_117+m319_117+m320_117+m321_117+m322_117+m323_117+m324_117+m325_117+m326_117+m327_117+m328_117+m329_117+m330_117+m331_117+m332_117+m333_117+m334_117+m335_117+m336_117+m337_117+m338_117+m339_117+m340_117+m341_117+m342_117+m343_117+m344_117+m345_117+m346_117+m347_117+m348_117+m349_117+m350_117+m351_117+m352_117+m353_117+m354_117+m355_117+m356_117+m357_117+m358_117+m359_117+m360_117+m361_117+m362_117+m363_117+m364_117+m365_117+m366_117+m367_117+m368_117+m369_117+m370_117+m371_117+m372_117+m373_117+m374_117+m375_117+m376_117+m377_117+m378_117+m379_117+m380_117+m381_117+b117;
endmodule