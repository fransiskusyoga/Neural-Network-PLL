module lenet300_top(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   input [14:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598;
   output [15:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   wire signed [14:0] s2_1,s2_2,s2_3,s2_4,s2_5,s2_6,s2_7,s2_8,s2_9,s2_10,s2_11,s2_12,s2_13,s2_14,s2_15,s2_16,s2_17,s2_18,s2_19,s2_20,s2_21,s2_22,s2_23,s2_24,s2_25,s2_26,s2_27,s2_28,s2_29,s2_30,s2_31,s2_32,s2_33,s2_34,s2_35,s2_36,s2_37,s2_38,s2_39,s2_40,s2_41,s2_42,s2_43,s2_44,s2_45,s2_46,s2_47,s2_48,s2_49,s2_50,s2_51,s2_52,s2_53,s2_54,s2_55,s2_56,s2_57,s2_58,s2_59,s2_60,s2_61,s2_62,s2_63,s2_64,s2_65,s2_66,s2_67,s2_68,s2_69,s2_70,s2_71,s2_72,s2_73,s2_74,s2_75,s2_76,s2_77,s2_78,s2_79,s2_80,s2_81,s2_82,s2_83,s2_84,s2_85,s2_86,s2_87,s2_88,s2_89,s2_90,s2_91,s2_92,s2_93,s2_94,s2_95,s2_96,s2_97,s2_98,s2_99,s2_100,s2_101,s2_102,s2_103,s2_104,s2_105,s2_106,s2_107,s2_108,s2_109,s2_110,s2_111,s2_112,s2_113,s2_114,s2_115,s2_116,s2_117,s2_118,s2_119,s2_120,s2_121,s2_122,s2_123,s2_124,s2_125,s2_126,s2_127,s2_128,s2_129,s2_130,s2_131,s2_132,s2_133,s2_134,s2_135,s2_136,s2_137,s2_138,s2_139,s2_140,s2_141,s2_142,s2_143,s2_144,s2_145,s2_146,s2_147,s2_148,s2_149,s2_150,s2_151,s2_152,s2_153,s2_154,s2_155,s2_156,s2_157,s2_158,s2_159,s2_160,s2_161,s2_162,s2_163,s2_164,s2_165,s2_166,s2_167,s2_168,s2_169,s2_170,s2_171,s2_172,s2_173,s2_174,s2_175,s2_176,s2_177,s2_178,s2_179,s2_180,s2_181,s2_182,s2_183,s2_184,s2_185,s2_186,s2_187,s2_188,s2_189,s2_190,s2_191,s2_192,s2_193,s2_194,s2_195,s2_196,s2_197,s2_198,s2_199,s2_200,s2_201,s2_202,s2_203,s2_204,s2_205,s2_206,s2_207,s2_208,s2_209,s2_210,s2_211,s2_212,s2_213,s2_214,s2_215,s2_216,s2_217,s2_218,s2_219,s2_220,s2_221,s2_222,s2_223,s2_224,s2_225,s2_226,s2_227,s2_228,s2_229,s2_230,s2_231,s2_232,s2_233,s2_234,s2_235,s2_236,s2_237,s2_238,s2_239,s2_240,s2_241,s2_242,s2_243,s2_244,s2_245,s2_246,s2_247,s2_248,s2_249,s2_250,s2_251,s2_252,s2_253,s2_254,s2_255,s2_256,s2_257,s2_258,s2_259,s2_260,s2_261,s2_262,s2_263;
   wire signed [14:0] s3_1,s3_2,s3_3,s3_4,s3_5,s3_6,s3_7,s3_8,s3_9,s3_10,s3_11,s3_12,s3_13,s3_14,s3_15,s3_16,s3_17,s3_18,s3_19,s3_20,s3_21,s3_22,s3_23,s3_24,s3_25,s3_26,s3_27,s3_28,s3_29,s3_30,s3_31,s3_32,s3_33,s3_34,s3_35,s3_36,s3_37,s3_38,s3_39,s3_40,s3_41,s3_42,s3_43,s3_44,s3_45,s3_46,s3_47,s3_48,s3_49,s3_50,s3_51,s3_52,s3_53,s3_54,s3_55,s3_56,s3_57,s3_58,s3_59,s3_60,s3_61,s3_62,s3_63,s3_64,s3_65,s3_66,s3_67,s3_68,s3_69,s3_70,s3_71,s3_72,s3_73,s3_74,s3_75,s3_76,s3_77,s3_78,s3_79,s3_80,s3_81,s3_82,s3_83,s3_84,s3_85,s3_86,s3_87,s3_88,s3_89,s3_90,s3_91,s3_92,s3_93,s3_94,s3_95,s3_96,s3_97,s3_98,s3_99,s3_100;
   wire signed [14:0] h2_1,h2_2,h2_3,h2_4,h2_5,h2_6,h2_7,h2_8,h2_9,h2_10,h2_11,h2_12,h2_13,h2_14,h2_15,h2_16,h2_17,h2_18,h2_19,h2_20,h2_21,h2_22,h2_23,h2_24,h2_25,h2_26,h2_27,h2_28,h2_29,h2_30,h2_31,h2_32,h2_33,h2_34,h2_35,h2_36,h2_37,h2_38,h2_39,h2_40,h2_41,h2_42,h2_43,h2_44,h2_45,h2_46,h2_47,h2_48,h2_49,h2_50,h2_51,h2_52,h2_53,h2_54,h2_55,h2_56,h2_57,h2_58,h2_59,h2_60,h2_61,h2_62,h2_63,h2_64,h2_65,h2_66,h2_67,h2_68,h2_69,h2_70,h2_71,h2_72,h2_73,h2_74,h2_75,h2_76,h2_77,h2_78,h2_79,h2_80,h2_81,h2_82,h2_83,h2_84,h2_85,h2_86,h2_87,h2_88,h2_89,h2_90,h2_91,h2_92,h2_93,h2_94,h2_95,h2_96,h2_97,h2_98,h2_99,h2_100,h2_101,h2_102,h2_103,h2_104,h2_105,h2_106,h2_107,h2_108,h2_109,h2_110,h2_111,h2_112,h2_113,h2_114,h2_115,h2_116,h2_117,h2_118,h2_119,h2_120,h2_121,h2_122,h2_123,h2_124,h2_125,h2_126,h2_127,h2_128,h2_129,h2_130,h2_131,h2_132,h2_133,h2_134,h2_135,h2_136,h2_137,h2_138,h2_139,h2_140,h2_141,h2_142,h2_143,h2_144,h2_145,h2_146,h2_147,h2_148,h2_149,h2_150,h2_151,h2_152,h2_153,h2_154,h2_155,h2_156,h2_157,h2_158,h2_159,h2_160,h2_161,h2_162,h2_163,h2_164,h2_165,h2_166,h2_167,h2_168,h2_169,h2_170,h2_171,h2_172,h2_173,h2_174,h2_175,h2_176,h2_177,h2_178,h2_179,h2_180,h2_181,h2_182,h2_183,h2_184,h2_185,h2_186,h2_187,h2_188,h2_189,h2_190,h2_191,h2_192,h2_193,h2_194,h2_195,h2_196,h2_197,h2_198,h2_199,h2_200,h2_201,h2_202,h2_203,h2_204,h2_205,h2_206,h2_207,h2_208,h2_209,h2_210,h2_211,h2_212,h2_213,h2_214,h2_215,h2_216,h2_217,h2_218,h2_219,h2_220,h2_221,h2_222,h2_223,h2_224,h2_225,h2_226,h2_227,h2_228,h2_229,h2_230,h2_231,h2_232,h2_233,h2_234,h2_235,h2_236,h2_237,h2_238,h2_239,h2_240,h2_241,h2_242,h2_243,h2_244,h2_245,h2_246,h2_247,h2_248,h2_249,h2_250,h2_251,h2_252,h2_253,h2_254,h2_255,h2_256,h2_257,h2_258,h2_259,h2_260,h2_261,h2_262,h2_263;
   wire signed [14:0] h3_1,h3_2,h3_3,h3_4,h3_5,h3_6,h3_7,h3_8,h3_9,h3_10,h3_11,h3_12,h3_13,h3_14,h3_15,h3_16,h3_17,h3_18,h3_19,h3_20,h3_21,h3_22,h3_23,h3_24,h3_25,h3_26,h3_27,h3_28,h3_29,h3_30,h3_31,h3_32,h3_33,h3_34,h3_35,h3_36,h3_37,h3_38,h3_39,h3_40,h3_41,h3_42,h3_43,h3_44,h3_45,h3_46,h3_47,h3_48,h3_49,h3_50,h3_51,h3_52,h3_53,h3_54,h3_55,h3_56,h3_57,h3_58,h3_59,h3_60,h3_61,h3_62,h3_63,h3_64,h3_65,h3_66,h3_67,h3_68,h3_69,h3_70,h3_71,h3_72,h3_73,h3_74,h3_75,h3_76,h3_77,h3_78,h3_79,h3_80,h3_81,h3_82,h3_83,h3_84,h3_85,h3_86,h3_87,h3_88,h3_89,h3_90,h3_91,h3_92,h3_93,h3_94,h3_95,h3_96,h3_97,h3_98,h3_99,h3_100;
   lenet300_layer_1 L1(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598,s2_1,s2_2,s2_3,s2_4,s2_5,s2_6,s2_7,s2_8,s2_9,s2_10,s2_11,s2_12,s2_13,s2_14,s2_15,s2_16,s2_17,s2_18,s2_19,s2_20,s2_21,s2_22,s2_23,s2_24,s2_25,s2_26,s2_27,s2_28,s2_29,s2_30,s2_31,s2_32,s2_33,s2_34,s2_35,s2_36,s2_37,s2_38,s2_39,s2_40,s2_41,s2_42,s2_43,s2_44,s2_45,s2_46,s2_47,s2_48,s2_49,s2_50,s2_51,s2_52,s2_53,s2_54,s2_55,s2_56,s2_57,s2_58,s2_59,s2_60,s2_61,s2_62,s2_63,s2_64,s2_65,s2_66,s2_67,s2_68,s2_69,s2_70,s2_71,s2_72,s2_73,s2_74,s2_75,s2_76,s2_77,s2_78,s2_79,s2_80,s2_81,s2_82,s2_83,s2_84,s2_85,s2_86,s2_87,s2_88,s2_89,s2_90,s2_91,s2_92,s2_93,s2_94,s2_95,s2_96,s2_97,s2_98,s2_99,s2_100,s2_101,s2_102,s2_103,s2_104,s2_105,s2_106,s2_107,s2_108,s2_109,s2_110,s2_111,s2_112,s2_113,s2_114,s2_115,s2_116,s2_117,s2_118,s2_119,s2_120,s2_121,s2_122,s2_123,s2_124,s2_125,s2_126,s2_127,s2_128,s2_129,s2_130,s2_131,s2_132,s2_133,s2_134,s2_135,s2_136,s2_137,s2_138,s2_139,s2_140,s2_141,s2_142,s2_143,s2_144,s2_145,s2_146,s2_147,s2_148,s2_149,s2_150,s2_151,s2_152,s2_153,s2_154,s2_155,s2_156,s2_157,s2_158,s2_159,s2_160,s2_161,s2_162,s2_163,s2_164,s2_165,s2_166,s2_167,s2_168,s2_169,s2_170,s2_171,s2_172,s2_173,s2_174,s2_175,s2_176,s2_177,s2_178,s2_179,s2_180,s2_181,s2_182,s2_183,s2_184,s2_185,s2_186,s2_187,s2_188,s2_189,s2_190,s2_191,s2_192,s2_193,s2_194,s2_195,s2_196,s2_197,s2_198,s2_199,s2_200,s2_201,s2_202,s2_203,s2_204,s2_205,s2_206,s2_207,s2_208,s2_209,s2_210,s2_211,s2_212,s2_213,s2_214,s2_215,s2_216,s2_217,s2_218,s2_219,s2_220,s2_221,s2_222,s2_223,s2_224,s2_225,s2_226,s2_227,s2_228,s2_229,s2_230,s2_231,s2_232,s2_233,s2_234,s2_235,s2_236,s2_237,s2_238,s2_239,s2_240,s2_241,s2_242,s2_243,s2_244,s2_245,s2_246,s2_247,s2_248,s2_249,s2_250,s2_251,s2_252,s2_253,s2_254,s2_255,s2_256,s2_257,s2_258,s2_259,s2_260,s2_261,s2_262,s2_263);
   actifunc #(15) AF2_1(s2_1,h2_1);
   actifunc #(15) AF2_2(s2_2,h2_2);
   actifunc #(15) AF2_3(s2_3,h2_3);
   actifunc #(15) AF2_4(s2_4,h2_4);
   actifunc #(15) AF2_5(s2_5,h2_5);
   actifunc #(15) AF2_6(s2_6,h2_6);
   actifunc #(15) AF2_7(s2_7,h2_7);
   actifunc #(15) AF2_8(s2_8,h2_8);
   actifunc #(15) AF2_9(s2_9,h2_9);
   actifunc #(15) AF2_10(s2_10,h2_10);
   actifunc #(15) AF2_11(s2_11,h2_11);
   actifunc #(15) AF2_12(s2_12,h2_12);
   actifunc #(15) AF2_13(s2_13,h2_13);
   actifunc #(15) AF2_14(s2_14,h2_14);
   actifunc #(15) AF2_15(s2_15,h2_15);
   actifunc #(15) AF2_16(s2_16,h2_16);
   actifunc #(15) AF2_17(s2_17,h2_17);
   actifunc #(15) AF2_18(s2_18,h2_18);
   actifunc #(15) AF2_19(s2_19,h2_19);
   actifunc #(15) AF2_20(s2_20,h2_20);
   actifunc #(15) AF2_21(s2_21,h2_21);
   actifunc #(15) AF2_22(s2_22,h2_22);
   actifunc #(15) AF2_23(s2_23,h2_23);
   actifunc #(15) AF2_24(s2_24,h2_24);
   actifunc #(15) AF2_25(s2_25,h2_25);
   actifunc #(15) AF2_26(s2_26,h2_26);
   actifunc #(15) AF2_27(s2_27,h2_27);
   actifunc #(15) AF2_28(s2_28,h2_28);
   actifunc #(15) AF2_29(s2_29,h2_29);
   actifunc #(15) AF2_30(s2_30,h2_30);
   actifunc #(15) AF2_31(s2_31,h2_31);
   actifunc #(15) AF2_32(s2_32,h2_32);
   actifunc #(15) AF2_33(s2_33,h2_33);
   actifunc #(15) AF2_34(s2_34,h2_34);
   actifunc #(15) AF2_35(s2_35,h2_35);
   actifunc #(15) AF2_36(s2_36,h2_36);
   actifunc #(15) AF2_37(s2_37,h2_37);
   actifunc #(15) AF2_38(s2_38,h2_38);
   actifunc #(15) AF2_39(s2_39,h2_39);
   actifunc #(15) AF2_40(s2_40,h2_40);
   actifunc #(15) AF2_41(s2_41,h2_41);
   actifunc #(15) AF2_42(s2_42,h2_42);
   actifunc #(15) AF2_43(s2_43,h2_43);
   actifunc #(15) AF2_44(s2_44,h2_44);
   actifunc #(15) AF2_45(s2_45,h2_45);
   actifunc #(15) AF2_46(s2_46,h2_46);
   actifunc #(15) AF2_47(s2_47,h2_47);
   actifunc #(15) AF2_48(s2_48,h2_48);
   actifunc #(15) AF2_49(s2_49,h2_49);
   actifunc #(15) AF2_50(s2_50,h2_50);
   actifunc #(15) AF2_51(s2_51,h2_51);
   actifunc #(15) AF2_52(s2_52,h2_52);
   actifunc #(15) AF2_53(s2_53,h2_53);
   actifunc #(15) AF2_54(s2_54,h2_54);
   actifunc #(15) AF2_55(s2_55,h2_55);
   actifunc #(15) AF2_56(s2_56,h2_56);
   actifunc #(15) AF2_57(s2_57,h2_57);
   actifunc #(15) AF2_58(s2_58,h2_58);
   actifunc #(15) AF2_59(s2_59,h2_59);
   actifunc #(15) AF2_60(s2_60,h2_60);
   actifunc #(15) AF2_61(s2_61,h2_61);
   actifunc #(15) AF2_62(s2_62,h2_62);
   actifunc #(15) AF2_63(s2_63,h2_63);
   actifunc #(15) AF2_64(s2_64,h2_64);
   actifunc #(15) AF2_65(s2_65,h2_65);
   actifunc #(15) AF2_66(s2_66,h2_66);
   actifunc #(15) AF2_67(s2_67,h2_67);
   actifunc #(15) AF2_68(s2_68,h2_68);
   actifunc #(15) AF2_69(s2_69,h2_69);
   actifunc #(15) AF2_70(s2_70,h2_70);
   actifunc #(15) AF2_71(s2_71,h2_71);
   actifunc #(15) AF2_72(s2_72,h2_72);
   actifunc #(15) AF2_73(s2_73,h2_73);
   actifunc #(15) AF2_74(s2_74,h2_74);
   actifunc #(15) AF2_75(s2_75,h2_75);
   actifunc #(15) AF2_76(s2_76,h2_76);
   actifunc #(15) AF2_77(s2_77,h2_77);
   actifunc #(15) AF2_78(s2_78,h2_78);
   actifunc #(15) AF2_79(s2_79,h2_79);
   actifunc #(15) AF2_80(s2_80,h2_80);
   actifunc #(15) AF2_81(s2_81,h2_81);
   actifunc #(15) AF2_82(s2_82,h2_82);
   actifunc #(15) AF2_83(s2_83,h2_83);
   actifunc #(15) AF2_84(s2_84,h2_84);
   actifunc #(15) AF2_85(s2_85,h2_85);
   actifunc #(15) AF2_86(s2_86,h2_86);
   actifunc #(15) AF2_87(s2_87,h2_87);
   actifunc #(15) AF2_88(s2_88,h2_88);
   actifunc #(15) AF2_89(s2_89,h2_89);
   actifunc #(15) AF2_90(s2_90,h2_90);
   actifunc #(15) AF2_91(s2_91,h2_91);
   actifunc #(15) AF2_92(s2_92,h2_92);
   actifunc #(15) AF2_93(s2_93,h2_93);
   actifunc #(15) AF2_94(s2_94,h2_94);
   actifunc #(15) AF2_95(s2_95,h2_95);
   actifunc #(15) AF2_96(s2_96,h2_96);
   actifunc #(15) AF2_97(s2_97,h2_97);
   actifunc #(15) AF2_98(s2_98,h2_98);
   actifunc #(15) AF2_99(s2_99,h2_99);
   actifunc #(15) AF2_100(s2_100,h2_100);
   actifunc #(15) AF2_101(s2_101,h2_101);
   actifunc #(15) AF2_102(s2_102,h2_102);
   actifunc #(15) AF2_103(s2_103,h2_103);
   actifunc #(15) AF2_104(s2_104,h2_104);
   actifunc #(15) AF2_105(s2_105,h2_105);
   actifunc #(15) AF2_106(s2_106,h2_106);
   actifunc #(15) AF2_107(s2_107,h2_107);
   actifunc #(15) AF2_108(s2_108,h2_108);
   actifunc #(15) AF2_109(s2_109,h2_109);
   actifunc #(15) AF2_110(s2_110,h2_110);
   actifunc #(15) AF2_111(s2_111,h2_111);
   actifunc #(15) AF2_112(s2_112,h2_112);
   actifunc #(15) AF2_113(s2_113,h2_113);
   actifunc #(15) AF2_114(s2_114,h2_114);
   actifunc #(15) AF2_115(s2_115,h2_115);
   actifunc #(15) AF2_116(s2_116,h2_116);
   actifunc #(15) AF2_117(s2_117,h2_117);
   actifunc #(15) AF2_118(s2_118,h2_118);
   actifunc #(15) AF2_119(s2_119,h2_119);
   actifunc #(15) AF2_120(s2_120,h2_120);
   actifunc #(15) AF2_121(s2_121,h2_121);
   actifunc #(15) AF2_122(s2_122,h2_122);
   actifunc #(15) AF2_123(s2_123,h2_123);
   actifunc #(15) AF2_124(s2_124,h2_124);
   actifunc #(15) AF2_125(s2_125,h2_125);
   actifunc #(15) AF2_126(s2_126,h2_126);
   actifunc #(15) AF2_127(s2_127,h2_127);
   actifunc #(15) AF2_128(s2_128,h2_128);
   actifunc #(15) AF2_129(s2_129,h2_129);
   actifunc #(15) AF2_130(s2_130,h2_130);
   actifunc #(15) AF2_131(s2_131,h2_131);
   actifunc #(15) AF2_132(s2_132,h2_132);
   actifunc #(15) AF2_133(s2_133,h2_133);
   actifunc #(15) AF2_134(s2_134,h2_134);
   actifunc #(15) AF2_135(s2_135,h2_135);
   actifunc #(15) AF2_136(s2_136,h2_136);
   actifunc #(15) AF2_137(s2_137,h2_137);
   actifunc #(15) AF2_138(s2_138,h2_138);
   actifunc #(15) AF2_139(s2_139,h2_139);
   actifunc #(15) AF2_140(s2_140,h2_140);
   actifunc #(15) AF2_141(s2_141,h2_141);
   actifunc #(15) AF2_142(s2_142,h2_142);
   actifunc #(15) AF2_143(s2_143,h2_143);
   actifunc #(15) AF2_144(s2_144,h2_144);
   actifunc #(15) AF2_145(s2_145,h2_145);
   actifunc #(15) AF2_146(s2_146,h2_146);
   actifunc #(15) AF2_147(s2_147,h2_147);
   actifunc #(15) AF2_148(s2_148,h2_148);
   actifunc #(15) AF2_149(s2_149,h2_149);
   actifunc #(15) AF2_150(s2_150,h2_150);
   actifunc #(15) AF2_151(s2_151,h2_151);
   actifunc #(15) AF2_152(s2_152,h2_152);
   actifunc #(15) AF2_153(s2_153,h2_153);
   actifunc #(15) AF2_154(s2_154,h2_154);
   actifunc #(15) AF2_155(s2_155,h2_155);
   actifunc #(15) AF2_156(s2_156,h2_156);
   actifunc #(15) AF2_157(s2_157,h2_157);
   actifunc #(15) AF2_158(s2_158,h2_158);
   actifunc #(15) AF2_159(s2_159,h2_159);
   actifunc #(15) AF2_160(s2_160,h2_160);
   actifunc #(15) AF2_161(s2_161,h2_161);
   actifunc #(15) AF2_162(s2_162,h2_162);
   actifunc #(15) AF2_163(s2_163,h2_163);
   actifunc #(15) AF2_164(s2_164,h2_164);
   actifunc #(15) AF2_165(s2_165,h2_165);
   actifunc #(15) AF2_166(s2_166,h2_166);
   actifunc #(15) AF2_167(s2_167,h2_167);
   actifunc #(15) AF2_168(s2_168,h2_168);
   actifunc #(15) AF2_169(s2_169,h2_169);
   actifunc #(15) AF2_170(s2_170,h2_170);
   actifunc #(15) AF2_171(s2_171,h2_171);
   actifunc #(15) AF2_172(s2_172,h2_172);
   actifunc #(15) AF2_173(s2_173,h2_173);
   actifunc #(15) AF2_174(s2_174,h2_174);
   actifunc #(15) AF2_175(s2_175,h2_175);
   actifunc #(15) AF2_176(s2_176,h2_176);
   actifunc #(15) AF2_177(s2_177,h2_177);
   actifunc #(15) AF2_178(s2_178,h2_178);
   actifunc #(15) AF2_179(s2_179,h2_179);
   actifunc #(15) AF2_180(s2_180,h2_180);
   actifunc #(15) AF2_181(s2_181,h2_181);
   actifunc #(15) AF2_182(s2_182,h2_182);
   actifunc #(15) AF2_183(s2_183,h2_183);
   actifunc #(15) AF2_184(s2_184,h2_184);
   actifunc #(15) AF2_185(s2_185,h2_185);
   actifunc #(15) AF2_186(s2_186,h2_186);
   actifunc #(15) AF2_187(s2_187,h2_187);
   actifunc #(15) AF2_188(s2_188,h2_188);
   actifunc #(15) AF2_189(s2_189,h2_189);
   actifunc #(15) AF2_190(s2_190,h2_190);
   actifunc #(15) AF2_191(s2_191,h2_191);
   actifunc #(15) AF2_192(s2_192,h2_192);
   actifunc #(15) AF2_193(s2_193,h2_193);
   actifunc #(15) AF2_194(s2_194,h2_194);
   actifunc #(15) AF2_195(s2_195,h2_195);
   actifunc #(15) AF2_196(s2_196,h2_196);
   actifunc #(15) AF2_197(s2_197,h2_197);
   actifunc #(15) AF2_198(s2_198,h2_198);
   actifunc #(15) AF2_199(s2_199,h2_199);
   actifunc #(15) AF2_200(s2_200,h2_200);
   actifunc #(15) AF2_201(s2_201,h2_201);
   actifunc #(15) AF2_202(s2_202,h2_202);
   actifunc #(15) AF2_203(s2_203,h2_203);
   actifunc #(15) AF2_204(s2_204,h2_204);
   actifunc #(15) AF2_205(s2_205,h2_205);
   actifunc #(15) AF2_206(s2_206,h2_206);
   actifunc #(15) AF2_207(s2_207,h2_207);
   actifunc #(15) AF2_208(s2_208,h2_208);
   actifunc #(15) AF2_209(s2_209,h2_209);
   actifunc #(15) AF2_210(s2_210,h2_210);
   actifunc #(15) AF2_211(s2_211,h2_211);
   actifunc #(15) AF2_212(s2_212,h2_212);
   actifunc #(15) AF2_213(s2_213,h2_213);
   actifunc #(15) AF2_214(s2_214,h2_214);
   actifunc #(15) AF2_215(s2_215,h2_215);
   actifunc #(15) AF2_216(s2_216,h2_216);
   actifunc #(15) AF2_217(s2_217,h2_217);
   actifunc #(15) AF2_218(s2_218,h2_218);
   actifunc #(15) AF2_219(s2_219,h2_219);
   actifunc #(15) AF2_220(s2_220,h2_220);
   actifunc #(15) AF2_221(s2_221,h2_221);
   actifunc #(15) AF2_222(s2_222,h2_222);
   actifunc #(15) AF2_223(s2_223,h2_223);
   actifunc #(15) AF2_224(s2_224,h2_224);
   actifunc #(15) AF2_225(s2_225,h2_225);
   actifunc #(15) AF2_226(s2_226,h2_226);
   actifunc #(15) AF2_227(s2_227,h2_227);
   actifunc #(15) AF2_228(s2_228,h2_228);
   actifunc #(15) AF2_229(s2_229,h2_229);
   actifunc #(15) AF2_230(s2_230,h2_230);
   actifunc #(15) AF2_231(s2_231,h2_231);
   actifunc #(15) AF2_232(s2_232,h2_232);
   actifunc #(15) AF2_233(s2_233,h2_233);
   actifunc #(15) AF2_234(s2_234,h2_234);
   actifunc #(15) AF2_235(s2_235,h2_235);
   actifunc #(15) AF2_236(s2_236,h2_236);
   actifunc #(15) AF2_237(s2_237,h2_237);
   actifunc #(15) AF2_238(s2_238,h2_238);
   actifunc #(15) AF2_239(s2_239,h2_239);
   actifunc #(15) AF2_240(s2_240,h2_240);
   actifunc #(15) AF2_241(s2_241,h2_241);
   actifunc #(15) AF2_242(s2_242,h2_242);
   actifunc #(15) AF2_243(s2_243,h2_243);
   actifunc #(15) AF2_244(s2_244,h2_244);
   actifunc #(15) AF2_245(s2_245,h2_245);
   actifunc #(15) AF2_246(s2_246,h2_246);
   actifunc #(15) AF2_247(s2_247,h2_247);
   actifunc #(15) AF2_248(s2_248,h2_248);
   actifunc #(15) AF2_249(s2_249,h2_249);
   actifunc #(15) AF2_250(s2_250,h2_250);
   actifunc #(15) AF2_251(s2_251,h2_251);
   actifunc #(15) AF2_252(s2_252,h2_252);
   actifunc #(15) AF2_253(s2_253,h2_253);
   actifunc #(15) AF2_254(s2_254,h2_254);
   actifunc #(15) AF2_255(s2_255,h2_255);
   actifunc #(15) AF2_256(s2_256,h2_256);
   actifunc #(15) AF2_257(s2_257,h2_257);
   actifunc #(15) AF2_258(s2_258,h2_258);
   actifunc #(15) AF2_259(s2_259,h2_259);
   actifunc #(15) AF2_260(s2_260,h2_260);
   actifunc #(15) AF2_261(s2_261,h2_261);
   actifunc #(15) AF2_262(s2_262,h2_262);
   actifunc #(15) AF2_263(s2_263,h2_263);
   lenet300_layer_2 L2(h2_1[14:0],h2_2[14:0],h2_3[14:0],h2_4[14:0],h2_5[14:0],h2_6[14:0],h2_7[14:0],h2_8[14:0],h2_9[14:0],h2_10[14:0],h2_11[14:0],h2_12[14:0],h2_13[14:0],h2_14[14:0],h2_15[14:0],h2_16[14:0],h2_17[14:0],h2_18[14:0],h2_19[14:0],h2_20[14:0],h2_21[14:0],h2_22[14:0],h2_23[14:0],h2_24[14:0],h2_25[14:0],h2_26[14:0],h2_27[14:0],h2_28[14:0],h2_29[14:0],h2_30[14:0],h2_31[14:0],h2_32[14:0],h2_33[14:0],h2_34[14:0],h2_35[14:0],h2_36[14:0],h2_37[14:0],h2_38[14:0],h2_39[14:0],h2_40[14:0],h2_41[14:0],h2_42[14:0],h2_43[14:0],h2_44[14:0],h2_45[14:0],h2_46[14:0],h2_47[14:0],h2_48[14:0],h2_49[14:0],h2_50[14:0],h2_51[14:0],h2_52[14:0],h2_53[14:0],h2_54[14:0],h2_55[14:0],h2_56[14:0],h2_57[14:0],h2_58[14:0],h2_59[14:0],h2_60[14:0],h2_61[14:0],h2_62[14:0],h2_63[14:0],h2_64[14:0],h2_65[14:0],h2_66[14:0],h2_67[14:0],h2_68[14:0],h2_69[14:0],h2_70[14:0],h2_71[14:0],h2_72[14:0],h2_73[14:0],h2_74[14:0],h2_75[14:0],h2_76[14:0],h2_77[14:0],h2_78[14:0],h2_79[14:0],h2_80[14:0],h2_81[14:0],h2_82[14:0],h2_83[14:0],h2_84[14:0],h2_85[14:0],h2_86[14:0],h2_87[14:0],h2_88[14:0],h2_89[14:0],h2_90[14:0],h2_91[14:0],h2_92[14:0],h2_93[14:0],h2_94[14:0],h2_95[14:0],h2_96[14:0],h2_97[14:0],h2_98[14:0],h2_99[14:0],h2_100[14:0],h2_101[14:0],h2_102[14:0],h2_103[14:0],h2_104[14:0],h2_105[14:0],h2_106[14:0],h2_107[14:0],h2_108[14:0],h2_109[14:0],h2_110[14:0],h2_111[14:0],h2_112[14:0],h2_113[14:0],h2_114[14:0],h2_115[14:0],h2_116[14:0],h2_117[14:0],h2_118[14:0],h2_119[14:0],h2_120[14:0],h2_121[14:0],h2_122[14:0],h2_123[14:0],h2_124[14:0],h2_125[14:0],h2_126[14:0],h2_127[14:0],h2_128[14:0],h2_129[14:0],h2_130[14:0],h2_131[14:0],h2_132[14:0],h2_133[14:0],h2_134[14:0],h2_135[14:0],h2_136[14:0],h2_137[14:0],h2_138[14:0],h2_139[14:0],h2_140[14:0],h2_141[14:0],h2_142[14:0],h2_143[14:0],h2_144[14:0],h2_145[14:0],h2_146[14:0],h2_147[14:0],h2_148[14:0],h2_149[14:0],h2_150[14:0],h2_151[14:0],h2_152[14:0],h2_153[14:0],h2_154[14:0],h2_155[14:0],h2_156[14:0],h2_157[14:0],h2_158[14:0],h2_159[14:0],h2_160[14:0],h2_161[14:0],h2_162[14:0],h2_163[14:0],h2_164[14:0],h2_165[14:0],h2_166[14:0],h2_167[14:0],h2_168[14:0],h2_169[14:0],h2_170[14:0],h2_171[14:0],h2_172[14:0],h2_173[14:0],h2_174[14:0],h2_175[14:0],h2_176[14:0],h2_177[14:0],h2_178[14:0],h2_179[14:0],h2_180[14:0],h2_181[14:0],h2_182[14:0],h2_183[14:0],h2_184[14:0],h2_185[14:0],h2_186[14:0],h2_187[14:0],h2_188[14:0],h2_189[14:0],h2_190[14:0],h2_191[14:0],h2_192[14:0],h2_193[14:0],h2_194[14:0],h2_195[14:0],h2_196[14:0],h2_197[14:0],h2_198[14:0],h2_199[14:0],h2_200[14:0],h2_201[14:0],h2_202[14:0],h2_203[14:0],h2_204[14:0],h2_205[14:0],h2_206[14:0],h2_207[14:0],h2_208[14:0],h2_209[14:0],h2_210[14:0],h2_211[14:0],h2_212[14:0],h2_213[14:0],h2_214[14:0],h2_215[14:0],h2_216[14:0],h2_217[14:0],h2_218[14:0],h2_219[14:0],h2_220[14:0],h2_221[14:0],h2_222[14:0],h2_223[14:0],h2_224[14:0],h2_225[14:0],h2_226[14:0],h2_227[14:0],h2_228[14:0],h2_229[14:0],h2_230[14:0],h2_231[14:0],h2_232[14:0],h2_233[14:0],h2_234[14:0],h2_235[14:0],h2_236[14:0],h2_237[14:0],h2_238[14:0],h2_239[14:0],h2_240[14:0],h2_241[14:0],h2_242[14:0],h2_243[14:0],h2_244[14:0],h2_245[14:0],h2_246[14:0],h2_247[14:0],h2_248[14:0],h2_249[14:0],h2_250[14:0],h2_251[14:0],h2_252[14:0],h2_253[14:0],h2_254[14:0],h2_255[14:0],h2_256[14:0],h2_257[14:0],h2_258[14:0],h2_259[14:0],h2_260[14:0],h2_261[14:0],h2_262[14:0],h2_263[14:0],s3_1,s3_2,s3_3,s3_4,s3_5,s3_6,s3_7,s3_8,s3_9,s3_10,s3_11,s3_12,s3_13,s3_14,s3_15,s3_16,s3_17,s3_18,s3_19,s3_20,s3_21,s3_22,s3_23,s3_24,s3_25,s3_26,s3_27,s3_28,s3_29,s3_30,s3_31,s3_32,s3_33,s3_34,s3_35,s3_36,s3_37,s3_38,s3_39,s3_40,s3_41,s3_42,s3_43,s3_44,s3_45,s3_46,s3_47,s3_48,s3_49,s3_50,s3_51,s3_52,s3_53,s3_54,s3_55,s3_56,s3_57,s3_58,s3_59,s3_60,s3_61,s3_62,s3_63,s3_64,s3_65,s3_66,s3_67,s3_68,s3_69,s3_70,s3_71,s3_72,s3_73,s3_74,s3_75,s3_76,s3_77,s3_78,s3_79,s3_80,s3_81,s3_82,s3_83,s3_84,s3_85,s3_86,s3_87,s3_88,s3_89,s3_90,s3_91,s3_92,s3_93,s3_94,s3_95,s3_96,s3_97,s3_98,s3_99,s3_100);
   actifunc #(15) AF3_1(s3_1,h3_1);
   actifunc #(15) AF3_2(s3_2,h3_2);
   actifunc #(15) AF3_3(s3_3,h3_3);
   actifunc #(15) AF3_4(s3_4,h3_4);
   actifunc #(15) AF3_5(s3_5,h3_5);
   actifunc #(15) AF3_6(s3_6,h3_6);
   actifunc #(15) AF3_7(s3_7,h3_7);
   actifunc #(15) AF3_8(s3_8,h3_8);
   actifunc #(15) AF3_9(s3_9,h3_9);
   actifunc #(15) AF3_10(s3_10,h3_10);
   actifunc #(15) AF3_11(s3_11,h3_11);
   actifunc #(15) AF3_12(s3_12,h3_12);
   actifunc #(15) AF3_13(s3_13,h3_13);
   actifunc #(15) AF3_14(s3_14,h3_14);
   actifunc #(15) AF3_15(s3_15,h3_15);
   actifunc #(15) AF3_16(s3_16,h3_16);
   actifunc #(15) AF3_17(s3_17,h3_17);
   actifunc #(15) AF3_18(s3_18,h3_18);
   actifunc #(15) AF3_19(s3_19,h3_19);
   actifunc #(15) AF3_20(s3_20,h3_20);
   actifunc #(15) AF3_21(s3_21,h3_21);
   actifunc #(15) AF3_22(s3_22,h3_22);
   actifunc #(15) AF3_23(s3_23,h3_23);
   actifunc #(15) AF3_24(s3_24,h3_24);
   actifunc #(15) AF3_25(s3_25,h3_25);
   actifunc #(15) AF3_26(s3_26,h3_26);
   actifunc #(15) AF3_27(s3_27,h3_27);
   actifunc #(15) AF3_28(s3_28,h3_28);
   actifunc #(15) AF3_29(s3_29,h3_29);
   actifunc #(15) AF3_30(s3_30,h3_30);
   actifunc #(15) AF3_31(s3_31,h3_31);
   actifunc #(15) AF3_32(s3_32,h3_32);
   actifunc #(15) AF3_33(s3_33,h3_33);
   actifunc #(15) AF3_34(s3_34,h3_34);
   actifunc #(15) AF3_35(s3_35,h3_35);
   actifunc #(15) AF3_36(s3_36,h3_36);
   actifunc #(15) AF3_37(s3_37,h3_37);
   actifunc #(15) AF3_38(s3_38,h3_38);
   actifunc #(15) AF3_39(s3_39,h3_39);
   actifunc #(15) AF3_40(s3_40,h3_40);
   actifunc #(15) AF3_41(s3_41,h3_41);
   actifunc #(15) AF3_42(s3_42,h3_42);
   actifunc #(15) AF3_43(s3_43,h3_43);
   actifunc #(15) AF3_44(s3_44,h3_44);
   actifunc #(15) AF3_45(s3_45,h3_45);
   actifunc #(15) AF3_46(s3_46,h3_46);
   actifunc #(15) AF3_47(s3_47,h3_47);
   actifunc #(15) AF3_48(s3_48,h3_48);
   actifunc #(15) AF3_49(s3_49,h3_49);
   actifunc #(15) AF3_50(s3_50,h3_50);
   actifunc #(15) AF3_51(s3_51,h3_51);
   actifunc #(15) AF3_52(s3_52,h3_52);
   actifunc #(15) AF3_53(s3_53,h3_53);
   actifunc #(15) AF3_54(s3_54,h3_54);
   actifunc #(15) AF3_55(s3_55,h3_55);
   actifunc #(15) AF3_56(s3_56,h3_56);
   actifunc #(15) AF3_57(s3_57,h3_57);
   actifunc #(15) AF3_58(s3_58,h3_58);
   actifunc #(15) AF3_59(s3_59,h3_59);
   actifunc #(15) AF3_60(s3_60,h3_60);
   actifunc #(15) AF3_61(s3_61,h3_61);
   actifunc #(15) AF3_62(s3_62,h3_62);
   actifunc #(15) AF3_63(s3_63,h3_63);
   actifunc #(15) AF3_64(s3_64,h3_64);
   actifunc #(15) AF3_65(s3_65,h3_65);
   actifunc #(15) AF3_66(s3_66,h3_66);
   actifunc #(15) AF3_67(s3_67,h3_67);
   actifunc #(15) AF3_68(s3_68,h3_68);
   actifunc #(15) AF3_69(s3_69,h3_69);
   actifunc #(15) AF3_70(s3_70,h3_70);
   actifunc #(15) AF3_71(s3_71,h3_71);
   actifunc #(15) AF3_72(s3_72,h3_72);
   actifunc #(15) AF3_73(s3_73,h3_73);
   actifunc #(15) AF3_74(s3_74,h3_74);
   actifunc #(15) AF3_75(s3_75,h3_75);
   actifunc #(15) AF3_76(s3_76,h3_76);
   actifunc #(15) AF3_77(s3_77,h3_77);
   actifunc #(15) AF3_78(s3_78,h3_78);
   actifunc #(15) AF3_79(s3_79,h3_79);
   actifunc #(15) AF3_80(s3_80,h3_80);
   actifunc #(15) AF3_81(s3_81,h3_81);
   actifunc #(15) AF3_82(s3_82,h3_82);
   actifunc #(15) AF3_83(s3_83,h3_83);
   actifunc #(15) AF3_84(s3_84,h3_84);
   actifunc #(15) AF3_85(s3_85,h3_85);
   actifunc #(15) AF3_86(s3_86,h3_86);
   actifunc #(15) AF3_87(s3_87,h3_87);
   actifunc #(15) AF3_88(s3_88,h3_88);
   actifunc #(15) AF3_89(s3_89,h3_89);
   actifunc #(15) AF3_90(s3_90,h3_90);
   actifunc #(15) AF3_91(s3_91,h3_91);
   actifunc #(15) AF3_92(s3_92,h3_92);
   actifunc #(15) AF3_93(s3_93,h3_93);
   actifunc #(15) AF3_94(s3_94,h3_94);
   actifunc #(15) AF3_95(s3_95,h3_95);
   actifunc #(15) AF3_96(s3_96,h3_96);
   actifunc #(15) AF3_97(s3_97,h3_97);
   actifunc #(15) AF3_98(s3_98,h3_98);
   actifunc #(15) AF3_99(s3_99,h3_99);
   actifunc #(15) AF3_100(s3_100,h3_100);
   lenet300_layer_3 L3(h3_1[15:0],h3_2[15:0],h3_3[15:0],h3_4[15:0],h3_5[15:0],h3_6[15:0],h3_7[15:0],h3_8[15:0],h3_9[15:0],h3_10[15:0],h3_11[15:0],h3_12[15:0],h3_13[15:0],h3_14[15:0],h3_15[15:0],h3_16[15:0],h3_17[15:0],h3_18[15:0],h3_19[15:0],h3_20[15:0],h3_21[15:0],h3_22[15:0],h3_23[15:0],h3_24[15:0],h3_25[15:0],h3_26[15:0],h3_27[15:0],h3_28[15:0],h3_29[15:0],h3_30[15:0],h3_31[15:0],h3_32[15:0],h3_33[15:0],h3_34[15:0],h3_35[15:0],h3_36[15:0],h3_37[15:0],h3_38[15:0],h3_39[15:0],h3_40[15:0],h3_41[15:0],h3_42[15:0],h3_43[15:0],h3_44[15:0],h3_45[15:0],h3_46[15:0],h3_47[15:0],h3_48[15:0],h3_49[15:0],h3_50[15:0],h3_51[15:0],h3_52[15:0],h3_53[15:0],h3_54[15:0],h3_55[15:0],h3_56[15:0],h3_57[15:0],h3_58[15:0],h3_59[15:0],h3_60[15:0],h3_61[15:0],h3_62[15:0],h3_63[15:0],h3_64[15:0],h3_65[15:0],h3_66[15:0],h3_67[15:0],h3_68[15:0],h3_69[15:0],h3_70[15:0],h3_71[15:0],h3_72[15:0],h3_73[15:0],h3_74[15:0],h3_75[15:0],h3_76[15:0],h3_77[15:0],h3_78[15:0],h3_79[15:0],h3_80[15:0],h3_81[15:0],h3_82[15:0],h3_83[15:0],h3_84[15:0],h3_85[15:0],h3_86[15:0],h3_87[15:0],h3_88[15:0],h3_89[15:0],h3_90[15:0],h3_91[15:0],h3_92[15:0],h3_93[15:0],h3_94[15:0],h3_95[15:0],h3_96[15:0],h3_97[15:0],h3_98[15:0],h3_99[15:0],h3_100[15:0],out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
endmodule