module tanh(in,out);
   // 1 sign bit, 2 decimal, 13 fractional
   input signed [15:0] in;
   // 1 sign bit, 0 decimal, 7 fractional
   output [7:0] out;
   //not implemented yet
endmodule
