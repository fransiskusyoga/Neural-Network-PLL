module test_tb();
   reg [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80;
   wire [7:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   test_top TopModule(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   initial begin
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'hC; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h4; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h3; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h2; in23=6'h0; in24=6'h0; in25=6'h1; in26=6'h1; in27=6'h0; in28=6'h2; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h2; in34=6'h4; in35=6'h0; in36=6'h2; in37=6'h8; in38=6'h0; in39=6'h0; in40=6'h2; in41=6'h0; in42=6'h5; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h1; in51=6'h0; in52=6'h7; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h4; in65=6'h0; in66=6'h1; in67=6'h0; in68=6'h0; in69=6'h9; in70=6'h0; in71=6'hB; in72=6'h0; in73=6'h8; in74=6'h1; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h7; in79=6'hA; in80=6'h9;
      #50 in1=6'h0; in2=6'h0; in3=6'h2; in4=6'h0; in5=6'h2; in6=6'h0; in7=6'h0; in8=6'h2; in9=6'h3; in10=6'h0; in11=6'h0; in12=6'h1; in13=6'h0; in14=6'h2; in15=6'h0; in16=6'h0; in17=6'h9; in18=6'h7; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h3; in23=6'h1; in24=6'h0; in25=6'h7; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h2; in30=6'h9; in31=6'h0; in32=6'h0; in33=6'h3; in34=6'h9; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h3; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h5; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h6; in49=6'h0; in50=6'h0; in51=6'h9; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h5; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h1; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h8; in70=6'h0; in71=6'h9; in72=6'h3; in73=6'h0; in74=6'h0; in75=6'h6; in76=6'h0; in77=6'h0; in78=6'h2; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h1; in3=6'h0; in4=6'h0; in5=6'h3; in6=6'h0; in7=6'h7; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h3; in15=6'h0; in16=6'h3; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h3; in21=6'h2; in22=6'h0; in23=6'h3; in24=6'h5; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h7; in29=6'h0; in30=6'h1; in31=6'h0; in32=6'hC; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h2; in37=6'h8; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h4; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h8; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h1; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h4; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'hE; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'hA; in71=6'h0; in72=6'hC; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h2; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h2;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h5; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h2; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h5; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h1; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h3; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h5; in42=6'hC; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h2; in50=6'h0; in51=6'h0; in52=6'h6; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h1; in57=6'h0; in58=6'h0; in59=6'h1; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h8; in65=6'h2; in66=6'h3; in67=6'h0; in68=6'h0; in69=6'h3; in70=6'h0; in71=6'h4; in72=6'h0; in73=6'h6; in74=6'h2; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h1; in79=6'h6; in80=6'h6;
      #50 in1=6'h0; in2=6'h4; in3=6'h0; in4=6'h0; in5=6'h1; in6=6'h0; in7=6'h3; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h3; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h5; in21=6'h2; in22=6'h0; in23=6'h6; in24=6'h6; in25=6'h0; in26=6'h1; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h4; in31=6'h0; in32=6'h8; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h4; in38=6'h0; in39=6'h2; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h9; in47=6'h0; in48=6'h0; in49=6'h2; in50=6'h0; in51=6'h1; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h7; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h8; in71=6'h0; in72=6'h9; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h6; in3=6'h0; in4=6'h6; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h5; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h6; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h7; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h9; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h9; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h3; in42=6'h7; in43=6'h6; in44=6'h0; in45=6'h1; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h1; in53=6'h0; in54=6'h4; in55=6'h0; in56=6'h3; in57=6'h4; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h6; in62=6'h0; in63=6'h2; in64=6'h0; in65=6'h5; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h5; in6=6'h0; in7=6'h5; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h5; in21=6'h5; in22=6'h0; in23=6'h5; in24=6'h6; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h2; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h9; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h7; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h9; in47=6'h0; in48=6'h0; in49=6'h3; in50=6'h0; in51=6'h0; in52=6'h0; in53=6'h1; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h6; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'hA; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'hA; in71=6'h0; in72=6'hA; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h3; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h3;
      #50 in1=6'h0; in2=6'h0; in3=6'h7; in4=6'h0; in5=6'h4; in6=6'hD; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h1; in11=6'h5; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h2; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h9; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h5; in29=6'h3; in30=6'h2; in31=6'h1; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h4; in40=6'h0; in41=6'h1; in42=6'h0; in43=6'h2; in44=6'h8; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h1; in51=6'h0; in52=6'h0; in53=6'hA; in54=6'h1; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h2; in61=6'h0; in62=6'h6; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h5; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h1; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h5; in5=6'h7; in6=6'h2; in7=6'h0; in8=6'h9; in9=6'h0; in10=6'h4; in11=6'h0; in12=6'h0; in13=6'h7; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h1; in20=6'h8; in21=6'h0; in22=6'hA; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h8; in41=6'hC; in42=6'h0; in43=6'h0; in44=6'h4; in45=6'h0; in46=6'h1; in47=6'h2; in48=6'h0; in49=6'h5; in50=6'h0; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'hB; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h4; in62=6'h1; in63=6'h0; in64=6'hA; in65=6'h0; in66=6'h1; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h6; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h8; in3=6'h0; in4=6'h9; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h9; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h5; in16=6'h8; in17=6'h0; in18=6'h0; in19=6'h2; in20=6'h2; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h8; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'hA; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h7; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h1; in40=6'h0; in41=6'h3; in42=6'h4; in43=6'h8; in44=6'h0; in45=6'h4; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h5; in53=6'h2; in54=6'h6; in55=6'h0; in56=6'h5; in57=6'h2; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h4; in62=6'h0; in63=6'h7; in64=6'h0; in65=6'h5; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h6; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h2; in7=6'h0; in8=6'h0; in9=6'hB; in10=6'h0; in11=6'h6; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h6; in21=6'h4; in22=6'h3; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h8; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h9; in36=6'h0; in37=6'h4; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h1; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h5; in47=6'h0; in48=6'h0; in49=6'h2; in50=6'h3; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h8; in59=6'h7; in60=6'h0; in61=6'h0; in62=6'h1; in63=6'h0; in64=6'h0; in65=6'h1; in66=6'h1; in67=6'h0; in68=6'h6; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h9; in74=6'h6; in75=6'h0; in76=6'h0; in77=6'h2; in78=6'h7; in79=6'h0; in80=6'h4;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h8; in6=6'h0; in7=6'h4; in8=6'h0; in9=6'h3; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h5; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h7; in21=6'h3; in22=6'h0; in23=6'h5; in24=6'h8; in25=6'h0; in26=6'h2; in27=6'h0; in28=6'h1; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h7; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h6; in37=6'hD; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h5; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h9; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h0; in53=6'h1; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h4; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'hB; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'hC; in71=6'h0; in72=6'h4; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h3; in77=6'h0; in78=6'h1; in79=6'h0; in80=6'hB;
      #50 in1=6'h6; in2=6'h0; in3=6'h0; in4=6'h5; in5=6'h1; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h5; in17=6'h0; in18=6'h0; in19=6'h6; in20=6'h0; in21=6'h0; in22=6'h3; in23=6'h0; in24=6'h0; in25=6'h5; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h6; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h6; in39=6'h0; in40=6'h1; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h5; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h8; in56=6'h4; in57=6'h1; in58=6'h0; in59=6'h0; in60=6'h2; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h4; in66=6'h0; in67=6'h5; in68=6'h0; in69=6'h1; in70=6'h0; in71=6'h0; in72=6'h3; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h6; in77=6'h0; in78=6'h1; in79=6'h0; in80=6'h0;
      #50 in1=6'h2; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h1; in7=6'h0; in8=6'h2; in9=6'h4; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h1; in17=6'h1; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h2; in24=6'h0; in25=6'h2; in26=6'h0; in27=6'h2; in28=6'h0; in29=6'h1; in30=6'h3; in31=6'h0; in32=6'h0; in33=6'h2; in34=6'h4; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h1; in40=6'h1; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h2; in50=6'h2; in51=6'h3; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h1; in58=6'h0; in59=6'h0; in60=6'h2; in61=6'h0; in62=6'h3; in63=6'h0; in64=6'h2; in65=6'h0; in66=6'h0; in67=6'h1; in68=6'h1; in69=6'h4; in70=6'h0; in71=6'h4; in72=6'h0; in73=6'h1; in74=6'h0; in75=6'h4; in76=6'h0; in77=6'h0; in78=6'h2; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'hA; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h1; in10=6'hB; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h5; in17=6'h0; in18=6'h0; in19=6'h8; in20=6'h0; in21=6'h0; in22=6'h3; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h8; in42=6'h8; in43=6'h0; in44=6'h0; in45=6'h3; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h9; in53=6'h3; in54=6'hA; in55=6'h0; in56=6'h9; in57=6'h7; in58=6'h0; in59=6'h5; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h5; in64=6'h4; in65=6'h0; in66=6'h7; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h1; in72=6'h0; in73=6'h8; in74=6'h9; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h6; in80=6'h0;
      #50 in1=6'h7; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h2; in6=6'h0; in7=6'h4; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h1; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h2; in22=6'h1; in23=6'h0; in24=6'h0; in25=6'h5; in26=6'h0; in27=6'h0; in28=6'h1; in29=6'h3; in30=6'h5; in31=6'h5; in32=6'h0; in33=6'h0; in34=6'h5; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h6; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h7; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h4; in56=6'h0; in57=6'h1; in58=6'h0; in59=6'h0; in60=6'h6; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h3; in66=6'h0; in67=6'h5; in68=6'h0; in69=6'h1; in70=6'h0; in71=6'h0; in72=6'h7; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h3; in77=6'h0; in78=6'h3; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h5; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h7; in10=6'h0; in11=6'hA; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h5; in21=6'hC; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h5; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h6; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h6; in47=6'h0; in48=6'h0; in49=6'h1; in50=6'h1; in51=6'h0; in52=6'h0; in53=6'h1; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h3; in59=6'h4; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h6; in69=6'h0; in70=6'h0; in71=6'h1; in72=6'h0; in73=6'h3; in74=6'h3; in75=6'h0; in76=6'h0; in77=6'h5; in78=6'h5; in79=6'h0; in80=6'h4;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h4; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h2; in11=6'h0; in12=6'h0; in13=6'h1; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'hA; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h6; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h2; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h5; in47=6'h5; in48=6'h0; in49=6'h2; in50=6'h2; in51=6'h6; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h2; in58=6'h2; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h9; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h2; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h1; in72=6'h0; in73=6'h0; in74=6'h2; in75=6'h3; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h1; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h2; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h2; in13=6'h3; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h4; in18=6'h4; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h1; in23=6'h3; in24=6'h0; in25=6'h4; in26=6'h0; in27=6'h1; in28=6'h0; in29=6'h0; in30=6'h4; in31=6'h0; in32=6'h0; in33=6'h1; in34=6'h7; in35=6'h0; in36=6'h1; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h3; in45=6'h0; in46=6'h1; in47=6'h3; in48=6'h3; in49=6'h0; in50=6'h0; in51=6'h4; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h1; in58=6'h0; in59=6'h0; in60=6'h4; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h5; in70=6'h0; in71=6'h4; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h4; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h1; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h1; in9=6'h1; in10=6'h0; in11=6'h0; in12=6'h5; in13=6'h0; in14=6'h4; in15=6'h0; in16=6'h0; in17=6'hA; in18=6'h8; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h1; in23=6'h2; in24=6'h0; in25=6'h9; in26=6'h3; in27=6'h0; in28=6'h0; in29=6'h4; in30=6'h9; in31=6'h1; in32=6'h0; in33=6'h5; in34=6'h6; in35=6'h0; in36=6'h4; in37=6'h0; in38=6'h1; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h6; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h6; in49=6'h0; in50=6'h0; in51=6'hA; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h7; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'hA; in70=6'h0; in71=6'h8; in72=6'h3; in73=6'h0; in74=6'h0; in75=6'h9; in76=6'h0; in77=6'h0; in78=6'h1; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h5; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h8; in9=6'h0; in10=6'h3; in11=6'h0; in12=6'h0; in13=6'h3; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'hA; in21=6'h0; in22=6'h7; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h8; in41=6'h9; in42=6'h4; in43=6'h0; in44=6'h2; in45=6'h0; in46=6'h2; in47=6'h0; in48=6'h0; in49=6'h5; in50=6'h0; in51=6'h0; in52=6'h0; in53=6'h1; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h8; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'hC; in62=6'h0; in63=6'h0; in64=6'hB; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h4; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h6; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h6; in4=6'h0; in5=6'h3; in6=6'h9; in7=6'h1; in8=6'h0; in9=6'h0; in10=6'h1; in11=6'h1; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h4; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h6; in30=6'h2; in31=6'h6; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h1; in40=6'h0; in41=6'h1; in42=6'h0; in43=6'h3; in44=6'h5; in45=6'h3; in46=6'h2; in47=6'h0; in48=6'h0; in49=6'h1; in50=6'h3; in51=6'h0; in52=6'h0; in53=6'h5; in54=6'h2; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h5; in61=6'h0; in62=6'h6; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h5; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h7; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h7; in7=6'h0; in8=6'h6; in9=6'h0; in10=6'h2; in11=6'h0; in12=6'h0; in13=6'h5; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h2; in21=6'h0; in22=6'h0; in23=6'h6; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h5; in28=6'h0; in29=6'h1; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h1; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h1; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h4; in45=6'h5; in46=6'h4; in47=6'h4; in48=6'h0; in49=6'h4; in50=6'h5; in51=6'h4; in52=6'h0; in53=6'h0; in54=6'h3; in55=6'h0; in56=6'h0; in57=6'h6; in58=6'h2; in59=6'h0; in60=6'h5; in61=6'h0; in62=6'h9; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h4; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h5; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h6; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h9; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h7; in14=6'h0; in15=6'h1; in16=6'h1; in17=6'h1; in18=6'h0; in19=6'h0; in20=6'h7; in21=6'h0; in22=6'hA; in23=6'h2; in24=6'h1; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h1; in40=6'hA; in41=6'h8; in42=6'h8; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h1; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h2; in51=6'h2; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h4; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h6; in62=6'h0; in63=6'h0; in64=6'h6; in65=6'h2; in66=6'h4; in67=6'h0; in68=6'h6; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h8; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h5; in2=6'h1; in3=6'h0; in4=6'h3; in5=6'h1; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h1; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h3; in17=6'h0; in18=6'h0; in19=6'h6; in20=6'h0; in21=6'h2; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h2; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h2; in33=6'h0; in34=6'h1; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h2; in39=6'h2; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h1; in46=6'h1; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h5; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h5; in56=6'h2; in57=6'h1; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h5; in66=6'h0; in67=6'h4; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h5; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h2; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h1; in3=6'h0; in4=6'h0; in5=6'h2; in6=6'h0; in7=6'h8; in8=6'h0; in9=6'h2; in10=6'h0; in11=6'h0; in12=6'h3; in13=6'h0; in14=6'h5; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h2; in19=6'h0; in20=6'h4; in21=6'h0; in22=6'h0; in23=6'h4; in24=6'hC; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h3; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'hC; in33=6'h0; in34=6'h0; in35=6'h1; in36=6'hB; in37=6'hA; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h7; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h5; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h1; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h4; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'hD; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'hA; in71=6'h1; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h8;
      #50 in1=6'h0; in2=6'h0; in3=6'h2; in4=6'h0; in5=6'h0; in6=6'h1; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h9; in13=6'h0; in14=6'h7; in15=6'h0; in16=6'h0; in17=6'hA; in18=6'h9; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h5; in24=6'h0; in25=6'h7; in26=6'h0; in27=6'h2; in28=6'h0; in29=6'h3; in30=6'hA; in31=6'h0; in32=6'h0; in33=6'h6; in34=6'h4; in35=6'h0; in36=6'h9; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h6; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h8; in49=6'h0; in50=6'h0; in51=6'hA; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h9; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'hB; in70=6'h0; in71=6'h8; in72=6'h2; in73=6'h0; in74=6'h0; in75=6'hB; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'hC; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h6; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h2; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h7; in23=6'h0; in24=6'h0; in25=6'h3; in26=6'h1; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h2; in34=6'h5; in35=6'h0; in36=6'h0; in37=6'h7; in38=6'h0; in39=6'h0; in40=6'h1; in41=6'h0; in42=6'h6; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h6; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h5; in65=6'h1; in66=6'h2; in67=6'h0; in68=6'h0; in69=6'hA; in70=6'h0; in71=6'hB; in72=6'h0; in73=6'hA; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h8; in79=6'hA; in80=6'h7;
      #50 in1=6'h7; in2=6'h0; in3=6'h0; in4=6'h2; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h3; in17=6'h0; in18=6'h0; in19=6'h5; in20=6'h0; in21=6'h0; in22=6'h3; in23=6'h0; in24=6'h0; in25=6'h6; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h1; in30=6'h5; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h6; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h7; in39=6'h0; in40=6'h0; in41=6'h1; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h4; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h7; in56=6'h2; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h3; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h4; in66=6'h0; in67=6'h5; in68=6'h0; in69=6'h2; in70=6'h0; in71=6'h0; in72=6'h3; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h5; in77=6'h0; in78=6'h3; in79=6'h0; in80=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h9; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h4; in15=6'h2; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h3; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h2; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h6; in38=6'h0; in39=6'h0; in40=6'h1; in41=6'h0; in42=6'h8; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h9; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h7; in65=6'h1; in66=6'h5; in67=6'h0; in68=6'h0; in69=6'h7; in70=6'h0; in71=6'h8; in72=6'h0; in73=6'hC; in74=6'h3; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h4; in79=6'h9; in80=6'h7;
   end
endmodule