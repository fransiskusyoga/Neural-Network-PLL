module test_tb();
   reg [8:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36;
   wire [10:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   test_top TopModule(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   initial begin
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h1C; in15=9'h0; in16=9'hD; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h1E; in29=9'h0; in30=9'h0; in31=9'h44; in32=9'h0; in33=9'h0; in34=9'h39; in35=9'h4F; in36=9'h45;
      #50 in1=9'h15; in2=9'h0; in3=9'h14; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h6; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h48; in13=9'h0; in14=9'h48; in15=9'h0; in16=9'h16; in17=9'h0; in18=9'h2B; in19=9'h0; in20=9'h45; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'hB; in29=9'h0; in30=9'h0; in31=9'h41; in32=9'h34; in33=9'h0; in34=9'h12; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h49; in3=9'h0; in4=9'h60; in5=9'h38; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h27; in12=9'h4; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h7; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h1F; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h2; in35=9'h0; in36=9'h11;
      #50 in1=9'h0; in2=9'hA; in3=9'h0; in4=9'h14; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h1; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h8; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h43; in29=9'h0; in30=9'h0; in31=9'h18; in32=9'h0; in33=9'h0; in34=9'hA; in35=9'h32; in36=9'h31;
      #50 in1=9'h0; in2=9'h3E; in3=9'h0; in4=9'h32; in5=9'h18; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h30; in12=9'h1F; in13=9'h0; in14=9'h0; in15=9'hF; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h5; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'hF; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h2; in11=9'h4B; in12=9'h0; in13=9'h2D; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h31; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h1C; in22=9'h0; in23=9'h0; in24=9'h14; in25=9'h22; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h24; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h4A; in3=9'h0; in4=9'h51; in5=9'h25; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h32; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h14; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h3; in35=9'h0; in36=9'h17;
      #50 in1=9'h1E; in2=9'h14; in3=9'h3C; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h28; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h12; in13=9'h36; in14=9'h0; in15=9'h1F; in16=9'h0; in17=9'hD; in18=9'h3E; in19=9'h0; in20=9'h0; in21=9'hC; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h33; in28=9'h0; in29=9'h0; in30=9'h27; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h38; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h43; in17=9'h0; in18=9'h22; in19=9'h11; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h56; in26=9'h4; in27=9'hA; in28=9'h52; in29=9'h15; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h3A; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h2B; in11=9'h3E; in12=9'h0; in13=9'h30; in14=9'h0; in15=9'h7; in16=9'h0; in17=9'h3F; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h30; in22=9'h0; in23=9'h0; in24=9'h26; in25=9'hD; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h17; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h2C; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h3D; in27=9'h8; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'hE; in34=9'h36; in35=9'h0; in36=9'h21;
      #50 in1=9'h0; in2=9'h18; in3=9'h0; in4=9'h17; in5=9'h21; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h40; in12=9'h0; in13=9'h14; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h35; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'hC; in35=9'h0; in36=9'h56;
      #50 in1=9'h15; in2=9'h6; in3=9'h0; in4=9'h1C; in5=9'h0; in6=9'h3; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h28; in13=9'h0; in14=9'h32; in15=9'h0; in16=9'h6; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h40; in23=9'h0; in24=9'h1E; in25=9'h6; in26=9'h0; in27=9'h0; in28=9'h2; in29=9'h0; in30=9'h2B; in31=9'h6; in32=9'h0; in33=9'h0; in34=9'hB; in35=9'h0; in36=9'h0;
      #50 in1=9'h4; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h3; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h19; in13=9'h0; in14=9'h1D; in15=9'h7; in16=9'h8; in17=9'h0; in18=9'h3; in19=9'h0; in20=9'h16; in21=9'h0; in22=9'h0; in23=9'h2; in24=9'h0; in25=9'hC; in26=9'h0; in27=9'h17; in28=9'h13; in29=9'h0; in30=9'h6; in31=9'h21; in32=9'h1E; in33=9'h0; in34=9'hE; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h1; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h51; in22=9'h0; in23=9'h0; in24=9'h4A; in25=9'h3C; in26=9'h0; in27=9'h0; in28=9'h1D; in29=9'h0; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h32; in36=9'h0;
      #50 in1=9'h36; in2=9'h10; in3=9'h0; in4=9'h15; in5=9'h20; in6=9'h33; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h2A; in13=9'h0; in14=9'h29; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h20; in23=9'h0; in24=9'h0; in25=9'h5; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h2B; in31=9'h6; in32=9'h0; in33=9'h0; in34=9'h18; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h14; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h22; in7=9'h50; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h30; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h1A; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h25; in34=9'h25; in35=9'h0; in36=9'h1D;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h9; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h29; in20=9'h2D; in21=9'h1; in22=9'h0; in23=9'hF; in24=9'h0; in25=9'h12; in26=9'h11; in27=9'h4B; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h0; in32=9'h1C; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h15; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h14; in9=9'h18; in10=9'h0; in11=9'h0; in12=9'h22; in13=9'h0; in14=9'h35; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h17; in19=9'h15; in20=9'h1F; in21=9'h0; in22=9'h0; in23=9'h31; in24=9'h0; in25=9'hA; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h25; in32=9'h23; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h27; in2=9'h0; in3=9'hB; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h28; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h4C; in13=9'h0; in14=9'h33; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h31; in19=9'h0; in20=9'h54; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h52; in32=9'h4A; in33=9'h0; in34=9'h9; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h16; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'h42; in17=9'h0; in18=9'h13; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h41; in26=9'h0; in27=9'h0; in28=9'h54; in29=9'h44; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h24; in2=9'h2C; in3=9'h31; in4=9'h1; in5=9'hA; in6=9'h0; in7=9'h8; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h10; in13=9'h10; in14=9'h0; in15=9'h6; in16=9'h0; in17=9'h1A; in18=9'h27; in19=9'h0; in20=9'h0; in21=9'h11; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h4; in27=9'h33; in28=9'h0; in29=9'h0; in30=9'h29; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h2A; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h7; in16=9'h0; in17=9'h0; in18=9'h1E; in19=9'h1D; in20=9'h21; in21=9'h18; in22=9'h0; in23=9'h27; in24=9'h0; in25=9'h32; in26=9'h12; in27=9'h49; in28=9'h4; in29=9'h0; in30=9'h0; in31=9'h0; in32=9'h2B; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h38; in10=9'h6; in11=9'h6; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h4; in16=9'h50; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h13; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h23; in26=9'h0; in27=9'h0; in28=9'h30; in29=9'h54; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'hA; in2=9'h1F; in3=9'h0; in4=9'h29; in5=9'h0; in6=9'h2; in7=9'h2; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h1; in13=9'h0; in14=9'h6; in15=9'hD; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h24; in23=9'h0; in24=9'hF; in25=9'hC; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h22; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h11; in5=9'h3D; in6=9'h0; in7=9'h0; in8=9'h17; in9=9'h0; in10=9'h0; in11=9'h5E; in12=9'h0; in13=9'h2E; in14=9'h0; in15=9'h0; in16=9'h0; in17=9'h2; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h2B; in30=9'h0; in31=9'h0; in32=9'h0; in33=9'h0; in34=9'h2; in35=9'h0; in36=9'h3E;
      #50 in1=9'h2E; in2=9'h0; in3=9'h13; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h45; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h54; in13=9'h0; in14=9'h1C; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h32; in19=9'h0; in20=9'h50; in21=9'h0; in22=9'h0; in23=9'h11; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h0; in31=9'h59; in32=9'h55; in33=9'h0; in34=9'h0; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h25; in15=9'h0; in16=9'h9; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h2; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h2C; in29=9'h0; in30=9'h0; in31=9'h51; in32=9'h0; in33=9'h0; in34=9'h42; in35=9'h4E; in36=9'h38;
      #50 in1=9'h13; in2=9'h6; in3=9'h0; in4=9'h1F; in5=9'h0; in6=9'h12; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h0; in11=9'h0; in12=9'h28; in13=9'h0; in14=9'h32; in15=9'h0; in16=9'h0; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h3B; in23=9'h0; in24=9'h13; in25=9'h1; in26=9'h0; in27=9'h0; in28=9'h0; in29=9'h0; in30=9'h27; in31=9'hC; in32=9'h0; in33=9'h0; in34=9'h19; in35=9'h0; in36=9'h0;
      #50 in1=9'h0; in2=9'h0; in3=9'h0; in4=9'h0; in5=9'h0; in6=9'h0; in7=9'h0; in8=9'h0; in9=9'h0; in10=9'h12; in11=9'h0; in12=9'h0; in13=9'h0; in14=9'h0; in15=9'h0; in16=9'hA; in17=9'h0; in18=9'h0; in19=9'h0; in20=9'h0; in21=9'h0; in22=9'h0; in23=9'h0; in24=9'h0; in25=9'h0; in26=9'h0; in27=9'h0; in28=9'h39; in29=9'h0; in30=9'h0; in31=9'h36; in32=9'h0; in33=9'h0; in34=9'h24; in35=9'h45; in36=9'h3A;
   end
endmodule