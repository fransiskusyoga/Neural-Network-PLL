module lenet5_top(clk,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   input clk;
   input [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381;
   output [9:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   wire signed [9:0] s2_1,s2_2,s2_3,s2_4,s2_5,s2_6,s2_7,s2_8,s2_9,s2_10,s2_11,s2_12,s2_13,s2_14,s2_15,s2_16,s2_17,s2_18,s2_19,s2_20,s2_21,s2_22,s2_23,s2_24,s2_25,s2_26,s2_27,s2_28,s2_29,s2_30,s2_31,s2_32,s2_33,s2_34,s2_35,s2_36,s2_37,s2_38,s2_39,s2_40,s2_41,s2_42,s2_43,s2_44,s2_45,s2_46,s2_47,s2_48,s2_49,s2_50,s2_51,s2_52,s2_53,s2_54,s2_55,s2_56,s2_57,s2_58,s2_59,s2_60,s2_61,s2_62,s2_63,s2_64,s2_65,s2_66,s2_67,s2_68,s2_69,s2_70,s2_71,s2_72,s2_73,s2_74,s2_75,s2_76,s2_77,s2_78,s2_79,s2_80,s2_81,s2_82,s2_83,s2_84,s2_85,s2_86,s2_87,s2_88,s2_89,s2_90,s2_91,s2_92,s2_93,s2_94,s2_95,s2_96,s2_97,s2_98,s2_99,s2_100,s2_101,s2_102,s2_103,s2_104,s2_105,s2_106,s2_107,s2_108,s2_109,s2_110,s2_111,s2_112,s2_113,s2_114,s2_115,s2_116,s2_117;
   wire signed [9:0] s3_1,s3_2,s3_3,s3_4,s3_5,s3_6,s3_7,s3_8,s3_9,s3_10,s3_11,s3_12,s3_13,s3_14,s3_15,s3_16,s3_17,s3_18,s3_19,s3_20,s3_21,s3_22,s3_23,s3_24,s3_25,s3_26,s3_27,s3_28,s3_29,s3_30,s3_31,s3_32,s3_33,s3_34,s3_35,s3_36,s3_37,s3_38,s3_39,s3_40,s3_41,s3_42,s3_43,s3_44,s3_45,s3_46,s3_47,s3_48,s3_49,s3_50,s3_51,s3_52,s3_53,s3_54,s3_55,s3_56,s3_57,s3_58,s3_59,s3_60,s3_61,s3_62,s3_63,s3_64,s3_65,s3_66,s3_67,s3_68,s3_69,s3_70,s3_71,s3_72,s3_73,s3_74,s3_75,s3_76,s3_77,s3_78,s3_79,s3_80,s3_81;
   wire signed [9:0] h2_1,h2_2,h2_3,h2_4,h2_5,h2_6,h2_7,h2_8,h2_9,h2_10,h2_11,h2_12,h2_13,h2_14,h2_15,h2_16,h2_17,h2_18,h2_19,h2_20,h2_21,h2_22,h2_23,h2_24,h2_25,h2_26,h2_27,h2_28,h2_29,h2_30,h2_31,h2_32,h2_33,h2_34,h2_35,h2_36,h2_37,h2_38,h2_39,h2_40,h2_41,h2_42,h2_43,h2_44,h2_45,h2_46,h2_47,h2_48,h2_49,h2_50,h2_51,h2_52,h2_53,h2_54,h2_55,h2_56,h2_57,h2_58,h2_59,h2_60,h2_61,h2_62,h2_63,h2_64,h2_65,h2_66,h2_67,h2_68,h2_69,h2_70,h2_71,h2_72,h2_73,h2_74,h2_75,h2_76,h2_77,h2_78,h2_79,h2_80,h2_81,h2_82,h2_83,h2_84,h2_85,h2_86,h2_87,h2_88,h2_89,h2_90,h2_91,h2_92,h2_93,h2_94,h2_95,h2_96,h2_97,h2_98,h2_99,h2_100,h2_101,h2_102,h2_103,h2_104,h2_105,h2_106,h2_107,h2_108,h2_109,h2_110,h2_111,h2_112,h2_113,h2_114,h2_115,h2_116,h2_117;
   wire signed [9:0] h3_1,h3_2,h3_3,h3_4,h3_5,h3_6,h3_7,h3_8,h3_9,h3_10,h3_11,h3_12,h3_13,h3_14,h3_15,h3_16,h3_17,h3_18,h3_19,h3_20,h3_21,h3_22,h3_23,h3_24,h3_25,h3_26,h3_27,h3_28,h3_29,h3_30,h3_31,h3_32,h3_33,h3_34,h3_35,h3_36,h3_37,h3_38,h3_39,h3_40,h3_41,h3_42,h3_43,h3_44,h3_45,h3_46,h3_47,h3_48,h3_49,h3_50,h3_51,h3_52,h3_53,h3_54,h3_55,h3_56,h3_57,h3_58,h3_59,h3_60,h3_61,h3_62,h3_63,h3_64,h3_65,h3_66,h3_67,h3_68,h3_69,h3_70,h3_71,h3_72,h3_73,h3_74,h3_75,h3_76,h3_77,h3_78,h3_79,h3_80,h3_81;
   lenet5_layer_1 L1(clk,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,s2_1,s2_2,s2_3,s2_4,s2_5,s2_6,s2_7,s2_8,s2_9,s2_10,s2_11,s2_12,s2_13,s2_14,s2_15,s2_16,s2_17,s2_18,s2_19,s2_20,s2_21,s2_22,s2_23,s2_24,s2_25,s2_26,s2_27,s2_28,s2_29,s2_30,s2_31,s2_32,s2_33,s2_34,s2_35,s2_36,s2_37,s2_38,s2_39,s2_40,s2_41,s2_42,s2_43,s2_44,s2_45,s2_46,s2_47,s2_48,s2_49,s2_50,s2_51,s2_52,s2_53,s2_54,s2_55,s2_56,s2_57,s2_58,s2_59,s2_60,s2_61,s2_62,s2_63,s2_64,s2_65,s2_66,s2_67,s2_68,s2_69,s2_70,s2_71,s2_72,s2_73,s2_74,s2_75,s2_76,s2_77,s2_78,s2_79,s2_80,s2_81,s2_82,s2_83,s2_84,s2_85,s2_86,s2_87,s2_88,s2_89,s2_90,s2_91,s2_92,s2_93,s2_94,s2_95,s2_96,s2_97,s2_98,s2_99,s2_100,s2_101,s2_102,s2_103,s2_104,s2_105,s2_106,s2_107,s2_108,s2_109,s2_110,s2_111,s2_112,s2_113,s2_114,s2_115,s2_116,s2_117);
   actifunc #(10) AF2_1(s2_1,h2_1);
   actifunc #(10) AF2_2(s2_2,h2_2);
   actifunc #(10) AF2_3(s2_3,h2_3);
   actifunc #(10) AF2_4(s2_4,h2_4);
   actifunc #(10) AF2_5(s2_5,h2_5);
   actifunc #(10) AF2_6(s2_6,h2_6);
   actifunc #(10) AF2_7(s2_7,h2_7);
   actifunc #(10) AF2_8(s2_8,h2_8);
   actifunc #(10) AF2_9(s2_9,h2_9);
   actifunc #(10) AF2_10(s2_10,h2_10);
   actifunc #(10) AF2_11(s2_11,h2_11);
   actifunc #(10) AF2_12(s2_12,h2_12);
   actifunc #(10) AF2_13(s2_13,h2_13);
   actifunc #(10) AF2_14(s2_14,h2_14);
   actifunc #(10) AF2_15(s2_15,h2_15);
   actifunc #(10) AF2_16(s2_16,h2_16);
   actifunc #(10) AF2_17(s2_17,h2_17);
   actifunc #(10) AF2_18(s2_18,h2_18);
   actifunc #(10) AF2_19(s2_19,h2_19);
   actifunc #(10) AF2_20(s2_20,h2_20);
   actifunc #(10) AF2_21(s2_21,h2_21);
   actifunc #(10) AF2_22(s2_22,h2_22);
   actifunc #(10) AF2_23(s2_23,h2_23);
   actifunc #(10) AF2_24(s2_24,h2_24);
   actifunc #(10) AF2_25(s2_25,h2_25);
   actifunc #(10) AF2_26(s2_26,h2_26);
   actifunc #(10) AF2_27(s2_27,h2_27);
   actifunc #(10) AF2_28(s2_28,h2_28);
   actifunc #(10) AF2_29(s2_29,h2_29);
   actifunc #(10) AF2_30(s2_30,h2_30);
   actifunc #(10) AF2_31(s2_31,h2_31);
   actifunc #(10) AF2_32(s2_32,h2_32);
   actifunc #(10) AF2_33(s2_33,h2_33);
   actifunc #(10) AF2_34(s2_34,h2_34);
   actifunc #(10) AF2_35(s2_35,h2_35);
   actifunc #(10) AF2_36(s2_36,h2_36);
   actifunc #(10) AF2_37(s2_37,h2_37);
   actifunc #(10) AF2_38(s2_38,h2_38);
   actifunc #(10) AF2_39(s2_39,h2_39);
   actifunc #(10) AF2_40(s2_40,h2_40);
   actifunc #(10) AF2_41(s2_41,h2_41);
   actifunc #(10) AF2_42(s2_42,h2_42);
   actifunc #(10) AF2_43(s2_43,h2_43);
   actifunc #(10) AF2_44(s2_44,h2_44);
   actifunc #(10) AF2_45(s2_45,h2_45);
   actifunc #(10) AF2_46(s2_46,h2_46);
   actifunc #(10) AF2_47(s2_47,h2_47);
   actifunc #(10) AF2_48(s2_48,h2_48);
   actifunc #(10) AF2_49(s2_49,h2_49);
   actifunc #(10) AF2_50(s2_50,h2_50);
   actifunc #(10) AF2_51(s2_51,h2_51);
   actifunc #(10) AF2_52(s2_52,h2_52);
   actifunc #(10) AF2_53(s2_53,h2_53);
   actifunc #(10) AF2_54(s2_54,h2_54);
   actifunc #(10) AF2_55(s2_55,h2_55);
   actifunc #(10) AF2_56(s2_56,h2_56);
   actifunc #(10) AF2_57(s2_57,h2_57);
   actifunc #(10) AF2_58(s2_58,h2_58);
   actifunc #(10) AF2_59(s2_59,h2_59);
   actifunc #(10) AF2_60(s2_60,h2_60);
   actifunc #(10) AF2_61(s2_61,h2_61);
   actifunc #(10) AF2_62(s2_62,h2_62);
   actifunc #(10) AF2_63(s2_63,h2_63);
   actifunc #(10) AF2_64(s2_64,h2_64);
   actifunc #(10) AF2_65(s2_65,h2_65);
   actifunc #(10) AF2_66(s2_66,h2_66);
   actifunc #(10) AF2_67(s2_67,h2_67);
   actifunc #(10) AF2_68(s2_68,h2_68);
   actifunc #(10) AF2_69(s2_69,h2_69);
   actifunc #(10) AF2_70(s2_70,h2_70);
   actifunc #(10) AF2_71(s2_71,h2_71);
   actifunc #(10) AF2_72(s2_72,h2_72);
   actifunc #(10) AF2_73(s2_73,h2_73);
   actifunc #(10) AF2_74(s2_74,h2_74);
   actifunc #(10) AF2_75(s2_75,h2_75);
   actifunc #(10) AF2_76(s2_76,h2_76);
   actifunc #(10) AF2_77(s2_77,h2_77);
   actifunc #(10) AF2_78(s2_78,h2_78);
   actifunc #(10) AF2_79(s2_79,h2_79);
   actifunc #(10) AF2_80(s2_80,h2_80);
   actifunc #(10) AF2_81(s2_81,h2_81);
   actifunc #(10) AF2_82(s2_82,h2_82);
   actifunc #(10) AF2_83(s2_83,h2_83);
   actifunc #(10) AF2_84(s2_84,h2_84);
   actifunc #(10) AF2_85(s2_85,h2_85);
   actifunc #(10) AF2_86(s2_86,h2_86);
   actifunc #(10) AF2_87(s2_87,h2_87);
   actifunc #(10) AF2_88(s2_88,h2_88);
   actifunc #(10) AF2_89(s2_89,h2_89);
   actifunc #(10) AF2_90(s2_90,h2_90);
   actifunc #(10) AF2_91(s2_91,h2_91);
   actifunc #(10) AF2_92(s2_92,h2_92);
   actifunc #(10) AF2_93(s2_93,h2_93);
   actifunc #(10) AF2_94(s2_94,h2_94);
   actifunc #(10) AF2_95(s2_95,h2_95);
   actifunc #(10) AF2_96(s2_96,h2_96);
   actifunc #(10) AF2_97(s2_97,h2_97);
   actifunc #(10) AF2_98(s2_98,h2_98);
   actifunc #(10) AF2_99(s2_99,h2_99);
   actifunc #(10) AF2_100(s2_100,h2_100);
   actifunc #(10) AF2_101(s2_101,h2_101);
   actifunc #(10) AF2_102(s2_102,h2_102);
   actifunc #(10) AF2_103(s2_103,h2_103);
   actifunc #(10) AF2_104(s2_104,h2_104);
   actifunc #(10) AF2_105(s2_105,h2_105);
   actifunc #(10) AF2_106(s2_106,h2_106);
   actifunc #(10) AF2_107(s2_107,h2_107);
   actifunc #(10) AF2_108(s2_108,h2_108);
   actifunc #(10) AF2_109(s2_109,h2_109);
   actifunc #(10) AF2_110(s2_110,h2_110);
   actifunc #(10) AF2_111(s2_111,h2_111);
   actifunc #(10) AF2_112(s2_112,h2_112);
   actifunc #(10) AF2_113(s2_113,h2_113);
   actifunc #(10) AF2_114(s2_114,h2_114);
   actifunc #(10) AF2_115(s2_115,h2_115);
   actifunc #(10) AF2_116(s2_116,h2_116);
   actifunc #(10) AF2_117(s2_117,h2_117);
   lenet5_layer_2 L2(clk,h2_1[9:4],h2_2[9:4],h2_3[9:4],h2_4[9:4],h2_5[9:4],h2_6[9:4],h2_7[9:4],h2_8[9:4],h2_9[9:4],h2_10[9:4],h2_11[9:4],h2_12[9:4],h2_13[9:4],h2_14[9:4],h2_15[9:4],h2_16[9:4],h2_17[9:4],h2_18[9:4],h2_19[9:4],h2_20[9:4],h2_21[9:4],h2_22[9:4],h2_23[9:4],h2_24[9:4],h2_25[9:4],h2_26[9:4],h2_27[9:4],h2_28[9:4],h2_29[9:4],h2_30[9:4],h2_31[9:4],h2_32[9:4],h2_33[9:4],h2_34[9:4],h2_35[9:4],h2_36[9:4],h2_37[9:4],h2_38[9:4],h2_39[9:4],h2_40[9:4],h2_41[9:4],h2_42[9:4],h2_43[9:4],h2_44[9:4],h2_45[9:4],h2_46[9:4],h2_47[9:4],h2_48[9:4],h2_49[9:4],h2_50[9:4],h2_51[9:4],h2_52[9:4],h2_53[9:4],h2_54[9:4],h2_55[9:4],h2_56[9:4],h2_57[9:4],h2_58[9:4],h2_59[9:4],h2_60[9:4],h2_61[9:4],h2_62[9:4],h2_63[9:4],h2_64[9:4],h2_65[9:4],h2_66[9:4],h2_67[9:4],h2_68[9:4],h2_69[9:4],h2_70[9:4],h2_71[9:4],h2_72[9:4],h2_73[9:4],h2_74[9:4],h2_75[9:4],h2_76[9:4],h2_77[9:4],h2_78[9:4],h2_79[9:4],h2_80[9:4],h2_81[9:4],h2_82[9:4],h2_83[9:4],h2_84[9:4],h2_85[9:4],h2_86[9:4],h2_87[9:4],h2_88[9:4],h2_89[9:4],h2_90[9:4],h2_91[9:4],h2_92[9:4],h2_93[9:4],h2_94[9:4],h2_95[9:4],h2_96[9:4],h2_97[9:4],h2_98[9:4],h2_99[9:4],h2_100[9:4],h2_101[9:4],h2_102[9:4],h2_103[9:4],h2_104[9:4],h2_105[9:4],h2_106[9:4],h2_107[9:4],h2_108[9:4],h2_109[9:4],h2_110[9:4],h2_111[9:4],h2_112[9:4],h2_113[9:4],h2_114[9:4],h2_115[9:4],h2_116[9:4],h2_117[9:4],s3_1,s3_2,s3_3,s3_4,s3_5,s3_6,s3_7,s3_8,s3_9,s3_10,s3_11,s3_12,s3_13,s3_14,s3_15,s3_16,s3_17,s3_18,s3_19,s3_20,s3_21,s3_22,s3_23,s3_24,s3_25,s3_26,s3_27,s3_28,s3_29,s3_30,s3_31,s3_32,s3_33,s3_34,s3_35,s3_36,s3_37,s3_38,s3_39,s3_40,s3_41,s3_42,s3_43,s3_44,s3_45,s3_46,s3_47,s3_48,s3_49,s3_50,s3_51,s3_52,s3_53,s3_54,s3_55,s3_56,s3_57,s3_58,s3_59,s3_60,s3_61,s3_62,s3_63,s3_64,s3_65,s3_66,s3_67,s3_68,s3_69,s3_70,s3_71,s3_72,s3_73,s3_74,s3_75,s3_76,s3_77,s3_78,s3_79,s3_80,s3_81);
   actifunc #(10) AF3_1(s3_1,h3_1);
   actifunc #(10) AF3_2(s3_2,h3_2);
   actifunc #(10) AF3_3(s3_3,h3_3);
   actifunc #(10) AF3_4(s3_4,h3_4);
   actifunc #(10) AF3_5(s3_5,h3_5);
   actifunc #(10) AF3_6(s3_6,h3_6);
   actifunc #(10) AF3_7(s3_7,h3_7);
   actifunc #(10) AF3_8(s3_8,h3_8);
   actifunc #(10) AF3_9(s3_9,h3_9);
   actifunc #(10) AF3_10(s3_10,h3_10);
   actifunc #(10) AF3_11(s3_11,h3_11);
   actifunc #(10) AF3_12(s3_12,h3_12);
   actifunc #(10) AF3_13(s3_13,h3_13);
   actifunc #(10) AF3_14(s3_14,h3_14);
   actifunc #(10) AF3_15(s3_15,h3_15);
   actifunc #(10) AF3_16(s3_16,h3_16);
   actifunc #(10) AF3_17(s3_17,h3_17);
   actifunc #(10) AF3_18(s3_18,h3_18);
   actifunc #(10) AF3_19(s3_19,h3_19);
   actifunc #(10) AF3_20(s3_20,h3_20);
   actifunc #(10) AF3_21(s3_21,h3_21);
   actifunc #(10) AF3_22(s3_22,h3_22);
   actifunc #(10) AF3_23(s3_23,h3_23);
   actifunc #(10) AF3_24(s3_24,h3_24);
   actifunc #(10) AF3_25(s3_25,h3_25);
   actifunc #(10) AF3_26(s3_26,h3_26);
   actifunc #(10) AF3_27(s3_27,h3_27);
   actifunc #(10) AF3_28(s3_28,h3_28);
   actifunc #(10) AF3_29(s3_29,h3_29);
   actifunc #(10) AF3_30(s3_30,h3_30);
   actifunc #(10) AF3_31(s3_31,h3_31);
   actifunc #(10) AF3_32(s3_32,h3_32);
   actifunc #(10) AF3_33(s3_33,h3_33);
   actifunc #(10) AF3_34(s3_34,h3_34);
   actifunc #(10) AF3_35(s3_35,h3_35);
   actifunc #(10) AF3_36(s3_36,h3_36);
   actifunc #(10) AF3_37(s3_37,h3_37);
   actifunc #(10) AF3_38(s3_38,h3_38);
   actifunc #(10) AF3_39(s3_39,h3_39);
   actifunc #(10) AF3_40(s3_40,h3_40);
   actifunc #(10) AF3_41(s3_41,h3_41);
   actifunc #(10) AF3_42(s3_42,h3_42);
   actifunc #(10) AF3_43(s3_43,h3_43);
   actifunc #(10) AF3_44(s3_44,h3_44);
   actifunc #(10) AF3_45(s3_45,h3_45);
   actifunc #(10) AF3_46(s3_46,h3_46);
   actifunc #(10) AF3_47(s3_47,h3_47);
   actifunc #(10) AF3_48(s3_48,h3_48);
   actifunc #(10) AF3_49(s3_49,h3_49);
   actifunc #(10) AF3_50(s3_50,h3_50);
   actifunc #(10) AF3_51(s3_51,h3_51);
   actifunc #(10) AF3_52(s3_52,h3_52);
   actifunc #(10) AF3_53(s3_53,h3_53);
   actifunc #(10) AF3_54(s3_54,h3_54);
   actifunc #(10) AF3_55(s3_55,h3_55);
   actifunc #(10) AF3_56(s3_56,h3_56);
   actifunc #(10) AF3_57(s3_57,h3_57);
   actifunc #(10) AF3_58(s3_58,h3_58);
   actifunc #(10) AF3_59(s3_59,h3_59);
   actifunc #(10) AF3_60(s3_60,h3_60);
   actifunc #(10) AF3_61(s3_61,h3_61);
   actifunc #(10) AF3_62(s3_62,h3_62);
   actifunc #(10) AF3_63(s3_63,h3_63);
   actifunc #(10) AF3_64(s3_64,h3_64);
   actifunc #(10) AF3_65(s3_65,h3_65);
   actifunc #(10) AF3_66(s3_66,h3_66);
   actifunc #(10) AF3_67(s3_67,h3_67);
   actifunc #(10) AF3_68(s3_68,h3_68);
   actifunc #(10) AF3_69(s3_69,h3_69);
   actifunc #(10) AF3_70(s3_70,h3_70);
   actifunc #(10) AF3_71(s3_71,h3_71);
   actifunc #(10) AF3_72(s3_72,h3_72);
   actifunc #(10) AF3_73(s3_73,h3_73);
   actifunc #(10) AF3_74(s3_74,h3_74);
   actifunc #(10) AF3_75(s3_75,h3_75);
   actifunc #(10) AF3_76(s3_76,h3_76);
   actifunc #(10) AF3_77(s3_77,h3_77);
   actifunc #(10) AF3_78(s3_78,h3_78);
   actifunc #(10) AF3_79(s3_79,h3_79);
   actifunc #(10) AF3_80(s3_80,h3_80);
   actifunc #(10) AF3_81(s3_81,h3_81);
   lenet5_layer_3 L3(clk,h3_1[9:4],h3_2[9:4],h3_3[9:4],h3_4[9:4],h3_5[9:4],h3_6[9:4],h3_7[9:4],h3_8[9:4],h3_9[9:4],h3_10[9:4],h3_11[9:4],h3_12[9:4],h3_13[9:4],h3_14[9:4],h3_15[9:4],h3_16[9:4],h3_17[9:4],h3_18[9:4],h3_19[9:4],h3_20[9:4],h3_21[9:4],h3_22[9:4],h3_23[9:4],h3_24[9:4],h3_25[9:4],h3_26[9:4],h3_27[9:4],h3_28[9:4],h3_29[9:4],h3_30[9:4],h3_31[9:4],h3_32[9:4],h3_33[9:4],h3_34[9:4],h3_35[9:4],h3_36[9:4],h3_37[9:4],h3_38[9:4],h3_39[9:4],h3_40[9:4],h3_41[9:4],h3_42[9:4],h3_43[9:4],h3_44[9:4],h3_45[9:4],h3_46[9:4],h3_47[9:4],h3_48[9:4],h3_49[9:4],h3_50[9:4],h3_51[9:4],h3_52[9:4],h3_53[9:4],h3_54[9:4],h3_55[9:4],h3_56[9:4],h3_57[9:4],h3_58[9:4],h3_59[9:4],h3_60[9:4],h3_61[9:4],h3_62[9:4],h3_63[9:4],h3_64[9:4],h3_65[9:4],h3_66[9:4],h3_67[9:4],h3_68[9:4],h3_69[9:4],h3_70[9:4],h3_71[9:4],h3_72[9:4],h3_73[9:4],h3_74[9:4],h3_75[9:4],h3_76[9:4],h3_77[9:4],h3_78[9:4],h3_79[9:4],h3_80[9:4],h3_81[9:4],out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
endmodule