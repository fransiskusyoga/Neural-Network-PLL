module lenet5_tb();
   reg [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381;
   wire [9:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   lenet5_top TopModule(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   initial begin
      #50 in1=6'h0; in2=6'h0; in3=6'h9; in4=6'h12; in5=6'hF; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h2; in14=6'h0; in15=6'h0; in16=6'h3; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h1; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h6; in31=6'h1; in32=6'h2; in33=6'h6; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h2; in41=6'h2; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'hC; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h1; in57=6'h0; in58=6'hA; in59=6'hB; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'hA; in65=6'h3; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h1; in70=6'h0; in71=6'h0; in72=6'h3; in73=6'h3; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h6; in78=6'h0; in79=6'h8; in80=6'h0; in81=6'h0; in82=6'h8; in83=6'hA; in84=6'h0; in85=6'h0; in86=6'h4; in87=6'h6; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h4; in92=6'h9; in93=6'h0; in94=6'h0; in95=6'h4; in96=6'h0; in97=6'h5; in98=6'h0; in99=6'h2; in100=6'h3; in101=6'h9; in102=6'h5; in103=6'h0; in104=6'h0; in105=6'h1; in106=6'h2; in107=6'h0; in108=6'h2; in109=6'h0; in110=6'h1; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h2; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h3; in120=6'h0; in121=6'h1; in122=6'hE; in123=6'h5; in124=6'h0; in125=6'h0; in126=6'hA; in127=6'h9; in128=6'hA; in129=6'h3; in130=6'h1; in131=6'h0; in132=6'h5; in133=6'hD; in134=6'h0; in135=6'h0; in136=6'h8; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h1; in141=6'h4; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h8; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h5; in159=6'h1; in160=6'h5; in161=6'h9; in162=6'h2; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h3; in167=6'h1; in168=6'h0; in169=6'h3; in170=6'h0; in171=6'hD; in172=6'h0; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'hE; in177=6'h2; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'h6; in182=6'h4; in183=6'h0; in184=6'h0; in185=6'h4; in186=6'hA; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h2; in191=6'h0; in192=6'h0; in193=6'h6; in194=6'h8; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h2; in199=6'h1; in200=6'h5; in201=6'h0; in202=6'h0; in203=6'h1; in204=6'h1; in205=6'h0; in206=6'h5; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h3; in211=6'h2; in212=6'h3; in213=6'h3; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'hF; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h3; in225=6'h0; in226=6'h4; in227=6'h0; in228=6'h0; in229=6'h4; in230=6'hB; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h2; in236=6'h8; in237=6'h10; in238=6'h5; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h5; in246=6'h1; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h7; in251=6'h3; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h2; in256=6'h4; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h6; in262=6'h5; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h3; in270=6'h2; in271=6'h2; in272=6'h3; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h3; in280=6'hE; in281=6'hD; in282=6'h3; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h8; in292=6'h7; in293=6'h2; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h2; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h2; in316=6'h0; in317=6'h0; in318=6'h2; in319=6'h0; in320=6'h7; in321=6'h3; in322=6'h5; in323=6'h8; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h2; in328=6'h0; in329=6'h0; in330=6'h1; in331=6'h0; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h1; in336=6'h0; in337=6'h0; in338=6'h3; in339=6'h0; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h9; in344=6'h4; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h3; in349=6'h6; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h4; in354=6'h3; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h0; in363=6'h2; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h1; in369=6'h0; in370=6'h6; in371=6'h4; in372=6'h2; in373=6'h0; in374=6'h2; in375=6'h3; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h0; in380=6'h1; in381=6'h1;
      #50 in1=6'h2; in2=6'h3; in3=6'hC; in4=6'h14; in5=6'hC; in6=6'h1; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h2; in13=6'h9; in14=6'h8; in15=6'h2; in16=6'h1; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h1; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h5; in31=6'h0; in32=6'h2; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h2; in42=6'h4; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'hB; in51=6'h9; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h2; in56=6'hA; in57=6'h0; in58=6'h4; in59=6'h0; in60=6'h7; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h4; in66=6'h1; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h3; in73=6'h4; in74=6'h0; in75=6'h0; in76=6'h6; in77=6'hB; in78=6'h0; in79=6'h2; in80=6'h0; in81=6'h3; in82=6'h1; in83=6'h6; in84=6'h3; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h5; in89=6'h0; in90=6'h0; in91=6'h1; in92=6'hA; in93=6'h5; in94=6'h0; in95=6'h2; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h0; in101=6'h5; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h0; in106=6'h2; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h3; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h1; in116=6'h6; in117=6'h5; in118=6'h0; in119=6'h1; in120=6'h0; in121=6'h2; in122=6'hB; in123=6'h0; in124=6'h0; in125=6'h3; in126=6'h13; in127=6'hC; in128=6'h4; in129=6'h0; in130=6'h2; in131=6'h0; in132=6'h0; in133=6'h4; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h9; in138=6'h6; in139=6'h0; in140=6'h0; in141=6'hE; in142=6'hE; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h3; in151=6'h0; in152=6'h6; in153=6'hA; in154=6'h3; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h1; in160=6'h2; in161=6'h1; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h1; in169=6'h0; in170=6'h7; in171=6'hE; in172=6'h0; in173=6'h1; in174=6'h0; in175=6'h7; in176=6'h6; in177=6'h4; in178=6'h8; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h0; in183=6'h1; in184=6'h0; in185=6'h0; in186=6'h2; in187=6'h1; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'hA; in194=6'h6; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h3; in208=6'h0; in209=6'h0; in210=6'h1; in211=6'h0; in212=6'h8; in213=6'h0; in214=6'h5; in215=6'h7; in216=6'h0; in217=6'h6; in218=6'h0; in219=6'h0; in220=6'h12; in221=6'h7; in222=6'h4; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h2; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h3; in237=6'h7; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'hA; in242=6'hD; in243=6'h2; in244=6'h0; in245=6'hE; in246=6'h10; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h6; in251=6'hA; in252=6'h3; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h9; in262=6'h7; in263=6'h2; in264=6'h0; in265=6'h0; in266=6'h1; in267=6'h0; in268=6'h0; in269=6'h2; in270=6'hD; in271=6'hD; in272=6'h1; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h7; in281=6'h1; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h3; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'hA; in301=6'hD; in302=6'h2; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h5; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h3; in321=6'h0; in322=6'h0; in323=6'h1; in324=6'h5; in325=6'h4; in326=6'h0; in327=6'h4; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'h9; in332=6'hA; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h7; in339=6'h0; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h6; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h2; in358=6'h3; in359=6'h1; in360=6'h5; in361=6'h2; in362=6'h0; in363=6'h3; in364=6'h6; in365=6'h1; in366=6'h0; in367=6'h1; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h5; in373=6'h5; in374=6'h3; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h2; in380=6'h2; in381=6'h1;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h3; in5=6'h1; in6=6'h1; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h6; in12=6'h10; in13=6'hE; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h9; in19=6'h2; in20=6'h1; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h1; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h1; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h2; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h1; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h10; in51=6'h7; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h6; in56=6'h8; in57=6'h2; in58=6'h5; in59=6'h8; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h5; in65=6'h6; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h5; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h4; in84=6'h0; in85=6'h0; in86=6'h4; in87=6'hC; in88=6'h8; in89=6'h0; in90=6'h0; in91=6'h5; in92=6'h8; in93=6'h0; in94=6'h0; in95=6'h2; in96=6'h2; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h3; in101=6'h3; in102=6'h0; in103=6'h3; in104=6'h5; in105=6'h0; in106=6'h2; in107=6'h0; in108=6'h7; in109=6'h5; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h1; in120=6'h0; in121=6'h0; in122=6'h3; in123=6'h0; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h7; in132=6'h1; in133=6'h9; in134=6'h0; in135=6'h7; in136=6'h4; in137=6'h6; in138=6'h1; in139=6'h0; in140=6'h1; in141=6'h0; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h1; in146=6'h2; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h1; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h1; in156=6'h0; in157=6'h5; in158=6'h8; in159=6'h2; in160=6'h0; in161=6'h2; in162=6'h3; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h0; in169=6'h0; in170=6'h2; in171=6'h0; in172=6'h0; in173=6'h5; in174=6'h0; in175=6'h7; in176=6'h4; in177=6'h0; in178=6'h5; in179=6'h0; in180=6'h9; in181=6'h1; in182=6'h3; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h3; in199=6'h1; in200=6'h2; in201=6'h0; in202=6'h0; in203=6'h2; in204=6'h0; in205=6'h4; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h0; in212=6'hE; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h3; in218=6'h0; in219=6'h4; in220=6'h1; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h4; in225=6'hA; in226=6'hB; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h3; in232=6'h4; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h2; in237=6'h5; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h1; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h3; in250=6'h7; in251=6'h4; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h6; in256=6'h3; in257=6'h5; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h3; in262=6'h1; in263=6'h0; in264=6'h0; in265=6'h1; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'hA; in276=6'h5; in277=6'h1; in278=6'h0; in279=6'h1; in280=6'h1; in281=6'h2; in282=6'h3; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h1; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h7; in306=6'h3; in307=6'h3; in308=6'h0; in309=6'h3; in310=6'h3; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h4; in315=6'h3; in316=6'h0; in317=6'h2; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h1; in323=6'h5; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h1; in329=6'h1; in330=6'h3; in331=6'h2; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h6; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h6; in341=6'h2; in342=6'h0; in343=6'h2; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h7; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h7; in363=6'h8; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h3; in368=6'hA; in369=6'h3; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h1; in376=6'h0; in377=6'h5; in378=6'h9; in379=6'h9; in380=6'h5; in381=6'h3;
      #50 in1=6'h4; in2=6'hA; in3=6'hC; in4=6'hE; in5=6'hE; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h3; in12=6'hC; in13=6'h12; in14=6'h9; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h9; in19=6'hC; in20=6'h4; in21=6'h0; in22=6'h4; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'hB; in30=6'h9; in31=6'h3; in32=6'h1; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h2; in40=6'h5; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h6; in49=6'h0; in50=6'h0; in51=6'h3; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h1; in58=6'h4; in59=6'hC; in60=6'h5; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h4; in65=6'h15; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h4; in70=6'h2; in71=6'h1; in72=6'h0; in73=6'h7; in74=6'hA; in75=6'h0; in76=6'hC; in77=6'hC; in78=6'hB; in79=6'h5; in80=6'h0; in81=6'h5; in82=6'h4; in83=6'h0; in84=6'h0; in85=6'h4; in86=6'h7; in87=6'h9; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'hA; in93=6'hE; in94=6'h0; in95=6'h0; in96=6'h5; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h0; in101=6'h4; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h2; in106=6'h0; in107=6'h0; in108=6'h0; in109=6'h2; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h1; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h1; in121=6'h7; in122=6'h5; in123=6'hA; in124=6'h6; in125=6'h8; in126=6'hB; in127=6'h2; in128=6'h0; in129=6'h0; in130=6'h2; in131=6'h0; in132=6'h0; in133=6'h0; in134=6'h0; in135=6'h4; in136=6'h0; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h1; in141=6'h4; in142=6'h2; in143=6'h5; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h6; in149=6'h6; in150=6'h1; in151=6'h0; in152=6'h8; in153=6'h5; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h4; in158=6'h3; in159=6'h4; in160=6'h0; in161=6'h7; in162=6'h5; in163=6'h0; in164=6'h0; in165=6'h8; in166=6'h4; in167=6'h0; in168=6'h0; in169=6'h0; in170=6'hF; in171=6'h0; in172=6'h0; in173=6'h0; in174=6'h0; in175=6'hD; in176=6'h0; in177=6'h0; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h0; in183=6'h1; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h3; in190=6'h1; in191=6'h0; in192=6'h3; in193=6'h7; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h2; in198=6'h3; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h6; in210=6'h6; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'hA; in220=6'h5; in221=6'h9; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h3; in226=6'hE; in227=6'h8; in228=6'h0; in229=6'h0; in230=6'hD; in231=6'h9; in232=6'h0; in233=6'h0; in234=6'h2; in235=6'h3; in236=6'h5; in237=6'h9; in238=6'h8; in239=6'h0; in240=6'h8; in241=6'hB; in242=6'h9; in243=6'h5; in244=6'h3; in245=6'h5; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h6; in250=6'hA; in251=6'h7; in252=6'h1; in253=6'h0; in254=6'h0; in255=6'h5; in256=6'h4; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h1; in261=6'h6; in262=6'h9; in263=6'h7; in264=6'h0; in265=6'h7; in266=6'hC; in267=6'h4; in268=6'h0; in269=6'h7; in270=6'hA; in271=6'h4; in272=6'h0; in273=6'h0; in274=6'h2; in275=6'h2; in276=6'h4; in277=6'h3; in278=6'h0; in279=6'h2; in280=6'h5; in281=6'hB; in282=6'h5; in283=6'h2; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h2; in291=6'hB; in292=6'h9; in293=6'h6; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h6; in300=6'h6; in301=6'h4; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h0; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h3; in315=6'h2; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h0; in323=6'h0; in324=6'h1; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'h1; in330=6'h0; in331=6'h0; in332=6'h0; in333=6'h0; in334=6'h3; in335=6'h0; in336=6'h0; in337=6'h5; in338=6'h3; in339=6'h0; in340=6'h0; in341=6'h0; in342=6'hA; in343=6'h8; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h4; in349=6'h0; in350=6'h6; in351=6'h0; in352=6'h0; in353=6'h5; in354=6'h1; in355=6'h1; in356=6'h0; in357=6'h0; in358=6'h1; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h5; in363=6'hB; in364=6'h11; in365=6'hD; in366=6'h9; in367=6'h0; in368=6'h5; in369=6'hF; in370=6'h6; in371=6'h0; in372=6'h4; in373=6'h9; in374=6'h6; in375=6'h3; in376=6'h1; in377=6'h1; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h1; in2=6'h3; in3=6'h1; in4=6'h2; in5=6'h1; in6=6'h0; in7=6'h0; in8=6'h1; in9=6'h0; in10=6'h0; in11=6'h2; in12=6'hE; in13=6'h10; in14=6'h8; in15=6'h2; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h8; in30=6'h4; in31=6'h0; in32=6'h2; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h1; in41=6'h4; in42=6'hC; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h3; in47=6'h6; in48=6'h7; in49=6'h0; in50=6'hB; in51=6'h9; in52=6'h1; in53=6'h2; in54=6'h0; in55=6'h4; in56=6'h8; in57=6'h0; in58=6'h6; in59=6'h0; in60=6'h0; in61=6'h3; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h1; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h2; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h3; in81=6'h3; in82=6'h0; in83=6'h5; in84=6'h3; in85=6'h2; in86=6'h3; in87=6'h2; in88=6'h5; in89=6'h1; in90=6'h0; in91=6'h0; in92=6'h0; in93=6'h1; in94=6'h0; in95=6'h0; in96=6'hA; in97=6'h2; in98=6'h3; in99=6'hB; in100=6'h4; in101=6'hF; in102=6'h0; in103=6'h7; in104=6'hE; in105=6'h0; in106=6'h0; in107=6'h0; in108=6'h3; in109=6'h5; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h1; in114=6'h0; in115=6'h2; in116=6'h2; in117=6'h3; in118=6'hB; in119=6'h0; in120=6'h0; in121=6'h2; in122=6'h0; in123=6'h0; in124=6'h2; in125=6'h4; in126=6'h6; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h2; in131=6'h0; in132=6'h0; in133=6'h2; in134=6'h0; in135=6'h1; in136=6'h0; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h0; in142=6'h5; in143=6'h4; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h4; in151=6'h1; in152=6'hB; in153=6'hA; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h2; in158=6'h4; in159=6'h0; in160=6'h0; in161=6'h0; in162=6'h2; in163=6'h2; in164=6'h0; in165=6'h5; in166=6'h0; in167=6'h0; in168=6'h8; in169=6'h0; in170=6'h10; in171=6'h0; in172=6'h0; in173=6'hB; in174=6'h0; in175=6'hB; in176=6'h0; in177=6'h0; in178=6'h9; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h0; in183=6'hB; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'hA; in188=6'h4; in189=6'h2; in190=6'h0; in191=6'h0; in192=6'h3; in193=6'h6; in194=6'h0; in195=6'h0; in196=6'h1; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h1; in201=6'h1; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h3; in210=6'h0; in211=6'h0; in212=6'h5; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h4; in218=6'h0; in219=6'h11; in220=6'hA; in221=6'h2; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h1; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h1; in235=6'h0; in236=6'h0; in237=6'h1; in238=6'h0; in239=6'h1; in240=6'h0; in241=6'h0; in242=6'h2; in243=6'h0; in244=6'h7; in245=6'hB; in246=6'h2; in247=6'h2; in248=6'h0; in249=6'h5; in250=6'hE; in251=6'hE; in252=6'h7; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h2; in267=6'h0; in268=6'h0; in269=6'h6; in270=6'hD; in271=6'hB; in272=6'h5; in273=6'h2; in274=6'h0; in275=6'h5; in276=6'h5; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h0; in281=6'h2; in282=6'h1; in283=6'h2; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h3; in300=6'h9; in301=6'hE; in302=6'h7; in303=6'h1; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h0; in311=6'h0; in312=6'h3; in313=6'h0; in314=6'h4; in315=6'h5; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h0; in323=6'h1; in324=6'h3; in325=6'h1; in326=6'h0; in327=6'h3; in328=6'h3; in329=6'h5; in330=6'h7; in331=6'h1; in332=6'hA; in333=6'h3; in334=6'h0; in335=6'h0; in336=6'h2; in337=6'h7; in338=6'h7; in339=6'h0; in340=6'h4; in341=6'h5; in342=6'h5; in343=6'hA; in344=6'h0; in345=6'h4; in346=6'h5; in347=6'h0; in348=6'h0; in349=6'h0; in350=6'h3; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h3; in356=6'h0; in357=6'h5; in358=6'h5; in359=6'h0; in360=6'h5; in361=6'h3; in362=6'h0; in363=6'h2; in364=6'h1; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h5; in373=6'h5; in374=6'h7; in375=6'h4; in376=6'h0; in377=6'h4; in378=6'h4; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h4; in2=6'h12; in3=6'h15; in4=6'hC; in5=6'h3; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h3; in10=6'h1; in11=6'h0; in12=6'h3; in13=6'h7; in14=6'h6; in15=6'hA; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h1; in30=6'h1; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h6; in41=6'h0; in42=6'hB; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h9; in50=6'h11; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'hF; in56=6'h2; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h3; in61=6'h7; in62=6'h0; in63=6'h2; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h2; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h6; in72=6'h4; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h4; in83=6'h6; in84=6'h6; in85=6'h0; in86=6'h5; in87=6'h1; in88=6'h5; in89=6'h6; in90=6'h0; in91=6'h5; in92=6'h8; in93=6'h5; in94=6'h0; in95=6'h0; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h1; in100=6'h1; in101=6'h0; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h1; in106=6'h6; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'h5; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h9; in121=6'h7; in122=6'h0; in123=6'h0; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'hE; in132=6'hC; in133=6'h4; in134=6'h0; in135=6'h1; in136=6'hA; in137=6'h5; in138=6'h7; in139=6'h0; in140=6'h1; in141=6'h0; in142=6'h5; in143=6'h0; in144=6'h0; in145=6'h2; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h3; in150=6'h2; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h2; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h2; in160=6'h5; in161=6'h9; in162=6'h1; in163=6'h0; in164=6'h0; in165=6'h1; in166=6'h0; in167=6'h1; in168=6'h2; in169=6'h0; in170=6'h1; in171=6'h0; in172=6'h0; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'h3; in177=6'h0; in178=6'h7; in179=6'h0; in180=6'hA; in181=6'hD; in182=6'h0; in183=6'h2; in184=6'h0; in185=6'h7; in186=6'h1; in187=6'h1; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h1; in197=6'h0; in198=6'h0; in199=6'h1; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h9; in204=6'h5; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h7; in211=6'h11; in212=6'h5; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'hD; in218=6'h0; in219=6'h0; in220=6'h3; in221=6'h0; in222=6'h5; in223=6'h2; in224=6'h5; in225=6'h8; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h10; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h7; in235=6'hA; in236=6'h8; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h8; in242=6'h4; in243=6'h0; in244=6'h0; in245=6'h1; in246=6'hA; in247=6'h8; in248=6'h4; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h3; in253=6'h6; in254=6'h0; in255=6'h9; in256=6'h3; in257=6'h0; in258=6'h0; in259=6'h3; in260=6'h3; in261=6'h3; in262=6'h2; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h1; in268=6'h0; in269=6'h0; in270=6'h4; in271=6'h3; in272=6'h0; in273=6'h5; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h4; in280=6'hA; in281=6'hA; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h3; in290=6'h4; in291=6'h3; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h1; in301=6'h3; in302=6'h3; in303=6'h5; in304=6'h0; in305=6'h3; in306=6'h2; in307=6'h0; in308=6'h0; in309=6'h0; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'hB; in315=6'h5; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h4; in320=6'h0; in321=6'h0; in322=6'h0; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h6; in328=6'h1; in329=6'h0; in330=6'h1; in331=6'h2; in332=6'hC; in333=6'h5; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'hA; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h3; in346=6'h0; in347=6'h0; in348=6'h8; in349=6'h0; in350=6'h1; in351=6'h0; in352=6'h0; in353=6'h7; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h4; in360=6'h3; in361=6'h0; in362=6'h7; in363=6'h6; in364=6'h3; in365=6'h4; in366=6'h4; in367=6'h2; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'hC; in380=6'h7; in381=6'h2;
      #50 in1=6'h0; in2=6'h0; in3=6'hD; in4=6'hA; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h2; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h2; in17=6'h4; in18=6'h7; in19=6'h11; in20=6'h10; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h2; in29=6'h0; in30=6'h2; in31=6'h0; in32=6'h6; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h7; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h4; in45=6'h1; in46=6'h1; in47=6'h0; in48=6'h0; in49=6'hA; in50=6'h13; in51=6'h0; in52=6'h0; in53=6'h1; in54=6'h0; in55=6'hA; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h2; in64=6'h0; in65=6'h3; in66=6'h4; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h2; in71=6'h0; in72=6'h5; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h2; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h1; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'hB; in88=6'hD; in89=6'h0; in90=6'h0; in91=6'h7; in92=6'h9; in93=6'h5; in94=6'h2; in95=6'h2; in96=6'h3; in97=6'h0; in98=6'h0; in99=6'h2; in100=6'h0; in101=6'h4; in102=6'h0; in103=6'h7; in104=6'h1; in105=6'h3; in106=6'h0; in107=6'h0; in108=6'h9; in109=6'h0; in110=6'h3; in111=6'h0; in112=6'h1; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h5; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h0; in121=6'hF; in122=6'h7; in123=6'h0; in124=6'h0; in125=6'h2; in126=6'h6; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h0; in133=6'h2; in134=6'h0; in135=6'h0; in136=6'h6; in137=6'hD; in138=6'h0; in139=6'h0; in140=6'h3; in141=6'h9; in142=6'h5; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h1; in148=6'h4; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h2; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h0; in160=6'h2; in161=6'h9; in162=6'h4; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h7; in167=6'h0; in168=6'h2; in169=6'h0; in170=6'h0; in171=6'hC; in172=6'h4; in173=6'h8; in174=6'h0; in175=6'h0; in176=6'h0; in177=6'h10; in178=6'hC; in179=6'h0; in180=6'h0; in181=6'h2; in182=6'h10; in183=6'h3; in184=6'h0; in185=6'h0; in186=6'h3; in187=6'h0; in188=6'h0; in189=6'h1; in190=6'h7; in191=6'h0; in192=6'h0; in193=6'h3; in194=6'h1; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h4; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h5; in205=6'h4; in206=6'h1; in207=6'h2; in208=6'h0; in209=6'h0; in210=6'h1; in211=6'h8; in212=6'h8; in213=6'h0; in214=6'h0; in215=6'h6; in216=6'h0; in217=6'h7; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h2; in226=6'h0; in227=6'h9; in228=6'h3; in229=6'h0; in230=6'h7; in231=6'h0; in232=6'h0; in233=6'h1; in234=6'h1; in235=6'h0; in236=6'h5; in237=6'h1; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h1; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h2; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h1; in252=6'h6; in253=6'h3; in254=6'h1; in255=6'h4; in256=6'h4; in257=6'hE; in258=6'hB; in259=6'h0; in260=6'h1; in261=6'h0; in262=6'h1; in263=6'h0; in264=6'h3; in265=6'h4; in266=6'h4; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h1; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h9; in278=6'hC; in279=6'h4; in280=6'h7; in281=6'h4; in282=6'h3; in283=6'h2; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h1; in295=6'h3; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h4; in306=6'h1; in307=6'h3; in308=6'h7; in309=6'h1; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h7; in316=6'h0; in317=6'h1; in318=6'h0; in319=6'h5; in320=6'h8; in321=6'h0; in322=6'h5; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h3; in331=6'h7; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h3; in337=6'h0; in338=6'h3; in339=6'h0; in340=6'h8; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h7; in346=6'h0; in347=6'h0; in348=6'h3; in349=6'h0; in350=6'h5; in351=6'h0; in352=6'h0; in353=6'h3; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h0; in363=6'h1; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h7; in368=6'h9; in369=6'h3; in370=6'h5; in371=6'h0; in372=6'h2; in373=6'h2; in374=6'h0; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h2; in379=6'h3; in380=6'h6; in381=6'h8;
      #50 in1=6'h0; in2=6'h4; in3=6'hB; in4=6'hD; in5=6'h9; in6=6'h1; in7=6'h1; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h5; in12=6'h0; in13=6'h2; in14=6'hC; in15=6'h8; in16=6'hF; in17=6'h10; in18=6'h6; in19=6'h0; in20=6'h2; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h7; in32=6'hB; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h2; in45=6'h2; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h3; in50=6'h6; in51=6'h6; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h2; in57=6'h4; in58=6'h0; in59=6'h0; in60=6'hE; in61=6'h1; in62=6'h5; in63=6'h5; in64=6'h0; in65=6'h7; in66=6'h5; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h2; in74=6'h1; in75=6'h0; in76=6'h0; in77=6'h1; in78=6'hA; in79=6'h5; in80=6'h0; in81=6'h2; in82=6'hA; in83=6'h8; in84=6'h0; in85=6'h1; in86=6'h3; in87=6'h0; in88=6'h7; in89=6'h3; in90=6'h1; in91=6'h6; in92=6'hC; in93=6'hD; in94=6'h0; in95=6'h2; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h1; in100=6'h2; in101=6'h0; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h0; in106=6'h0; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h0; in121=6'h1; in122=6'h8; in123=6'h3; in124=6'h1; in125=6'h0; in126=6'h7; in127=6'h2; in128=6'h5; in129=6'h0; in130=6'h0; in131=6'h8; in132=6'h6; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h1; in138=6'h8; in139=6'h0; in140=6'h1; in141=6'h0; in142=6'h5; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h1; in149=6'h6; in150=6'h3; in151=6'h0; in152=6'h0; in153=6'h7; in154=6'hB; in155=6'h7; in156=6'h0; in157=6'h4; in158=6'h0; in159=6'h5; in160=6'h4; in161=6'h3; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h3; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'h0; in173=6'h1; in174=6'h0; in175=6'h0; in176=6'h0; in177=6'h3; in178=6'h0; in179=6'h0; in180=6'h1; in181=6'h0; in182=6'h0; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h1; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h2; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h3; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h3; in221=6'h8; in222=6'h12; in223=6'h0; in224=6'h13; in225=6'h7; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h7; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h1; in236=6'hC; in237=6'h9; in238=6'h0; in239=6'h0; in240=6'h5; in241=6'hA; in242=6'h5; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h3; in247=6'h1; in248=6'h0; in249=6'h2; in250=6'h0; in251=6'h6; in252=6'h7; in253=6'h1; in254=6'hA; in255=6'hC; in256=6'h6; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h6; in261=6'hB; in262=6'h1; in263=6'h0; in264=6'h0; in265=6'h3; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'hA; in271=6'hD; in272=6'h4; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h3; in280=6'hC; in281=6'hB; in282=6'h1; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h2; in290=6'h5; in291=6'h3; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h3; in301=6'h8; in302=6'h0; in303=6'h1; in304=6'h2; in305=6'hE; in306=6'hE; in307=6'h4; in308=6'h1; in309=6'h2; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h2; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'h0; in332=6'h7; in333=6'h2; in334=6'h0; in335=6'h1; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h2; in340=6'h2; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h1; in348=6'h0; in349=6'h0; in350=6'h3; in351=6'h0; in352=6'h0; in353=6'h1; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h0; in363=6'h7; in364=6'h7; in365=6'h0; in366=6'h0; in367=6'h7; in368=6'h0; in369=6'h0; in370=6'h6; in371=6'h1; in372=6'h1; in373=6'hC; in374=6'hB; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h3; in379=6'hF; in380=6'hE; in381=6'h3;
      #50 in1=6'h0; in2=6'h0; in3=6'hA; in4=6'hD; in5=6'h4; in6=6'h0; in7=6'h0; in8=6'h4; in9=6'h0; in10=6'h6; in11=6'h4; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h2; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h4; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h6; in31=6'h7; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h7; in37=6'h4; in38=6'h0; in39=6'h0; in40=6'h3; in41=6'h9; in42=6'h3; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h8; in51=6'h6; in52=6'h0; in53=6'h0; in54=6'hB; in55=6'h0; in56=6'h7; in57=6'h0; in58=6'h0; in59=6'h6; in60=6'h1; in61=6'h0; in62=6'h0; in63=6'h5; in64=6'h4; in65=6'hB; in66=6'h0; in67=6'h1; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'hE; in73=6'h4; in74=6'h0; in75=6'h0; in76=6'h3; in77=6'h4; in78=6'h0; in79=6'h2; in80=6'h0; in81=6'h0; in82=6'h9; in83=6'h10; in84=6'hD; in85=6'h0; in86=6'h5; in87=6'h5; in88=6'h0; in89=6'h0; in90=6'h1; in91=6'h5; in92=6'hA; in93=6'h3; in94=6'h0; in95=6'h2; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h1; in101=6'h0; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h1; in106=6'h0; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'hA; in112=6'h0; in113=6'h2; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h2; in120=6'h0; in121=6'hA; in122=6'hB; in123=6'h0; in124=6'h0; in125=6'h2; in126=6'h3; in127=6'h0; in128=6'h8; in129=6'hD; in130=6'h0; in131=6'hC; in132=6'h5; in133=6'hB; in134=6'h1; in135=6'h2; in136=6'hB; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h1; in141=6'h0; in142=6'h3; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h9; in149=6'h3; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h2; in155=6'h0; in156=6'h0; in157=6'h1; in158=6'h0; in159=6'h7; in160=6'h8; in161=6'hA; in162=6'h4; in163=6'h2; in164=6'h0; in165=6'h0; in166=6'hC; in167=6'h0; in168=6'h0; in169=6'h4; in170=6'h0; in171=6'hA; in172=6'h0; in173=6'h0; in174=6'h2; in175=6'h1; in176=6'h2; in177=6'h3; in178=6'h0; in179=6'h0; in180=6'h10; in181=6'hA; in182=6'h5; in183=6'h0; in184=6'h0; in185=6'h9; in186=6'h0; in187=6'h4; in188=6'h0; in189=6'h0; in190=6'h7; in191=6'h0; in192=6'h0; in193=6'h1; in194=6'h1; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h1; in199=6'h1; in200=6'h1; in201=6'h0; in202=6'h1; in203=6'h9; in204=6'h1; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h3; in211=6'h2; in212=6'h4; in213=6'h0; in214=6'h0; in215=6'h12; in216=6'hA; in217=6'h0; in218=6'h0; in219=6'h1; in220=6'h0; in221=6'h4; in222=6'h0; in223=6'h0; in224=6'h8; in225=6'h7; in226=6'h6; in227=6'h0; in228=6'h0; in229=6'h3; in230=6'h13; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h1; in236=6'h0; in237=6'h2; in238=6'h0; in239=6'h0; in240=6'h1; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h4; in247=6'h2; in248=6'h2; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h2; in255=6'h8; in256=6'h6; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h1; in262=6'h6; in263=6'h0; in264=6'h2; in265=6'h1; in266=6'h0; in267=6'h0; in268=6'h2; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h2; in273=6'h2; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h6; in280=6'hE; in281=6'hC; in282=6'h4; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h1; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h4; in298=6'h5; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h0; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h1; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h0; in323=6'h1; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h4; in328=6'h3; in329=6'h0; in330=6'h0; in331=6'h2; in332=6'h7; in333=6'h0; in334=6'h6; in335=6'h1; in336=6'h0; in337=6'h0; in338=6'h5; in339=6'hC; in340=6'h0; in341=6'h1; in342=6'h0; in343=6'h0; in344=6'hA; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'hA; in349=6'h8; in350=6'h8; in351=6'h0; in352=6'h0; in353=6'h9; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h4; in361=6'h9; in362=6'h0; in363=6'h3; in364=6'h5; in365=6'h5; in366=6'h0; in367=6'h1; in368=6'h0; in369=6'h0; in370=6'hA; in371=6'hA; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h3; in376=6'h2; in377=6'h0; in378=6'h0; in379=6'h4; in380=6'h0; in381=6'h1;
      #50 in1=6'h0; in2=6'h0; in3=6'h8; in4=6'h11; in5=6'hF; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h1; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h1; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h4; in32=6'h0; in33=6'h3; in34=6'h0; in35=6'h3; in36=6'h0; in37=6'h0; in38=6'h1; in39=6'h9; in40=6'h4; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h2; in50=6'h6; in51=6'h11; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h10; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h1; in62=6'h3; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h1; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h7; in74=6'h1; in75=6'h0; in76=6'h0; in77=6'h7; in78=6'h5; in79=6'h0; in80=6'h0; in81=6'h4; in82=6'h4; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h3; in87=6'h0; in88=6'h7; in89=6'h6; in90=6'h3; in91=6'h7; in92=6'hE; in93=6'h9; in94=6'h0; in95=6'h4; in96=6'h2; in97=6'h5; in98=6'h2; in99=6'h0; in100=6'h4; in101=6'h6; in102=6'hB; in103=6'h0; in104=6'h3; in105=6'h0; in106=6'h10; in107=6'hA; in108=6'h0; in109=6'h8; in110=6'hB; in111=6'h13; in112=6'h0; in113=6'h7; in114=6'h7; in115=6'h4; in116=6'h0; in117=6'h0; in118=6'h2; in119=6'h0; in120=6'h0; in121=6'h0; in122=6'hE; in123=6'hD; in124=6'h1; in125=6'h0; in126=6'h7; in127=6'hB; in128=6'h1; in129=6'h0; in130=6'h0; in131=6'h8; in132=6'h0; in133=6'h1; in134=6'h8; in135=6'h4; in136=6'h3; in137=6'h4; in138=6'hE; in139=6'h3; in140=6'h1; in141=6'h4; in142=6'hF; in143=6'h0; in144=6'h0; in145=6'h1; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h1; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h1; in160=6'hE; in161=6'hA; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h5; in168=6'h0; in169=6'h3; in170=6'h0; in171=6'h9; in172=6'h8; in173=6'h0; in174=6'h4; in175=6'h6; in176=6'hB; in177=6'h0; in178=6'h5; in179=6'h9; in180=6'h11; in181=6'h7; in182=6'h0; in183=6'h7; in184=6'h0; in185=6'hE; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h1; in191=6'h4; in192=6'h0; in193=6'h0; in194=6'h6; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h7; in199=6'h5; in200=6'h0; in201=6'h2; in202=6'h3; in203=6'h7; in204=6'h0; in205=6'h4; in206=6'h2; in207=6'h0; in208=6'h2; in209=6'h0; in210=6'h0; in211=6'h4; in212=6'h4; in213=6'h9; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'hF; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'hB; in230=6'h6; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h3; in236=6'h5; in237=6'h6; in238=6'h1; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'hB; in243=6'h5; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h2; in255=6'h7; in256=6'h1; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h3; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h9; in280=6'h11; in281=6'h9; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h1; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h3; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'hA; in317=6'h6; in318=6'h0; in319=6'h0; in320=6'h9; in321=6'h11; in322=6'h3; in323=6'h6; in324=6'h6; in325=6'hC; in326=6'h3; in327=6'h1; in328=6'hB; in329=6'h2; in330=6'h0; in331=6'h0; in332=6'h9; in333=6'h8; in334=6'h0; in335=6'h1; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h0; in341=6'h6; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h3; in347=6'h6; in348=6'h1; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h9; in353=6'h9; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h2; in362=6'h0; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h1; in370=6'h0; in371=6'h0; in372=6'h2; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h5; in380=6'h8; in381=6'h2;
      #50 in1=6'h1; in2=6'h7; in3=6'h15; in4=6'h10; in5=6'h3; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h1; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h1; in31=6'h1; in32=6'h8; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h4; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h4; in42=6'h2; in43=6'h0; in44=6'h0; in45=6'h4; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h5; in50=6'hE; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h10; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h5; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h2; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h2; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h4; in77=6'h4; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h3; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h2; in93=6'h1; in94=6'h0; in95=6'h0; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h2; in100=6'h0; in101=6'h0; in102=6'h0; in103=6'h3; in104=6'h1; in105=6'h2; in106=6'h2; in107=6'h0; in108=6'hC; in109=6'h0; in110=6'h4; in111=6'h4; in112=6'hE; in113=6'hE; in114=6'h0; in115=6'h4; in116=6'h0; in117=6'hE; in118=6'h3; in119=6'h2; in120=6'h0; in121=6'h9; in122=6'h7; in123=6'h0; in124=6'h0; in125=6'h4; in126=6'hB; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h0; in133=6'h3; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h6; in138=6'h3; in139=6'h0; in140=6'h0; in141=6'h0; in142=6'h5; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h1; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h0; in160=6'h0; in161=6'h4; in162=6'h4; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'h0; in173=6'h6; in174=6'h0; in175=6'h0; in176=6'h0; in177=6'hB; in178=6'h9; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'hE; in183=6'h5; in184=6'h0; in185=6'h0; in186=6'h5; in187=6'hF; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h1; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h2; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h2; in205=6'h5; in206=6'h0; in207=6'h6; in208=6'h3; in209=6'h3; in210=6'h0; in211=6'h7; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h3; in217=6'hA; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h2; in231=6'h5; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h3; in237=6'h0; in238=6'h0; in239=6'h2; in240=6'h9; in241=6'hD; in242=6'h4; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h5; in261=6'h5; in262=6'h1; in263=6'h0; in264=6'h5; in265=6'h8; in266=6'h3; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h0; in281=6'h2; in282=6'h1; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h4; in290=6'h9; in291=6'h7; in292=6'h3; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h1; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h1; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h4; in320=6'hA; in321=6'h0; in322=6'h5; in323=6'h2; in324=6'h1; in325=6'h1; in326=6'h0; in327=6'h8; in328=6'h2; in329=6'h0; in330=6'h0; in331=6'hB; in332=6'h8; in333=6'h0; in334=6'h1; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h6; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h4; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h2; in355=6'h0; in356=6'h0; in357=6'h2; in358=6'h3; in359=6'h6; in360=6'h4; in361=6'h0; in362=6'h0; in363=6'h5; in364=6'h0; in365=6'h1; in366=6'h0; in367=6'h8; in368=6'h9; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h1; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h0; in377=6'h1; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h1;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h1; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h1; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h4; in32=6'h4; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h5; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h3; in41=6'h5; in42=6'h0; in43=6'h0; in44=6'h4; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h8; in51=6'h1; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h3; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h2; in83=6'h2; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h1; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h3; in92=6'h1; in93=6'h0; in94=6'h0; in95=6'h2; in96=6'h4; in97=6'h0; in98=6'hC; in99=6'h2; in100=6'h4; in101=6'h4; in102=6'hE; in103=6'hE; in104=6'h0; in105=6'h4; in106=6'h0; in107=6'h11; in108=6'h7; in109=6'h2; in110=6'h4; in111=6'h7; in112=6'h10; in113=6'h0; in114=6'h3; in115=6'h1; in116=6'hA; in117=6'h8; in118=6'h1; in119=6'h3; in120=6'h0; in121=6'h0; in122=6'h0; in123=6'h7; in124=6'h1; in125=6'h0; in126=6'h0; in127=6'h5; in128=6'h5; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h4; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h3; in137=6'h3; in138=6'h0; in139=6'h0; in140=6'h1; in141=6'h5; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h0; in160=6'h0; in161=6'h8; in162=6'h6; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h5; in168=6'h9; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'hE; in173=6'h7; in174=6'h0; in175=6'h0; in176=6'h5; in177=6'hF; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'hF; in182=6'hB; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'hA; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h5; in192=6'h0; in193=6'h0; in194=6'h1; in195=6'h6; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h5; in200=6'h3; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h6; in205=6'h0; in206=6'h0; in207=6'h2; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h2; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h1; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h1; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h4; in280=6'h6; in281=6'h5; in282=6'h1; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h1; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h3; in311=6'h1; in312=6'h0; in313=6'h1; in314=6'h1; in315=6'h0; in316=6'h0; in317=6'hA; in318=6'h3; in319=6'h0; in320=6'h0; in321=6'hA; in322=6'hB; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'hB; in327=6'h7; in328=6'h0; in329=6'h0; in330=6'h8; in331=6'hB; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h1; in349=6'h2; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h2; in354=6'h1; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h1; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h1; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h1; in377=6'h0; in378=6'h1; in379=6'h0; in380=6'h1; in381=6'h1;
      #50 in1=6'h1; in2=6'h2; in3=6'h8; in4=6'hC; in5=6'h5; in6=6'h2; in7=6'h0; in8=6'h0; in9=6'h3; in10=6'h4; in11=6'h0; in12=6'h0; in13=6'h2; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h4; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h2; in31=6'h0; in32=6'h1; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'hB; in42=6'h5; in43=6'h0; in44=6'h0; in45=6'h4; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'hC; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'hF; in56=6'h7; in57=6'h0; in58=6'h0; in59=6'h2; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h2; in65=6'h1; in66=6'h0; in67=6'h0; in68=6'h2; in69=6'h1; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h8; in77=6'h9; in78=6'h5; in79=6'h0; in80=6'h3; in81=6'h3; in82=6'h3; in83=6'h9; in84=6'h3; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h3; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h4; in93=6'h0; in94=6'h0; in95=6'h3; in96=6'h0; in97=6'h0; in98=6'h1; in99=6'h0; in100=6'h0; in101=6'h3; in102=6'h1; in103=6'h0; in104=6'h0; in105=6'h0; in106=6'h2; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'h0; in112=6'h1; in113=6'h1; in114=6'h0; in115=6'h1; in116=6'h0; in117=6'h5; in118=6'h0; in119=6'h2; in120=6'h0; in121=6'h0; in122=6'hA; in123=6'h7; in124=6'h2; in125=6'h0; in126=6'hE; in127=6'h10; in128=6'h0; in129=6'h0; in130=6'h6; in131=6'h1; in132=6'h0; in133=6'h9; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h1; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h2; in142=6'h5; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h2; in150=6'h4; in151=6'h0; in152=6'h8; in153=6'h9; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h1; in158=6'h3; in159=6'h2; in160=6'h0; in161=6'h6; in162=6'hC; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h7; in169=6'h0; in170=6'h5; in171=6'h8; in172=6'h0; in173=6'h4; in174=6'h0; in175=6'hC; in176=6'h7; in177=6'h5; in178=6'h6; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h7; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h5; in187=6'hD; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h1; in192=6'h0; in193=6'hA; in194=6'h6; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h5; in199=6'h0; in200=6'h1; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h3; in208=6'h0; in209=6'h0; in210=6'h3; in211=6'h0; in212=6'h4; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'hA; in218=6'h0; in219=6'hB; in220=6'h8; in221=6'h2; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h2; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h9; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h1; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h8; in242=6'h2; in243=6'h2; in244=6'h1; in245=6'hB; in246=6'hA; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h10; in251=6'h6; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h1; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h2; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h4; in266=6'h7; in267=6'h0; in268=6'h0; in269=6'h4; in270=6'hF; in271=6'hA; in272=6'h0; in273=6'h0; in274=6'h1; in275=6'h3; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h4; in281=6'hB; in282=6'h9; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h2; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h3; in300=6'hB; in301=6'h6; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h5; in310=6'h5; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h2; in323=6'h3; in324=6'h2; in325=6'h0; in326=6'h4; in327=6'h7; in328=6'h4; in329=6'h2; in330=6'h0; in331=6'h9; in332=6'h3; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h1; in337=6'h1; in338=6'h1; in339=6'h0; in340=6'h4; in341=6'h0; in342=6'h0; in343=6'h6; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h5; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h7; in355=6'h0; in356=6'h0; in357=6'h2; in358=6'h5; in359=6'h1; in360=6'h3; in361=6'h0; in362=6'h0; in363=6'h0; in364=6'h7; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h3; in373=6'h2; in374=6'h4; in375=6'h0; in376=6'h0; in377=6'h2; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h3; in4=6'h4; in5=6'h1; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h1; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h7; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h8; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h9; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h6; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'hA; in50=6'h8; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h3; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h6; in60=6'h1; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h3; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h3; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h1; in78=6'h3; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h2; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h2; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h1; in92=6'h2; in93=6'h0; in94=6'h0; in95=6'h3; in96=6'h3; in97=6'h8; in98=6'hE; in99=6'h2; in100=6'h4; in101=6'h0; in102=6'hE; in103=6'h9; in104=6'h2; in105=6'h3; in106=6'h0; in107=6'hE; in108=6'h2; in109=6'h3; in110=6'h2; in111=6'h0; in112=6'hB; in113=6'h0; in114=6'h3; in115=6'h2; in116=6'h0; in117=6'h7; in118=6'h0; in119=6'h3; in120=6'h0; in121=6'h0; in122=6'h6; in123=6'h5; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h5; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h1; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h1; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h1; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h1; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h3; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h3; in160=6'h0; in161=6'h8; in162=6'h9; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h9; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h2; in172=6'h11; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'h9; in177=6'h11; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'hE; in182=6'hF; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'hC; in187=6'h4; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h4; in192=6'h0; in193=6'h0; in194=6'h4; in195=6'h5; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h4; in200=6'h1; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h3; in205=6'h0; in206=6'h0; in207=6'h1; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h4; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h2; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h1; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h2; in231=6'h4; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h1; in236=6'h4; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h2; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h6; in281=6'h7; in282=6'h4; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h3; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h7; in317=6'h5; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h9; in322=6'h4; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'hA; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'hA; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h2; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h6; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h6; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h8; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h8; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h1; in362=6'h1; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h1; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h1; in377=6'h0; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h2; in2=6'h7; in3=6'h14; in4=6'h13; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h2; in9=6'h9; in10=6'h4; in11=6'h1; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h2; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h3; in31=6'h0; in32=6'h2; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h4; in37=6'h7; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h9; in42=6'h7; in43=6'h0; in44=6'h0; in45=6'h4; in46=6'h0; in47=6'h0; in48=6'h1; in49=6'h2; in50=6'hA; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'hC; in56=6'h3; in57=6'h0; in58=6'h0; in59=6'h4; in60=6'h2; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h3; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h6; in78=6'h1; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h2; in83=6'h7; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h1; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h4; in93=6'h1; in94=6'h0; in95=6'h4; in96=6'h0; in97=6'h1; in98=6'h0; in99=6'h1; in100=6'h2; in101=6'h0; in102=6'h0; in103=6'h1; in104=6'h0; in105=6'h1; in106=6'h0; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h4; in111=6'h0; in112=6'h8; in113=6'h6; in114=6'h1; in115=6'h3; in116=6'h0; in117=6'hD; in118=6'h4; in119=6'h2; in120=6'h0; in121=6'h0; in122=6'h3; in123=6'h2; in124=6'h0; in125=6'h0; in126=6'h9; in127=6'h10; in128=6'h0; in129=6'h0; in130=6'h2; in131=6'h2; in132=6'h0; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h5; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h2; in142=6'h7; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h2; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'hB; in154=6'h8; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h1; in160=6'h0; in161=6'h1; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h1; in167=6'h0; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h9; in172=6'h0; in173=6'h1; in174=6'h0; in175=6'h0; in176=6'h4; in177=6'h5; in178=6'h4; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h9; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h8; in187=6'hB; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h2; in194=6'h7; in195=6'h1; in196=6'h2; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h1; in206=6'h0; in207=6'h5; in208=6'h1; in209=6'h0; in210=6'h2; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h9; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'hB; in221=6'hB; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h1; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h0; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h1; in241=6'h8; in242=6'h3; in243=6'h0; in244=6'h0; in245=6'h8; in246=6'h10; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h1; in270=6'h5; in271=6'h9; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h0; in281=6'h0; in282=6'h1; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h6; in296=6'h7; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h4; in301=6'h3; in302=6'h3; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h5; in310=6'h5; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h3; in321=6'h1; in322=6'h0; in323=6'h0; in324=6'h2; in325=6'h2; in326=6'h5; in327=6'h9; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'hB; in332=6'hB; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h6; in339=6'h3; in340=6'h1; in341=6'h0; in342=6'h0; in343=6'h2; in344=6'h3; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h4; in350=6'h4; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h1; in355=6'h0; in356=6'h0; in357=6'h2; in358=6'h8; in359=6'hD; in360=6'hC; in361=6'h1; in362=6'h0; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h3; in369=6'h1; in370=6'h1; in371=6'h0; in372=6'h2; in373=6'h3; in374=6'h2; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h1;
      #50 in1=6'h3; in2=6'hD; in3=6'h14; in4=6'hF; in5=6'h5; in6=6'h0; in7=6'h0; in8=6'h3; in9=6'h7; in10=6'h5; in11=6'h1; in12=6'h4; in13=6'h2; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h6; in30=6'h0; in31=6'h0; in32=6'h3; in33=6'h0; in34=6'h5; in35=6'h0; in36=6'h0; in37=6'h2; in38=6'h0; in39=6'h0; in40=6'h1; in41=6'h3; in42=6'hA; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h5; in47=6'h0; in48=6'h0; in49=6'h1; in50=6'h7; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'hA; in56=6'h2; in57=6'h5; in58=6'h5; in59=6'h0; in60=6'h3; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h6; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h4; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'hB; in77=6'h5; in78=6'h0; in79=6'h1; in80=6'h1; in81=6'h0; in82=6'h1; in83=6'h5; in84=6'h1; in85=6'h2; in86=6'h3; in87=6'h3; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h0; in93=6'h0; in94=6'h0; in95=6'h1; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h1; in100=6'h6; in101=6'h1; in102=6'h0; in103=6'h3; in104=6'h1; in105=6'h2; in106=6'h0; in107=6'h0; in108=6'h3; in109=6'h0; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h2; in114=6'h0; in115=6'h1; in116=6'h0; in117=6'h0; in118=6'h4; in119=6'h0; in120=6'h0; in121=6'h6; in122=6'h7; in123=6'h0; in124=6'h0; in125=6'hD; in126=6'h11; in127=6'h2; in128=6'h3; in129=6'h0; in130=6'h3; in131=6'h0; in132=6'h8; in133=6'h9; in134=6'h0; in135=6'h1; in136=6'h4; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h0; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h7; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h7; in158=6'h4; in159=6'h0; in160=6'h0; in161=6'h0; in162=6'h3; in163=6'h4; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h0; in169=6'h0; in170=6'h8; in171=6'h0; in172=6'h0; in173=6'h6; in174=6'h0; in175=6'hE; in176=6'h0; in177=6'h6; in178=6'h9; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h6; in183=6'h7; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h8; in188=6'h7; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h3; in193=6'h9; in194=6'h0; in195=6'h0; in196=6'h2; in197=6'h5; in198=6'h3; in199=6'h0; in200=6'h2; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h1; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h1; in215=6'h0; in216=6'h1; in217=6'h6; in218=6'h0; in219=6'h13; in220=6'h2; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h3; in225=6'h3; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h5; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h0; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h6; in241=6'hD; in242=6'h5; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'hA; in250=6'hC; in251=6'h4; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h1; in261=6'h6; in262=6'h1; in263=6'h0; in264=6'h2; in265=6'h6; in266=6'h6; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h5; in271=6'h6; in272=6'h0; in273=6'h0; in274=6'h8; in275=6'hE; in276=6'h4; in277=6'h0; in278=6'h0; in279=6'h0; in280=6'h0; in281=6'h0; in282=6'h0; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h3; in291=6'h7; in292=6'h0; in293=6'h0; in294=6'h1; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h6; in300=6'hE; in301=6'h9; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h5; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h4; in320=6'h2; in321=6'h0; in322=6'h5; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h9; in328=6'h0; in329=6'h5; in330=6'h7; in331=6'h1; in332=6'h9; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h4; in338=6'h0; in339=6'h0; in340=6'h2; in341=6'h0; in342=6'h9; in343=6'h5; in344=6'h0; in345=6'h3; in346=6'h0; in347=6'h2; in348=6'h1; in349=6'h0; in350=6'h6; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h8; in356=6'h0; in357=6'h4; in358=6'h7; in359=6'h9; in360=6'h5; in361=6'h2; in362=6'h0; in363=6'h1; in364=6'h2; in365=6'h1; in366=6'h0; in367=6'h9; in368=6'h9; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h2; in373=6'h6; in374=6'h5; in375=6'h3; in376=6'h0; in377=6'h6; in378=6'h8; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h1; in2=6'h0; in3=6'h5; in4=6'h4; in5=6'h1; in6=6'h0; in7=6'h1; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'hD; in13=6'hC; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h6; in30=6'h2; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h5; in38=6'h0; in39=6'h1; in40=6'h3; in41=6'h2; in42=6'hB; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h2; in47=6'hA; in48=6'h8; in49=6'h8; in50=6'h10; in51=6'h0; in52=6'h3; in53=6'h4; in54=6'h0; in55=6'h11; in56=6'h0; in57=6'h0; in58=6'h1; in59=6'h0; in60=6'h6; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'hC; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h8; in70=6'h3; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h4; in81=6'h3; in82=6'h6; in83=6'h5; in84=6'h0; in85=6'h2; in86=6'h2; in87=6'h0; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h0; in93=6'h1; in94=6'h0; in95=6'h5; in96=6'hF; in97=6'h0; in98=6'h6; in99=6'h3; in100=6'h8; in101=6'hE; in102=6'h0; in103=6'h7; in104=6'h2; in105=6'h2; in106=6'h0; in107=6'h0; in108=6'h1; in109=6'h0; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h1; in114=6'h0; in115=6'h2; in116=6'h2; in117=6'h0; in118=6'h4; in119=6'h0; in120=6'h0; in121=6'h1; in122=6'h0; in123=6'h0; in124=6'h0; in125=6'h2; in126=6'h1; in127=6'h0; in128=6'h1; in129=6'h0; in130=6'h4; in131=6'h0; in132=6'h6; in133=6'h2; in134=6'h0; in135=6'h1; in136=6'h0; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h0; in142=6'h1; in143=6'h2; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h4; in150=6'h1; in151=6'h0; in152=6'hB; in153=6'h9; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h2; in158=6'h4; in159=6'h4; in160=6'h0; in161=6'h0; in162=6'h2; in163=6'h7; in164=6'h0; in165=6'hA; in166=6'h0; in167=6'h7; in168=6'h1; in169=6'h0; in170=6'hF; in171=6'h0; in172=6'h7; in173=6'h3; in174=6'h0; in175=6'hB; in176=6'h0; in177=6'h9; in178=6'h9; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h0; in183=6'h9; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'hB; in189=6'h2; in190=6'h0; in191=6'h2; in192=6'h3; in193=6'h5; in194=6'h0; in195=6'h1; in196=6'h1; in197=6'h0; in198=6'h0; in199=6'h2; in200=6'h3; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h5; in210=6'h0; in211=6'hA; in212=6'h0; in213=6'h0; in214=6'h2; in215=6'h0; in216=6'h4; in217=6'h6; in218=6'h0; in219=6'hF; in220=6'h4; in221=6'h2; in222=6'h3; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h1; in227=6'hB; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h4; in233=6'h0; in234=6'h2; in235=6'h0; in236=6'h0; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h1; in242=6'h0; in243=6'h0; in244=6'hA; in245=6'hF; in246=6'h5; in247=6'h0; in248=6'h0; in249=6'h2; in250=6'h8; in251=6'h5; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h1; in258=6'h1; in259=6'h0; in260=6'h0; in261=6'h2; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h2; in267=6'h0; in268=6'h0; in269=6'h7; in270=6'hC; in271=6'h7; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h1; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h1; in281=6'h2; in282=6'h5; in283=6'h6; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h8; in300=6'hC; in301=6'hB; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h0; in311=6'h3; in312=6'h2; in313=6'h0; in314=6'h6; in315=6'h4; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h3; in323=6'h0; in324=6'h6; in325=6'h5; in326=6'h0; in327=6'h6; in328=6'h0; in329=6'h6; in330=6'h7; in331=6'h0; in332=6'h5; in333=6'h0; in334=6'h2; in335=6'h0; in336=6'h6; in337=6'h8; in338=6'h7; in339=6'h0; in340=6'hA; in341=6'h0; in342=6'h7; in343=6'h8; in344=6'h0; in345=6'h4; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h0; in350=6'hC; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'hD; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h5; in360=6'h5; in361=6'h0; in362=6'h0; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h7; in373=6'h8; in374=6'h3; in375=6'h2; in376=6'h0; in377=6'h3; in378=6'h3; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h9; in2=6'hF; in3=6'h12; in4=6'h12; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h4; in14=6'h8; in15=6'h2; in16=6'h7; in17=6'h5; in18=6'h0; in19=6'hF; in20=6'h9; in21=6'hA; in22=6'hE; in23=6'hA; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h1; in30=6'h1; in31=6'h4; in32=6'h6; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h1; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h1; in50=6'h9; in51=6'h6; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h2; in57=6'h0; in58=6'h0; in59=6'h3; in60=6'hB; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h12; in66=6'hA; in67=6'h2; in68=6'h0; in69=6'h0; in70=6'h3; in71=6'h9; in72=6'h2; in73=6'h0; in74=6'h0; in75=6'h8; in76=6'h3; in77=6'h0; in78=6'hB; in79=6'h2; in80=6'h0; in81=6'h0; in82=6'h6; in83=6'hA; in84=6'h0; in85=6'h0; in86=6'h3; in87=6'h4; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h1; in92=6'hA; in93=6'hF; in94=6'h4; in95=6'h0; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h0; in101=6'h0; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h0; in106=6'h0; in107=6'h3; in108=6'h0; in109=6'h0; in110=6'h2; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'hC; in121=6'h9; in122=6'h1; in123=6'h0; in124=6'h0; in125=6'h6; in126=6'h0; in127=6'h7; in128=6'hB; in129=6'h0; in130=6'h0; in131=6'h7; in132=6'h9; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h2; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h4; in141=6'h3; in142=6'h6; in143=6'h8; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h3; in148=6'h0; in149=6'h1; in150=6'h1; in151=6'h0; in152=6'h0; in153=6'h7; in154=6'h6; in155=6'h0; in156=6'h1; in157=6'h0; in158=6'h7; in159=6'hE; in160=6'h4; in161=6'h5; in162=6'h0; in163=6'h2; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h6; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'h1; in173=6'h2; in174=6'h0; in175=6'h0; in176=6'h5; in177=6'h8; in178=6'h0; in179=6'h0; in180=6'h1; in181=6'h0; in182=6'h0; in183=6'h0; in184=6'h0; in185=6'h1; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h6; in200=6'h7; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h1; in210=6'h0; in211=6'h1; in212=6'h4; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h5; in221=6'hA; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h7; in227=6'h10; in228=6'h0; in229=6'h9; in230=6'h6; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h8; in235=6'hC; in236=6'h11; in237=6'hA; in238=6'h0; in239=6'h6; in240=6'h4; in241=6'h7; in242=6'h5; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'hA; in252=6'h8; in253=6'h0; in254=6'h5; in255=6'h8; in256=6'h3; in257=6'h0; in258=6'h0; in259=6'hA; in260=6'hC; in261=6'hB; in262=6'h0; in263=6'h0; in264=6'h4; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h3; in271=6'h1; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h7; in276=6'hC; in277=6'h6; in278=6'h0; in279=6'h7; in280=6'hB; in281=6'hB; in282=6'h7; in283=6'h2; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h8; in290=6'hC; in291=6'hD; in292=6'h2; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h1; in300=6'h2; in301=6'h5; in302=6'h1; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h0; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h6; in315=6'h2; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h8; in320=6'h0; in321=6'h1; in322=6'h6; in323=6'h0; in324=6'h2; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'h0; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h1; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h1; in345=6'h1; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h0; in350=6'h5; in351=6'h0; in352=6'h0; in353=6'h2; in354=6'h0; in355=6'h2; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h1; in362=6'hC; in363=6'h8; in364=6'h4; in365=6'h0; in366=6'h0; in367=6'h4; in368=6'h0; in369=6'h0; in370=6'h5; in371=6'h1; in372=6'h8; in373=6'h11; in374=6'hB; in375=6'h1; in376=6'h3; in377=6'h0; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h0; in2=6'h3; in3=6'hF; in4=6'hF; in5=6'h4; in6=6'h1; in7=6'h0; in8=6'h0; in9=6'hC; in10=6'h7; in11=6'hD; in12=6'h13; in13=6'h6; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h6; in20=6'hA; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h4; in38=6'h0; in39=6'h6; in40=6'h5; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h2; in45=6'h0; in46=6'h1; in47=6'h0; in48=6'h2; in49=6'h5; in50=6'hC; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h10; in56=6'h7; in57=6'h5; in58=6'h3; in59=6'h0; in60=6'h5; in61=6'h6; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h9; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h2; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h4; in78=6'h4; in79=6'h1; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h5; in84=6'h1; in85=6'h7; in86=6'hE; in87=6'hC; in88=6'hA; in89=6'h3; in90=6'h4; in91=6'h5; in92=6'h0; in93=6'h0; in94=6'h0; in95=6'h3; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h3; in101=6'h0; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h1; in106=6'h0; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h0; in121=6'h0; in122=6'h3; in123=6'h1; in124=6'h0; in125=6'h0; in126=6'h3; in127=6'h7; in128=6'h0; in129=6'h0; in130=6'h9; in131=6'h9; in132=6'h6; in133=6'h6; in134=6'h0; in135=6'h8; in136=6'h6; in137=6'h7; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h0; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h7; in149=6'h8; in150=6'h4; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'hB; in158=6'h7; in159=6'h2; in160=6'h8; in161=6'h5; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h1; in167=6'h3; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h2; in172=6'h1; in173=6'h0; in174=6'h0; in175=6'h5; in176=6'h4; in177=6'h0; in178=6'h7; in179=6'h0; in180=6'h9; in181=6'h0; in182=6'h0; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h2; in191=6'h3; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h3; in198=6'h7; in199=6'h3; in200=6'h2; in201=6'h0; in202=6'h6; in203=6'h6; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h4; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h2; in217=6'h8; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h8; in225=6'h0; in226=6'h0; in227=6'hF; in228=6'hC; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h0; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h3; in241=6'h6; in242=6'h3; in243=6'h0; in244=6'h2; in245=6'h1; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h2; in250=6'h1; in251=6'h2; in252=6'hC; in253=6'hA; in254=6'h6; in255=6'h6; in256=6'h0; in257=6'h4; in258=6'h7; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h2; in265=6'h7; in266=6'hA; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h8; in275=6'hB; in276=6'h5; in277=6'h6; in278=6'h8; in279=6'h6; in280=6'h5; in281=6'h0; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h3; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h1; in302=6'h0; in303=6'h0; in304=6'h9; in305=6'hB; in306=6'h5; in307=6'h6; in308=6'h8; in309=6'h2; in310=6'h1; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h4; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h0; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'hA; in330=6'h9; in331=6'h6; in332=6'h3; in333=6'h1; in334=6'h0; in335=6'h3; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h1; in340=6'h2; in341=6'h0; in342=6'h3; in343=6'h0; in344=6'h0; in345=6'h9; in346=6'h4; in347=6'h7; in348=6'h2; in349=6'h0; in350=6'h0; in351=6'h3; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h5; in359=6'hB; in360=6'h9; in361=6'h0; in362=6'h7; in363=6'h9; in364=6'h3; in365=6'h0; in366=6'h1; in367=6'h2; in368=6'h7; in369=6'h7; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h0; in374=6'h2; in375=6'h0; in376=6'h0; in377=6'hC; in378=6'hF; in379=6'hF; in380=6'h9; in381=6'h6;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h4; in5=6'h1; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h2; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h3; in24=6'h8; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h7; in32=6'h6; in33=6'h0; in34=6'h0; in35=6'h3; in36=6'h6; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h7; in41=6'h8; in42=6'h0; in43=6'h0; in44=6'h4; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h2; in50=6'hB; in51=6'h2; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h1; in57=6'h0; in58=6'h2; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h4; in64=6'h5; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h2; in69=6'h1; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h2; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h6; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h7; in83=6'h3; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h5; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h7; in92=6'h7; in93=6'h0; in94=6'h0; in95=6'h3; in96=6'h4; in97=6'h0; in98=6'hC; in99=6'h0; in100=6'h4; in101=6'h1; in102=6'hC; in103=6'h9; in104=6'h0; in105=6'h4; in106=6'h5; in107=6'hE; in108=6'h3; in109=6'h1; in110=6'h2; in111=6'h9; in112=6'hC; in113=6'h0; in114=6'h2; in115=6'h1; in116=6'h1; in117=6'h0; in118=6'h0; in119=6'h2; in120=6'h0; in121=6'h0; in122=6'h5; in123=6'h7; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h6; in128=6'h4; in129=6'h0; in130=6'h0; in131=6'h2; in132=6'h6; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h1; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h2; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h1; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h1; in150=6'h1; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h1; in155=6'h1; in156=6'h0; in157=6'h0; in158=6'h4; in159=6'h0; in160=6'h0; in161=6'hD; in162=6'hB; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'hA; in168=6'h6; in169=6'h0; in170=6'h0; in171=6'h1; in172=6'hE; in173=6'h2; in174=6'h0; in175=6'h0; in176=6'hC; in177=6'hD; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'h10; in182=6'h9; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h7; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h5; in192=6'h0; in193=6'h0; in194=6'h6; in195=6'h6; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h6; in200=6'h1; in201=6'h0; in202=6'h0; in203=6'h2; in204=6'h7; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h3; in212=6'h2; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h1; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h3; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h6; in231=6'h1; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h5; in237=6'h1; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h4; in256=6'hA; in257=6'h3; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h1; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h3; in280=6'hA; in281=6'hC; in282=6'h3; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h1; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h3; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h2; in317=6'h9; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h8; in322=6'hB; in323=6'h0; in324=6'h0; in325=6'h3; in326=6'h9; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h4; in331=6'h5; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h1; in336=6'h4; in337=6'h0; in338=6'h0; in339=6'h2; in340=6'h2; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h2; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'hA; in349=6'h9; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h8; in354=6'h8; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h0; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h1; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h1; in376=6'h1; in377=6'h0; in378=6'h0; in379=6'h0; in380=6'h2; in381=6'h1;
      #50 in1=6'h0; in2=6'h0; in3=6'h9; in4=6'h10; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h2; in12=6'h1; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h2; in19=6'h1; in20=6'h0; in21=6'h0; in22=6'h4; in23=6'h5; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h6; in32=6'h0; in33=6'h2; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h1; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'hA; in51=6'h11; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'hB; in57=6'h4; in58=6'h2; in59=6'h0; in60=6'h0; in61=6'h3; in62=6'h4; in63=6'h5; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h1; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h3; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h1; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h1; in87=6'h0; in88=6'h7; in89=6'h4; in90=6'h5; in91=6'h7; in92=6'hB; in93=6'hA; in94=6'h0; in95=6'h1; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h2; in101=6'h0; in102=6'h3; in103=6'h0; in104=6'h4; in105=6'h1; in106=6'h8; in107=6'h5; in108=6'h0; in109=6'h6; in110=6'h0; in111=6'hE; in112=6'h0; in113=6'h5; in114=6'h7; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h0; in121=6'h5; in122=6'h6; in123=6'h1; in124=6'h0; in125=6'h1; in126=6'h0; in127=6'h2; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h3; in132=6'h0; in133=6'h0; in134=6'h6; in135=6'h1; in136=6'h5; in137=6'h4; in138=6'hE; in139=6'h4; in140=6'h2; in141=6'h0; in142=6'hC; in143=6'h1; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h2; in149=6'h1; in150=6'h0; in151=6'h1; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h2; in160=6'h9; in161=6'hB; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h2; in168=6'h1; in169=6'h2; in170=6'h0; in171=6'h0; in172=6'h3; in173=6'h0; in174=6'h3; in175=6'h2; in176=6'h4; in177=6'h0; in178=6'h4; in179=6'h6; in180=6'h11; in181=6'h6; in182=6'h0; in183=6'h6; in184=6'h0; in185=6'hB; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h3; in199=6'h1; in200=6'h0; in201=6'h1; in202=6'h2; in203=6'h6; in204=6'h0; in205=6'h3; in206=6'h0; in207=6'h0; in208=6'h1; in209=6'h0; in210=6'h0; in211=6'h2; in212=6'h8; in213=6'h7; in214=6'h0; in215=6'h2; in216=6'h1; in217=6'h0; in218=6'hB; in219=6'h2; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h6; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'hD; in230=6'hC; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h8; in236=6'h6; in237=6'h5; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h3; in243=6'h2; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h6; in255=6'hC; in256=6'h6; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h3; in261=6'h5; in262=6'h2; in263=6'h0; in264=6'h0; in265=6'h3; in266=6'h2; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h1; in278=6'h0; in279=6'hA; in280=6'hF; in281=6'h8; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h2; in286=6'h1; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h1; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h1; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h1; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h1; in315=6'h0; in316=6'h8; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h1; in321=6'h9; in322=6'h0; in323=6'h3; in324=6'h1; in325=6'h2; in326=6'h0; in327=6'h0; in328=6'h8; in329=6'h0; in330=6'h0; in331=6'h0; in332=6'h7; in333=6'h6; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h2; in340=6'h0; in341=6'h5; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h2; in348=6'h9; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h1; in353=6'hB; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h3; in362=6'h1; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h2; in368=6'h3; in369=6'h5; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h2; in374=6'h0; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h9; in380=6'hA; in381=6'h3;
      #50 in1=6'h0; in2=6'h0; in3=6'h1; in4=6'h0; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h1; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h4; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h2; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h1; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'hB; in50=6'h6; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h1; in55=6'h3; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h3; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h5; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h4; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h0; in93=6'h0; in94=6'h0; in95=6'h2; in96=6'h3; in97=6'h9; in98=6'hA; in99=6'h3; in100=6'h2; in101=6'h3; in102=6'hA; in103=6'h7; in104=6'h3; in105=6'h2; in106=6'h3; in107=6'h7; in108=6'h1; in109=6'h3; in110=6'h2; in111=6'h3; in112=6'h8; in113=6'h1; in114=6'h3; in115=6'h2; in116=6'h2; in117=6'h8; in118=6'h1; in119=6'h3; in120=6'h0; in121=6'h0; in122=6'h2; in123=6'h1; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h1; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h0; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h1; in142=6'h2; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h1; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h0; in160=6'h0; in161=6'h1; in162=6'h4; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h5; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'hA; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'h0; in177=6'hA; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'hA; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'hA; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h2; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h1; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h3; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h1; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h1; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h2; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h1; in236=6'h2; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h4; in281=6'h4; in282=6'h4; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h1; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h2; in311=6'h2; in312=6'h0; in313=6'h1; in314=6'h0; in315=6'h0; in316=6'h6; in317=6'h3; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h8; in322=6'h3; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h4; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'h5; in332=6'h2; in333=6'h0; in334=6'h0; in335=6'h4; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h5; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h4; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h5; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h6; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h1; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h1; in367=6'h1; in368=6'h0; in369=6'h2; in370=6'h0; in371=6'h1; in372=6'h1; in373=6'h0; in374=6'h2; in375=6'h1; in376=6'h1; in377=6'h1; in378=6'h0; in379=6'h0; in380=6'h0; in381=6'h0;
      #50 in1=6'h0; in2=6'h0; in3=6'h4; in4=6'h2; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h2; in15=6'h1; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h2; in25=6'h1; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'hB; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h7; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h8; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h4; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'hE; in50=6'h5; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h9; in55=6'h3; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'hA; in60=6'h8; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h3; in65=6'h5; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h1; in70=6'h0; in71=6'h0; in72=6'h2; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h2; in78=6'h2; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h1; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h1; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h5; in93=6'h3; in94=6'h0; in95=6'h2; in96=6'h0; in97=6'hA; in98=6'h0; in99=6'h3; in100=6'h2; in101=6'h0; in102=6'h7; in103=6'h0; in104=6'h3; in105=6'h3; in106=6'h0; in107=6'h7; in108=6'h1; in109=6'h3; in110=6'h3; in111=6'h0; in112=6'h5; in113=6'h1; in114=6'h2; in115=6'h2; in116=6'h0; in117=6'h3; in118=6'h0; in119=6'h0; in120=6'h0; in121=6'h1; in122=6'h4; in123=6'h0; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h0; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h0; in142=6'h1; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h2; in149=6'h4; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h5; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h5; in160=6'h0; in161=6'h4; in162=6'hA; in163=6'h4; in164=6'h0; in165=6'h0; in166=6'h6; in167=6'hB; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h6; in172=6'hD; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'h6; in177=6'hD; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'h6; in182=6'hD; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h4; in187=6'h8; in188=6'h0; in189=6'h0; in190=6'h3; in191=6'h2; in192=6'h0; in193=6'h0; in194=6'h1; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h2; in205=6'h1; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h1; in211=6'h3; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h4; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h3; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h1; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h4; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h5; in236=6'h1; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h2; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h2; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h6; in257=6'h5; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h5; in281=6'h9; in282=6'h5; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h2; in307=6'h0; in308=6'h0; in309=6'h2; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h1; in314=6'h0; in315=6'h0; in316=6'h9; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h9; in322=6'h0; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h6; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'hA; in332=6'h4; in333=6'h0; in334=6'h0; in335=6'h7; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'hA; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'hA; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'hB; in350=6'h3; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h7; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h0; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h1; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h1; in372=6'h1; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h0; in377=6'h1; in378=6'h0; in379=6'h1; in380=6'h2; in381=6'h2;
      #50 in1=6'h0; in2=6'h9; in3=6'h9; in4=6'hE; in5=6'hA; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h3; in17=6'h7; in18=6'h4; in19=6'h1; in20=6'h0; in21=6'h6; in22=6'hA; in23=6'h7; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h4; in30=6'h0; in31=6'h1; in32=6'h0; in33=6'h3; in34=6'h6; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h2; in39=6'h8; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h5; in51=6'h11; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'hE; in57=6'h4; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h3; in62=6'h7; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h6; in72=6'h6; in73=6'h5; in74=6'h0; in75=6'h2; in76=6'h7; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h1; in81=6'h0; in82=6'h0; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h5; in89=6'h4; in90=6'h4; in91=6'h9; in92=6'hB; in93=6'hA; in94=6'h0; in95=6'h0; in96=6'h2; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'hE; in101=6'h7; in102=6'h0; in103=6'h0; in104=6'h7; in105=6'hD; in106=6'h0; in107=6'h2; in108=6'h0; in109=6'hB; in110=6'h8; in111=6'h0; in112=6'h0; in113=6'h7; in114=6'h9; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h1; in119=6'h0; in120=6'h0; in121=6'hF; in122=6'h4; in123=6'h2; in124=6'h0; in125=6'hB; in126=6'hB; in127=6'h0; in128=6'h0; in129=6'h0; in130=6'h2; in131=6'h0; in132=6'h0; in133=6'h0; in134=6'h5; in135=6'h0; in136=6'h0; in137=6'h2; in138=6'hC; in139=6'h5; in140=6'h0; in141=6'h3; in142=6'hE; in143=6'h5; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h1; in156=6'h2; in157=6'h1; in158=6'h0; in159=6'h2; in160=6'h9; in161=6'h4; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h0; in169=6'h1; in170=6'hA; in171=6'h1; in172=6'h0; in173=6'h0; in174=6'h9; in175=6'hE; in176=6'h0; in177=6'h0; in178=6'h7; in179=6'hC; in180=6'hC; in181=6'h0; in182=6'h0; in183=6'h8; in184=6'h2; in185=6'h4; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h1; in190=6'h0; in191=6'h0; in192=6'h5; in193=6'h6; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h4; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h2; in202=6'h2; in203=6'h0; in204=6'h0; in205=6'h3; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h1; in210=6'h0; in211=6'h0; in212=6'h8; in213=6'hD; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h8; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'hC; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'hD; in230=6'h1; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h7; in236=6'h8; in237=6'h9; in238=6'h4; in239=6'h1; in240=6'h0; in241=6'h0; in242=6'h4; in243=6'h3; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'hC; in255=6'hE; in256=6'h7; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h4; in261=6'h3; in262=6'h5; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h1; in271=6'h1; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h2; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'hC; in280=6'h10; in281=6'h8; in282=6'h2; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h4; in291=6'h7; in292=6'h8; in293=6'h1; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h1; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h8; in316=6'h3; in317=6'h0; in318=6'h0; in319=6'hA; in320=6'hA; in321=6'h3; in322=6'h0; in323=6'h5; in324=6'hC; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'hA; in329=6'h0; in330=6'h0; in331=6'h0; in332=6'h8; in333=6'h9; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h1; in338=6'h0; in339=6'h0; in340=6'h0; in341=6'h6; in342=6'h4; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h3; in347=6'h8; in348=6'h0; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h9; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h0; in363=6'h3; in364=6'h4; in365=6'h0; in366=6'h0; in367=6'h1; in368=6'h0; in369=6'h1; in370=6'h0; in371=6'h0; in372=6'h3; in373=6'h2; in374=6'h1; in375=6'h0; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h8; in380=6'hC; in381=6'h3;
      #50 in1=6'h0; in2=6'h1; in3=6'h8; in4=6'hD; in5=6'h8; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h1; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h3; in31=6'h2; in32=6'h5; in33=6'h0; in34=6'h0; in35=6'h4; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h4; in41=6'hA; in42=6'h0; in43=6'h0; in44=6'h4; in45=6'h4; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h1; in50=6'h8; in51=6'h1; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h4; in56=6'h1; in57=6'h0; in58=6'h2; in59=6'h6; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h3; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h4; in78=6'h4; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h6; in83=6'h7; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h3; in88=6'h3; in89=6'h0; in90=6'h0; in91=6'h0; in92=6'h4; in93=6'h0; in94=6'h0; in95=6'h4; in96=6'h2; in97=6'h0; in98=6'h2; in99=6'h0; in100=6'h4; in101=6'h1; in102=6'h4; in103=6'h0; in104=6'h0; in105=6'h1; in106=6'h3; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h4; in111=6'h0; in112=6'h6; in113=6'h0; in114=6'h2; in115=6'h3; in116=6'hA; in117=6'hB; in118=6'h0; in119=6'h3; in120=6'h0; in121=6'h0; in122=6'h7; in123=6'h7; in124=6'h0; in125=6'h0; in126=6'h8; in127=6'hF; in128=6'h0; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h0; in133=6'h2; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'h0; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h6; in142=6'h4; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'hA; in154=6'h5; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h8; in159=6'h7; in160=6'h1; in161=6'h4; in162=6'h2; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h2; in168=6'h1; in169=6'h0; in170=6'h0; in171=6'hE; in172=6'h5; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'hC; in177=6'h2; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'h6; in182=6'h5; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'hC; in187=6'h2; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h1; in192=6'h0; in193=6'h1; in194=6'hA; in195=6'h3; in196=6'h0; in197=6'h0; in198=6'h3; in199=6'h5; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h3; in208=6'h0; in209=6'h0; in210=6'h1; in211=6'h0; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'hE; in221=6'h4; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h2; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h3; in237=6'h2; in238=6'h0; in239=6'h0; in240=6'h1; in241=6'h7; in242=6'h2; in243=6'h0; in244=6'h0; in245=6'h5; in246=6'h6; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h7; in251=6'h5; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h1; in270=6'h6; in271=6'h6; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h1; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h0; in280=6'h5; in281=6'h2; in282=6'h1; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h5; in301=6'h3; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h4; in310=6'h5; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h2; in321=6'h2; in322=6'h4; in323=6'h1; in324=6'h0; in325=6'h3; in326=6'h6; in327=6'h5; in328=6'h0; in329=6'h0; in330=6'h4; in331=6'hD; in332=6'h3; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h3; in339=6'h1; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h8; in344=6'h7; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h1; in349=6'h7; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h1; in354=6'h3; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h2; in359=6'h3; in360=6'h6; in361=6'h1; in362=6'h0; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h3; in374=6'h0; in375=6'h0; in376=6'h1; in377=6'h0; in378=6'h0; in379=6'h0; in380=6'h1; in381=6'h1;
      #50 in1=6'h0; in2=6'h2; in3=6'h8; in4=6'hB; in5=6'hA; in6=6'h2; in7=6'h4; in8=6'hB; in9=6'hF; in10=6'hE; in11=6'h0; in12=6'h0; in13=6'h5; in14=6'h7; in15=6'h0; in16=6'hB; in17=6'hB; in18=6'h1; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h2; in45=6'h1; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h0; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h4; in60=6'h12; in61=6'h0; in62=6'h1; in63=6'h1; in64=6'h0; in65=6'h7; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h5; in78=6'hA; in79=6'h7; in80=6'h0; in81=6'h6; in82=6'h9; in83=6'h6; in84=6'h1; in85=6'h0; in86=6'h0; in87=6'h5; in88=6'hA; in89=6'h0; in90=6'h2; in91=6'h6; in92=6'hA; in93=6'h2; in94=6'h0; in95=6'h4; in96=6'h3; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h3; in101=6'h0; in102=6'h2; in103=6'h0; in104=6'h0; in105=6'h1; in106=6'h0; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h0; in121=6'h0; in122=6'h0; in123=6'h0; in124=6'h0; in125=6'h0; in126=6'h4; in127=6'hD; in128=6'h8; in129=6'h4; in130=6'h2; in131=6'h9; in132=6'h1; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h0; in137=6'hB; in138=6'h4; in139=6'h0; in140=6'h3; in141=6'h0; in142=6'h1; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h2; in151=6'h0; in152=6'h2; in153=6'h8; in154=6'hC; in155=6'h0; in156=6'h0; in157=6'h3; in158=6'h0; in159=6'h0; in160=6'h2; in161=6'h1; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h0; in169=6'h0; in170=6'h0; in171=6'h6; in172=6'h4; in173=6'h0; in174=6'h0; in175=6'h2; in176=6'h8; in177=6'h0; in178=6'h0; in179=6'h0; in180=6'h4; in181=6'h0; in182=6'h0; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h8; in195=6'h2; in196=6'h0; in197=6'h0; in198=6'h1; in199=6'h3; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h3; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h1; in211=6'h2; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h1; in216=6'h0; in217=6'h1; in218=6'h0; in219=6'h0; in220=6'h5; in221=6'hC; in222=6'h3; in223=6'h0; in224=6'hF; in225=6'h5; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h0; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h8; in243=6'h9; in244=6'h0; in245=6'h2; in246=6'hB; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h1; in252=6'h1; in253=6'h0; in254=6'hA; in255=6'hE; in256=6'h6; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h2; in267=6'hD; in268=6'hE; in269=6'h0; in270=6'h8; in271=6'h7; in272=6'h0; in273=6'h0; in274=6'h2; in275=6'h5; in276=6'h5; in277=6'h0; in278=6'h0; in279=6'h5; in280=6'h9; in281=6'h3; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h1; in287=6'h0; in288=6'h0; in289=6'h1; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h4; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h7; in299=6'h1; in300=6'h6; in301=6'h5; in302=6'h0; in303=6'h0; in304=6'h5; in305=6'hE; in306=6'hB; in307=6'h1; in308=6'h1; in309=6'h3; in310=6'h7; in311=6'h7; in312=6'h1; in313=6'h0; in314=6'h1; in315=6'h0; in316=6'h0; in317=6'h0; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h0; in322=6'h0; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h0; in331=6'h4; in332=6'h6; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h1; in339=6'h2; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h1; in344=6'h1; in345=6'h2; in346=6'h0; in347=6'h3; in348=6'h0; in349=6'h3; in350=6'h6; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h4; in359=6'h7; in360=6'h7; in361=6'h5; in362=6'h1; in363=6'h1; in364=6'h0; in365=6'h0; in366=6'h3; in367=6'h3; in368=6'h0; in369=6'h0; in370=6'h8; in371=6'h9; in372=6'h5; in373=6'hC; in374=6'h1; in375=6'h0; in376=6'h0; in377=6'h4; in378=6'hB; in379=6'h10; in380=6'h9; in381=6'h2;
      #50 in1=6'h0; in2=6'h4; in3=6'hD; in4=6'hF; in5=6'h7; in6=6'h4; in7=6'h1; in8=6'h0; in9=6'h0; in10=6'h1; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h2; in16=6'h3; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h8; in22=6'h7; in23=6'h2; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h7; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h6; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h2; in43=6'h0; in44=6'h0; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'hB; in51=6'h2; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'hA; in56=6'h1; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'hB; in61=6'h7; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h0; in74=6'h2; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h7; in79=6'h3; in80=6'h0; in81=6'h5; in82=6'h7; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h4; in89=6'h0; in90=6'h0; in91=6'h7; in92=6'hC; in93=6'h6; in94=6'h0; in95=6'h2; in96=6'h0; in97=6'h0; in98=6'h3; in99=6'h1; in100=6'h2; in101=6'h0; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h0; in106=6'h2; in107=6'h0; in108=6'h0; in109=6'h0; in110=6'h0; in111=6'h1; in112=6'h0; in113=6'h7; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h5; in118=6'h1; in119=6'h1; in120=6'h0; in121=6'h6; in122=6'h2; in123=6'h0; in124=6'h1; in125=6'h0; in126=6'h0; in127=6'hB; in128=6'h1; in129=6'h0; in130=6'h5; in131=6'hE; in132=6'hC; in133=6'h0; in134=6'h0; in135=6'h1; in136=6'h0; in137=6'h8; in138=6'h9; in139=6'h0; in140=6'h1; in141=6'hB; in142=6'hC; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h1; in154=6'h2; in155=6'h4; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h0; in160=6'h5; in161=6'h0; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h6; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'h0; in173=6'h7; in174=6'h0; in175=6'h0; in176=6'h0; in177=6'h0; in178=6'h5; in179=6'h0; in180=6'h0; in181=6'h0; in182=6'h3; in183=6'h7; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h3; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h1; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h1; in203=6'h0; in204=6'h0; in205=6'h1; in206=6'h0; in207=6'h1; in208=6'h1; in209=6'h0; in210=6'h5; in211=6'h0; in212=6'h4; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h3; in218=6'h0; in219=6'h2; in220=6'h0; in221=6'h0; in222=6'h6; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'hA; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h7; in236=6'hE; in237=6'h7; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h1; in245=6'h2; in246=6'h7; in247=6'h6; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h3; in255=6'h4; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h2; in260=6'h7; in261=6'h8; in262=6'h2; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h4; in270=6'h9; in271=6'h6; in272=6'h0; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'hE; in280=6'h11; in281=6'h6; in282=6'h0; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h1; in290=6'h9; in291=6'h8; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h7; in296=6'h7; in297=6'h0; in298=6'h0; in299=6'h2; in300=6'h5; in301=6'h1; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h0; in306=6'h0; in307=6'h0; in308=6'h0; in309=6'h1; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h0; in317=6'h1; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'h1; in322=6'h1; in323=6'h0; in324=6'h3; in325=6'h7; in326=6'h1; in327=6'h9; in328=6'h6; in329=6'h0; in330=6'h0; in331=6'h4; in332=6'hA; in333=6'h3; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h6; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h6; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h0; in350=6'h2; in351=6'h0; in352=6'h1; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h1; in363=6'h4; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h0; in368=6'h1; in369=6'h6; in370=6'h0; in371=6'h0; in372=6'hC; in373=6'hB; in374=6'h3; in375=6'h0; in376=6'h0; in377=6'h2; in378=6'h0; in379=6'h7; in380=6'h6; in381=6'h1;
      #50 in1=6'h0; in2=6'h0; in3=6'h0; in4=6'h1; in5=6'h0; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h0; in17=6'h0; in18=6'h0; in19=6'h0; in20=6'h0; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h1; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h5; in32=6'h0; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h7; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h7; in42=6'h0; in43=6'h0; in44=6'h0; in45=6'h2; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h9; in51=6'h0; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h0; in57=6'h0; in58=6'h0; in59=6'h5; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h5; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h1; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h4; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h2; in83=6'h0; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h0; in88=6'h0; in89=6'h0; in90=6'h0; in91=6'h3; in92=6'h3; in93=6'h0; in94=6'h0; in95=6'h3; in96=6'h4; in97=6'h0; in98=6'hD; in99=6'h0; in100=6'h4; in101=6'h3; in102=6'h10; in103=6'hB; in104=6'h0; in105=6'h4; in106=6'h0; in107=6'h10; in108=6'h2; in109=6'h3; in110=6'h3; in111=6'h0; in112=6'hD; in113=6'h0; in114=6'h3; in115=6'h1; in116=6'h0; in117=6'h7; in118=6'h0; in119=6'h3; in120=6'h0; in121=6'h0; in122=6'h3; in123=6'h6; in124=6'h0; in125=6'h0; in126=6'h0; in127=6'h6; in128=6'h2; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'h1; in133=6'h0; in134=6'h0; in135=6'h0; in136=6'h2; in137=6'h2; in138=6'h0; in139=6'h0; in140=6'h0; in141=6'h5; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h0; in146=6'h0; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h1; in155=6'h0; in156=6'h0; in157=6'h0; in158=6'h1; in159=6'h1; in160=6'h0; in161=6'h7; in162=6'h8; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h9; in168=6'h3; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'hE; in173=6'h0; in174=6'h0; in175=6'h0; in176=6'hA; in177=6'h12; in178=6'h0; in179=6'h0; in180=6'h0; in181=6'hF; in182=6'hC; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h9; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h3; in192=6'h0; in193=6'h0; in194=6'h4; in195=6'h6; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h5; in200=6'h1; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h4; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h1; in212=6'h0; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h0; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h3; in231=6'h2; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h2; in237=6'h0; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h0; in254=6'h0; in255=6'h0; in256=6'h3; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h0; in261=6'h0; in262=6'h0; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h1; in273=6'h0; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h0; in278=6'h0; in279=6'h1; in280=6'h5; in281=6'h5; in282=6'h3; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h0; in291=6'h0; in292=6'h0; in293=6'h0; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h1; in306=6'h2; in307=6'h0; in308=6'h0; in309=6'h3; in310=6'h3; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h0; in315=6'h0; in316=6'h4; in317=6'h8; in318=6'h0; in319=6'h0; in320=6'h0; in321=6'hA; in322=6'h7; in323=6'h0; in324=6'h0; in325=6'h0; in326=6'h8; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h2; in331=6'h9; in332=6'h0; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h1; in337=6'h0; in338=6'h0; in339=6'h2; in340=6'h0; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h4; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h0; in349=6'h8; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h5; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h1; in363=6'h0; in364=6'h0; in365=6'h0; in366=6'h0; in367=6'h1; in368=6'h0; in369=6'h0; in370=6'h0; in371=6'h1; in372=6'h0; in373=6'h0; in374=6'h0; in375=6'h0; in376=6'h1; in377=6'h0; in378=6'h3; in379=6'h1; in380=6'h1; in381=6'h1;
      #50 in1=6'h0; in2=6'h0; in3=6'h3; in4=6'hE; in5=6'hB; in6=6'h0; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h4; in12=6'hA; in13=6'hB; in14=6'h9; in15=6'h0; in16=6'h6; in17=6'h6; in18=6'h9; in19=6'h9; in20=6'h2; in21=6'h0; in22=6'h0; in23=6'h0; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h0; in32=6'h0; in33=6'h3; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h2; in45=6'h1; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'h4; in51=6'hC; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h7; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h1; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h0; in72=6'h0; in73=6'h4; in74=6'h0; in75=6'h0; in76=6'h0; in77=6'h0; in78=6'h0; in79=6'h0; in80=6'h0; in81=6'h0; in82=6'h0; in83=6'h1; in84=6'h0; in85=6'h0; in86=6'hC; in87=6'hC; in88=6'h7; in89=6'h0; in90=6'h6; in91=6'h8; in92=6'h0; in93=6'h0; in94=6'h0; in95=6'h2; in96=6'h2; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h3; in101=6'h3; in102=6'h0; in103=6'h0; in104=6'h0; in105=6'h3; in106=6'h1; in107=6'h0; in108=6'h0; in109=6'h1; in110=6'h0; in111=6'h0; in112=6'h0; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h0; in117=6'h0; in118=6'h0; in119=6'h2; in120=6'h0; in121=6'h0; in122=6'h9; in123=6'h6; in124=6'h1; in125=6'h0; in126=6'h1; in127=6'h3; in128=6'h0; in129=6'h1; in130=6'h0; in131=6'h0; in132=6'h2; in133=6'h7; in134=6'h2; in135=6'h8; in136=6'hB; in137=6'hD; in138=6'h1; in139=6'h0; in140=6'h6; in141=6'h0; in142=6'h0; in143=6'h0; in144=6'h0; in145=6'h1; in146=6'h1; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h0; in156=6'h0; in157=6'h3; in158=6'h0; in159=6'h0; in160=6'h3; in161=6'h3; in162=6'h0; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h0; in169=6'h1; in170=6'h0; in171=6'h0; in172=6'h0; in173=6'h0; in174=6'h0; in175=6'h2; in176=6'h0; in177=6'h0; in178=6'h0; in179=6'h0; in180=6'h2; in181=6'h0; in182=6'h0; in183=6'h0; in184=6'h0; in185=6'h0; in186=6'h0; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h0; in200=6'h0; in201=6'h0; in202=6'h0; in203=6'h0; in204=6'h0; in205=6'h0; in206=6'h0; in207=6'h0; in208=6'h0; in209=6'h0; in210=6'h0; in211=6'h5; in212=6'h4; in213=6'h6; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h3; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h5; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h0; in230=6'h0; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h0; in235=6'h0; in236=6'h7; in237=6'hC; in238=6'h4; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h5; in243=6'h2; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h6; in250=6'h9; in251=6'h7; in252=6'h4; in253=6'h0; in254=6'h6; in255=6'h5; in256=6'h0; in257=6'h0; in258=6'h0; in259=6'h0; in260=6'h2; in261=6'h9; in262=6'hA; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h0; in274=6'hA; in275=6'hC; in276=6'h7; in277=6'h4; in278=6'h0; in279=6'h3; in280=6'h2; in281=6'h0; in282=6'h0; in283=6'h1; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h0; in290=6'h1; in291=6'h9; in292=6'hA; in293=6'h4; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h3; in302=6'h4; in303=6'h1; in304=6'h8; in305=6'hB; in306=6'h5; in307=6'h1; in308=6'h1; in309=6'h3; in310=6'h2; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h2; in315=6'h3; in316=6'h5; in317=6'h0; in318=6'h0; in319=6'h5; in320=6'h3; in321=6'h0; in322=6'h0; in323=6'h1; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h1; in329=6'h4; in330=6'h9; in331=6'h6; in332=6'h1; in333=6'h0; in334=6'h0; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h0; in341=6'h1; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h4; in348=6'h2; in349=6'h0; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h0; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h1; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h1; in363=6'h3; in364=6'h7; in365=6'h2; in366=6'h1; in367=6'h8; in368=6'h7; in369=6'h9; in370=6'h0; in371=6'h0; in372=6'h0; in373=6'h0; in374=6'h5; in375=6'h9; in376=6'h3; in377=6'hC; in378=6'hC; in379=6'hC; in380=6'h5; in381=6'h1;
      #50 in1=6'h1; in2=6'h4; in3=6'h10; in4=6'h11; in5=6'h8; in6=6'h1; in7=6'h0; in8=6'h0; in9=6'h0; in10=6'h0; in11=6'h0; in12=6'h0; in13=6'h0; in14=6'h0; in15=6'h0; in16=6'h1; in17=6'h1; in18=6'h3; in19=6'h9; in20=6'h9; in21=6'h0; in22=6'h0; in23=6'h1; in24=6'h0; in25=6'h0; in26=6'h0; in27=6'h0; in28=6'h0; in29=6'h0; in30=6'h0; in31=6'h3; in32=6'h7; in33=6'h0; in34=6'h0; in35=6'h0; in36=6'h0; in37=6'h0; in38=6'h0; in39=6'h0; in40=6'h0; in41=6'h0; in42=6'h0; in43=6'h0; in44=6'h2; in45=6'h0; in46=6'h0; in47=6'h0; in48=6'h0; in49=6'h0; in50=6'hE; in51=6'h7; in52=6'h0; in53=6'h0; in54=6'h0; in55=6'h0; in56=6'h2; in57=6'h0; in58=6'h0; in59=6'h0; in60=6'h0; in61=6'h0; in62=6'h0; in63=6'h0; in64=6'h0; in65=6'h0; in66=6'h0; in67=6'h0; in68=6'h0; in69=6'h0; in70=6'h0; in71=6'h6; in72=6'h4; in73=6'h1; in74=6'h0; in75=6'h0; in76=6'h2; in77=6'h0; in78=6'h6; in79=6'h1; in80=6'h0; in81=6'h0; in82=6'h4; in83=6'h5; in84=6'h0; in85=6'h0; in86=6'h0; in87=6'h4; in88=6'h0; in89=6'h1; in90=6'h2; in91=6'hA; in92=6'hB; in93=6'hA; in94=6'h0; in95=6'h0; in96=6'h0; in97=6'h0; in98=6'h0; in99=6'h0; in100=6'h0; in101=6'h0; in102=6'h0; in103=6'h1; in104=6'h0; in105=6'h4; in106=6'h0; in107=6'hC; in108=6'hA; in109=6'h0; in110=6'h2; in111=6'h6; in112=6'h8; in113=6'h0; in114=6'h0; in115=6'h0; in116=6'h3; in117=6'h0; in118=6'h0; in119=6'h0; in120=6'h4; in121=6'hA; in122=6'h8; in123=6'h0; in124=6'h0; in125=6'h4; in126=6'h0; in127=6'h0; in128=6'h9; in129=6'h0; in130=6'h0; in131=6'h0; in132=6'hA; in133=6'h4; in134=6'h0; in135=6'h0; in136=6'hA; in137=6'h8; in138=6'h8; in139=6'h4; in140=6'h4; in141=6'h5; in142=6'h7; in143=6'h6; in144=6'h0; in145=6'h0; in146=6'h1; in147=6'h0; in148=6'h0; in149=6'h0; in150=6'h0; in151=6'h0; in152=6'h0; in153=6'h0; in154=6'h0; in155=6'h1; in156=6'h0; in157=6'h0; in158=6'h0; in159=6'h0; in160=6'h5; in161=6'hB; in162=6'h4; in163=6'h0; in164=6'h0; in165=6'h0; in166=6'h0; in167=6'h0; in168=6'h2; in169=6'h0; in170=6'h0; in171=6'h0; in172=6'h0; in173=6'h5; in174=6'h0; in175=6'h0; in176=6'h0; in177=6'h8; in178=6'h1; in179=6'h0; in180=6'h1; in181=6'hC; in182=6'h6; in183=6'h0; in184=6'h0; in185=6'h4; in186=6'hA; in187=6'h0; in188=6'h0; in189=6'h0; in190=6'h0; in191=6'h0; in192=6'h0; in193=6'h0; in194=6'h0; in195=6'h0; in196=6'h0; in197=6'h0; in198=6'h0; in199=6'h6; in200=6'h4; in201=6'h0; in202=6'h0; in203=6'h9; in204=6'h9; in205=6'h0; in206=6'h2; in207=6'h0; in208=6'h0; in209=6'h6; in210=6'h2; in211=6'h2; in212=6'h8; in213=6'h0; in214=6'h0; in215=6'h0; in216=6'h0; in217=6'h0; in218=6'h0; in219=6'h0; in220=6'h0; in221=6'h0; in222=6'h0; in223=6'h0; in224=6'h1; in225=6'h0; in226=6'h0; in227=6'h0; in228=6'h0; in229=6'h4; in230=6'h8; in231=6'h0; in232=6'h0; in233=6'h0; in234=6'h3; in235=6'hA; in236=6'h11; in237=6'hC; in238=6'h0; in239=6'h0; in240=6'h0; in241=6'h0; in242=6'h0; in243=6'h0; in244=6'h0; in245=6'h0; in246=6'h0; in247=6'h0; in248=6'h0; in249=6'h0; in250=6'h0; in251=6'h0; in252=6'h0; in253=6'h1; in254=6'h0; in255=6'hB; in256=6'hB; in257=6'hA; in258=6'h1; in259=6'h7; in260=6'hB; in261=6'h7; in262=6'h4; in263=6'h0; in264=6'h0; in265=6'h0; in266=6'h0; in267=6'h0; in268=6'h0; in269=6'h0; in270=6'h0; in271=6'h0; in272=6'h0; in273=6'h1; in274=6'h0; in275=6'h0; in276=6'h0; in277=6'h4; in278=6'h1; in279=6'h7; in280=6'hC; in281=6'hC; in282=6'h7; in283=6'h0; in284=6'h0; in285=6'h0; in286=6'h0; in287=6'h0; in288=6'h0; in289=6'h5; in290=6'hB; in291=6'hB; in292=6'h3; in293=6'h2; in294=6'h0; in295=6'h0; in296=6'h0; in297=6'h0; in298=6'h0; in299=6'h0; in300=6'h0; in301=6'h0; in302=6'h0; in303=6'h0; in304=6'h0; in305=6'h1; in306=6'h4; in307=6'h4; in308=6'h1; in309=6'h0; in310=6'h0; in311=6'h0; in312=6'h0; in313=6'h0; in314=6'h3; in315=6'h9; in316=6'h0; in317=6'h5; in318=6'h4; in319=6'h5; in320=6'h5; in321=6'h3; in322=6'hE; in323=6'h5; in324=6'h0; in325=6'h0; in326=6'h0; in327=6'h0; in328=6'h0; in329=6'h0; in330=6'h3; in331=6'h0; in332=6'h0; in333=6'h1; in334=6'h1; in335=6'h0; in336=6'h0; in337=6'h0; in338=6'h0; in339=6'h0; in340=6'h2; in341=6'h0; in342=6'h0; in343=6'h0; in344=6'h0; in345=6'h0; in346=6'h0; in347=6'h0; in348=6'h4; in349=6'h1; in350=6'h0; in351=6'h0; in352=6'h0; in353=6'h5; in354=6'h0; in355=6'h0; in356=6'h0; in357=6'h0; in358=6'h0; in359=6'h0; in360=6'h0; in361=6'h0; in362=6'h7; in363=6'h8; in364=6'h4; in365=6'h0; in366=6'h0; in367=6'h2; in368=6'h0; in369=6'h3; in370=6'h4; in371=6'h4; in372=6'h0; in373=6'h0; in374=6'h8; in375=6'h4; in376=6'h0; in377=6'h0; in378=6'h0; in379=6'h7; in380=6'hC; in381=6'h5;
   end
endmodule