module upcount3rst(clk,out);
   input in,clk;
   output out;
   
endmodule
