module test_top(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
   input [9:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12;
   output [11:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10;
   wire signed [10:0] s2_1,s2_2,s2_3,s2_4,s2_5,s2_6,s2_7,s2_8,s2_9,s2_10,s2_11,s2_12,s2_13,s2_14,s2_15;
   wire signed [10:0] h2_1,h2_2,h2_3,h2_4,h2_5,h2_6,h2_7,h2_8,h2_9,h2_10,h2_11,h2_12,h2_13,h2_14,h2_15;
   test_layer_1 L1(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,s2_1,s2_2,s2_3,s2_4,s2_5,s2_6,s2_7,s2_8,s2_9,s2_10,s2_11,s2_12,s2_13,s2_14,s2_15);
   actifunc #(11) AF2_1(s2_1,h2_1);
   actifunc #(11) AF2_2(s2_2,h2_2);
   actifunc #(11) AF2_3(s2_3,h2_3);
   actifunc #(11) AF2_4(s2_4,h2_4);
   actifunc #(11) AF2_5(s2_5,h2_5);
   actifunc #(11) AF2_6(s2_6,h2_6);
   actifunc #(11) AF2_7(s2_7,h2_7);
   actifunc #(11) AF2_8(s2_8,h2_8);
   actifunc #(11) AF2_9(s2_9,h2_9);
   actifunc #(11) AF2_10(s2_10,h2_10);
   actifunc #(11) AF2_11(s2_11,h2_11);
   actifunc #(11) AF2_12(s2_12,h2_12);
   actifunc #(11) AF2_13(s2_13,h2_13);
   actifunc #(11) AF2_14(s2_14,h2_14);
   actifunc #(11) AF2_15(s2_15,h2_15);
   test_layer_2 L2(h2_1[10:0],h2_2[10:0],h2_3[10:0],h2_4[10:0],h2_5[10:0],h2_6[10:0],h2_7[10:0],h2_8[10:0],h2_9[10:0],h2_10[10:0],h2_11[10:0],h2_12[10:0],h2_13[10:0],h2_14[10:0],h2_15[10:0],out1,out2,out3,out4,out5,out6,out7,out8,out9,out10);
endmodule