module lenet300_layer_2(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81,out82,out83,out84,out85,out86,out87,out88,out89,out90,out91,out92,out93,out94,out95,out96,out97,out98,out99,out100);
   input signed [14:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263;
   output signed [14:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81,out82,out83,out84,out85,out86,out87,out88,out89,out90,out91,out92,out93,out94,out95,out96,out97,out98,out99,out100;
   wire signed [14:0] neg1,neg2,neg3,neg4,neg5,neg6,neg7,neg8,neg9,neg10,neg11,neg12,neg13,neg14,neg15,neg16,neg17,neg18,neg19,neg20,neg21,neg22,neg23,neg24,neg25,neg26,neg27,neg28,neg29,neg30,neg31,neg32,neg33,neg34,neg35,neg36,neg37,neg38,neg39,neg40,neg41,neg42,neg43,neg44,neg45,neg46,neg47,neg48,neg49,neg50,neg51,neg52,neg53,neg54,neg55,neg56,neg57,neg58,neg59,neg60,neg61,neg62,neg63,neg64,neg65,neg66,neg67,neg68,neg69,neg70,neg71,neg72,neg73,neg74,neg75,neg76,neg77,neg78,neg79,neg80,neg81,neg82,neg83,neg84,neg85,neg86,neg87,neg88,neg89,neg90,neg91,neg92,neg93,neg94,neg95,neg96,neg97,neg98,neg99,neg100,neg101,neg102,neg103,neg104,neg105,neg106,neg107,neg108,neg109,neg110,neg111,neg112,neg113,neg114,neg115,neg116,neg117,neg118,neg119,neg120,neg121,neg122,neg123,neg124,neg125,neg126,neg127,neg128,neg129,neg130,neg131,neg132,neg133,neg134,neg135,neg136,neg137,neg138,neg139,neg140,neg141,neg142,neg143,neg144,neg145,neg146,neg147,neg148,neg149,neg150,neg151,neg152,neg153,neg154,neg155,neg156,neg157,neg158,neg159,neg160,neg161,neg162,neg163,neg164,neg165,neg166,neg167,neg168,neg169,neg170,neg171,neg172,neg173,neg174,neg175,neg176,neg177,neg178,neg179,neg180,neg181,neg182,neg183,neg184,neg185,neg186,neg187,neg188,neg189,neg190,neg191,neg192,neg193,neg194,neg195,neg196,neg197,neg198,neg199,neg200,neg201,neg202,neg203,neg204,neg205,neg206,neg207,neg208,neg209,neg210,neg211,neg212,neg213,neg214,neg215,neg216,neg217,neg218,neg219,neg220,neg221,neg222,neg223,neg224,neg225,neg226,neg227,neg228,neg229,neg230,neg231,neg232,neg233,neg234,neg235,neg236,neg237,neg238,neg239,neg240,neg241,neg242,neg243,neg244,neg245,neg246,neg247,neg248,neg249,neg250,neg251,neg252,neg253,neg254,neg255,neg256,neg257,neg258,neg259,neg260,neg261,neg262,neg263;

   //Bias value
   wire signed [14:0] b1 = $signed(15'h161);
   wire signed [14:0] b2 = $signed(15'h227);
   wire signed [14:0] b3 = $signed(15'h7E8F);
   wire signed [14:0] b4 = $signed(15'h7B);
   wire signed [14:0] b5 = $signed(15'h190);
   wire signed [14:0] b6 = $signed(15'h7DDE);
   wire signed [14:0] b7 = $signed(15'h7A);
   wire signed [14:0] b8 = $signed(15'h7F14);
   wire signed [14:0] b9 = $signed(15'h7FC8);
   wire signed [14:0] b10 = $signed(15'h26D);
   wire signed [14:0] b11 = $signed(15'h46);
   wire signed [14:0] b12 = $signed(15'h9F);
   wire signed [14:0] b13 = $signed(15'h13C);
   wire signed [14:0] b14 = $signed(15'hDD);
   wire signed [14:0] b15 = $signed(15'h80);
   wire signed [14:0] b16 = $signed(15'h1E7);
   wire signed [14:0] b17 = $signed(15'h7F4D);
   wire signed [14:0] b18 = $signed(15'h7F80);
   wire signed [14:0] b19 = $signed(15'h18A);
   wire signed [14:0] b20 = $signed(15'h7EE8);
   wire signed [14:0] b21 = $signed(15'h7F71);
   wire signed [14:0] b22 = $signed(15'h11D);
   wire signed [14:0] b23 = $signed(15'h7E6A);
   wire signed [14:0] b24 = $signed(15'h7F94);
   wire signed [14:0] b25 = $signed(15'h55);
   wire signed [14:0] b26 = $signed(15'h124);
   wire signed [14:0] b27 = $signed(15'h28A);
   wire signed [14:0] b28 = $signed(15'h7F3F);
   wire signed [14:0] b29 = $signed(15'hCE);
   wire signed [14:0] b30 = $signed(15'h1D1);
   wire signed [14:0] b31 = $signed(15'h2B);
   wire signed [14:0] b32 = $signed(15'h1FB);
   wire signed [14:0] b33 = $signed(15'h1D0);
   wire signed [14:0] b34 = $signed(15'h19);
   wire signed [14:0] b35 = $signed(15'h94);
   wire signed [14:0] b36 = $signed(15'h2D);
   wire signed [14:0] b37 = $signed(15'h7DFD);
   wire signed [14:0] b38 = $signed(15'h18C);
   wire signed [14:0] b39 = $signed(15'h1D3);
   wire signed [14:0] b40 = $signed(15'h7FCF);
   wire signed [14:0] b41 = $signed(15'h7E5B);
   wire signed [14:0] b42 = $signed(15'hCC);
   wire signed [14:0] b43 = $signed(15'h2AE);
   wire signed [14:0] b44 = $signed(15'h9C);
   wire signed [14:0] b45 = $signed(15'h7E80);
   wire signed [14:0] b46 = $signed(15'h215);
   wire signed [14:0] b47 = $signed(15'h16);
   wire signed [14:0] b48 = $signed(15'h7F5E);
   wire signed [14:0] b49 = $signed(15'h7F64);
   wire signed [14:0] b50 = $signed(15'h7FDB);
   wire signed [14:0] b51 = $signed(15'h7DE6);
   wire signed [14:0] b52 = $signed(15'h7E0D);
   wire signed [14:0] b53 = $signed(15'h7F25);
   wire signed [14:0] b54 = $signed(15'h7FC6);
   wire signed [14:0] b55 = $signed(15'h7FA8);
   wire signed [14:0] b56 = $signed(15'h7EEF);
   wire signed [14:0] b57 = $signed(15'hBD);
   wire signed [14:0] b58 = $signed(15'h7ED2);
   wire signed [14:0] b59 = $signed(15'h25);
   wire signed [14:0] b60 = $signed(15'h7EA2);
   wire signed [14:0] b61 = $signed(15'h12);
   wire signed [14:0] b62 = $signed(15'h7F30);
   wire signed [14:0] b63 = $signed(15'h1AF);
   wire signed [14:0] b64 = $signed(15'h7FAE);
   wire signed [14:0] b65 = $signed(15'h233);
   wire signed [14:0] b66 = $signed(15'h1AD);
   wire signed [14:0] b67 = $signed(15'hF0);
   wire signed [14:0] b68 = $signed(15'h7F9A);
   wire signed [14:0] b69 = $signed(15'h9B);
   wire signed [14:0] b70 = $signed(15'h7EC0);
   wire signed [14:0] b71 = $signed(15'h7E3A);
   wire signed [14:0] b72 = $signed(15'h7FF2);
   wire signed [14:0] b73 = $signed(15'h7FB7);
   wire signed [14:0] b74 = $signed(15'h7FB0);
   wire signed [14:0] b75 = $signed(15'h7FC1);
   wire signed [14:0] b76 = $signed(15'h146);
   wire signed [14:0] b77 = $signed(15'h7F4B);
   wire signed [14:0] b78 = $signed(15'h7EF6);
   wire signed [14:0] b79 = $signed(15'hD1);
   wire signed [14:0] b80 = $signed(15'h135);
   wire signed [14:0] b81 = $signed(15'h7FEE);
   wire signed [14:0] b82 = $signed(15'h252);
   wire signed [14:0] b83 = $signed(15'h9A);
   wire signed [14:0] b84 = $signed(15'h13C);
   wire signed [14:0] b85 = $signed(15'h7FD8);
   wire signed [14:0] b86 = $signed(15'hD0);
   wire signed [14:0] b87 = $signed(15'h7F67);
   wire signed [14:0] b88 = $signed(15'h7DB5);
   wire signed [14:0] b89 = $signed(15'h7E5A);
   wire signed [14:0] b90 = $signed(15'h196);
   wire signed [14:0] b91 = $signed(15'h7DFA);
   wire signed [14:0] b92 = $signed(15'hD4);
   wire signed [14:0] b93 = $signed(15'h7EFB);
   wire signed [14:0] b94 = $signed(15'h1A4);
   wire signed [14:0] b95 = $signed(15'h3A);
   wire signed [14:0] b96 = $signed(15'h7D76);
   wire signed [14:0] b97 = $signed(15'h359);
   wire signed [14:0] b98 = $signed(15'h7F3A);
   wire signed [14:0] b99 = $signed(15'h7F50);
   wire signed [14:0] b100 = $signed(15'h120);

   //Negation modules
   negate #(15) N1(in1,neg1);
   negate #(15) N2(in2,neg2);
   negate #(15) N3(in3,neg3);
   negate #(15) N4(in4,neg4);
   negate #(15) N5(in5,neg5);
   negate #(15) N6(in6,neg6);
   negate #(15) N7(in7,neg7);
   negate #(15) N8(in8,neg8);
   negate #(15) N9(in9,neg9);
   negate #(15) N10(in10,neg10);
   negate #(15) N11(in11,neg11);
   negate #(15) N12(in12,neg12);
   negate #(15) N13(in13,neg13);
   negate #(15) N14(in14,neg14);
   negate #(15) N15(in15,neg15);
   negate #(15) N16(in16,neg16);
   negate #(15) N17(in17,neg17);
   negate #(15) N18(in18,neg18);
   negate #(15) N19(in19,neg19);
   negate #(15) N20(in20,neg20);
   negate #(15) N21(in21,neg21);
   negate #(15) N22(in22,neg22);
   negate #(15) N23(in23,neg23);
   negate #(15) N24(in24,neg24);
   negate #(15) N25(in25,neg25);
   negate #(15) N26(in26,neg26);
   negate #(15) N27(in27,neg27);
   negate #(15) N28(in28,neg28);
   negate #(15) N29(in29,neg29);
   negate #(15) N30(in30,neg30);
   negate #(15) N31(in31,neg31);
   negate #(15) N32(in32,neg32);
   negate #(15) N33(in33,neg33);
   negate #(15) N34(in34,neg34);
   negate #(15) N35(in35,neg35);
   negate #(15) N36(in36,neg36);
   negate #(15) N37(in37,neg37);
   negate #(15) N38(in38,neg38);
   negate #(15) N39(in39,neg39);
   negate #(15) N40(in40,neg40);
   negate #(15) N41(in41,neg41);
   negate #(15) N42(in42,neg42);
   negate #(15) N43(in43,neg43);
   negate #(15) N44(in44,neg44);
   negate #(15) N45(in45,neg45);
   negate #(15) N46(in46,neg46);
   negate #(15) N47(in47,neg47);
   negate #(15) N48(in48,neg48);
   negate #(15) N49(in49,neg49);
   negate #(15) N50(in50,neg50);
   negate #(15) N51(in51,neg51);
   negate #(15) N52(in52,neg52);
   negate #(15) N53(in53,neg53);
   negate #(15) N54(in54,neg54);
   negate #(15) N55(in55,neg55);
   negate #(15) N56(in56,neg56);
   negate #(15) N57(in57,neg57);
   negate #(15) N58(in58,neg58);
   negate #(15) N59(in59,neg59);
   negate #(15) N60(in60,neg60);
   negate #(15) N61(in61,neg61);
   negate #(15) N62(in62,neg62);
   negate #(15) N63(in63,neg63);
   negate #(15) N64(in64,neg64);
   negate #(15) N65(in65,neg65);
   negate #(15) N66(in66,neg66);
   negate #(15) N67(in67,neg67);
   negate #(15) N68(in68,neg68);
   negate #(15) N69(in69,neg69);
   negate #(15) N70(in70,neg70);
   negate #(15) N71(in71,neg71);
   negate #(15) N72(in72,neg72);
   negate #(15) N73(in73,neg73);
   negate #(15) N74(in74,neg74);
   negate #(15) N75(in75,neg75);
   negate #(15) N76(in76,neg76);
   negate #(15) N77(in77,neg77);
   negate #(15) N78(in78,neg78);
   negate #(15) N79(in79,neg79);
   negate #(15) N80(in80,neg80);
   negate #(15) N81(in81,neg81);
   negate #(15) N82(in82,neg82);
   negate #(15) N83(in83,neg83);
   negate #(15) N84(in84,neg84);
   negate #(15) N85(in85,neg85);
   negate #(15) N86(in86,neg86);
   negate #(15) N87(in87,neg87);
   negate #(15) N88(in88,neg88);
   negate #(15) N89(in89,neg89);
   negate #(15) N90(in90,neg90);
   negate #(15) N91(in91,neg91);
   negate #(15) N92(in92,neg92);
   negate #(15) N93(in93,neg93);
   negate #(15) N94(in94,neg94);
   negate #(15) N95(in95,neg95);
   negate #(15) N96(in96,neg96);
   negate #(15) N97(in97,neg97);
   negate #(15) N98(in98,neg98);
   negate #(15) N99(in99,neg99);
   negate #(15) N100(in100,neg100);
   negate #(15) N101(in101,neg101);
   negate #(15) N102(in102,neg102);
   negate #(15) N103(in103,neg103);
   negate #(15) N104(in104,neg104);
   negate #(15) N105(in105,neg105);
   negate #(15) N106(in106,neg106);
   negate #(15) N107(in107,neg107);
   negate #(15) N108(in108,neg108);
   negate #(15) N109(in109,neg109);
   negate #(15) N110(in110,neg110);
   negate #(15) N111(in111,neg111);
   negate #(15) N112(in112,neg112);
   negate #(15) N113(in113,neg113);
   negate #(15) N114(in114,neg114);
   negate #(15) N115(in115,neg115);
   negate #(15) N116(in116,neg116);
   negate #(15) N117(in117,neg117);
   negate #(15) N118(in118,neg118);
   negate #(15) N119(in119,neg119);
   negate #(15) N120(in120,neg120);
   negate #(15) N121(in121,neg121);
   negate #(15) N122(in122,neg122);
   negate #(15) N123(in123,neg123);
   negate #(15) N124(in124,neg124);
   negate #(15) N125(in125,neg125);
   negate #(15) N126(in126,neg126);
   negate #(15) N127(in127,neg127);
   negate #(15) N128(in128,neg128);
   negate #(15) N129(in129,neg129);
   negate #(15) N130(in130,neg130);
   negate #(15) N131(in131,neg131);
   negate #(15) N132(in132,neg132);
   negate #(15) N133(in133,neg133);
   negate #(15) N134(in134,neg134);
   negate #(15) N135(in135,neg135);
   negate #(15) N136(in136,neg136);
   negate #(15) N137(in137,neg137);
   negate #(15) N138(in138,neg138);
   negate #(15) N139(in139,neg139);
   negate #(15) N140(in140,neg140);
   negate #(15) N141(in141,neg141);
   negate #(15) N142(in142,neg142);
   negate #(15) N143(in143,neg143);
   negate #(15) N144(in144,neg144);
   negate #(15) N145(in145,neg145);
   negate #(15) N146(in146,neg146);
   negate #(15) N147(in147,neg147);
   negate #(15) N148(in148,neg148);
   negate #(15) N149(in149,neg149);
   negate #(15) N150(in150,neg150);
   negate #(15) N151(in151,neg151);
   negate #(15) N152(in152,neg152);
   negate #(15) N153(in153,neg153);
   negate #(15) N154(in154,neg154);
   negate #(15) N155(in155,neg155);
   negate #(15) N156(in156,neg156);
   negate #(15) N157(in157,neg157);
   negate #(15) N158(in158,neg158);
   negate #(15) N159(in159,neg159);
   negate #(15) N160(in160,neg160);
   negate #(15) N161(in161,neg161);
   negate #(15) N162(in162,neg162);
   negate #(15) N163(in163,neg163);
   negate #(15) N164(in164,neg164);
   negate #(15) N165(in165,neg165);
   negate #(15) N166(in166,neg166);
   negate #(15) N167(in167,neg167);
   negate #(15) N168(in168,neg168);
   negate #(15) N169(in169,neg169);
   negate #(15) N170(in170,neg170);
   negate #(15) N171(in171,neg171);
   negate #(15) N172(in172,neg172);
   negate #(15) N173(in173,neg173);
   negate #(15) N174(in174,neg174);
   negate #(15) N175(in175,neg175);
   negate #(15) N176(in176,neg176);
   negate #(15) N177(in177,neg177);
   negate #(15) N178(in178,neg178);
   negate #(15) N179(in179,neg179);
   negate #(15) N180(in180,neg180);
   negate #(15) N181(in181,neg181);
   negate #(15) N182(in182,neg182);
   negate #(15) N183(in183,neg183);
   negate #(15) N184(in184,neg184);
   negate #(15) N185(in185,neg185);
   negate #(15) N186(in186,neg186);
   negate #(15) N187(in187,neg187);
   negate #(15) N188(in188,neg188);
   negate #(15) N189(in189,neg189);
   negate #(15) N190(in190,neg190);
   negate #(15) N191(in191,neg191);
   negate #(15) N192(in192,neg192);
   negate #(15) N193(in193,neg193);
   negate #(15) N194(in194,neg194);
   negate #(15) N195(in195,neg195);
   negate #(15) N196(in196,neg196);
   negate #(15) N197(in197,neg197);
   negate #(15) N198(in198,neg198);
   negate #(15) N199(in199,neg199);
   negate #(15) N200(in200,neg200);
   negate #(15) N201(in201,neg201);
   negate #(15) N202(in202,neg202);
   negate #(15) N203(in203,neg203);
   negate #(15) N204(in204,neg204);
   negate #(15) N205(in205,neg205);
   negate #(15) N206(in206,neg206);
   negate #(15) N207(in207,neg207);
   negate #(15) N208(in208,neg208);
   negate #(15) N209(in209,neg209);
   negate #(15) N210(in210,neg210);
   negate #(15) N211(in211,neg211);
   negate #(15) N212(in212,neg212);
   negate #(15) N213(in213,neg213);
   negate #(15) N214(in214,neg214);
   negate #(15) N215(in215,neg215);
   negate #(15) N216(in216,neg216);
   negate #(15) N217(in217,neg217);
   negate #(15) N218(in218,neg218);
   negate #(15) N219(in219,neg219);
   negate #(15) N220(in220,neg220);
   negate #(15) N221(in221,neg221);
   negate #(15) N222(in222,neg222);
   negate #(15) N223(in223,neg223);
   negate #(15) N224(in224,neg224);
   negate #(15) N225(in225,neg225);
   negate #(15) N226(in226,neg226);
   negate #(15) N227(in227,neg227);
   negate #(15) N228(in228,neg228);
   negate #(15) N229(in229,neg229);
   negate #(15) N230(in230,neg230);
   negate #(15) N231(in231,neg231);
   negate #(15) N232(in232,neg232);
   negate #(15) N233(in233,neg233);
   negate #(15) N234(in234,neg234);
   negate #(15) N235(in235,neg235);
   negate #(15) N236(in236,neg236);
   negate #(15) N237(in237,neg237);
   negate #(15) N238(in238,neg238);
   negate #(15) N239(in239,neg239);
   negate #(15) N240(in240,neg240);
   negate #(15) N241(in241,neg241);
   negate #(15) N242(in242,neg242);
   negate #(15) N243(in243,neg243);
   negate #(15) N244(in244,neg244);
   negate #(15) N245(in245,neg245);
   negate #(15) N246(in246,neg246);
   negate #(15) N247(in247,neg247);
   negate #(15) N248(in248,neg248);
   negate #(15) N249(in249,neg249);
   negate #(15) N250(in250,neg250);
   negate #(15) N251(in251,neg251);
   negate #(15) N252(in252,neg252);
   negate #(15) N253(in253,neg253);
   negate #(15) N254(in254,neg254);
   negate #(15) N255(in255,neg255);
   negate #(15) N256(in256,neg256);
   negate #(15) N257(in257,neg257);
   negate #(15) N258(in258,neg258);
   negate #(15) N259(in259,neg259);
   negate #(15) N260(in260,neg260);
   negate #(15) N261(in261,neg261);
   negate #(15) N262(in262,neg262);
   negate #(15) N263(in263,neg263);

   // m1_1 = W*in
   wire signed [14:0] m1_1;
   assign m1_1 =15'b0;

   // m1_2 = W*in
   wire signed [14:0] m1_2;
   assign m1_2 =15'b0;

   // m1_3 = W*in
   wire signed [14:0] m1_3;
   assign m1_3 =15'b0;

   // m1_4 = W*in
   wire signed [14:0] m1_4;
   assign m1_4 =15'b0;

   // m1_5 = W*in
   wire signed [14:0] m1_5;
   assign m1_5 =15'b0;

   // m1_6 = W*in
   wire signed [14:0] m1_6;
   assign m1_6 =15'b0;

   // m1_7 = W*in
   wire signed [14:0] m1_7;
   assign m1_7 ={ {3{in1[14]}} , in1[14:3] };

   // m1_8 = W*in
   wire signed [14:0] m1_8;
   assign m1_8 =15'b0;

   // m1_9 = W*in
   wire signed [14:0] m1_9;
   assign m1_9 =15'b0;

   // m1_10 = W*in
   wire signed [14:0] m1_10;
   assign m1_10 =15'b0;

   // m1_11 = W*in
   wire signed [14:0] m1_11;
   assign m1_11 =15'b0;

   // m1_12 = W*in
   wire signed [14:0] m1_12;
   assign m1_12 =15'b0;

   // m1_13 = W*in
   wire signed [14:0] m1_13;
   assign m1_13 =15'b0;

   // m1_14 = W*in
   wire signed [14:0] m1_14;
   assign m1_14 =15'b0;

   // m1_15 = W*in
   wire signed [14:0] m1_15;
   assign m1_15 =15'b0;

   // m1_16 = W*in
   wire signed [14:0] m1_16;
   assign m1_16 =15'b0;

   // m1_17 = W*in
   wire signed [14:0] m1_17;
   assign m1_17 =15'b0;

   // m1_18 = W*in
   wire signed [14:0] m1_18;
   assign m1_18 =15'b0;

   // m1_19 = W*in
   wire signed [14:0] m1_19;
   assign m1_19 ={ {4{in1[14]}} , in1[14:4] };

   // m1_20 = W*in
   wire signed [14:0] m1_20;
   assign m1_20 =15'b0;

   // m1_21 = W*in
   wire signed [14:0] m1_21;
   assign m1_21 =15'b0;

   // m1_22 = W*in
   wire signed [14:0] m1_22;
   assign m1_22 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_23 = W*in
   wire signed [14:0] m1_23;
   assign m1_23 =15'b0;

   // m1_24 = W*in
   wire signed [14:0] m1_24;
   assign m1_24 =15'b0;

   // m1_25 = W*in
   wire signed [14:0] m1_25;
   assign m1_25 ={ {3{neg1[14]}} , neg1[14:3] };

   // m1_26 = W*in
   wire signed [14:0] m1_26;
   assign m1_26 =15'b0;

   // m1_27 = W*in
   wire signed [14:0] m1_27;
   assign m1_27 =15'b0;

   // m1_28 = W*in
   wire signed [14:0] m1_28;
   assign m1_28 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_29 = W*in
   wire signed [14:0] m1_29;
   assign m1_29 =15'b0;

   // m1_30 = W*in
   wire signed [14:0] m1_30;
   assign m1_30 =15'b0;

   // m1_31 = W*in
   wire signed [14:0] m1_31;
   assign m1_31 =15'b0;

   // m1_32 = W*in
   wire signed [14:0] m1_32;
   assign m1_32 ={ {3{in1[14]}} , in1[14:3] };

   // m1_33 = W*in
   wire signed [14:0] m1_33;
   assign m1_33 ={ {4{in1[14]}} , in1[14:4] };

   // m1_34 = W*in
   wire signed [14:0] m1_34;
   assign m1_34 =15'b0;

   // m1_35 = W*in
   wire signed [14:0] m1_35;
   assign m1_35 ={ {3{in1[14]}} , in1[14:3] };

   // m1_36 = W*in
   wire signed [14:0] m1_36;
   assign m1_36 =15'b0;

   // m1_37 = W*in
   wire signed [14:0] m1_37;
   assign m1_37 =15'b0;

   // m1_38 = W*in
   wire signed [14:0] m1_38;
   assign m1_38 =15'b0;

   // m1_39 = W*in
   wire signed [14:0] m1_39;
   assign m1_39 =15'b0;

   // m1_40 = W*in
   wire signed [14:0] m1_40;
   assign m1_40 =15'b0;

   // m1_41 = W*in
   wire signed [14:0] m1_41;
   assign m1_41 =15'b0;

   // m1_42 = W*in
   wire signed [14:0] m1_42;
   assign m1_42 ={ {3{in1[14]}} , in1[14:3] };

   // m1_43 = W*in
   wire signed [14:0] m1_43;
   assign m1_43 =15'b0;

   // m1_44 = W*in
   wire signed [14:0] m1_44;
   assign m1_44 =15'b0;

   // m1_45 = W*in
   wire signed [14:0] m1_45;
   assign m1_45 =15'b0;

   // m1_46 = W*in
   wire signed [14:0] m1_46;
   assign m1_46 =15'b0;

   // m1_47 = W*in
   wire signed [14:0] m1_47;
   assign m1_47 ={ {4{in1[14]}} , in1[14:4] };

   // m1_48 = W*in
   wire signed [14:0] m1_48;
   assign m1_48 =15'b0;

   // m1_49 = W*in
   wire signed [14:0] m1_49;
   assign m1_49 ={ {3{neg1[14]}} , neg1[14:3] };

   // m1_50 = W*in
   wire signed [14:0] m1_50;
   assign m1_50 =15'b0;

   // m1_51 = W*in
   wire signed [14:0] m1_51;
   assign m1_51 =15'b0;

   // m1_52 = W*in
   wire signed [14:0] m1_52;
   assign m1_52 =15'b0;

   // m1_53 = W*in
   wire signed [14:0] m1_53;
   assign m1_53 =15'b0;

   // m1_54 = W*in
   wire signed [14:0] m1_54;
   assign m1_54 =15'b0;

   // m1_55 = W*in
   wire signed [14:0] m1_55;
   assign m1_55 =15'b0;

   // m1_56 = W*in
   wire signed [14:0] m1_56;
   assign m1_56 ={ {3{in1[14]}} , in1[14:3] };

   // m1_57 = W*in
   wire signed [14:0] m1_57;
   assign m1_57 =15'b0;

   // m1_58 = W*in
   wire signed [14:0] m1_58;
   assign m1_58 ={ {3{neg1[14]}} , neg1[14:3] };

   // m1_59 = W*in
   wire signed [14:0] m1_59;
   assign m1_59 =15'b0;

   // m1_60 = W*in
   wire signed [14:0] m1_60;
   assign m1_60 =15'b0;

   // m1_61 = W*in
   wire signed [14:0] m1_61;
   assign m1_61 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_62 = W*in
   wire signed [14:0] m1_62;
   assign m1_62 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_63 = W*in
   wire signed [14:0] m1_63;
   assign m1_63 =15'b0;

   // m1_64 = W*in
   wire signed [14:0] m1_64;
   assign m1_64 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_65 = W*in
   wire signed [14:0] m1_65;
   assign m1_65 ={ {3{neg1[14]}} , neg1[14:3] };

   // m1_66 = W*in
   wire signed [14:0] m1_66;
   assign m1_66 ={ {4{in1[14]}} , in1[14:4] };

   // m1_67 = W*in
   wire signed [14:0] m1_67;
   assign m1_67 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_68 = W*in
   wire signed [14:0] m1_68;
   assign m1_68 =15'b0;

   // m1_69 = W*in
   wire signed [14:0] m1_69;
   assign m1_69 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_70 = W*in
   wire signed [14:0] m1_70;
   assign m1_70 ={ {3{in1[14]}} , in1[14:3] };

   // m1_71 = W*in
   wire signed [14:0] m1_71;
   assign m1_71 =15'b0;

   // m1_72 = W*in
   wire signed [14:0] m1_72;
   assign m1_72 =15'b0;

   // m1_73 = W*in
   wire signed [14:0] m1_73;
   assign m1_73 =15'b0;

   // m1_74 = W*in
   wire signed [14:0] m1_74;
   assign m1_74 =15'b0;

   // m1_75 = W*in
   wire signed [14:0] m1_75;
   assign m1_75 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_76 = W*in
   wire signed [14:0] m1_76;
   assign m1_76 =15'b0;

   // m1_77 = W*in
   wire signed [14:0] m1_77;
   assign m1_77 ={ {4{neg1[14]}} , neg1[14:4] };

   // m1_78 = W*in
   wire signed [14:0] m1_78;
   assign m1_78 =15'b0;

   // m1_79 = W*in
   wire signed [14:0] m1_79;
   assign m1_79 ={ {4{in1[14]}} , in1[14:4] };

   // m1_80 = W*in
   wire signed [14:0] m1_80;
   assign m1_80 =15'b0;

   // m1_81 = W*in
   wire signed [14:0] m1_81;
   assign m1_81 =15'b0;

   // m1_82 = W*in
   wire signed [14:0] m1_82;
   assign m1_82 =15'b0;

   // m1_83 = W*in
   wire signed [14:0] m1_83;
   assign m1_83 =15'b0;

   // m1_84 = W*in
   wire signed [14:0] m1_84;
   assign m1_84 =15'b0;

   // m1_85 = W*in
   wire signed [14:0] m1_85;
   assign m1_85 =15'b0;

   // m1_86 = W*in
   wire signed [14:0] m1_86;
   assign m1_86 =15'b0;

   // m1_87 = W*in
   wire signed [14:0] m1_87;
   assign m1_87 =15'b0;

   // m1_88 = W*in
   wire signed [14:0] m1_88;
   assign m1_88 =15'b0;

   // m1_89 = W*in
   wire signed [14:0] m1_89;
   assign m1_89 =15'b0;

   // m1_90 = W*in
   wire signed [14:0] m1_90;
   assign m1_90 =15'b0;

   // m1_91 = W*in
   wire signed [14:0] m1_91;
   assign m1_91 =15'b0;

   // m1_92 = W*in
   wire signed [14:0] m1_92;
   assign m1_92 =15'b0;

   // m1_93 = W*in
   wire signed [14:0] m1_93;
   assign m1_93 =15'b0;

   // m1_94 = W*in
   wire signed [14:0] m1_94;
   assign m1_94 ={ {4{in1[14]}} , in1[14:4] };

   // m1_95 = W*in
   wire signed [14:0] m1_95;
   assign m1_95 =15'b0;

   // m1_96 = W*in
   wire signed [14:0] m1_96;
   assign m1_96 =15'b0;

   // m1_97 = W*in
   wire signed [14:0] m1_97;
   assign m1_97 =15'b0;

   // m1_98 = W*in
   wire signed [14:0] m1_98;
   assign m1_98 =15'b0;

   // m1_99 = W*in
   wire signed [14:0] m1_99;
   assign m1_99 =15'b0;

   // m1_100 = W*in
   wire signed [14:0] m1_100;
   assign m1_100 =15'b0;

   // m2_1 = W*in
   wire signed [14:0] m2_1;
   assign m2_1 =15'b0;

   // m2_2 = W*in
   wire signed [14:0] m2_2;
   assign m2_2 =15'b0;

   // m2_3 = W*in
   wire signed [14:0] m2_3;
   assign m2_3 =15'b0;

   // m2_4 = W*in
   wire signed [14:0] m2_4;
   assign m2_4 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_5 = W*in
   wire signed [14:0] m2_5;
   assign m2_5 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_6 = W*in
   wire signed [14:0] m2_6;
   assign m2_6 =15'b0;

   // m2_7 = W*in
   wire signed [14:0] m2_7;
   assign m2_7 =15'b0;

   // m2_8 = W*in
   wire signed [14:0] m2_8;
   assign m2_8 ={ {3{in2[14]}} , in2[14:3] };

   // m2_9 = W*in
   wire signed [14:0] m2_9;
   assign m2_9 ={ {3{in2[14]}} , in2[14:3] };

   // m2_10 = W*in
   wire signed [14:0] m2_10;
   assign m2_10 =15'b0;

   // m2_11 = W*in
   wire signed [14:0] m2_11;
   assign m2_11 =15'b0;

   // m2_12 = W*in
   wire signed [14:0] m2_12;
   assign m2_12 =15'b0;

   // m2_13 = W*in
   wire signed [14:0] m2_13;
   assign m2_13 =15'b0;

   // m2_14 = W*in
   wire signed [14:0] m2_14;
   assign m2_14 =15'b0;

   // m2_15 = W*in
   wire signed [14:0] m2_15;
   assign m2_15 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_16 = W*in
   wire signed [14:0] m2_16;
   assign m2_16 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_17 = W*in
   wire signed [14:0] m2_17;
   assign m2_17 =15'b0;

   // m2_18 = W*in
   wire signed [14:0] m2_18;
   assign m2_18 =15'b0;

   // m2_19 = W*in
   wire signed [14:0] m2_19;
   assign m2_19 ={ {4{in2[14]}} , in2[14:4] };

   // m2_20 = W*in
   wire signed [14:0] m2_20;
   assign m2_20 ={ {3{in2[14]}} , in2[14:3] };

   // m2_21 = W*in
   wire signed [14:0] m2_21;
   assign m2_21 ={ {3{in2[14]}} , in2[14:3] };

   // m2_22 = W*in
   wire signed [14:0] m2_22;
   assign m2_22 =15'b0;

   // m2_23 = W*in
   wire signed [14:0] m2_23;
   assign m2_23 ={ {3{in2[14]}} , in2[14:3] };

   // m2_24 = W*in
   wire signed [14:0] m2_24;
   assign m2_24 =15'b0;

   // m2_25 = W*in
   wire signed [14:0] m2_25;
   assign m2_25 =15'b0;

   // m2_26 = W*in
   wire signed [14:0] m2_26;
   assign m2_26 ={ {4{neg2[14]}} , neg2[14:4] };

   // m2_27 = W*in
   wire signed [14:0] m2_27;
   assign m2_27 ={ {4{neg2[14]}} , neg2[14:4] };

   // m2_28 = W*in
   wire signed [14:0] m2_28;
   assign m2_28 =15'b0;

   // m2_29 = W*in
   wire signed [14:0] m2_29;
   assign m2_29 ={ {4{neg2[14]}} , neg2[14:4] };

   // m2_30 = W*in
   wire signed [14:0] m2_30;
   assign m2_30 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_31 = W*in
   wire signed [14:0] m2_31;
   assign m2_31 =15'b0;

   // m2_32 = W*in
   wire signed [14:0] m2_32;
   assign m2_32 ={ {4{neg2[14]}} , neg2[14:4] };

   // m2_33 = W*in
   wire signed [14:0] m2_33;
   assign m2_33 =15'b0;

   // m2_34 = W*in
   wire signed [14:0] m2_34;
   assign m2_34 =15'b0;

   // m2_35 = W*in
   wire signed [14:0] m2_35;
   assign m2_35 =15'b0;

   // m2_36 = W*in
   wire signed [14:0] m2_36;
   assign m2_36 =15'b0;

   // m2_37 = W*in
   wire signed [14:0] m2_37;
   assign m2_37 ={ {2{in2[14]}} , in2[14:2] };

   // m2_38 = W*in
   wire signed [14:0] m2_38;
   assign m2_38 =15'b0;

   // m2_39 = W*in
   wire signed [14:0] m2_39;
   assign m2_39 =15'b0;

   // m2_40 = W*in
   wire signed [14:0] m2_40;
   assign m2_40 =15'b0;

   // m2_41 = W*in
   wire signed [14:0] m2_41;
   assign m2_41 ={ {4{in2[14]}} , in2[14:4] };

   // m2_42 = W*in
   wire signed [14:0] m2_42;
   assign m2_42 =15'b0;

   // m2_43 = W*in
   wire signed [14:0] m2_43;
   assign m2_43 =15'b0;

   // m2_44 = W*in
   wire signed [14:0] m2_44;
   assign m2_44 ={ {3{in2[14]}} , in2[14:3] };

   // m2_45 = W*in
   wire signed [14:0] m2_45;
   assign m2_45 ={ {3{in2[14]}} , in2[14:3] };

   // m2_46 = W*in
   wire signed [14:0] m2_46;
   assign m2_46 =15'b0;

   // m2_47 = W*in
   wire signed [14:0] m2_47;
   assign m2_47 ={ {3{in2[14]}} , in2[14:3] };

   // m2_48 = W*in
   wire signed [14:0] m2_48;
   assign m2_48 =15'b0;

   // m2_49 = W*in
   wire signed [14:0] m2_49;
   assign m2_49 =15'b0;

   // m2_50 = W*in
   wire signed [14:0] m2_50;
   assign m2_50 =15'b0;

   // m2_51 = W*in
   wire signed [14:0] m2_51;
   assign m2_51 ={ {3{in2[14]}} , in2[14:3] };

   // m2_52 = W*in
   wire signed [14:0] m2_52;
   assign m2_52 =15'b0;

   // m2_53 = W*in
   wire signed [14:0] m2_53;
   assign m2_53 ={ {3{in2[14]}} , in2[14:3] };

   // m2_54 = W*in
   wire signed [14:0] m2_54;
   assign m2_54 =15'b0;

   // m2_55 = W*in
   wire signed [14:0] m2_55;
   assign m2_55 =15'b0;

   // m2_56 = W*in
   wire signed [14:0] m2_56;
   assign m2_56 ={ {3{in2[14]}} , in2[14:3] };

   // m2_57 = W*in
   wire signed [14:0] m2_57;
   assign m2_57 =15'b0;

   // m2_58 = W*in
   wire signed [14:0] m2_58;
   assign m2_58 =15'b0;

   // m2_59 = W*in
   wire signed [14:0] m2_59;
   assign m2_59 ={ {3{in2[14]}} , in2[14:3] };

   // m2_60 = W*in
   wire signed [14:0] m2_60;
   assign m2_60 =15'b0;

   // m2_61 = W*in
   wire signed [14:0] m2_61;
   assign m2_61 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_62 = W*in
   wire signed [14:0] m2_62;
   assign m2_62 =15'b0;

   // m2_63 = W*in
   wire signed [14:0] m2_63;
   assign m2_63 =15'b0;

   // m2_64 = W*in
   wire signed [14:0] m2_64;
   assign m2_64 ={ {3{in2[14]}} , in2[14:3] };

   // m2_65 = W*in
   wire signed [14:0] m2_65;
   assign m2_65 =15'b0;

   // m2_66 = W*in
   wire signed [14:0] m2_66;
   assign m2_66 ={ {4{neg2[14]}} , neg2[14:4] };

   // m2_67 = W*in
   wire signed [14:0] m2_67;
   assign m2_67 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_68 = W*in
   wire signed [14:0] m2_68;
   assign m2_68 =15'b0;

   // m2_69 = W*in
   wire signed [14:0] m2_69;
   assign m2_69 =15'b0;

   // m2_70 = W*in
   wire signed [14:0] m2_70;
   assign m2_70 ={ {3{in2[14]}} , in2[14:3] };

   // m2_71 = W*in
   wire signed [14:0] m2_71;
   assign m2_71 ={ {4{in2[14]}} , in2[14:4] };

   // m2_72 = W*in
   wire signed [14:0] m2_72;
   assign m2_72 =15'b0;

   // m2_73 = W*in
   wire signed [14:0] m2_73;
   assign m2_73 =15'b0;

   // m2_74 = W*in
   wire signed [14:0] m2_74;
   assign m2_74 ={ {3{in2[14]}} , in2[14:3] };

   // m2_75 = W*in
   wire signed [14:0] m2_75;
   assign m2_75 ={ {3{in2[14]}} , in2[14:3] };

   // m2_76 = W*in
   wire signed [14:0] m2_76;
   assign m2_76 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_77 = W*in
   wire signed [14:0] m2_77;
   assign m2_77 =15'b0;

   // m2_78 = W*in
   wire signed [14:0] m2_78;
   assign m2_78 =15'b0;

   // m2_79 = W*in
   wire signed [14:0] m2_79;
   assign m2_79 =15'b0;

   // m2_80 = W*in
   wire signed [14:0] m2_80;
   assign m2_80 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_81 = W*in
   wire signed [14:0] m2_81;
   assign m2_81 =15'b0;

   // m2_82 = W*in
   wire signed [14:0] m2_82;
   assign m2_82 ={ {3{neg2[14]}} , neg2[14:3] };

   // m2_83 = W*in
   wire signed [14:0] m2_83;
   assign m2_83 =15'b0;

   // m2_84 = W*in
   wire signed [14:0] m2_84;
   assign m2_84 =15'b0;

   // m2_85 = W*in
   wire signed [14:0] m2_85;
   assign m2_85 =15'b0;

   // m2_86 = W*in
   wire signed [14:0] m2_86;
   assign m2_86 =15'b0;

   // m2_87 = W*in
   wire signed [14:0] m2_87;
   assign m2_87 =15'b0;

   // m2_88 = W*in
   wire signed [14:0] m2_88;
   assign m2_88 ={ {2{in2[14]}} , in2[14:2] };

   // m2_89 = W*in
   wire signed [14:0] m2_89;
   assign m2_89 ={ {3{in2[14]}} , in2[14:3] };

   // m2_90 = W*in
   wire signed [14:0] m2_90;
   assign m2_90 =15'b0;

   // m2_91 = W*in
   wire signed [14:0] m2_91;
   assign m2_91 =15'b0;

   // m2_92 = W*in
   wire signed [14:0] m2_92;
   assign m2_92 =15'b0;

   // m2_93 = W*in
   wire signed [14:0] m2_93;
   assign m2_93 =15'b0;

   // m2_94 = W*in
   wire signed [14:0] m2_94;
   assign m2_94 =15'b0;

   // m2_95 = W*in
   wire signed [14:0] m2_95;
   assign m2_95 =15'b0;

   // m2_96 = W*in
   wire signed [14:0] m2_96;
   assign m2_96 =15'b0;

   // m2_97 = W*in
   wire signed [14:0] m2_97;
   assign m2_97 =15'b0;

   // m2_98 = W*in
   wire signed [14:0] m2_98;
   assign m2_98 =15'b0;

   // m2_99 = W*in
   wire signed [14:0] m2_99;
   assign m2_99 ={ {3{in2[14]}} , in2[14:3] };

   // m2_100 = W*in
   wire signed [14:0] m2_100;
   assign m2_100 =15'b0;

   // m3_1 = W*in
   wire signed [14:0] m3_1;
   assign m3_1 =15'b0;

   // m3_2 = W*in
   wire signed [14:0] m3_2;
   assign m3_2 =15'b0;

   // m3_3 = W*in
   wire signed [14:0] m3_3;
   assign m3_3 =15'b0;

   // m3_4 = W*in
   wire signed [14:0] m3_4;
   assign m3_4 =15'b0;

   // m3_5 = W*in
   wire signed [14:0] m3_5;
   assign m3_5 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_6 = W*in
   wire signed [14:0] m3_6;
   assign m3_6 =15'b0;

   // m3_7 = W*in
   wire signed [14:0] m3_7;
   assign m3_7 =15'b0;

   // m3_8 = W*in
   wire signed [14:0] m3_8;
   assign m3_8 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_9 = W*in
   wire signed [14:0] m3_9;
   assign m3_9 =15'b0;

   // m3_10 = W*in
   wire signed [14:0] m3_10;
   assign m3_10 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_11 = W*in
   wire signed [14:0] m3_11;
   assign m3_11 =15'b0;

   // m3_12 = W*in
   wire signed [14:0] m3_12;
   assign m3_12 =15'b0;

   // m3_13 = W*in
   wire signed [14:0] m3_13;
   assign m3_13 ={ {3{in3[14]}} , in3[14:3] };

   // m3_14 = W*in
   wire signed [14:0] m3_14;
   assign m3_14 =15'b0;

   // m3_15 = W*in
   wire signed [14:0] m3_15;
   assign m3_15 =15'b0;

   // m3_16 = W*in
   wire signed [14:0] m3_16;
   assign m3_16 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_17 = W*in
   wire signed [14:0] m3_17;
   assign m3_17 =15'b0;

   // m3_18 = W*in
   wire signed [14:0] m3_18;
   assign m3_18 =15'b0;

   // m3_19 = W*in
   wire signed [14:0] m3_19;
   assign m3_19 =15'b0;

   // m3_20 = W*in
   wire signed [14:0] m3_20;
   assign m3_20 =15'b0;

   // m3_21 = W*in
   wire signed [14:0] m3_21;
   assign m3_21 =15'b0;

   // m3_22 = W*in
   wire signed [14:0] m3_22;
   assign m3_22 =15'b0;

   // m3_23 = W*in
   wire signed [14:0] m3_23;
   assign m3_23 =15'b0;

   // m3_24 = W*in
   wire signed [14:0] m3_24;
   assign m3_24 =15'b0;

   // m3_25 = W*in
   wire signed [14:0] m3_25;
   assign m3_25 =15'b0;

   // m3_26 = W*in
   wire signed [14:0] m3_26;
   assign m3_26 =15'b0;

   // m3_27 = W*in
   wire signed [14:0] m3_27;
   assign m3_27 =15'b0;

   // m3_28 = W*in
   wire signed [14:0] m3_28;
   assign m3_28 ={ {2{in3[14]}} , in3[14:2] };

   // m3_29 = W*in
   wire signed [14:0] m3_29;
   assign m3_29 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_30 = W*in
   wire signed [14:0] m3_30;
   assign m3_30 =15'b0;

   // m3_31 = W*in
   wire signed [14:0] m3_31;
   assign m3_31 =15'b0;

   // m3_32 = W*in
   wire signed [14:0] m3_32;
   assign m3_32 =15'b0;

   // m3_33 = W*in
   wire signed [14:0] m3_33;
   assign m3_33 =15'b0;

   // m3_34 = W*in
   wire signed [14:0] m3_34;
   assign m3_34 =15'b0;

   // m3_35 = W*in
   wire signed [14:0] m3_35;
   assign m3_35 =15'b0;

   // m3_36 = W*in
   wire signed [14:0] m3_36;
   assign m3_36 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_37 = W*in
   wire signed [14:0] m3_37;
   assign m3_37 =15'b0;

   // m3_38 = W*in
   wire signed [14:0] m3_38;
   assign m3_38 =15'b0;

   // m3_39 = W*in
   wire signed [14:0] m3_39;
   assign m3_39 ={ {3{in3[14]}} , in3[14:3] };

   // m3_40 = W*in
   wire signed [14:0] m3_40;
   assign m3_40 =15'b0;

   // m3_41 = W*in
   wire signed [14:0] m3_41;
   assign m3_41 ={ {3{in3[14]}} , in3[14:3] };

   // m3_42 = W*in
   wire signed [14:0] m3_42;
   assign m3_42 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_43 = W*in
   wire signed [14:0] m3_43;
   assign m3_43 =15'b0;

   // m3_44 = W*in
   wire signed [14:0] m3_44;
   assign m3_44 =15'b0;

   // m3_45 = W*in
   wire signed [14:0] m3_45;
   assign m3_45 ={ {3{in3[14]}} , in3[14:3] };

   // m3_46 = W*in
   wire signed [14:0] m3_46;
   assign m3_46 =15'b0;

   // m3_47 = W*in
   wire signed [14:0] m3_47;
   assign m3_47 =15'b0;

   // m3_48 = W*in
   wire signed [14:0] m3_48;
   assign m3_48 =15'b0;

   // m3_49 = W*in
   wire signed [14:0] m3_49;
   assign m3_49 =15'b0;

   // m3_50 = W*in
   wire signed [14:0] m3_50;
   assign m3_50 =15'b0;

   // m3_51 = W*in
   wire signed [14:0] m3_51;
   assign m3_51 =15'b0;

   // m3_52 = W*in
   wire signed [14:0] m3_52;
   assign m3_52 =15'b0;

   // m3_53 = W*in
   wire signed [14:0] m3_53;
   assign m3_53 =15'b0;

   // m3_54 = W*in
   wire signed [14:0] m3_54;
   assign m3_54 =15'b0;

   // m3_55 = W*in
   wire signed [14:0] m3_55;
   assign m3_55 =15'b0;

   // m3_56 = W*in
   wire signed [14:0] m3_56;
   assign m3_56 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_57 = W*in
   wire signed [14:0] m3_57;
   assign m3_57 =15'b0;

   // m3_58 = W*in
   wire signed [14:0] m3_58;
   assign m3_58 =15'b0;

   // m3_59 = W*in
   wire signed [14:0] m3_59;
   assign m3_59 =15'b0;

   // m3_60 = W*in
   wire signed [14:0] m3_60;
   assign m3_60 =15'b0;

   // m3_61 = W*in
   wire signed [14:0] m3_61;
   assign m3_61 =15'b0;

   // m3_62 = W*in
   wire signed [14:0] m3_62;
   assign m3_62 =15'b0;

   // m3_63 = W*in
   wire signed [14:0] m3_63;
   assign m3_63 =15'b0;

   // m3_64 = W*in
   wire signed [14:0] m3_64;
   assign m3_64 =15'b0;

   // m3_65 = W*in
   wire signed [14:0] m3_65;
   assign m3_65 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_66 = W*in
   wire signed [14:0] m3_66;
   assign m3_66 =15'b0;

   // m3_67 = W*in
   wire signed [14:0] m3_67;
   assign m3_67 =15'b0;

   // m3_68 = W*in
   wire signed [14:0] m3_68;
   assign m3_68 =15'b0;

   // m3_69 = W*in
   wire signed [14:0] m3_69;
   assign m3_69 =15'b0;

   // m3_70 = W*in
   wire signed [14:0] m3_70;
   assign m3_70 =15'b0;

   // m3_71 = W*in
   wire signed [14:0] m3_71;
   assign m3_71 =15'b0;

   // m3_72 = W*in
   wire signed [14:0] m3_72;
   assign m3_72 =15'b0;

   // m3_73 = W*in
   wire signed [14:0] m3_73;
   assign m3_73 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_74 = W*in
   wire signed [14:0] m3_74;
   assign m3_74 =15'b0;

   // m3_75 = W*in
   wire signed [14:0] m3_75;
   assign m3_75 =15'b0;

   // m3_76 = W*in
   wire signed [14:0] m3_76;
   assign m3_76 =15'b0;

   // m3_77 = W*in
   wire signed [14:0] m3_77;
   assign m3_77 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_78 = W*in
   wire signed [14:0] m3_78;
   assign m3_78 =15'b0;

   // m3_79 = W*in
   wire signed [14:0] m3_79;
   assign m3_79 ={ {3{neg3[14]}} , neg3[14:3] };

   // m3_80 = W*in
   wire signed [14:0] m3_80;
   assign m3_80 =15'b0;

   // m3_81 = W*in
   wire signed [14:0] m3_81;
   assign m3_81 =15'b0;

   // m3_82 = W*in
   wire signed [14:0] m3_82;
   assign m3_82 =15'b0;

   // m3_83 = W*in
   wire signed [14:0] m3_83;
   assign m3_83 =15'b0;

   // m3_84 = W*in
   wire signed [14:0] m3_84;
   assign m3_84 =15'b0;

   // m3_85 = W*in
   wire signed [14:0] m3_85;
   assign m3_85 =15'b0;

   // m3_86 = W*in
   wire signed [14:0] m3_86;
   assign m3_86 ={ {3{in3[14]}} , in3[14:3] };

   // m3_87 = W*in
   wire signed [14:0] m3_87;
   assign m3_87 =15'b0;

   // m3_88 = W*in
   wire signed [14:0] m3_88;
   assign m3_88 =15'b0;

   // m3_89 = W*in
   wire signed [14:0] m3_89;
   assign m3_89 =15'b0;

   // m3_90 = W*in
   wire signed [14:0] m3_90;
   assign m3_90 =15'b0;

   // m3_91 = W*in
   wire signed [14:0] m3_91;
   assign m3_91 =15'b0;

   // m3_92 = W*in
   wire signed [14:0] m3_92;
   assign m3_92 =15'b0;

   // m3_93 = W*in
   wire signed [14:0] m3_93;
   assign m3_93 =15'b0;

   // m3_94 = W*in
   wire signed [14:0] m3_94;
   assign m3_94 =15'b0;

   // m3_95 = W*in
   wire signed [14:0] m3_95;
   assign m3_95 =15'b0;

   // m3_96 = W*in
   wire signed [14:0] m3_96;
   assign m3_96 =15'b0;

   // m3_97 = W*in
   wire signed [14:0] m3_97;
   assign m3_97 =15'b0;

   // m3_98 = W*in
   wire signed [14:0] m3_98;
   assign m3_98 =15'b0;

   // m3_99 = W*in
   wire signed [14:0] m3_99;
   assign m3_99 =15'b0;

   // m3_100 = W*in
   wire signed [14:0] m3_100;
   assign m3_100 =15'b0;

   // m4_1 = W*in
   wire signed [14:0] m4_1;
   assign m4_1 =15'b0;

   // m4_2 = W*in
   wire signed [14:0] m4_2;
   assign m4_2 =15'b0;

   // m4_3 = W*in
   wire signed [14:0] m4_3;
   assign m4_3 =15'b0;

   // m4_4 = W*in
   wire signed [14:0] m4_4;
   assign m4_4 =15'b0;

   // m4_5 = W*in
   wire signed [14:0] m4_5;
   assign m4_5 ={ {3{neg4[14]}} , neg4[14:3] };

   // m4_6 = W*in
   wire signed [14:0] m4_6;
   assign m4_6 =15'b0;

   // m4_7 = W*in
   wire signed [14:0] m4_7;
   assign m4_7 =15'b0;

   // m4_8 = W*in
   wire signed [14:0] m4_8;
   assign m4_8 =15'b0;

   // m4_9 = W*in
   wire signed [14:0] m4_9;
   assign m4_9 =15'b0;

   // m4_10 = W*in
   wire signed [14:0] m4_10;
   assign m4_10 =15'b0;

   // m4_11 = W*in
   wire signed [14:0] m4_11;
   assign m4_11 =15'b0;

   // m4_12 = W*in
   wire signed [14:0] m4_12;
   assign m4_12 =15'b0;

   // m4_13 = W*in
   wire signed [14:0] m4_13;
   assign m4_13 =15'b0;

   // m4_14 = W*in
   wire signed [14:0] m4_14;
   assign m4_14 =15'b0;

   // m4_15 = W*in
   wire signed [14:0] m4_15;
   assign m4_15 =15'b0;

   // m4_16 = W*in
   wire signed [14:0] m4_16;
   assign m4_16 =15'b0;

   // m4_17 = W*in
   wire signed [14:0] m4_17;
   assign m4_17 =15'b0;

   // m4_18 = W*in
   wire signed [14:0] m4_18;
   assign m4_18 ={ {4{in4[14]}} , in4[14:4] };

   // m4_19 = W*in
   wire signed [14:0] m4_19;
   assign m4_19 =15'b0;

   // m4_20 = W*in
   wire signed [14:0] m4_20;
   assign m4_20 =15'b0;

   // m4_21 = W*in
   wire signed [14:0] m4_21;
   assign m4_21 ={ {3{in4[14]}} , in4[14:3] };

   // m4_22 = W*in
   wire signed [14:0] m4_22;
   assign m4_22 =15'b0;

   // m4_23 = W*in
   wire signed [14:0] m4_23;
   assign m4_23 =15'b0;

   // m4_24 = W*in
   wire signed [14:0] m4_24;
   assign m4_24 =15'b0;

   // m4_25 = W*in
   wire signed [14:0] m4_25;
   assign m4_25 =15'b0;

   // m4_26 = W*in
   wire signed [14:0] m4_26;
   assign m4_26 =15'b0;

   // m4_27 = W*in
   wire signed [14:0] m4_27;
   assign m4_27 =15'b0;

   // m4_28 = W*in
   wire signed [14:0] m4_28;
   assign m4_28 =15'b0;

   // m4_29 = W*in
   wire signed [14:0] m4_29;
   assign m4_29 =15'b0;

   // m4_30 = W*in
   wire signed [14:0] m4_30;
   assign m4_30 =15'b0;

   // m4_31 = W*in
   wire signed [14:0] m4_31;
   assign m4_31 =15'b0;

   // m4_32 = W*in
   wire signed [14:0] m4_32;
   assign m4_32 =15'b0;

   // m4_33 = W*in
   wire signed [14:0] m4_33;
   assign m4_33 =15'b0;

   // m4_34 = W*in
   wire signed [14:0] m4_34;
   assign m4_34 =15'b0;

   // m4_35 = W*in
   wire signed [14:0] m4_35;
   assign m4_35 =15'b0;

   // m4_36 = W*in
   wire signed [14:0] m4_36;
   assign m4_36 =15'b0;

   // m4_37 = W*in
   wire signed [14:0] m4_37;
   assign m4_37 =15'b0;

   // m4_38 = W*in
   wire signed [14:0] m4_38;
   assign m4_38 =15'b0;

   // m4_39 = W*in
   wire signed [14:0] m4_39;
   assign m4_39 =15'b0;

   // m4_40 = W*in
   wire signed [14:0] m4_40;
   assign m4_40 =15'b0;

   // m4_41 = W*in
   wire signed [14:0] m4_41;
   assign m4_41 =15'b0;

   // m4_42 = W*in
   wire signed [14:0] m4_42;
   assign m4_42 =15'b0;

   // m4_43 = W*in
   wire signed [14:0] m4_43;
   assign m4_43 =15'b0;

   // m4_44 = W*in
   wire signed [14:0] m4_44;
   assign m4_44 ={ {3{in4[14]}} , in4[14:3] };

   // m4_45 = W*in
   wire signed [14:0] m4_45;
   assign m4_45 =15'b0;

   // m4_46 = W*in
   wire signed [14:0] m4_46;
   assign m4_46 =15'b0;

   // m4_47 = W*in
   wire signed [14:0] m4_47;
   assign m4_47 =15'b0;

   // m4_48 = W*in
   wire signed [14:0] m4_48;
   assign m4_48 =15'b0;

   // m4_49 = W*in
   wire signed [14:0] m4_49;
   assign m4_49 =15'b0;

   // m4_50 = W*in
   wire signed [14:0] m4_50;
   assign m4_50 =15'b0;

   // m4_51 = W*in
   wire signed [14:0] m4_51;
   assign m4_51 =15'b0;

   // m4_52 = W*in
   wire signed [14:0] m4_52;
   assign m4_52 =15'b0;

   // m4_53 = W*in
   wire signed [14:0] m4_53;
   assign m4_53 =15'b0;

   // m4_54 = W*in
   wire signed [14:0] m4_54;
   assign m4_54 ={ {3{neg4[14]}} , neg4[14:3] };

   // m4_55 = W*in
   wire signed [14:0] m4_55;
   assign m4_55 =15'b0;

   // m4_56 = W*in
   wire signed [14:0] m4_56;
   assign m4_56 =15'b0;

   // m4_57 = W*in
   wire signed [14:0] m4_57;
   assign m4_57 =15'b0;

   // m4_58 = W*in
   wire signed [14:0] m4_58;
   assign m4_58 ={ {4{neg4[14]}} , neg4[14:4] };

   // m4_59 = W*in
   wire signed [14:0] m4_59;
   assign m4_59 =15'b0;

   // m4_60 = W*in
   wire signed [14:0] m4_60;
   assign m4_60 ={ {2{in4[14]}} , in4[14:2] };

   // m4_61 = W*in
   wire signed [14:0] m4_61;
   assign m4_61 ={ {3{neg4[14]}} , neg4[14:3] };

   // m4_62 = W*in
   wire signed [14:0] m4_62;
   assign m4_62 =15'b0;

   // m4_63 = W*in
   wire signed [14:0] m4_63;
   assign m4_63 =15'b0;

   // m4_64 = W*in
   wire signed [14:0] m4_64;
   assign m4_64 =15'b0;

   // m4_65 = W*in
   wire signed [14:0] m4_65;
   assign m4_65 =15'b0;

   // m4_66 = W*in
   wire signed [14:0] m4_66;
   assign m4_66 =15'b0;

   // m4_67 = W*in
   wire signed [14:0] m4_67;
   assign m4_67 ={ {3{in4[14]}} , in4[14:3] };

   // m4_68 = W*in
   wire signed [14:0] m4_68;
   assign m4_68 =15'b0;

   // m4_69 = W*in
   wire signed [14:0] m4_69;
   assign m4_69 =15'b0;

   // m4_70 = W*in
   wire signed [14:0] m4_70;
   assign m4_70 =15'b0;

   // m4_71 = W*in
   wire signed [14:0] m4_71;
   assign m4_71 =15'b0;

   // m4_72 = W*in
   wire signed [14:0] m4_72;
   assign m4_72 =15'b0;

   // m4_73 = W*in
   wire signed [14:0] m4_73;
   assign m4_73 =15'b0;

   // m4_74 = W*in
   wire signed [14:0] m4_74;
   assign m4_74 =15'b0;

   // m4_75 = W*in
   wire signed [14:0] m4_75;
   assign m4_75 =15'b0;

   // m4_76 = W*in
   wire signed [14:0] m4_76;
   assign m4_76 =15'b0;

   // m4_77 = W*in
   wire signed [14:0] m4_77;
   assign m4_77 =15'b0;

   // m4_78 = W*in
   wire signed [14:0] m4_78;
   assign m4_78 ={ {4{in4[14]}} , in4[14:4] };

   // m4_79 = W*in
   wire signed [14:0] m4_79;
   assign m4_79 =15'b0;

   // m4_80 = W*in
   wire signed [14:0] m4_80;
   assign m4_80 =15'b0;

   // m4_81 = W*in
   wire signed [14:0] m4_81;
   assign m4_81 =15'b0;

   // m4_82 = W*in
   wire signed [14:0] m4_82;
   assign m4_82 =15'b0;

   // m4_83 = W*in
   wire signed [14:0] m4_83;
   assign m4_83 =15'b0;

   // m4_84 = W*in
   wire signed [14:0] m4_84;
   assign m4_84 =15'b0;

   // m4_85 = W*in
   wire signed [14:0] m4_85;
   assign m4_85 =15'b0;

   // m4_86 = W*in
   wire signed [14:0] m4_86;
   assign m4_86 ={ {3{in4[14]}} , in4[14:3] };

   // m4_87 = W*in
   wire signed [14:0] m4_87;
   assign m4_87 =15'b0;

   // m4_88 = W*in
   wire signed [14:0] m4_88;
   assign m4_88 =15'b0;

   // m4_89 = W*in
   wire signed [14:0] m4_89;
   assign m4_89 =15'b0;

   // m4_90 = W*in
   wire signed [14:0] m4_90;
   assign m4_90 =15'b0;

   // m4_91 = W*in
   wire signed [14:0] m4_91;
   assign m4_91 =15'b0;

   // m4_92 = W*in
   wire signed [14:0] m4_92;
   assign m4_92 =15'b0;

   // m4_93 = W*in
   wire signed [14:0] m4_93;
   assign m4_93 =15'b0;

   // m4_94 = W*in
   wire signed [14:0] m4_94;
   assign m4_94 =15'b0;

   // m4_95 = W*in
   wire signed [14:0] m4_95;
   assign m4_95 ={ {3{in4[14]}} , in4[14:3] };

   // m4_96 = W*in
   wire signed [14:0] m4_96;
   assign m4_96 =15'b0;

   // m4_97 = W*in
   wire signed [14:0] m4_97;
   assign m4_97 =15'b0;

   // m4_98 = W*in
   wire signed [14:0] m4_98;
   assign m4_98 =15'b0;

   // m4_99 = W*in
   wire signed [14:0] m4_99;
   assign m4_99 =15'b0;

   // m4_100 = W*in
   wire signed [14:0] m4_100;
   assign m4_100 =15'b0;

   // m5_1 = W*in
   wire signed [14:0] m5_1;
   assign m5_1 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_2 = W*in
   wire signed [14:0] m5_2;
   assign m5_2 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_3 = W*in
   wire signed [14:0] m5_3;
   assign m5_3 ={ {3{in5[14]}} , in5[14:3] };

   // m5_4 = W*in
   wire signed [14:0] m5_4;
   assign m5_4 =15'b0;

   // m5_5 = W*in
   wire signed [14:0] m5_5;
   assign m5_5 =15'b0;

   // m5_6 = W*in
   wire signed [14:0] m5_6;
   assign m5_6 =15'b0;

   // m5_7 = W*in
   wire signed [14:0] m5_7;
   assign m5_7 =15'b0;

   // m5_8 = W*in
   wire signed [14:0] m5_8;
   assign m5_8 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_9 = W*in
   wire signed [14:0] m5_9;
   assign m5_9 =15'b0;

   // m5_10 = W*in
   wire signed [14:0] m5_10;
   assign m5_10 =15'b0;

   // m5_11 = W*in
   wire signed [14:0] m5_11;
   assign m5_11 =15'b0;

   // m5_12 = W*in
   wire signed [14:0] m5_12;
   assign m5_12 =15'b0;

   // m5_13 = W*in
   wire signed [14:0] m5_13;
   assign m5_13 =15'b0;

   // m5_14 = W*in
   wire signed [14:0] m5_14;
   assign m5_14 =15'b0;

   // m5_15 = W*in
   wire signed [14:0] m5_15;
   assign m5_15 =15'b0;

   // m5_16 = W*in
   wire signed [14:0] m5_16;
   assign m5_16 =15'b0;

   // m5_17 = W*in
   wire signed [14:0] m5_17;
   assign m5_17 ={ {3{in5[14]}} , in5[14:3] };

   // m5_18 = W*in
   wire signed [14:0] m5_18;
   assign m5_18 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_19 = W*in
   wire signed [14:0] m5_19;
   assign m5_19 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_20 = W*in
   wire signed [14:0] m5_20;
   assign m5_20 =15'b0;

   // m5_21 = W*in
   wire signed [14:0] m5_21;
   assign m5_21 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_22 = W*in
   wire signed [14:0] m5_22;
   assign m5_22 =15'b0;

   // m5_23 = W*in
   wire signed [14:0] m5_23;
   assign m5_23 =15'b0;

   // m5_24 = W*in
   wire signed [14:0] m5_24;
   assign m5_24 =15'b0;

   // m5_25 = W*in
   wire signed [14:0] m5_25;
   assign m5_25 =15'b0;

   // m5_26 = W*in
   wire signed [14:0] m5_26;
   assign m5_26 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_27 = W*in
   wire signed [14:0] m5_27;
   assign m5_27 =15'b0;

   // m5_28 = W*in
   wire signed [14:0] m5_28;
   assign m5_28 =15'b0;

   // m5_29 = W*in
   wire signed [14:0] m5_29;
   assign m5_29 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_30 = W*in
   wire signed [14:0] m5_30;
   assign m5_30 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_31 = W*in
   wire signed [14:0] m5_31;
   assign m5_31 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_32 = W*in
   wire signed [14:0] m5_32;
   assign m5_32 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_33 = W*in
   wire signed [14:0] m5_33;
   assign m5_33 =15'b0;

   // m5_34 = W*in
   wire signed [14:0] m5_34;
   assign m5_34 =15'b0;

   // m5_35 = W*in
   wire signed [14:0] m5_35;
   assign m5_35 =15'b0;

   // m5_36 = W*in
   wire signed [14:0] m5_36;
   assign m5_36 =15'b0;

   // m5_37 = W*in
   wire signed [14:0] m5_37;
   assign m5_37 =15'b0;

   // m5_38 = W*in
   wire signed [14:0] m5_38;
   assign m5_38 =15'b0;

   // m5_39 = W*in
   wire signed [14:0] m5_39;
   assign m5_39 ={ {3{in5[14]}} , in5[14:3] };

   // m5_40 = W*in
   wire signed [14:0] m5_40;
   assign m5_40 =15'b0;

   // m5_41 = W*in
   wire signed [14:0] m5_41;
   assign m5_41 =15'b0;

   // m5_42 = W*in
   wire signed [14:0] m5_42;
   assign m5_42 =15'b0;

   // m5_43 = W*in
   wire signed [14:0] m5_43;
   assign m5_43 =15'b0;

   // m5_44 = W*in
   wire signed [14:0] m5_44;
   assign m5_44 =15'b0;

   // m5_45 = W*in
   wire signed [14:0] m5_45;
   assign m5_45 ={ {3{in5[14]}} , in5[14:3] };

   // m5_46 = W*in
   wire signed [14:0] m5_46;
   assign m5_46 =15'b0;

   // m5_47 = W*in
   wire signed [14:0] m5_47;
   assign m5_47 =15'b0;

   // m5_48 = W*in
   wire signed [14:0] m5_48;
   assign m5_48 =15'b0;

   // m5_49 = W*in
   wire signed [14:0] m5_49;
   assign m5_49 ={ {3{in5[14]}} , in5[14:3] };

   // m5_50 = W*in
   wire signed [14:0] m5_50;
   assign m5_50 =15'b0;

   // m5_51 = W*in
   wire signed [14:0] m5_51;
   assign m5_51 =15'b0;

   // m5_52 = W*in
   wire signed [14:0] m5_52;
   assign m5_52 =15'b0;

   // m5_53 = W*in
   wire signed [14:0] m5_53;
   assign m5_53 =15'b0;

   // m5_54 = W*in
   wire signed [14:0] m5_54;
   assign m5_54 ={ {3{in5[14]}} , in5[14:3] };

   // m5_55 = W*in
   wire signed [14:0] m5_55;
   assign m5_55 =15'b0;

   // m5_56 = W*in
   wire signed [14:0] m5_56;
   assign m5_56 ={ {3{in5[14]}} , in5[14:3] };

   // m5_57 = W*in
   wire signed [14:0] m5_57;
   assign m5_57 =15'b0;

   // m5_58 = W*in
   wire signed [14:0] m5_58;
   assign m5_58 ={ {4{in5[14]}} , in5[14:4] };

   // m5_59 = W*in
   wire signed [14:0] m5_59;
   assign m5_59 =15'b0;

   // m5_60 = W*in
   wire signed [14:0] m5_60;
   assign m5_60 ={ {4{in5[14]}} , in5[14:4] };

   // m5_61 = W*in
   wire signed [14:0] m5_61;
   assign m5_61 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_62 = W*in
   wire signed [14:0] m5_62;
   assign m5_62 ={ {4{in5[14]}} , in5[14:4] };

   // m5_63 = W*in
   wire signed [14:0] m5_63;
   assign m5_63 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_64 = W*in
   wire signed [14:0] m5_64;
   assign m5_64 =15'b0;

   // m5_65 = W*in
   wire signed [14:0] m5_65;
   assign m5_65 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_66 = W*in
   wire signed [14:0] m5_66;
   assign m5_66 ={ {4{in5[14]}} , in5[14:4] };

   // m5_67 = W*in
   wire signed [14:0] m5_67;
   assign m5_67 =15'b0;

   // m5_68 = W*in
   wire signed [14:0] m5_68;
   assign m5_68 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_69 = W*in
   wire signed [14:0] m5_69;
   assign m5_69 =15'b0;

   // m5_70 = W*in
   wire signed [14:0] m5_70;
   assign m5_70 ={ {3{in5[14]}} , in5[14:3] };

   // m5_71 = W*in
   wire signed [14:0] m5_71;
   assign m5_71 =15'b0;

   // m5_72 = W*in
   wire signed [14:0] m5_72;
   assign m5_72 =15'b0;

   // m5_73 = W*in
   wire signed [14:0] m5_73;
   assign m5_73 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_74 = W*in
   wire signed [14:0] m5_74;
   assign m5_74 =15'b0;

   // m5_75 = W*in
   wire signed [14:0] m5_75;
   assign m5_75 ={ {4{in5[14]}} , in5[14:4] };

   // m5_76 = W*in
   wire signed [14:0] m5_76;
   assign m5_76 =15'b0;

   // m5_77 = W*in
   wire signed [14:0] m5_77;
   assign m5_77 =15'b0;

   // m5_78 = W*in
   wire signed [14:0] m5_78;
   assign m5_78 =15'b0;

   // m5_79 = W*in
   wire signed [14:0] m5_79;
   assign m5_79 ={ {4{neg5[14]}} , neg5[14:4] };

   // m5_80 = W*in
   wire signed [14:0] m5_80;
   assign m5_80 =15'b0;

   // m5_81 = W*in
   wire signed [14:0] m5_81;
   assign m5_81 =15'b0;

   // m5_82 = W*in
   wire signed [14:0] m5_82;
   assign m5_82 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_83 = W*in
   wire signed [14:0] m5_83;
   assign m5_83 =15'b0;

   // m5_84 = W*in
   wire signed [14:0] m5_84;
   assign m5_84 =15'b0;

   // m5_85 = W*in
   wire signed [14:0] m5_85;
   assign m5_85 =15'b0;

   // m5_86 = W*in
   wire signed [14:0] m5_86;
   assign m5_86 =15'b0;

   // m5_87 = W*in
   wire signed [14:0] m5_87;
   assign m5_87 =15'b0;

   // m5_88 = W*in
   wire signed [14:0] m5_88;
   assign m5_88 =15'b0;

   // m5_89 = W*in
   wire signed [14:0] m5_89;
   assign m5_89 =15'b0;

   // m5_90 = W*in
   wire signed [14:0] m5_90;
   assign m5_90 =15'b0;

   // m5_91 = W*in
   wire signed [14:0] m5_91;
   assign m5_91 =15'b0;

   // m5_92 = W*in
   wire signed [14:0] m5_92;
   assign m5_92 =15'b0;

   // m5_93 = W*in
   wire signed [14:0] m5_93;
   assign m5_93 =15'b0;

   // m5_94 = W*in
   wire signed [14:0] m5_94;
   assign m5_94 =15'b0;

   // m5_95 = W*in
   wire signed [14:0] m5_95;
   assign m5_95 =15'b0;

   // m5_96 = W*in
   wire signed [14:0] m5_96;
   assign m5_96 =15'b0;

   // m5_97 = W*in
   wire signed [14:0] m5_97;
   assign m5_97 ={ {3{neg5[14]}} , neg5[14:3] };

   // m5_98 = W*in
   wire signed [14:0] m5_98;
   assign m5_98 =15'b0;

   // m5_99 = W*in
   wire signed [14:0] m5_99;
   assign m5_99 =15'b0;

   // m5_100 = W*in
   wire signed [14:0] m5_100;
   assign m5_100 =15'b0;

   // m6_1 = W*in
   wire signed [14:0] m6_1;
   assign m6_1 =15'b0;

   // m6_2 = W*in
   wire signed [14:0] m6_2;
   assign m6_2 =15'b0;

   // m6_3 = W*in
   wire signed [14:0] m6_3;
   assign m6_3 =15'b0;

   // m6_4 = W*in
   wire signed [14:0] m6_4;
   assign m6_4 =15'b0;

   // m6_5 = W*in
   wire signed [14:0] m6_5;
   assign m6_5 =15'b0;

   // m6_6 = W*in
   wire signed [14:0] m6_6;
   assign m6_6 =15'b0;

   // m6_7 = W*in
   wire signed [14:0] m6_7;
   assign m6_7 =15'b0;

   // m6_8 = W*in
   wire signed [14:0] m6_8;
   assign m6_8 =15'b0;

   // m6_9 = W*in
   wire signed [14:0] m6_9;
   assign m6_9 =15'b0;

   // m6_10 = W*in
   wire signed [14:0] m6_10;
   assign m6_10 =15'b0;

   // m6_11 = W*in
   wire signed [14:0] m6_11;
   assign m6_11 =15'b0;

   // m6_12 = W*in
   wire signed [14:0] m6_12;
   assign m6_12 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_13 = W*in
   wire signed [14:0] m6_13;
   assign m6_13 =15'b0;

   // m6_14 = W*in
   wire signed [14:0] m6_14;
   assign m6_14 =15'b0;

   // m6_15 = W*in
   wire signed [14:0] m6_15;
   assign m6_15 =15'b0;

   // m6_16 = W*in
   wire signed [14:0] m6_16;
   assign m6_16 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_17 = W*in
   wire signed [14:0] m6_17;
   assign m6_17 =15'b0;

   // m6_18 = W*in
   wire signed [14:0] m6_18;
   assign m6_18 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_19 = W*in
   wire signed [14:0] m6_19;
   assign m6_19 =15'b0;

   // m6_20 = W*in
   wire signed [14:0] m6_20;
   assign m6_20 =15'b0;

   // m6_21 = W*in
   wire signed [14:0] m6_21;
   assign m6_21 =15'b0;

   // m6_22 = W*in
   wire signed [14:0] m6_22;
   assign m6_22 =15'b0;

   // m6_23 = W*in
   wire signed [14:0] m6_23;
   assign m6_23 =15'b0;

   // m6_24 = W*in
   wire signed [14:0] m6_24;
   assign m6_24 =15'b0;

   // m6_25 = W*in
   wire signed [14:0] m6_25;
   assign m6_25 =15'b0;

   // m6_26 = W*in
   wire signed [14:0] m6_26;
   assign m6_26 =15'b0;

   // m6_27 = W*in
   wire signed [14:0] m6_27;
   assign m6_27 =15'b0;

   // m6_28 = W*in
   wire signed [14:0] m6_28;
   assign m6_28 =15'b0;

   // m6_29 = W*in
   wire signed [14:0] m6_29;
   assign m6_29 =15'b0;

   // m6_30 = W*in
   wire signed [14:0] m6_30;
   assign m6_30 ={ {4{in6[14]}} , in6[14:4] };

   // m6_31 = W*in
   wire signed [14:0] m6_31;
   assign m6_31 =15'b0;

   // m6_32 = W*in
   wire signed [14:0] m6_32;
   assign m6_32 =15'b0;

   // m6_33 = W*in
   wire signed [14:0] m6_33;
   assign m6_33 =15'b0;

   // m6_34 = W*in
   wire signed [14:0] m6_34;
   assign m6_34 =15'b0;

   // m6_35 = W*in
   wire signed [14:0] m6_35;
   assign m6_35 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_36 = W*in
   wire signed [14:0] m6_36;
   assign m6_36 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_37 = W*in
   wire signed [14:0] m6_37;
   assign m6_37 =15'b0;

   // m6_38 = W*in
   wire signed [14:0] m6_38;
   assign m6_38 =15'b0;

   // m6_39 = W*in
   wire signed [14:0] m6_39;
   assign m6_39 =15'b0;

   // m6_40 = W*in
   wire signed [14:0] m6_40;
   assign m6_40 =15'b0;

   // m6_41 = W*in
   wire signed [14:0] m6_41;
   assign m6_41 =15'b0;

   // m6_42 = W*in
   wire signed [14:0] m6_42;
   assign m6_42 =15'b0;

   // m6_43 = W*in
   wire signed [14:0] m6_43;
   assign m6_43 =15'b0;

   // m6_44 = W*in
   wire signed [14:0] m6_44;
   assign m6_44 =15'b0;

   // m6_45 = W*in
   wire signed [14:0] m6_45;
   assign m6_45 ={ {3{in6[14]}} , in6[14:3] };

   // m6_46 = W*in
   wire signed [14:0] m6_46;
   assign m6_46 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_47 = W*in
   wire signed [14:0] m6_47;
   assign m6_47 =15'b0;

   // m6_48 = W*in
   wire signed [14:0] m6_48;
   assign m6_48 =15'b0;

   // m6_49 = W*in
   wire signed [14:0] m6_49;
   assign m6_49 ={ {3{in6[14]}} , in6[14:3] };

   // m6_50 = W*in
   wire signed [14:0] m6_50;
   assign m6_50 ={ {3{in6[14]}} , in6[14:3] };

   // m6_51 = W*in
   wire signed [14:0] m6_51;
   assign m6_51 =15'b0;

   // m6_52 = W*in
   wire signed [14:0] m6_52;
   assign m6_52 =15'b0;

   // m6_53 = W*in
   wire signed [14:0] m6_53;
   assign m6_53 =15'b0;

   // m6_54 = W*in
   wire signed [14:0] m6_54;
   assign m6_54 =15'b0;

   // m6_55 = W*in
   wire signed [14:0] m6_55;
   assign m6_55 ={ {3{in6[14]}} , in6[14:3] };

   // m6_56 = W*in
   wire signed [14:0] m6_56;
   assign m6_56 =15'b0;

   // m6_57 = W*in
   wire signed [14:0] m6_57;
   assign m6_57 =15'b0;

   // m6_58 = W*in
   wire signed [14:0] m6_58;
   assign m6_58 =15'b0;

   // m6_59 = W*in
   wire signed [14:0] m6_59;
   assign m6_59 =15'b0;

   // m6_60 = W*in
   wire signed [14:0] m6_60;
   assign m6_60 =15'b0;

   // m6_61 = W*in
   wire signed [14:0] m6_61;
   assign m6_61 =15'b0;

   // m6_62 = W*in
   wire signed [14:0] m6_62;
   assign m6_62 =15'b0;

   // m6_63 = W*in
   wire signed [14:0] m6_63;
   assign m6_63 =15'b0;

   // m6_64 = W*in
   wire signed [14:0] m6_64;
   assign m6_64 =15'b0;

   // m6_65 = W*in
   wire signed [14:0] m6_65;
   assign m6_65 =15'b0;

   // m6_66 = W*in
   wire signed [14:0] m6_66;
   assign m6_66 =15'b0;

   // m6_67 = W*in
   wire signed [14:0] m6_67;
   assign m6_67 =15'b0;

   // m6_68 = W*in
   wire signed [14:0] m6_68;
   assign m6_68 ={ {3{in6[14]}} , in6[14:3] };

   // m6_69 = W*in
   wire signed [14:0] m6_69;
   assign m6_69 =15'b0;

   // m6_70 = W*in
   wire signed [14:0] m6_70;
   assign m6_70 ={ {3{in6[14]}} , in6[14:3] };

   // m6_71 = W*in
   wire signed [14:0] m6_71;
   assign m6_71 =15'b0;

   // m6_72 = W*in
   wire signed [14:0] m6_72;
   assign m6_72 =15'b0;

   // m6_73 = W*in
   wire signed [14:0] m6_73;
   assign m6_73 =15'b0;

   // m6_74 = W*in
   wire signed [14:0] m6_74;
   assign m6_74 =15'b0;

   // m6_75 = W*in
   wire signed [14:0] m6_75;
   assign m6_75 =15'b0;

   // m6_76 = W*in
   wire signed [14:0] m6_76;
   assign m6_76 =15'b0;

   // m6_77 = W*in
   wire signed [14:0] m6_77;
   assign m6_77 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_78 = W*in
   wire signed [14:0] m6_78;
   assign m6_78 ={ {3{in6[14]}} , in6[14:3] };

   // m6_79 = W*in
   wire signed [14:0] m6_79;
   assign m6_79 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_80 = W*in
   wire signed [14:0] m6_80;
   assign m6_80 =15'b0;

   // m6_81 = W*in
   wire signed [14:0] m6_81;
   assign m6_81 =15'b0;

   // m6_82 = W*in
   wire signed [14:0] m6_82;
   assign m6_82 =15'b0;

   // m6_83 = W*in
   wire signed [14:0] m6_83;
   assign m6_83 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_84 = W*in
   wire signed [14:0] m6_84;
   assign m6_84 =15'b0;

   // m6_85 = W*in
   wire signed [14:0] m6_85;
   assign m6_85 ={ {3{in6[14]}} , in6[14:3] };

   // m6_86 = W*in
   wire signed [14:0] m6_86;
   assign m6_86 =15'b0;

   // m6_87 = W*in
   wire signed [14:0] m6_87;
   assign m6_87 =15'b0;

   // m6_88 = W*in
   wire signed [14:0] m6_88;
   assign m6_88 =15'b0;

   // m6_89 = W*in
   wire signed [14:0] m6_89;
   assign m6_89 =15'b0;

   // m6_90 = W*in
   wire signed [14:0] m6_90;
   assign m6_90 ={ {3{in6[14]}} , in6[14:3] };

   // m6_91 = W*in
   wire signed [14:0] m6_91;
   assign m6_91 =15'b0;

   // m6_92 = W*in
   wire signed [14:0] m6_92;
   assign m6_92 =15'b0;

   // m6_93 = W*in
   wire signed [14:0] m6_93;
   assign m6_93 =15'b0;

   // m6_94 = W*in
   wire signed [14:0] m6_94;
   assign m6_94 =15'b0;

   // m6_95 = W*in
   wire signed [14:0] m6_95;
   assign m6_95 =15'b0;

   // m6_96 = W*in
   wire signed [14:0] m6_96;
   assign m6_96 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_97 = W*in
   wire signed [14:0] m6_97;
   assign m6_97 =15'b0;

   // m6_98 = W*in
   wire signed [14:0] m6_98;
   assign m6_98 =15'b0;

   // m6_99 = W*in
   wire signed [14:0] m6_99;
   assign m6_99 ={ {3{neg6[14]}} , neg6[14:3] };

   // m6_100 = W*in
   wire signed [14:0] m6_100;
   assign m6_100 ={ {3{neg6[14]}} , neg6[14:3] };

   // m7_1 = W*in
   wire signed [14:0] m7_1;
   assign m7_1 =15'b0;

   // m7_2 = W*in
   wire signed [14:0] m7_2;
   assign m7_2 =15'b0;

   // m7_3 = W*in
   wire signed [14:0] m7_3;
   assign m7_3 =15'b0;

   // m7_4 = W*in
   wire signed [14:0] m7_4;
   assign m7_4 =15'b0;

   // m7_5 = W*in
   wire signed [14:0] m7_5;
   assign m7_5 =15'b0;

   // m7_6 = W*in
   wire signed [14:0] m7_6;
   assign m7_6 =15'b0;

   // m7_7 = W*in
   wire signed [14:0] m7_7;
   assign m7_7 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_8 = W*in
   wire signed [14:0] m7_8;
   assign m7_8 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_9 = W*in
   wire signed [14:0] m7_9;
   assign m7_9 =15'b0;

   // m7_10 = W*in
   wire signed [14:0] m7_10;
   assign m7_10 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_11 = W*in
   wire signed [14:0] m7_11;
   assign m7_11 =15'b0;

   // m7_12 = W*in
   wire signed [14:0] m7_12;
   assign m7_12 =15'b0;

   // m7_13 = W*in
   wire signed [14:0] m7_13;
   assign m7_13 =15'b0;

   // m7_14 = W*in
   wire signed [14:0] m7_14;
   assign m7_14 =15'b0;

   // m7_15 = W*in
   wire signed [14:0] m7_15;
   assign m7_15 =15'b0;

   // m7_16 = W*in
   wire signed [14:0] m7_16;
   assign m7_16 ={ {3{in7[14]}} , in7[14:3] };

   // m7_17 = W*in
   wire signed [14:0] m7_17;
   assign m7_17 =15'b0;

   // m7_18 = W*in
   wire signed [14:0] m7_18;
   assign m7_18 =15'b0;

   // m7_19 = W*in
   wire signed [14:0] m7_19;
   assign m7_19 =15'b0;

   // m7_20 = W*in
   wire signed [14:0] m7_20;
   assign m7_20 =15'b0;

   // m7_21 = W*in
   wire signed [14:0] m7_21;
   assign m7_21 ={ {4{neg7[14]}} , neg7[14:4] };

   // m7_22 = W*in
   wire signed [14:0] m7_22;
   assign m7_22 =15'b0;

   // m7_23 = W*in
   wire signed [14:0] m7_23;
   assign m7_23 =15'b0;

   // m7_24 = W*in
   wire signed [14:0] m7_24;
   assign m7_24 =15'b0;

   // m7_25 = W*in
   wire signed [14:0] m7_25;
   assign m7_25 ={ {4{neg7[14]}} , neg7[14:4] };

   // m7_26 = W*in
   wire signed [14:0] m7_26;
   assign m7_26 =15'b0;

   // m7_27 = W*in
   wire signed [14:0] m7_27;
   assign m7_27 =15'b0;

   // m7_28 = W*in
   wire signed [14:0] m7_28;
   assign m7_28 =15'b0;

   // m7_29 = W*in
   wire signed [14:0] m7_29;
   assign m7_29 =15'b0;

   // m7_30 = W*in
   wire signed [14:0] m7_30;
   assign m7_30 =15'b0;

   // m7_31 = W*in
   wire signed [14:0] m7_31;
   assign m7_31 =15'b0;

   // m7_32 = W*in
   wire signed [14:0] m7_32;
   assign m7_32 =15'b0;

   // m7_33 = W*in
   wire signed [14:0] m7_33;
   assign m7_33 =15'b0;

   // m7_34 = W*in
   wire signed [14:0] m7_34;
   assign m7_34 =15'b0;

   // m7_35 = W*in
   wire signed [14:0] m7_35;
   assign m7_35 =15'b0;

   // m7_36 = W*in
   wire signed [14:0] m7_36;
   assign m7_36 =15'b0;

   // m7_37 = W*in
   wire signed [14:0] m7_37;
   assign m7_37 =15'b0;

   // m7_38 = W*in
   wire signed [14:0] m7_38;
   assign m7_38 =15'b0;

   // m7_39 = W*in
   wire signed [14:0] m7_39;
   assign m7_39 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_40 = W*in
   wire signed [14:0] m7_40;
   assign m7_40 =15'b0;

   // m7_41 = W*in
   wire signed [14:0] m7_41;
   assign m7_41 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_42 = W*in
   wire signed [14:0] m7_42;
   assign m7_42 =15'b0;

   // m7_43 = W*in
   wire signed [14:0] m7_43;
   assign m7_43 =15'b0;

   // m7_44 = W*in
   wire signed [14:0] m7_44;
   assign m7_44 =15'b0;

   // m7_45 = W*in
   wire signed [14:0] m7_45;
   assign m7_45 =15'b0;

   // m7_46 = W*in
   wire signed [14:0] m7_46;
   assign m7_46 =15'b0;

   // m7_47 = W*in
   wire signed [14:0] m7_47;
   assign m7_47 =15'b0;

   // m7_48 = W*in
   wire signed [14:0] m7_48;
   assign m7_48 ={ {4{in7[14]}} , in7[14:4] };

   // m7_49 = W*in
   wire signed [14:0] m7_49;
   assign m7_49 =15'b0;

   // m7_50 = W*in
   wire signed [14:0] m7_50;
   assign m7_50 =15'b0;

   // m7_51 = W*in
   wire signed [14:0] m7_51;
   assign m7_51 =15'b0;

   // m7_52 = W*in
   wire signed [14:0] m7_52;
   assign m7_52 =15'b0;

   // m7_53 = W*in
   wire signed [14:0] m7_53;
   assign m7_53 =15'b0;

   // m7_54 = W*in
   wire signed [14:0] m7_54;
   assign m7_54 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_55 = W*in
   wire signed [14:0] m7_55;
   assign m7_55 =15'b0;

   // m7_56 = W*in
   wire signed [14:0] m7_56;
   assign m7_56 ={ {3{in7[14]}} , in7[14:3] };

   // m7_57 = W*in
   wire signed [14:0] m7_57;
   assign m7_57 ={ {3{in7[14]}} , in7[14:3] };

   // m7_58 = W*in
   wire signed [14:0] m7_58;
   assign m7_58 ={ {3{in7[14]}} , in7[14:3] };

   // m7_59 = W*in
   wire signed [14:0] m7_59;
   assign m7_59 =15'b0;

   // m7_60 = W*in
   wire signed [14:0] m7_60;
   assign m7_60 =15'b0;

   // m7_61 = W*in
   wire signed [14:0] m7_61;
   assign m7_61 ={ {4{neg7[14]}} , neg7[14:4] };

   // m7_62 = W*in
   wire signed [14:0] m7_62;
   assign m7_62 ={ {3{in7[14]}} , in7[14:3] };

   // m7_63 = W*in
   wire signed [14:0] m7_63;
   assign m7_63 =15'b0;

   // m7_64 = W*in
   wire signed [14:0] m7_64;
   assign m7_64 ={ {3{in7[14]}} , in7[14:3] };

   // m7_65 = W*in
   wire signed [14:0] m7_65;
   assign m7_65 =15'b0;

   // m7_66 = W*in
   wire signed [14:0] m7_66;
   assign m7_66 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_67 = W*in
   wire signed [14:0] m7_67;
   assign m7_67 =15'b0;

   // m7_68 = W*in
   wire signed [14:0] m7_68;
   assign m7_68 =15'b0;

   // m7_69 = W*in
   wire signed [14:0] m7_69;
   assign m7_69 ={ {4{neg7[14]}} , neg7[14:4] };

   // m7_70 = W*in
   wire signed [14:0] m7_70;
   assign m7_70 =15'b0;

   // m7_71 = W*in
   wire signed [14:0] m7_71;
   assign m7_71 =15'b0;

   // m7_72 = W*in
   wire signed [14:0] m7_72;
   assign m7_72 =15'b0;

   // m7_73 = W*in
   wire signed [14:0] m7_73;
   assign m7_73 =15'b0;

   // m7_74 = W*in
   wire signed [14:0] m7_74;
   assign m7_74 =15'b0;

   // m7_75 = W*in
   wire signed [14:0] m7_75;
   assign m7_75 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_76 = W*in
   wire signed [14:0] m7_76;
   assign m7_76 =15'b0;

   // m7_77 = W*in
   wire signed [14:0] m7_77;
   assign m7_77 =15'b0;

   // m7_78 = W*in
   wire signed [14:0] m7_78;
   assign m7_78 =15'b0;

   // m7_79 = W*in
   wire signed [14:0] m7_79;
   assign m7_79 =15'b0;

   // m7_80 = W*in
   wire signed [14:0] m7_80;
   assign m7_80 =15'b0;

   // m7_81 = W*in
   wire signed [14:0] m7_81;
   assign m7_81 =15'b0;

   // m7_82 = W*in
   wire signed [14:0] m7_82;
   assign m7_82 =15'b0;

   // m7_83 = W*in
   wire signed [14:0] m7_83;
   assign m7_83 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_84 = W*in
   wire signed [14:0] m7_84;
   assign m7_84 =15'b0;

   // m7_85 = W*in
   wire signed [14:0] m7_85;
   assign m7_85 =15'b0;

   // m7_86 = W*in
   wire signed [14:0] m7_86;
   assign m7_86 =15'b0;

   // m7_87 = W*in
   wire signed [14:0] m7_87;
   assign m7_87 =15'b0;

   // m7_88 = W*in
   wire signed [14:0] m7_88;
   assign m7_88 =15'b0;

   // m7_89 = W*in
   wire signed [14:0] m7_89;
   assign m7_89 =15'b0;

   // m7_90 = W*in
   wire signed [14:0] m7_90;
   assign m7_90 =15'b0;

   // m7_91 = W*in
   wire signed [14:0] m7_91;
   assign m7_91 =15'b0;

   // m7_92 = W*in
   wire signed [14:0] m7_92;
   assign m7_92 ={ {3{in7[14]}} , in7[14:3] };

   // m7_93 = W*in
   wire signed [14:0] m7_93;
   assign m7_93 =15'b0;

   // m7_94 = W*in
   wire signed [14:0] m7_94;
   assign m7_94 ={ {3{neg7[14]}} , neg7[14:3] };

   // m7_95 = W*in
   wire signed [14:0] m7_95;
   assign m7_95 =15'b0;

   // m7_96 = W*in
   wire signed [14:0] m7_96;
   assign m7_96 =15'b0;

   // m7_97 = W*in
   wire signed [14:0] m7_97;
   assign m7_97 =15'b0;

   // m7_98 = W*in
   wire signed [14:0] m7_98;
   assign m7_98 =15'b0;

   // m7_99 = W*in
   wire signed [14:0] m7_99;
   assign m7_99 =15'b0;

   // m7_100 = W*in
   wire signed [14:0] m7_100;
   assign m7_100 =15'b0;

   // m8_1 = W*in
   wire signed [14:0] m8_1;
   assign m8_1 =15'b0;

   // m8_2 = W*in
   wire signed [14:0] m8_2;
   assign m8_2 ={ {3{neg8[14]}} , neg8[14:3] };

   // m8_3 = W*in
   wire signed [14:0] m8_3;
   assign m8_3 =15'b0;

   // m8_4 = W*in
   wire signed [14:0] m8_4;
   assign m8_4 =15'b0;

   // m8_5 = W*in
   wire signed [14:0] m8_5;
   assign m8_5 =15'b0;

   // m8_6 = W*in
   wire signed [14:0] m8_6;
   assign m8_6 =15'b0;

   // m8_7 = W*in
   wire signed [14:0] m8_7;
   assign m8_7 =15'b0;

   // m8_8 = W*in
   wire signed [14:0] m8_8;
   assign m8_8 =15'b0;

   // m8_9 = W*in
   wire signed [14:0] m8_9;
   assign m8_9 =15'b0;

   // m8_10 = W*in
   wire signed [14:0] m8_10;
   assign m8_10 =15'b0;

   // m8_11 = W*in
   wire signed [14:0] m8_11;
   assign m8_11 =15'b0;

   // m8_12 = W*in
   wire signed [14:0] m8_12;
   assign m8_12 =15'b0;

   // m8_13 = W*in
   wire signed [14:0] m8_13;
   assign m8_13 =15'b0;

   // m8_14 = W*in
   wire signed [14:0] m8_14;
   assign m8_14 =15'b0;

   // m8_15 = W*in
   wire signed [14:0] m8_15;
   assign m8_15 =15'b0;

   // m8_16 = W*in
   wire signed [14:0] m8_16;
   assign m8_16 =15'b0;

   // m8_17 = W*in
   wire signed [14:0] m8_17;
   assign m8_17 ={ {3{in8[14]}} , in8[14:3] };

   // m8_18 = W*in
   wire signed [14:0] m8_18;
   assign m8_18 =15'b0;

   // m8_19 = W*in
   wire signed [14:0] m8_19;
   assign m8_19 =15'b0;

   // m8_20 = W*in
   wire signed [14:0] m8_20;
   assign m8_20 =15'b0;

   // m8_21 = W*in
   wire signed [14:0] m8_21;
   assign m8_21 =15'b0;

   // m8_22 = W*in
   wire signed [14:0] m8_22;
   assign m8_22 =15'b0;

   // m8_23 = W*in
   wire signed [14:0] m8_23;
   assign m8_23 =15'b0;

   // m8_24 = W*in
   wire signed [14:0] m8_24;
   assign m8_24 =15'b0;

   // m8_25 = W*in
   wire signed [14:0] m8_25;
   assign m8_25 =15'b0;

   // m8_26 = W*in
   wire signed [14:0] m8_26;
   assign m8_26 =15'b0;

   // m8_27 = W*in
   wire signed [14:0] m8_27;
   assign m8_27 =15'b0;

   // m8_28 = W*in
   wire signed [14:0] m8_28;
   assign m8_28 =15'b0;

   // m8_29 = W*in
   wire signed [14:0] m8_29;
   assign m8_29 =15'b0;

   // m8_30 = W*in
   wire signed [14:0] m8_30;
   assign m8_30 ={ {4{in8[14]}} , in8[14:4] };

   // m8_31 = W*in
   wire signed [14:0] m8_31;
   assign m8_31 =15'b0;

   // m8_32 = W*in
   wire signed [14:0] m8_32;
   assign m8_32 =15'b0;

   // m8_33 = W*in
   wire signed [14:0] m8_33;
   assign m8_33 =15'b0;

   // m8_34 = W*in
   wire signed [14:0] m8_34;
   assign m8_34 =15'b0;

   // m8_35 = W*in
   wire signed [14:0] m8_35;
   assign m8_35 ={ {3{neg8[14]}} , neg8[14:3] };

   // m8_36 = W*in
   wire signed [14:0] m8_36;
   assign m8_36 =15'b0;

   // m8_37 = W*in
   wire signed [14:0] m8_37;
   assign m8_37 =15'b0;

   // m8_38 = W*in
   wire signed [14:0] m8_38;
   assign m8_38 ={ {3{neg8[14]}} , neg8[14:3] };

   // m8_39 = W*in
   wire signed [14:0] m8_39;
   assign m8_39 =15'b0;

   // m8_40 = W*in
   wire signed [14:0] m8_40;
   assign m8_40 =15'b0;

   // m8_41 = W*in
   wire signed [14:0] m8_41;
   assign m8_41 =15'b0;

   // m8_42 = W*in
   wire signed [14:0] m8_42;
   assign m8_42 =15'b0;

   // m8_43 = W*in
   wire signed [14:0] m8_43;
   assign m8_43 =15'b0;

   // m8_44 = W*in
   wire signed [14:0] m8_44;
   assign m8_44 =15'b0;

   // m8_45 = W*in
   wire signed [14:0] m8_45;
   assign m8_45 =15'b0;

   // m8_46 = W*in
   wire signed [14:0] m8_46;
   assign m8_46 =15'b0;

   // m8_47 = W*in
   wire signed [14:0] m8_47;
   assign m8_47 =15'b0;

   // m8_48 = W*in
   wire signed [14:0] m8_48;
   assign m8_48 =15'b0;

   // m8_49 = W*in
   wire signed [14:0] m8_49;
   assign m8_49 =15'b0;

   // m8_50 = W*in
   wire signed [14:0] m8_50;
   assign m8_50 =15'b0;

   // m8_51 = W*in
   wire signed [14:0] m8_51;
   assign m8_51 =15'b0;

   // m8_52 = W*in
   wire signed [14:0] m8_52;
   assign m8_52 =15'b0;

   // m8_53 = W*in
   wire signed [14:0] m8_53;
   assign m8_53 ={ {3{in8[14]}} , in8[14:3] };

   // m8_54 = W*in
   wire signed [14:0] m8_54;
   assign m8_54 =15'b0;

   // m8_55 = W*in
   wire signed [14:0] m8_55;
   assign m8_55 =15'b0;

   // m8_56 = W*in
   wire signed [14:0] m8_56;
   assign m8_56 ={ {4{in8[14]}} , in8[14:4] };

   // m8_57 = W*in
   wire signed [14:0] m8_57;
   assign m8_57 =15'b0;

   // m8_58 = W*in
   wire signed [14:0] m8_58;
   assign m8_58 =15'b0;

   // m8_59 = W*in
   wire signed [14:0] m8_59;
   assign m8_59 =15'b0;

   // m8_60 = W*in
   wire signed [14:0] m8_60;
   assign m8_60 ={ {3{neg8[14]}} , neg8[14:3] };

   // m8_61 = W*in
   wire signed [14:0] m8_61;
   assign m8_61 =15'b0;

   // m8_62 = W*in
   wire signed [14:0] m8_62;
   assign m8_62 =15'b0;

   // m8_63 = W*in
   wire signed [14:0] m8_63;
   assign m8_63 =15'b0;

   // m8_64 = W*in
   wire signed [14:0] m8_64;
   assign m8_64 ={ {3{in8[14]}} , in8[14:3] };

   // m8_65 = W*in
   wire signed [14:0] m8_65;
   assign m8_65 ={ {4{in8[14]}} , in8[14:4] };

   // m8_66 = W*in
   wire signed [14:0] m8_66;
   assign m8_66 =15'b0;

   // m8_67 = W*in
   wire signed [14:0] m8_67;
   assign m8_67 =15'b0;

   // m8_68 = W*in
   wire signed [14:0] m8_68;
   assign m8_68 =15'b0;

   // m8_69 = W*in
   wire signed [14:0] m8_69;
   assign m8_69 =15'b0;

   // m8_70 = W*in
   wire signed [14:0] m8_70;
   assign m8_70 =15'b0;

   // m8_71 = W*in
   wire signed [14:0] m8_71;
   assign m8_71 =15'b0;

   // m8_72 = W*in
   wire signed [14:0] m8_72;
   assign m8_72 =15'b0;

   // m8_73 = W*in
   wire signed [14:0] m8_73;
   assign m8_73 =15'b0;

   // m8_74 = W*in
   wire signed [14:0] m8_74;
   assign m8_74 =15'b0;

   // m8_75 = W*in
   wire signed [14:0] m8_75;
   assign m8_75 =15'b0;

   // m8_76 = W*in
   wire signed [14:0] m8_76;
   assign m8_76 =15'b0;

   // m8_77 = W*in
   wire signed [14:0] m8_77;
   assign m8_77 =15'b0;

   // m8_78 = W*in
   wire signed [14:0] m8_78;
   assign m8_78 =15'b0;

   // m8_79 = W*in
   wire signed [14:0] m8_79;
   assign m8_79 =15'b0;

   // m8_80 = W*in
   wire signed [14:0] m8_80;
   assign m8_80 =15'b0;

   // m8_81 = W*in
   wire signed [14:0] m8_81;
   assign m8_81 =15'b0;

   // m8_82 = W*in
   wire signed [14:0] m8_82;
   assign m8_82 =15'b0;

   // m8_83 = W*in
   wire signed [14:0] m8_83;
   assign m8_83 =15'b0;

   // m8_84 = W*in
   wire signed [14:0] m8_84;
   assign m8_84 =15'b0;

   // m8_85 = W*in
   wire signed [14:0] m8_85;
   assign m8_85 ={ {3{in8[14]}} , in8[14:3] };

   // m8_86 = W*in
   wire signed [14:0] m8_86;
   assign m8_86 =15'b0;

   // m8_87 = W*in
   wire signed [14:0] m8_87;
   assign m8_87 =15'b0;

   // m8_88 = W*in
   wire signed [14:0] m8_88;
   assign m8_88 =15'b0;

   // m8_89 = W*in
   wire signed [14:0] m8_89;
   assign m8_89 =15'b0;

   // m8_90 = W*in
   wire signed [14:0] m8_90;
   assign m8_90 =15'b0;

   // m8_91 = W*in
   wire signed [14:0] m8_91;
   assign m8_91 ={ {3{neg8[14]}} , neg8[14:3] };

   // m8_92 = W*in
   wire signed [14:0] m8_92;
   assign m8_92 =15'b0;

   // m8_93 = W*in
   wire signed [14:0] m8_93;
   assign m8_93 =15'b0;

   // m8_94 = W*in
   wire signed [14:0] m8_94;
   assign m8_94 =15'b0;

   // m8_95 = W*in
   wire signed [14:0] m8_95;
   assign m8_95 =15'b0;

   // m8_96 = W*in
   wire signed [14:0] m8_96;
   assign m8_96 =15'b0;

   // m8_97 = W*in
   wire signed [14:0] m8_97;
   assign m8_97 =15'b0;

   // m8_98 = W*in
   wire signed [14:0] m8_98;
   assign m8_98 =15'b0;

   // m8_99 = W*in
   wire signed [14:0] m8_99;
   assign m8_99 =15'b0;

   // m8_100 = W*in
   wire signed [14:0] m8_100;
   assign m8_100 =15'b0;

   // m9_1 = W*in
   wire signed [14:0] m9_1;
   assign m9_1 =15'b0;

   // m9_2 = W*in
   wire signed [14:0] m9_2;
   assign m9_2 =15'b0;

   // m9_3 = W*in
   wire signed [14:0] m9_3;
   assign m9_3 =15'b0;

   // m9_4 = W*in
   wire signed [14:0] m9_4;
   assign m9_4 =15'b0;

   // m9_5 = W*in
   wire signed [14:0] m9_5;
   assign m9_5 =15'b0;

   // m9_6 = W*in
   wire signed [14:0] m9_6;
   assign m9_6 =15'b0;

   // m9_7 = W*in
   wire signed [14:0] m9_7;
   assign m9_7 =15'b0;

   // m9_8 = W*in
   wire signed [14:0] m9_8;
   assign m9_8 =15'b0;

   // m9_9 = W*in
   wire signed [14:0] m9_9;
   assign m9_9 =15'b0;

   // m9_10 = W*in
   wire signed [14:0] m9_10;
   assign m9_10 =15'b0;

   // m9_11 = W*in
   wire signed [14:0] m9_11;
   assign m9_11 ={ {4{neg9[14]}} , neg9[14:4] };

   // m9_12 = W*in
   wire signed [14:0] m9_12;
   assign m9_12 =15'b0;

   // m9_13 = W*in
   wire signed [14:0] m9_13;
   assign m9_13 =15'b0;

   // m9_14 = W*in
   wire signed [14:0] m9_14;
   assign m9_14 =15'b0;

   // m9_15 = W*in
   wire signed [14:0] m9_15;
   assign m9_15 =15'b0;

   // m9_16 = W*in
   wire signed [14:0] m9_16;
   assign m9_16 =15'b0;

   // m9_17 = W*in
   wire signed [14:0] m9_17;
   assign m9_17 =15'b0;

   // m9_18 = W*in
   wire signed [14:0] m9_18;
   assign m9_18 =15'b0;

   // m9_19 = W*in
   wire signed [14:0] m9_19;
   assign m9_19 =15'b0;

   // m9_20 = W*in
   wire signed [14:0] m9_20;
   assign m9_20 =15'b0;

   // m9_21 = W*in
   wire signed [14:0] m9_21;
   assign m9_21 =15'b0;

   // m9_22 = W*in
   wire signed [14:0] m9_22;
   assign m9_22 =15'b0;

   // m9_23 = W*in
   wire signed [14:0] m9_23;
   assign m9_23 =15'b0;

   // m9_24 = W*in
   wire signed [14:0] m9_24;
   assign m9_24 ={ {3{neg9[14]}} , neg9[14:3] };

   // m9_25 = W*in
   wire signed [14:0] m9_25;
   assign m9_25 =15'b0;

   // m9_26 = W*in
   wire signed [14:0] m9_26;
   assign m9_26 =15'b0;

   // m9_27 = W*in
   wire signed [14:0] m9_27;
   assign m9_27 =15'b0;

   // m9_28 = W*in
   wire signed [14:0] m9_28;
   assign m9_28 =15'b0;

   // m9_29 = W*in
   wire signed [14:0] m9_29;
   assign m9_29 =15'b0;

   // m9_30 = W*in
   wire signed [14:0] m9_30;
   assign m9_30 =15'b0;

   // m9_31 = W*in
   wire signed [14:0] m9_31;
   assign m9_31 =15'b0;

   // m9_32 = W*in
   wire signed [14:0] m9_32;
   assign m9_32 =15'b0;

   // m9_33 = W*in
   wire signed [14:0] m9_33;
   assign m9_33 ={ {3{neg9[14]}} , neg9[14:3] };

   // m9_34 = W*in
   wire signed [14:0] m9_34;
   assign m9_34 =15'b0;

   // m9_35 = W*in
   wire signed [14:0] m9_35;
   assign m9_35 =15'b0;

   // m9_36 = W*in
   wire signed [14:0] m9_36;
   assign m9_36 =15'b0;

   // m9_37 = W*in
   wire signed [14:0] m9_37;
   assign m9_37 =15'b0;

   // m9_38 = W*in
   wire signed [14:0] m9_38;
   assign m9_38 =15'b0;

   // m9_39 = W*in
   wire signed [14:0] m9_39;
   assign m9_39 ={ {3{in9[14]}} , in9[14:3] };

   // m9_40 = W*in
   wire signed [14:0] m9_40;
   assign m9_40 ={ {3{in9[14]}} , in9[14:3] };

   // m9_41 = W*in
   wire signed [14:0] m9_41;
   assign m9_41 =15'b0;

   // m9_42 = W*in
   wire signed [14:0] m9_42;
   assign m9_42 ={ {3{in9[14]}} , in9[14:3] };

   // m9_43 = W*in
   wire signed [14:0] m9_43;
   assign m9_43 =15'b0;

   // m9_44 = W*in
   wire signed [14:0] m9_44;
   assign m9_44 ={ {4{neg9[14]}} , neg9[14:4] };

   // m9_45 = W*in
   wire signed [14:0] m9_45;
   assign m9_45 =15'b0;

   // m9_46 = W*in
   wire signed [14:0] m9_46;
   assign m9_46 ={ {4{neg9[14]}} , neg9[14:4] };

   // m9_47 = W*in
   wire signed [14:0] m9_47;
   assign m9_47 =15'b0;

   // m9_48 = W*in
   wire signed [14:0] m9_48;
   assign m9_48 ={ {3{in9[14]}} , in9[14:3] };

   // m9_49 = W*in
   wire signed [14:0] m9_49;
   assign m9_49 =15'b0;

   // m9_50 = W*in
   wire signed [14:0] m9_50;
   assign m9_50 =15'b0;

   // m9_51 = W*in
   wire signed [14:0] m9_51;
   assign m9_51 =15'b0;

   // m9_52 = W*in
   wire signed [14:0] m9_52;
   assign m9_52 =15'b0;

   // m9_53 = W*in
   wire signed [14:0] m9_53;
   assign m9_53 =15'b0;

   // m9_54 = W*in
   wire signed [14:0] m9_54;
   assign m9_54 =15'b0;

   // m9_55 = W*in
   wire signed [14:0] m9_55;
   assign m9_55 =15'b0;

   // m9_56 = W*in
   wire signed [14:0] m9_56;
   assign m9_56 ={ {4{in9[14]}} , in9[14:4] };

   // m9_57 = W*in
   wire signed [14:0] m9_57;
   assign m9_57 =15'b0;

   // m9_58 = W*in
   wire signed [14:0] m9_58;
   assign m9_58 =15'b0;

   // m9_59 = W*in
   wire signed [14:0] m9_59;
   assign m9_59 =15'b0;

   // m9_60 = W*in
   wire signed [14:0] m9_60;
   assign m9_60 =15'b0;

   // m9_61 = W*in
   wire signed [14:0] m9_61;
   assign m9_61 =15'b0;

   // m9_62 = W*in
   wire signed [14:0] m9_62;
   assign m9_62 =15'b0;

   // m9_63 = W*in
   wire signed [14:0] m9_63;
   assign m9_63 =15'b0;

   // m9_64 = W*in
   wire signed [14:0] m9_64;
   assign m9_64 =15'b0;

   // m9_65 = W*in
   wire signed [14:0] m9_65;
   assign m9_65 =15'b0;

   // m9_66 = W*in
   wire signed [14:0] m9_66;
   assign m9_66 =15'b0;

   // m9_67 = W*in
   wire signed [14:0] m9_67;
   assign m9_67 =15'b0;

   // m9_68 = W*in
   wire signed [14:0] m9_68;
   assign m9_68 =15'b0;

   // m9_69 = W*in
   wire signed [14:0] m9_69;
   assign m9_69 =15'b0;

   // m9_70 = W*in
   wire signed [14:0] m9_70;
   assign m9_70 =15'b0;

   // m9_71 = W*in
   wire signed [14:0] m9_71;
   assign m9_71 =15'b0;

   // m9_72 = W*in
   wire signed [14:0] m9_72;
   assign m9_72 =15'b0;

   // m9_73 = W*in
   wire signed [14:0] m9_73;
   assign m9_73 =15'b0;

   // m9_74 = W*in
   wire signed [14:0] m9_74;
   assign m9_74 =15'b0;

   // m9_75 = W*in
   wire signed [14:0] m9_75;
   assign m9_75 =15'b0;

   // m9_76 = W*in
   wire signed [14:0] m9_76;
   assign m9_76 =15'b0;

   // m9_77 = W*in
   wire signed [14:0] m9_77;
   assign m9_77 =15'b0;

   // m9_78 = W*in
   wire signed [14:0] m9_78;
   assign m9_78 =15'b0;

   // m9_79 = W*in
   wire signed [14:0] m9_79;
   assign m9_79 =15'b0;

   // m9_80 = W*in
   wire signed [14:0] m9_80;
   assign m9_80 =15'b0;

   // m9_81 = W*in
   wire signed [14:0] m9_81;
   assign m9_81 =15'b0;

   // m9_82 = W*in
   wire signed [14:0] m9_82;
   assign m9_82 =15'b0;

   // m9_83 = W*in
   wire signed [14:0] m9_83;
   assign m9_83 =15'b0;

   // m9_84 = W*in
   wire signed [14:0] m9_84;
   assign m9_84 =15'b0;

   // m9_85 = W*in
   wire signed [14:0] m9_85;
   assign m9_85 =15'b0;

   // m9_86 = W*in
   wire signed [14:0] m9_86;
   assign m9_86 =15'b0;

   // m9_87 = W*in
   wire signed [14:0] m9_87;
   assign m9_87 =15'b0;

   // m9_88 = W*in
   wire signed [14:0] m9_88;
   assign m9_88 =15'b0;

   // m9_89 = W*in
   wire signed [14:0] m9_89;
   assign m9_89 =15'b0;

   // m9_90 = W*in
   wire signed [14:0] m9_90;
   assign m9_90 ={ {4{in9[14]}} , in9[14:4] };

   // m9_91 = W*in
   wire signed [14:0] m9_91;
   assign m9_91 =15'b0;

   // m9_92 = W*in
   wire signed [14:0] m9_92;
   assign m9_92 =15'b0;

   // m9_93 = W*in
   wire signed [14:0] m9_93;
   assign m9_93 =15'b0;

   // m9_94 = W*in
   wire signed [14:0] m9_94;
   assign m9_94 =15'b0;

   // m9_95 = W*in
   wire signed [14:0] m9_95;
   assign m9_95 =15'b0;

   // m9_96 = W*in
   wire signed [14:0] m9_96;
   assign m9_96 =15'b0;

   // m9_97 = W*in
   wire signed [14:0] m9_97;
   assign m9_97 =15'b0;

   // m9_98 = W*in
   wire signed [14:0] m9_98;
   assign m9_98 =15'b0;

   // m9_99 = W*in
   wire signed [14:0] m9_99;
   assign m9_99 =15'b0;

   // m9_100 = W*in
   wire signed [14:0] m9_100;
   assign m9_100 ={ {4{neg9[14]}} , neg9[14:4] };

   // m10_1 = W*in
   wire signed [14:0] m10_1;
   assign m10_1 =15'b0;

   // m10_2 = W*in
   wire signed [14:0] m10_2;
   assign m10_2 =15'b0;

   // m10_3 = W*in
   wire signed [14:0] m10_3;
   assign m10_3 =15'b0;

   // m10_4 = W*in
   wire signed [14:0] m10_4;
   assign m10_4 =15'b0;

   // m10_5 = W*in
   wire signed [14:0] m10_5;
   assign m10_5 =15'b0;

   // m10_6 = W*in
   wire signed [14:0] m10_6;
   assign m10_6 =15'b0;

   // m10_7 = W*in
   wire signed [14:0] m10_7;
   assign m10_7 ={ {3{neg10[14]}} , neg10[14:3] };

   // m10_8 = W*in
   wire signed [14:0] m10_8;
   assign m10_8 ={ {3{neg10[14]}} , neg10[14:3] };

   // m10_9 = W*in
   wire signed [14:0] m10_9;
   assign m10_9 =15'b0;

   // m10_10 = W*in
   wire signed [14:0] m10_10;
   assign m10_10 =15'b0;

   // m10_11 = W*in
   wire signed [14:0] m10_11;
   assign m10_11 =15'b0;

   // m10_12 = W*in
   wire signed [14:0] m10_12;
   assign m10_12 =15'b0;

   // m10_13 = W*in
   wire signed [14:0] m10_13;
   assign m10_13 =15'b0;

   // m10_14 = W*in
   wire signed [14:0] m10_14;
   assign m10_14 ={ {3{neg10[14]}} , neg10[14:3] };

   // m10_15 = W*in
   wire signed [14:0] m10_15;
   assign m10_15 =15'b0;

   // m10_16 = W*in
   wire signed [14:0] m10_16;
   assign m10_16 =15'b0;

   // m10_17 = W*in
   wire signed [14:0] m10_17;
   assign m10_17 =15'b0;

   // m10_18 = W*in
   wire signed [14:0] m10_18;
   assign m10_18 =15'b0;

   // m10_19 = W*in
   wire signed [14:0] m10_19;
   assign m10_19 =15'b0;

   // m10_20 = W*in
   wire signed [14:0] m10_20;
   assign m10_20 =15'b0;

   // m10_21 = W*in
   wire signed [14:0] m10_21;
   assign m10_21 ={ {4{in10[14]}} , in10[14:4] };

   // m10_22 = W*in
   wire signed [14:0] m10_22;
   assign m10_22 =15'b0;

   // m10_23 = W*in
   wire signed [14:0] m10_23;
   assign m10_23 =15'b0;

   // m10_24 = W*in
   wire signed [14:0] m10_24;
   assign m10_24 =15'b0;

   // m10_25 = W*in
   wire signed [14:0] m10_25;
   assign m10_25 ={ {4{in10[14]}} , in10[14:4] };

   // m10_26 = W*in
   wire signed [14:0] m10_26;
   assign m10_26 =15'b0;

   // m10_27 = W*in
   wire signed [14:0] m10_27;
   assign m10_27 =15'b0;

   // m10_28 = W*in
   wire signed [14:0] m10_28;
   assign m10_28 =15'b0;

   // m10_29 = W*in
   wire signed [14:0] m10_29;
   assign m10_29 ={ {4{neg10[14]}} , neg10[14:4] };

   // m10_30 = W*in
   wire signed [14:0] m10_30;
   assign m10_30 =15'b0;

   // m10_31 = W*in
   wire signed [14:0] m10_31;
   assign m10_31 =15'b0;

   // m10_32 = W*in
   wire signed [14:0] m10_32;
   assign m10_32 =15'b0;

   // m10_33 = W*in
   wire signed [14:0] m10_33;
   assign m10_33 =15'b0;

   // m10_34 = W*in
   wire signed [14:0] m10_34;
   assign m10_34 =15'b0;

   // m10_35 = W*in
   wire signed [14:0] m10_35;
   assign m10_35 =15'b0;

   // m10_36 = W*in
   wire signed [14:0] m10_36;
   assign m10_36 =15'b0;

   // m10_37 = W*in
   wire signed [14:0] m10_37;
   assign m10_37 =15'b0;

   // m10_38 = W*in
   wire signed [14:0] m10_38;
   assign m10_38 =15'b0;

   // m10_39 = W*in
   wire signed [14:0] m10_39;
   assign m10_39 =15'b0;

   // m10_40 = W*in
   wire signed [14:0] m10_40;
   assign m10_40 =15'b0;

   // m10_41 = W*in
   wire signed [14:0] m10_41;
   assign m10_41 ={ {4{neg10[14]}} , neg10[14:4] };

   // m10_42 = W*in
   wire signed [14:0] m10_42;
   assign m10_42 =15'b0;

   // m10_43 = W*in
   wire signed [14:0] m10_43;
   assign m10_43 =15'b0;

   // m10_44 = W*in
   wire signed [14:0] m10_44;
   assign m10_44 =15'b0;

   // m10_45 = W*in
   wire signed [14:0] m10_45;
   assign m10_45 =15'b0;

   // m10_46 = W*in
   wire signed [14:0] m10_46;
   assign m10_46 =15'b0;

   // m10_47 = W*in
   wire signed [14:0] m10_47;
   assign m10_47 =15'b0;

   // m10_48 = W*in
   wire signed [14:0] m10_48;
   assign m10_48 =15'b0;

   // m10_49 = W*in
   wire signed [14:0] m10_49;
   assign m10_49 =15'b0;

   // m10_50 = W*in
   wire signed [14:0] m10_50;
   assign m10_50 =15'b0;

   // m10_51 = W*in
   wire signed [14:0] m10_51;
   assign m10_51 =15'b0;

   // m10_52 = W*in
   wire signed [14:0] m10_52;
   assign m10_52 =15'b0;

   // m10_53 = W*in
   wire signed [14:0] m10_53;
   assign m10_53 =15'b0;

   // m10_54 = W*in
   wire signed [14:0] m10_54;
   assign m10_54 ={ {3{neg10[14]}} , neg10[14:3] };

   // m10_55 = W*in
   wire signed [14:0] m10_55;
   assign m10_55 =15'b0;

   // m10_56 = W*in
   wire signed [14:0] m10_56;
   assign m10_56 =15'b0;

   // m10_57 = W*in
   wire signed [14:0] m10_57;
   assign m10_57 =15'b0;

   // m10_58 = W*in
   wire signed [14:0] m10_58;
   assign m10_58 =15'b0;

   // m10_59 = W*in
   wire signed [14:0] m10_59;
   assign m10_59 ={ {4{in10[14]}} , in10[14:4] };

   // m10_60 = W*in
   wire signed [14:0] m10_60;
   assign m10_60 =15'b0;

   // m10_61 = W*in
   wire signed [14:0] m10_61;
   assign m10_61 ={ {4{in10[14]}} , in10[14:4] };

   // m10_62 = W*in
   wire signed [14:0] m10_62;
   assign m10_62 =15'b0;

   // m10_63 = W*in
   wire signed [14:0] m10_63;
   assign m10_63 =15'b0;

   // m10_64 = W*in
   wire signed [14:0] m10_64;
   assign m10_64 ={ {4{in10[14]}} , in10[14:4] };

   // m10_65 = W*in
   wire signed [14:0] m10_65;
   assign m10_65 ={ {4{in10[14]}} , in10[14:4] };

   // m10_66 = W*in
   wire signed [14:0] m10_66;
   assign m10_66 ={ {4{neg10[14]}} , neg10[14:4] };

   // m10_67 = W*in
   wire signed [14:0] m10_67;
   assign m10_67 ={ {4{in10[14]}} , in10[14:4] };

   // m10_68 = W*in
   wire signed [14:0] m10_68;
   assign m10_68 =15'b0;

   // m10_69 = W*in
   wire signed [14:0] m10_69;
   assign m10_69 ={ {4{in10[14]}} , in10[14:4] };

   // m10_70 = W*in
   wire signed [14:0] m10_70;
   assign m10_70 =15'b0;

   // m10_71 = W*in
   wire signed [14:0] m10_71;
   assign m10_71 =15'b0;

   // m10_72 = W*in
   wire signed [14:0] m10_72;
   assign m10_72 =15'b0;

   // m10_73 = W*in
   wire signed [14:0] m10_73;
   assign m10_73 =15'b0;

   // m10_74 = W*in
   wire signed [14:0] m10_74;
   assign m10_74 =15'b0;

   // m10_75 = W*in
   wire signed [14:0] m10_75;
   assign m10_75 ={ {4{in10[14]}} , in10[14:4] };

   // m10_76 = W*in
   wire signed [14:0] m10_76;
   assign m10_76 =15'b0;

   // m10_77 = W*in
   wire signed [14:0] m10_77;
   assign m10_77 =15'b0;

   // m10_78 = W*in
   wire signed [14:0] m10_78;
   assign m10_78 =15'b0;

   // m10_79 = W*in
   wire signed [14:0] m10_79;
   assign m10_79 =15'b0;

   // m10_80 = W*in
   wire signed [14:0] m10_80;
   assign m10_80 =15'b0;

   // m10_81 = W*in
   wire signed [14:0] m10_81;
   assign m10_81 =15'b0;

   // m10_82 = W*in
   wire signed [14:0] m10_82;
   assign m10_82 =15'b0;

   // m10_83 = W*in
   wire signed [14:0] m10_83;
   assign m10_83 =15'b0;

   // m10_84 = W*in
   wire signed [14:0] m10_84;
   assign m10_84 =15'b0;

   // m10_85 = W*in
   wire signed [14:0] m10_85;
   assign m10_85 =15'b0;

   // m10_86 = W*in
   wire signed [14:0] m10_86;
   assign m10_86 =15'b0;

   // m10_87 = W*in
   wire signed [14:0] m10_87;
   assign m10_87 =15'b0;

   // m10_88 = W*in
   wire signed [14:0] m10_88;
   assign m10_88 =15'b0;

   // m10_89 = W*in
   wire signed [14:0] m10_89;
   assign m10_89 =15'b0;

   // m10_90 = W*in
   wire signed [14:0] m10_90;
   assign m10_90 =15'b0;

   // m10_91 = W*in
   wire signed [14:0] m10_91;
   assign m10_91 =15'b0;

   // m10_92 = W*in
   wire signed [14:0] m10_92;
   assign m10_92 ={ {3{in10[14]}} , in10[14:3] };

   // m10_93 = W*in
   wire signed [14:0] m10_93;
   assign m10_93 =15'b0;

   // m10_94 = W*in
   wire signed [14:0] m10_94;
   assign m10_94 =15'b0;

   // m10_95 = W*in
   wire signed [14:0] m10_95;
   assign m10_95 =15'b0;

   // m10_96 = W*in
   wire signed [14:0] m10_96;
   assign m10_96 =15'b0;

   // m10_97 = W*in
   wire signed [14:0] m10_97;
   assign m10_97 =15'b0;

   // m10_98 = W*in
   wire signed [14:0] m10_98;
   assign m10_98 =15'b0;

   // m10_99 = W*in
   wire signed [14:0] m10_99;
   assign m10_99 =15'b0;

   // m10_100 = W*in
   wire signed [14:0] m10_100;
   assign m10_100 =15'b0;

   // m11_1 = W*in
   wire signed [14:0] m11_1;
   assign m11_1 =15'b0;

   // m11_2 = W*in
   wire signed [14:0] m11_2;
   assign m11_2 =15'b0;

   // m11_3 = W*in
   wire signed [14:0] m11_3;
   assign m11_3 =15'b0;

   // m11_4 = W*in
   wire signed [14:0] m11_4;
   assign m11_4 =15'b0;

   // m11_5 = W*in
   wire signed [14:0] m11_5;
   assign m11_5 =15'b0;

   // m11_6 = W*in
   wire signed [14:0] m11_6;
   assign m11_6 =15'b0;

   // m11_7 = W*in
   wire signed [14:0] m11_7;
   assign m11_7 =15'b0;

   // m11_8 = W*in
   wire signed [14:0] m11_8;
   assign m11_8 =15'b0;

   // m11_9 = W*in
   wire signed [14:0] m11_9;
   assign m11_9 =15'b0;

   // m11_10 = W*in
   wire signed [14:0] m11_10;
   assign m11_10 =15'b0;

   // m11_11 = W*in
   wire signed [14:0] m11_11;
   assign m11_11 =15'b0;

   // m11_12 = W*in
   wire signed [14:0] m11_12;
   assign m11_12 =15'b0;

   // m11_13 = W*in
   wire signed [14:0] m11_13;
   assign m11_13 =15'b0;

   // m11_14 = W*in
   wire signed [14:0] m11_14;
   assign m11_14 =15'b0;

   // m11_15 = W*in
   wire signed [14:0] m11_15;
   assign m11_15 =15'b0;

   // m11_16 = W*in
   wire signed [14:0] m11_16;
   assign m11_16 =15'b0;

   // m11_17 = W*in
   wire signed [14:0] m11_17;
   assign m11_17 =15'b0;

   // m11_18 = W*in
   wire signed [14:0] m11_18;
   assign m11_18 =15'b0;

   // m11_19 = W*in
   wire signed [14:0] m11_19;
   assign m11_19 =15'b0;

   // m11_20 = W*in
   wire signed [14:0] m11_20;
   assign m11_20 =15'b0;

   // m11_21 = W*in
   wire signed [14:0] m11_21;
   assign m11_21 =15'b0;

   // m11_22 = W*in
   wire signed [14:0] m11_22;
   assign m11_22 =15'b0;

   // m11_23 = W*in
   wire signed [14:0] m11_23;
   assign m11_23 =15'b0;

   // m11_24 = W*in
   wire signed [14:0] m11_24;
   assign m11_24 =15'b0;

   // m11_25 = W*in
   wire signed [14:0] m11_25;
   assign m11_25 =15'b0;

   // m11_26 = W*in
   wire signed [14:0] m11_26;
   assign m11_26 =15'b0;

   // m11_27 = W*in
   wire signed [14:0] m11_27;
   assign m11_27 =15'b0;

   // m11_28 = W*in
   wire signed [14:0] m11_28;
   assign m11_28 =15'b0;

   // m11_29 = W*in
   wire signed [14:0] m11_29;
   assign m11_29 =15'b0;

   // m11_30 = W*in
   wire signed [14:0] m11_30;
   assign m11_30 =15'b0;

   // m11_31 = W*in
   wire signed [14:0] m11_31;
   assign m11_31 =15'b0;

   // m11_32 = W*in
   wire signed [14:0] m11_32;
   assign m11_32 =15'b0;

   // m11_33 = W*in
   wire signed [14:0] m11_33;
   assign m11_33 =15'b0;

   // m11_34 = W*in
   wire signed [14:0] m11_34;
   assign m11_34 =15'b0;

   // m11_35 = W*in
   wire signed [14:0] m11_35;
   assign m11_35 =15'b0;

   // m11_36 = W*in
   wire signed [14:0] m11_36;
   assign m11_36 =15'b0;

   // m11_37 = W*in
   wire signed [14:0] m11_37;
   assign m11_37 =15'b0;

   // m11_38 = W*in
   wire signed [14:0] m11_38;
   assign m11_38 =15'b0;

   // m11_39 = W*in
   wire signed [14:0] m11_39;
   assign m11_39 =15'b0;

   // m11_40 = W*in
   wire signed [14:0] m11_40;
   assign m11_40 =15'b0;

   // m11_41 = W*in
   wire signed [14:0] m11_41;
   assign m11_41 =15'b0;

   // m11_42 = W*in
   wire signed [14:0] m11_42;
   assign m11_42 =15'b0;

   // m11_43 = W*in
   wire signed [14:0] m11_43;
   assign m11_43 =15'b0;

   // m11_44 = W*in
   wire signed [14:0] m11_44;
   assign m11_44 =15'b0;

   // m11_45 = W*in
   wire signed [14:0] m11_45;
   assign m11_45 =15'b0;

   // m11_46 = W*in
   wire signed [14:0] m11_46;
   assign m11_46 =15'b0;

   // m11_47 = W*in
   wire signed [14:0] m11_47;
   assign m11_47 =15'b0;

   // m11_48 = W*in
   wire signed [14:0] m11_48;
   assign m11_48 =15'b0;

   // m11_49 = W*in
   wire signed [14:0] m11_49;
   assign m11_49 =15'b0;

   // m11_50 = W*in
   wire signed [14:0] m11_50;
   assign m11_50 =15'b0;

   // m11_51 = W*in
   wire signed [14:0] m11_51;
   assign m11_51 =15'b0;

   // m11_52 = W*in
   wire signed [14:0] m11_52;
   assign m11_52 =15'b0;

   // m11_53 = W*in
   wire signed [14:0] m11_53;
   assign m11_53 =15'b0;

   // m11_54 = W*in
   wire signed [14:0] m11_54;
   assign m11_54 =15'b0;

   // m11_55 = W*in
   wire signed [14:0] m11_55;
   assign m11_55 =15'b0;

   // m11_56 = W*in
   wire signed [14:0] m11_56;
   assign m11_56 =15'b0;

   // m11_57 = W*in
   wire signed [14:0] m11_57;
   assign m11_57 =15'b0;

   // m11_58 = W*in
   wire signed [14:0] m11_58;
   assign m11_58 =15'b0;

   // m11_59 = W*in
   wire signed [14:0] m11_59;
   assign m11_59 =15'b0;

   // m11_60 = W*in
   wire signed [14:0] m11_60;
   assign m11_60 =15'b0;

   // m11_61 = W*in
   wire signed [14:0] m11_61;
   assign m11_61 =15'b0;

   // m11_62 = W*in
   wire signed [14:0] m11_62;
   assign m11_62 =15'b0;

   // m11_63 = W*in
   wire signed [14:0] m11_63;
   assign m11_63 =15'b0;

   // m11_64 = W*in
   wire signed [14:0] m11_64;
   assign m11_64 =15'b0;

   // m11_65 = W*in
   wire signed [14:0] m11_65;
   assign m11_65 =15'b0;

   // m11_66 = W*in
   wire signed [14:0] m11_66;
   assign m11_66 =15'b0;

   // m11_67 = W*in
   wire signed [14:0] m11_67;
   assign m11_67 =15'b0;

   // m11_68 = W*in
   wire signed [14:0] m11_68;
   assign m11_68 =15'b0;

   // m11_69 = W*in
   wire signed [14:0] m11_69;
   assign m11_69 =15'b0;

   // m11_70 = W*in
   wire signed [14:0] m11_70;
   assign m11_70 =15'b0;

   // m11_71 = W*in
   wire signed [14:0] m11_71;
   assign m11_71 =15'b0;

   // m11_72 = W*in
   wire signed [14:0] m11_72;
   assign m11_72 =15'b0;

   // m11_73 = W*in
   wire signed [14:0] m11_73;
   assign m11_73 =15'b0;

   // m11_74 = W*in
   wire signed [14:0] m11_74;
   assign m11_74 =15'b0;

   // m11_75 = W*in
   wire signed [14:0] m11_75;
   assign m11_75 ={ {4{neg11[14]}} , neg11[14:4] };

   // m11_76 = W*in
   wire signed [14:0] m11_76;
   assign m11_76 =15'b0;

   // m11_77 = W*in
   wire signed [14:0] m11_77;
   assign m11_77 =15'b0;

   // m11_78 = W*in
   wire signed [14:0] m11_78;
   assign m11_78 =15'b0;

   // m11_79 = W*in
   wire signed [14:0] m11_79;
   assign m11_79 =15'b0;

   // m11_80 = W*in
   wire signed [14:0] m11_80;
   assign m11_80 =15'b0;

   // m11_81 = W*in
   wire signed [14:0] m11_81;
   assign m11_81 =15'b0;

   // m11_82 = W*in
   wire signed [14:0] m11_82;
   assign m11_82 =15'b0;

   // m11_83 = W*in
   wire signed [14:0] m11_83;
   assign m11_83 =15'b0;

   // m11_84 = W*in
   wire signed [14:0] m11_84;
   assign m11_84 =15'b0;

   // m11_85 = W*in
   wire signed [14:0] m11_85;
   assign m11_85 =15'b0;

   // m11_86 = W*in
   wire signed [14:0] m11_86;
   assign m11_86 =15'b0;

   // m11_87 = W*in
   wire signed [14:0] m11_87;
   assign m11_87 =15'b0;

   // m11_88 = W*in
   wire signed [14:0] m11_88;
   assign m11_88 =15'b0;

   // m11_89 = W*in
   wire signed [14:0] m11_89;
   assign m11_89 =15'b0;

   // m11_90 = W*in
   wire signed [14:0] m11_90;
   assign m11_90 =15'b0;

   // m11_91 = W*in
   wire signed [14:0] m11_91;
   assign m11_91 =15'b0;

   // m11_92 = W*in
   wire signed [14:0] m11_92;
   assign m11_92 =15'b0;

   // m11_93 = W*in
   wire signed [14:0] m11_93;
   assign m11_93 =15'b0;

   // m11_94 = W*in
   wire signed [14:0] m11_94;
   assign m11_94 =15'b0;

   // m11_95 = W*in
   wire signed [14:0] m11_95;
   assign m11_95 =15'b0;

   // m11_96 = W*in
   wire signed [14:0] m11_96;
   assign m11_96 =15'b0;

   // m11_97 = W*in
   wire signed [14:0] m11_97;
   assign m11_97 =15'b0;

   // m11_98 = W*in
   wire signed [14:0] m11_98;
   assign m11_98 =15'b0;

   // m11_99 = W*in
   wire signed [14:0] m11_99;
   assign m11_99 =15'b0;

   // m11_100 = W*in
   wire signed [14:0] m11_100;
   assign m11_100 =15'b0;

   // m12_1 = W*in
   wire signed [14:0] m12_1;
   assign m12_1 =15'b0;

   // m12_2 = W*in
   wire signed [14:0] m12_2;
   assign m12_2 =15'b0;

   // m12_3 = W*in
   wire signed [14:0] m12_3;
   assign m12_3 =15'b0;

   // m12_4 = W*in
   wire signed [14:0] m12_4;
   assign m12_4 =15'b0;

   // m12_5 = W*in
   wire signed [14:0] m12_5;
   assign m12_5 =15'b0;

   // m12_6 = W*in
   wire signed [14:0] m12_6;
   assign m12_6 =15'b0;

   // m12_7 = W*in
   wire signed [14:0] m12_7;
   assign m12_7 =15'b0;

   // m12_8 = W*in
   wire signed [14:0] m12_8;
   assign m12_8 =15'b0;

   // m12_9 = W*in
   wire signed [14:0] m12_9;
   assign m12_9 =15'b0;

   // m12_10 = W*in
   wire signed [14:0] m12_10;
   assign m12_10 =15'b0;

   // m12_11 = W*in
   wire signed [14:0] m12_11;
   assign m12_11 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_12 = W*in
   wire signed [14:0] m12_12;
   assign m12_12 =15'b0;

   // m12_13 = W*in
   wire signed [14:0] m12_13;
   assign m12_13 =15'b0;

   // m12_14 = W*in
   wire signed [14:0] m12_14;
   assign m12_14 =15'b0;

   // m12_15 = W*in
   wire signed [14:0] m12_15;
   assign m12_15 ={ {3{in12[14]}} , in12[14:3] };

   // m12_16 = W*in
   wire signed [14:0] m12_16;
   assign m12_16 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_17 = W*in
   wire signed [14:0] m12_17;
   assign m12_17 =15'b0;

   // m12_18 = W*in
   wire signed [14:0] m12_18;
   assign m12_18 =15'b0;

   // m12_19 = W*in
   wire signed [14:0] m12_19;
   assign m12_19 =15'b0;

   // m12_20 = W*in
   wire signed [14:0] m12_20;
   assign m12_20 =15'b0;

   // m12_21 = W*in
   wire signed [14:0] m12_21;
   assign m12_21 =15'b0;

   // m12_22 = W*in
   wire signed [14:0] m12_22;
   assign m12_22 =15'b0;

   // m12_23 = W*in
   wire signed [14:0] m12_23;
   assign m12_23 =15'b0;

   // m12_24 = W*in
   wire signed [14:0] m12_24;
   assign m12_24 ={ {3{in12[14]}} , in12[14:3] };

   // m12_25 = W*in
   wire signed [14:0] m12_25;
   assign m12_25 =15'b0;

   // m12_26 = W*in
   wire signed [14:0] m12_26;
   assign m12_26 =15'b0;

   // m12_27 = W*in
   wire signed [14:0] m12_27;
   assign m12_27 =15'b0;

   // m12_28 = W*in
   wire signed [14:0] m12_28;
   assign m12_28 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_29 = W*in
   wire signed [14:0] m12_29;
   assign m12_29 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_30 = W*in
   wire signed [14:0] m12_30;
   assign m12_30 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_31 = W*in
   wire signed [14:0] m12_31;
   assign m12_31 =15'b0;

   // m12_32 = W*in
   wire signed [14:0] m12_32;
   assign m12_32 ={ {4{in12[14]}} , in12[14:4] };

   // m12_33 = W*in
   wire signed [14:0] m12_33;
   assign m12_33 =15'b0;

   // m12_34 = W*in
   wire signed [14:0] m12_34;
   assign m12_34 =15'b0;

   // m12_35 = W*in
   wire signed [14:0] m12_35;
   assign m12_35 ={ {3{in12[14]}} , in12[14:3] };

   // m12_36 = W*in
   wire signed [14:0] m12_36;
   assign m12_36 =15'b0;

   // m12_37 = W*in
   wire signed [14:0] m12_37;
   assign m12_37 =15'b0;

   // m12_38 = W*in
   wire signed [14:0] m12_38;
   assign m12_38 ={ {3{neg12[14]}} , neg12[14:3] };

   // m12_39 = W*in
   wire signed [14:0] m12_39;
   assign m12_39 ={ {3{in12[14]}} , in12[14:3] };

   // m12_40 = W*in
   wire signed [14:0] m12_40;
   assign m12_40 =15'b0;

   // m12_41 = W*in
   wire signed [14:0] m12_41;
   assign m12_41 =15'b0;

   // m12_42 = W*in
   wire signed [14:0] m12_42;
   assign m12_42 ={ {3{in12[14]}} , in12[14:3] };

   // m12_43 = W*in
   wire signed [14:0] m12_43;
   assign m12_43 =15'b0;

   // m12_44 = W*in
   wire signed [14:0] m12_44;
   assign m12_44 =15'b0;

   // m12_45 = W*in
   wire signed [14:0] m12_45;
   assign m12_45 =15'b0;

   // m12_46 = W*in
   wire signed [14:0] m12_46;
   assign m12_46 =15'b0;

   // m12_47 = W*in
   wire signed [14:0] m12_47;
   assign m12_47 =15'b0;

   // m12_48 = W*in
   wire signed [14:0] m12_48;
   assign m12_48 =15'b0;

   // m12_49 = W*in
   wire signed [14:0] m12_49;
   assign m12_49 =15'b0;

   // m12_50 = W*in
   wire signed [14:0] m12_50;
   assign m12_50 =15'b0;

   // m12_51 = W*in
   wire signed [14:0] m12_51;
   assign m12_51 =15'b0;

   // m12_52 = W*in
   wire signed [14:0] m12_52;
   assign m12_52 =15'b0;

   // m12_53 = W*in
   wire signed [14:0] m12_53;
   assign m12_53 =15'b0;

   // m12_54 = W*in
   wire signed [14:0] m12_54;
   assign m12_54 =15'b0;

   // m12_55 = W*in
   wire signed [14:0] m12_55;
   assign m12_55 =15'b0;

   // m12_56 = W*in
   wire signed [14:0] m12_56;
   assign m12_56 =15'b0;

   // m12_57 = W*in
   wire signed [14:0] m12_57;
   assign m12_57 =15'b0;

   // m12_58 = W*in
   wire signed [14:0] m12_58;
   assign m12_58 =15'b0;

   // m12_59 = W*in
   wire signed [14:0] m12_59;
   assign m12_59 =15'b0;

   // m12_60 = W*in
   wire signed [14:0] m12_60;
   assign m12_60 =15'b0;

   // m12_61 = W*in
   wire signed [14:0] m12_61;
   assign m12_61 =15'b0;

   // m12_62 = W*in
   wire signed [14:0] m12_62;
   assign m12_62 =15'b0;

   // m12_63 = W*in
   wire signed [14:0] m12_63;
   assign m12_63 ={ {4{in12[14]}} , in12[14:4] };

   // m12_64 = W*in
   wire signed [14:0] m12_64;
   assign m12_64 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_65 = W*in
   wire signed [14:0] m12_65;
   assign m12_65 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_66 = W*in
   wire signed [14:0] m12_66;
   assign m12_66 =15'b0;

   // m12_67 = W*in
   wire signed [14:0] m12_67;
   assign m12_67 =15'b0;

   // m12_68 = W*in
   wire signed [14:0] m12_68;
   assign m12_68 =15'b0;

   // m12_69 = W*in
   wire signed [14:0] m12_69;
   assign m12_69 =15'b0;

   // m12_70 = W*in
   wire signed [14:0] m12_70;
   assign m12_70 =15'b0;

   // m12_71 = W*in
   wire signed [14:0] m12_71;
   assign m12_71 =15'b0;

   // m12_72 = W*in
   wire signed [14:0] m12_72;
   assign m12_72 =15'b0;

   // m12_73 = W*in
   wire signed [14:0] m12_73;
   assign m12_73 =15'b0;

   // m12_74 = W*in
   wire signed [14:0] m12_74;
   assign m12_74 =15'b0;

   // m12_75 = W*in
   wire signed [14:0] m12_75;
   assign m12_75 =15'b0;

   // m12_76 = W*in
   wire signed [14:0] m12_76;
   assign m12_76 =15'b0;

   // m12_77 = W*in
   wire signed [14:0] m12_77;
   assign m12_77 ={ {3{neg12[14]}} , neg12[14:3] };

   // m12_78 = W*in
   wire signed [14:0] m12_78;
   assign m12_78 =15'b0;

   // m12_79 = W*in
   wire signed [14:0] m12_79;
   assign m12_79 =15'b0;

   // m12_80 = W*in
   wire signed [14:0] m12_80;
   assign m12_80 =15'b0;

   // m12_81 = W*in
   wire signed [14:0] m12_81;
   assign m12_81 =15'b0;

   // m12_82 = W*in
   wire signed [14:0] m12_82;
   assign m12_82 =15'b0;

   // m12_83 = W*in
   wire signed [14:0] m12_83;
   assign m12_83 =15'b0;

   // m12_84 = W*in
   wire signed [14:0] m12_84;
   assign m12_84 =15'b0;

   // m12_85 = W*in
   wire signed [14:0] m12_85;
   assign m12_85 =15'b0;

   // m12_86 = W*in
   wire signed [14:0] m12_86;
   assign m12_86 =15'b0;

   // m12_87 = W*in
   wire signed [14:0] m12_87;
   assign m12_87 =15'b0;

   // m12_88 = W*in
   wire signed [14:0] m12_88;
   assign m12_88 =15'b0;

   // m12_89 = W*in
   wire signed [14:0] m12_89;
   assign m12_89 =15'b0;

   // m12_90 = W*in
   wire signed [14:0] m12_90;
   assign m12_90 =15'b0;

   // m12_91 = W*in
   wire signed [14:0] m12_91;
   assign m12_91 =15'b0;

   // m12_92 = W*in
   wire signed [14:0] m12_92;
   assign m12_92 ={ {3{neg12[14]}} , neg12[14:3] };

   // m12_93 = W*in
   wire signed [14:0] m12_93;
   assign m12_93 =15'b0;

   // m12_94 = W*in
   wire signed [14:0] m12_94;
   assign m12_94 ={ {3{in12[14]}} , in12[14:3] };

   // m12_95 = W*in
   wire signed [14:0] m12_95;
   assign m12_95 =15'b0;

   // m12_96 = W*in
   wire signed [14:0] m12_96;
   assign m12_96 =15'b0;

   // m12_97 = W*in
   wire signed [14:0] m12_97;
   assign m12_97 ={ {4{neg12[14]}} , neg12[14:4] };

   // m12_98 = W*in
   wire signed [14:0] m12_98;
   assign m12_98 ={ {4{in12[14]}} , in12[14:4] };

   // m12_99 = W*in
   wire signed [14:0] m12_99;
   assign m12_99 ={ {3{neg12[14]}} , neg12[14:3] };

   // m12_100 = W*in
   wire signed [14:0] m12_100;
   assign m12_100 =15'b0;

   // m13_1 = W*in
   wire signed [14:0] m13_1;
   assign m13_1 =15'b0;

   // m13_2 = W*in
   wire signed [14:0] m13_2;
   assign m13_2 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_3 = W*in
   wire signed [14:0] m13_3;
   assign m13_3 =15'b0;

   // m13_4 = W*in
   wire signed [14:0] m13_4;
   assign m13_4 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_5 = W*in
   wire signed [14:0] m13_5;
   assign m13_5 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_6 = W*in
   wire signed [14:0] m13_6;
   assign m13_6 =15'b0;

   // m13_7 = W*in
   wire signed [14:0] m13_7;
   assign m13_7 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_8 = W*in
   wire signed [14:0] m13_8;
   assign m13_8 =15'b0;

   // m13_9 = W*in
   wire signed [14:0] m13_9;
   assign m13_9 =15'b0;

   // m13_10 = W*in
   wire signed [14:0] m13_10;
   assign m13_10 =15'b0;

   // m13_11 = W*in
   wire signed [14:0] m13_11;
   assign m13_11 =15'b0;

   // m13_12 = W*in
   wire signed [14:0] m13_12;
   assign m13_12 =15'b0;

   // m13_13 = W*in
   wire signed [14:0] m13_13;
   assign m13_13 =15'b0;

   // m13_14 = W*in
   wire signed [14:0] m13_14;
   assign m13_14 =15'b0;

   // m13_15 = W*in
   wire signed [14:0] m13_15;
   assign m13_15 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_16 = W*in
   wire signed [14:0] m13_16;
   assign m13_16 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_17 = W*in
   wire signed [14:0] m13_17;
   assign m13_17 ={ {3{in13[14]}} , in13[14:3] };

   // m13_18 = W*in
   wire signed [14:0] m13_18;
   assign m13_18 =15'b0;

   // m13_19 = W*in
   wire signed [14:0] m13_19;
   assign m13_19 =15'b0;

   // m13_20 = W*in
   wire signed [14:0] m13_20;
   assign m13_20 ={ {4{in13[14]}} , in13[14:4] };

   // m13_21 = W*in
   wire signed [14:0] m13_21;
   assign m13_21 ={ {3{in13[14]}} , in13[14:3] };

   // m13_22 = W*in
   wire signed [14:0] m13_22;
   assign m13_22 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_23 = W*in
   wire signed [14:0] m13_23;
   assign m13_23 =15'b0;

   // m13_24 = W*in
   wire signed [14:0] m13_24;
   assign m13_24 =15'b0;

   // m13_25 = W*in
   wire signed [14:0] m13_25;
   assign m13_25 =15'b0;

   // m13_26 = W*in
   wire signed [14:0] m13_26;
   assign m13_26 ={ {4{neg13[14]}} , neg13[14:4] };

   // m13_27 = W*in
   wire signed [14:0] m13_27;
   assign m13_27 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_28 = W*in
   wire signed [14:0] m13_28;
   assign m13_28 =15'b0;

   // m13_29 = W*in
   wire signed [14:0] m13_29;
   assign m13_29 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_30 = W*in
   wire signed [14:0] m13_30;
   assign m13_30 =15'b0;

   // m13_31 = W*in
   wire signed [14:0] m13_31;
   assign m13_31 =15'b0;

   // m13_32 = W*in
   wire signed [14:0] m13_32;
   assign m13_32 =15'b0;

   // m13_33 = W*in
   wire signed [14:0] m13_33;
   assign m13_33 ={ {4{neg13[14]}} , neg13[14:4] };

   // m13_34 = W*in
   wire signed [14:0] m13_34;
   assign m13_34 =15'b0;

   // m13_35 = W*in
   wire signed [14:0] m13_35;
   assign m13_35 =15'b0;

   // m13_36 = W*in
   wire signed [14:0] m13_36;
   assign m13_36 =15'b0;

   // m13_37 = W*in
   wire signed [14:0] m13_37;
   assign m13_37 =15'b0;

   // m13_38 = W*in
   wire signed [14:0] m13_38;
   assign m13_38 =15'b0;

   // m13_39 = W*in
   wire signed [14:0] m13_39;
   assign m13_39 ={ {4{in13[14]}} , in13[14:4] };

   // m13_40 = W*in
   wire signed [14:0] m13_40;
   assign m13_40 =15'b0;

   // m13_41 = W*in
   wire signed [14:0] m13_41;
   assign m13_41 =15'b0;

   // m13_42 = W*in
   wire signed [14:0] m13_42;
   assign m13_42 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_43 = W*in
   wire signed [14:0] m13_43;
   assign m13_43 =15'b0;

   // m13_44 = W*in
   wire signed [14:0] m13_44;
   assign m13_44 ={ {2{in13[14]}} , in13[14:2] };

   // m13_45 = W*in
   wire signed [14:0] m13_45;
   assign m13_45 ={ {3{in13[14]}} , in13[14:3] };

   // m13_46 = W*in
   wire signed [14:0] m13_46;
   assign m13_46 =15'b0;

   // m13_47 = W*in
   wire signed [14:0] m13_47;
   assign m13_47 =15'b0;

   // m13_48 = W*in
   wire signed [14:0] m13_48;
   assign m13_48 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_49 = W*in
   wire signed [14:0] m13_49;
   assign m13_49 =15'b0;

   // m13_50 = W*in
   wire signed [14:0] m13_50;
   assign m13_50 =15'b0;

   // m13_51 = W*in
   wire signed [14:0] m13_51;
   assign m13_51 =15'b0;

   // m13_52 = W*in
   wire signed [14:0] m13_52;
   assign m13_52 =15'b0;

   // m13_53 = W*in
   wire signed [14:0] m13_53;
   assign m13_53 =15'b0;

   // m13_54 = W*in
   wire signed [14:0] m13_54;
   assign m13_54 =15'b0;

   // m13_55 = W*in
   wire signed [14:0] m13_55;
   assign m13_55 =15'b0;

   // m13_56 = W*in
   wire signed [14:0] m13_56;
   assign m13_56 =15'b0;

   // m13_57 = W*in
   wire signed [14:0] m13_57;
   assign m13_57 =15'b0;

   // m13_58 = W*in
   wire signed [14:0] m13_58;
   assign m13_58 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_59 = W*in
   wire signed [14:0] m13_59;
   assign m13_59 =15'b0;

   // m13_60 = W*in
   wire signed [14:0] m13_60;
   assign m13_60 ={ {4{neg13[14]}} , neg13[14:4] };

   // m13_61 = W*in
   wire signed [14:0] m13_61;
   assign m13_61 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_62 = W*in
   wire signed [14:0] m13_62;
   assign m13_62 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_63 = W*in
   wire signed [14:0] m13_63;
   assign m13_63 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_64 = W*in
   wire signed [14:0] m13_64;
   assign m13_64 =15'b0;

   // m13_65 = W*in
   wire signed [14:0] m13_65;
   assign m13_65 =15'b0;

   // m13_66 = W*in
   wire signed [14:0] m13_66;
   assign m13_66 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_67 = W*in
   wire signed [14:0] m13_67;
   assign m13_67 =15'b0;

   // m13_68 = W*in
   wire signed [14:0] m13_68;
   assign m13_68 ={ {4{neg13[14]}} , neg13[14:4] };

   // m13_69 = W*in
   wire signed [14:0] m13_69;
   assign m13_69 =15'b0;

   // m13_70 = W*in
   wire signed [14:0] m13_70;
   assign m13_70 =15'b0;

   // m13_71 = W*in
   wire signed [14:0] m13_71;
   assign m13_71 =15'b0;

   // m13_72 = W*in
   wire signed [14:0] m13_72;
   assign m13_72 =15'b0;

   // m13_73 = W*in
   wire signed [14:0] m13_73;
   assign m13_73 =15'b0;

   // m13_74 = W*in
   wire signed [14:0] m13_74;
   assign m13_74 =15'b0;

   // m13_75 = W*in
   wire signed [14:0] m13_75;
   assign m13_75 ={ {3{in13[14]}} , in13[14:3] };

   // m13_76 = W*in
   wire signed [14:0] m13_76;
   assign m13_76 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_77 = W*in
   wire signed [14:0] m13_77;
   assign m13_77 =15'b0;

   // m13_78 = W*in
   wire signed [14:0] m13_78;
   assign m13_78 ={ {3{in13[14]}} , in13[14:3] };

   // m13_79 = W*in
   wire signed [14:0] m13_79;
   assign m13_79 =15'b0;

   // m13_80 = W*in
   wire signed [14:0] m13_80;
   assign m13_80 =15'b0;

   // m13_81 = W*in
   wire signed [14:0] m13_81;
   assign m13_81 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_82 = W*in
   wire signed [14:0] m13_82;
   assign m13_82 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_83 = W*in
   wire signed [14:0] m13_83;
   assign m13_83 =15'b0;

   // m13_84 = W*in
   wire signed [14:0] m13_84;
   assign m13_84 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_85 = W*in
   wire signed [14:0] m13_85;
   assign m13_85 ={ {3{neg13[14]}} , neg13[14:3] };

   // m13_86 = W*in
   wire signed [14:0] m13_86;
   assign m13_86 =15'b0;

   // m13_87 = W*in
   wire signed [14:0] m13_87;
   assign m13_87 =15'b0;

   // m13_88 = W*in
   wire signed [14:0] m13_88;
   assign m13_88 =15'b0;

   // m13_89 = W*in
   wire signed [14:0] m13_89;
   assign m13_89 =15'b0;

   // m13_90 = W*in
   wire signed [14:0] m13_90;
   assign m13_90 =15'b0;

   // m13_91 = W*in
   wire signed [14:0] m13_91;
   assign m13_91 =15'b0;

   // m13_92 = W*in
   wire signed [14:0] m13_92;
   assign m13_92 =15'b0;

   // m13_93 = W*in
   wire signed [14:0] m13_93;
   assign m13_93 =15'b0;

   // m13_94 = W*in
   wire signed [14:0] m13_94;
   assign m13_94 =15'b0;

   // m13_95 = W*in
   wire signed [14:0] m13_95;
   assign m13_95 =15'b0;

   // m13_96 = W*in
   wire signed [14:0] m13_96;
   assign m13_96 ={ {3{in13[14]}} , in13[14:3] };

   // m13_97 = W*in
   wire signed [14:0] m13_97;
   assign m13_97 =15'b0;

   // m13_98 = W*in
   wire signed [14:0] m13_98;
   assign m13_98 =15'b0;

   // m13_99 = W*in
   wire signed [14:0] m13_99;
   assign m13_99 =15'b0;

   // m13_100 = W*in
   wire signed [14:0] m13_100;
   assign m13_100 ={ {3{neg13[14]}} , neg13[14:3] };

   // m14_1 = W*in
   wire signed [14:0] m14_1;
   assign m14_1 ={ {3{in14[14]}} , in14[14:3] };

   // m14_2 = W*in
   wire signed [14:0] m14_2;
   assign m14_2 =15'b0;

   // m14_3 = W*in
   wire signed [14:0] m14_3;
   assign m14_3 =15'b0;

   // m14_4 = W*in
   wire signed [14:0] m14_4;
   assign m14_4 ={ {4{neg14[14]}} , neg14[14:4] };

   // m14_5 = W*in
   wire signed [14:0] m14_5;
   assign m14_5 =15'b0;

   // m14_6 = W*in
   wire signed [14:0] m14_6;
   assign m14_6 =15'b0;

   // m14_7 = W*in
   wire signed [14:0] m14_7;
   assign m14_7 =15'b0;

   // m14_8 = W*in
   wire signed [14:0] m14_8;
   assign m14_8 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_9 = W*in
   wire signed [14:0] m14_9;
   assign m14_9 =15'b0;

   // m14_10 = W*in
   wire signed [14:0] m14_10;
   assign m14_10 =15'b0;

   // m14_11 = W*in
   wire signed [14:0] m14_11;
   assign m14_11 =15'b0;

   // m14_12 = W*in
   wire signed [14:0] m14_12;
   assign m14_12 ={ {4{in14[14]}} , in14[14:4] };

   // m14_13 = W*in
   wire signed [14:0] m14_13;
   assign m14_13 =15'b0;

   // m14_14 = W*in
   wire signed [14:0] m14_14;
   assign m14_14 =15'b0;

   // m14_15 = W*in
   wire signed [14:0] m14_15;
   assign m14_15 =15'b0;

   // m14_16 = W*in
   wire signed [14:0] m14_16;
   assign m14_16 =15'b0;

   // m14_17 = W*in
   wire signed [14:0] m14_17;
   assign m14_17 =15'b0;

   // m14_18 = W*in
   wire signed [14:0] m14_18;
   assign m14_18 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_19 = W*in
   wire signed [14:0] m14_19;
   assign m14_19 ={ {4{neg14[14]}} , neg14[14:4] };

   // m14_20 = W*in
   wire signed [14:0] m14_20;
   assign m14_20 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_21 = W*in
   wire signed [14:0] m14_21;
   assign m14_21 =15'b0;

   // m14_22 = W*in
   wire signed [14:0] m14_22;
   assign m14_22 =15'b0;

   // m14_23 = W*in
   wire signed [14:0] m14_23;
   assign m14_23 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_24 = W*in
   wire signed [14:0] m14_24;
   assign m14_24 =15'b0;

   // m14_25 = W*in
   wire signed [14:0] m14_25;
   assign m14_25 ={ {3{in14[14]}} , in14[14:3] };

   // m14_26 = W*in
   wire signed [14:0] m14_26;
   assign m14_26 ={ {4{in14[14]}} , in14[14:4] };

   // m14_27 = W*in
   wire signed [14:0] m14_27;
   assign m14_27 =15'b0;

   // m14_28 = W*in
   wire signed [14:0] m14_28;
   assign m14_28 =15'b0;

   // m14_29 = W*in
   wire signed [14:0] m14_29;
   assign m14_29 ={ {4{in14[14]}} , in14[14:4] };

   // m14_30 = W*in
   wire signed [14:0] m14_30;
   assign m14_30 =15'b0;

   // m14_31 = W*in
   wire signed [14:0] m14_31;
   assign m14_31 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_32 = W*in
   wire signed [14:0] m14_32;
   assign m14_32 =15'b0;

   // m14_33 = W*in
   wire signed [14:0] m14_33;
   assign m14_33 =15'b0;

   // m14_34 = W*in
   wire signed [14:0] m14_34;
   assign m14_34 =15'b0;

   // m14_35 = W*in
   wire signed [14:0] m14_35;
   assign m14_35 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_36 = W*in
   wire signed [14:0] m14_36;
   assign m14_36 =15'b0;

   // m14_37 = W*in
   wire signed [14:0] m14_37;
   assign m14_37 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_38 = W*in
   wire signed [14:0] m14_38;
   assign m14_38 =15'b0;

   // m14_39 = W*in
   wire signed [14:0] m14_39;
   assign m14_39 =15'b0;

   // m14_40 = W*in
   wire signed [14:0] m14_40;
   assign m14_40 =15'b0;

   // m14_41 = W*in
   wire signed [14:0] m14_41;
   assign m14_41 =15'b0;

   // m14_42 = W*in
   wire signed [14:0] m14_42;
   assign m14_42 =15'b0;

   // m14_43 = W*in
   wire signed [14:0] m14_43;
   assign m14_43 ={ {3{in14[14]}} , in14[14:3] };

   // m14_44 = W*in
   wire signed [14:0] m14_44;
   assign m14_44 =15'b0;

   // m14_45 = W*in
   wire signed [14:0] m14_45;
   assign m14_45 =15'b0;

   // m14_46 = W*in
   wire signed [14:0] m14_46;
   assign m14_46 =15'b0;

   // m14_47 = W*in
   wire signed [14:0] m14_47;
   assign m14_47 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_48 = W*in
   wire signed [14:0] m14_48;
   assign m14_48 =15'b0;

   // m14_49 = W*in
   wire signed [14:0] m14_49;
   assign m14_49 =15'b0;

   // m14_50 = W*in
   wire signed [14:0] m14_50;
   assign m14_50 ={ {3{in14[14]}} , in14[14:3] };

   // m14_51 = W*in
   wire signed [14:0] m14_51;
   assign m14_51 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_52 = W*in
   wire signed [14:0] m14_52;
   assign m14_52 =15'b0;

   // m14_53 = W*in
   wire signed [14:0] m14_53;
   assign m14_53 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_54 = W*in
   wire signed [14:0] m14_54;
   assign m14_54 =15'b0;

   // m14_55 = W*in
   wire signed [14:0] m14_55;
   assign m14_55 =15'b0;

   // m14_56 = W*in
   wire signed [14:0] m14_56;
   assign m14_56 =15'b0;

   // m14_57 = W*in
   wire signed [14:0] m14_57;
   assign m14_57 =15'b0;

   // m14_58 = W*in
   wire signed [14:0] m14_58;
   assign m14_58 =15'b0;

   // m14_59 = W*in
   wire signed [14:0] m14_59;
   assign m14_59 =15'b0;

   // m14_60 = W*in
   wire signed [14:0] m14_60;
   assign m14_60 =15'b0;

   // m14_61 = W*in
   wire signed [14:0] m14_61;
   assign m14_61 =15'b0;

   // m14_62 = W*in
   wire signed [14:0] m14_62;
   assign m14_62 =15'b0;

   // m14_63 = W*in
   wire signed [14:0] m14_63;
   assign m14_63 ={ {4{neg14[14]}} , neg14[14:4] };

   // m14_64 = W*in
   wire signed [14:0] m14_64;
   assign m14_64 =15'b0;

   // m14_65 = W*in
   wire signed [14:0] m14_65;
   assign m14_65 =15'b0;

   // m14_66 = W*in
   wire signed [14:0] m14_66;
   assign m14_66 =15'b0;

   // m14_67 = W*in
   wire signed [14:0] m14_67;
   assign m14_67 =15'b0;

   // m14_68 = W*in
   wire signed [14:0] m14_68;
   assign m14_68 =15'b0;

   // m14_69 = W*in
   wire signed [14:0] m14_69;
   assign m14_69 =15'b0;

   // m14_70 = W*in
   wire signed [14:0] m14_70;
   assign m14_70 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_71 = W*in
   wire signed [14:0] m14_71;
   assign m14_71 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_72 = W*in
   wire signed [14:0] m14_72;
   assign m14_72 =15'b0;

   // m14_73 = W*in
   wire signed [14:0] m14_73;
   assign m14_73 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_74 = W*in
   wire signed [14:0] m14_74;
   assign m14_74 ={ {4{neg14[14]}} , neg14[14:4] };

   // m14_75 = W*in
   wire signed [14:0] m14_75;
   assign m14_75 =15'b0;

   // m14_76 = W*in
   wire signed [14:0] m14_76;
   assign m14_76 =15'b0;

   // m14_77 = W*in
   wire signed [14:0] m14_77;
   assign m14_77 =15'b0;

   // m14_78 = W*in
   wire signed [14:0] m14_78;
   assign m14_78 =15'b0;

   // m14_79 = W*in
   wire signed [14:0] m14_79;
   assign m14_79 ={ {3{in14[14]}} , in14[14:3] };

   // m14_80 = W*in
   wire signed [14:0] m14_80;
   assign m14_80 ={ {3{in14[14]}} , in14[14:3] };

   // m14_81 = W*in
   wire signed [14:0] m14_81;
   assign m14_81 =15'b0;

   // m14_82 = W*in
   wire signed [14:0] m14_82;
   assign m14_82 =15'b0;

   // m14_83 = W*in
   wire signed [14:0] m14_83;
   assign m14_83 ={ {4{neg14[14]}} , neg14[14:4] };

   // m14_84 = W*in
   wire signed [14:0] m14_84;
   assign m14_84 ={ {3{in14[14]}} , in14[14:3] };

   // m14_85 = W*in
   wire signed [14:0] m14_85;
   assign m14_85 =15'b0;

   // m14_86 = W*in
   wire signed [14:0] m14_86;
   assign m14_86 ={ {3{in14[14]}} , in14[14:3] };

   // m14_87 = W*in
   wire signed [14:0] m14_87;
   assign m14_87 =15'b0;

   // m14_88 = W*in
   wire signed [14:0] m14_88;
   assign m14_88 =15'b0;

   // m14_89 = W*in
   wire signed [14:0] m14_89;
   assign m14_89 ={ {3{neg14[14]}} , neg14[14:3] };

   // m14_90 = W*in
   wire signed [14:0] m14_90;
   assign m14_90 =15'b0;

   // m14_91 = W*in
   wire signed [14:0] m14_91;
   assign m14_91 =15'b0;

   // m14_92 = W*in
   wire signed [14:0] m14_92;
   assign m14_92 =15'b0;

   // m14_93 = W*in
   wire signed [14:0] m14_93;
   assign m14_93 =15'b0;

   // m14_94 = W*in
   wire signed [14:0] m14_94;
   assign m14_94 ={ {3{in14[14]}} , in14[14:3] };

   // m14_95 = W*in
   wire signed [14:0] m14_95;
   assign m14_95 ={ {4{in14[14]}} , in14[14:4] };

   // m14_96 = W*in
   wire signed [14:0] m14_96;
   assign m14_96 =15'b0;

   // m14_97 = W*in
   wire signed [14:0] m14_97;
   assign m14_97 =15'b0;

   // m14_98 = W*in
   wire signed [14:0] m14_98;
   assign m14_98 =15'b0;

   // m14_99 = W*in
   wire signed [14:0] m14_99;
   assign m14_99 =15'b0;

   // m14_100 = W*in
   wire signed [14:0] m14_100;
   assign m14_100 ={ {4{neg14[14]}} , neg14[14:4] };

   // m15_1 = W*in
   wire signed [14:0] m15_1;
   assign m15_1 =15'b0;

   // m15_2 = W*in
   wire signed [14:0] m15_2;
   assign m15_2 =15'b0;

   // m15_3 = W*in
   wire signed [14:0] m15_3;
   assign m15_3 =15'b0;

   // m15_4 = W*in
   wire signed [14:0] m15_4;
   assign m15_4 =15'b0;

   // m15_5 = W*in
   wire signed [14:0] m15_5;
   assign m15_5 =15'b0;

   // m15_6 = W*in
   wire signed [14:0] m15_6;
   assign m15_6 =15'b0;

   // m15_7 = W*in
   wire signed [14:0] m15_7;
   assign m15_7 =15'b0;

   // m15_8 = W*in
   wire signed [14:0] m15_8;
   assign m15_8 =15'b0;

   // m15_9 = W*in
   wire signed [14:0] m15_9;
   assign m15_9 =15'b0;

   // m15_10 = W*in
   wire signed [14:0] m15_10;
   assign m15_10 =15'b0;

   // m15_11 = W*in
   wire signed [14:0] m15_11;
   assign m15_11 =15'b0;

   // m15_12 = W*in
   wire signed [14:0] m15_12;
   assign m15_12 =15'b0;

   // m15_13 = W*in
   wire signed [14:0] m15_13;
   assign m15_13 =15'b0;

   // m15_14 = W*in
   wire signed [14:0] m15_14;
   assign m15_14 ={ {3{neg15[14]}} , neg15[14:3] };

   // m15_15 = W*in
   wire signed [14:0] m15_15;
   assign m15_15 =15'b0;

   // m15_16 = W*in
   wire signed [14:0] m15_16;
   assign m15_16 =15'b0;

   // m15_17 = W*in
   wire signed [14:0] m15_17;
   assign m15_17 =15'b0;

   // m15_18 = W*in
   wire signed [14:0] m15_18;
   assign m15_18 ={ {4{in15[14]}} , in15[14:4] };

   // m15_19 = W*in
   wire signed [14:0] m15_19;
   assign m15_19 =15'b0;

   // m15_20 = W*in
   wire signed [14:0] m15_20;
   assign m15_20 =15'b0;

   // m15_21 = W*in
   wire signed [14:0] m15_21;
   assign m15_21 =15'b0;

   // m15_22 = W*in
   wire signed [14:0] m15_22;
   assign m15_22 =15'b0;

   // m15_23 = W*in
   wire signed [14:0] m15_23;
   assign m15_23 =15'b0;

   // m15_24 = W*in
   wire signed [14:0] m15_24;
   assign m15_24 =15'b0;

   // m15_25 = W*in
   wire signed [14:0] m15_25;
   assign m15_25 =15'b0;

   // m15_26 = W*in
   wire signed [14:0] m15_26;
   assign m15_26 =15'b0;

   // m15_27 = W*in
   wire signed [14:0] m15_27;
   assign m15_27 =15'b0;

   // m15_28 = W*in
   wire signed [14:0] m15_28;
   assign m15_28 =15'b0;

   // m15_29 = W*in
   wire signed [14:0] m15_29;
   assign m15_29 ={ {4{neg15[14]}} , neg15[14:4] };

   // m15_30 = W*in
   wire signed [14:0] m15_30;
   assign m15_30 =15'b0;

   // m15_31 = W*in
   wire signed [14:0] m15_31;
   assign m15_31 =15'b0;

   // m15_32 = W*in
   wire signed [14:0] m15_32;
   assign m15_32 =15'b0;

   // m15_33 = W*in
   wire signed [14:0] m15_33;
   assign m15_33 =15'b0;

   // m15_34 = W*in
   wire signed [14:0] m15_34;
   assign m15_34 =15'b0;

   // m15_35 = W*in
   wire signed [14:0] m15_35;
   assign m15_35 =15'b0;

   // m15_36 = W*in
   wire signed [14:0] m15_36;
   assign m15_36 =15'b0;

   // m15_37 = W*in
   wire signed [14:0] m15_37;
   assign m15_37 ={ {3{neg15[14]}} , neg15[14:3] };

   // m15_38 = W*in
   wire signed [14:0] m15_38;
   assign m15_38 =15'b0;

   // m15_39 = W*in
   wire signed [14:0] m15_39;
   assign m15_39 ={ {3{neg15[14]}} , neg15[14:3] };

   // m15_40 = W*in
   wire signed [14:0] m15_40;
   assign m15_40 =15'b0;

   // m15_41 = W*in
   wire signed [14:0] m15_41;
   assign m15_41 =15'b0;

   // m15_42 = W*in
   wire signed [14:0] m15_42;
   assign m15_42 =15'b0;

   // m15_43 = W*in
   wire signed [14:0] m15_43;
   assign m15_43 =15'b0;

   // m15_44 = W*in
   wire signed [14:0] m15_44;
   assign m15_44 =15'b0;

   // m15_45 = W*in
   wire signed [14:0] m15_45;
   assign m15_45 =15'b0;

   // m15_46 = W*in
   wire signed [14:0] m15_46;
   assign m15_46 =15'b0;

   // m15_47 = W*in
   wire signed [14:0] m15_47;
   assign m15_47 =15'b0;

   // m15_48 = W*in
   wire signed [14:0] m15_48;
   assign m15_48 =15'b0;

   // m15_49 = W*in
   wire signed [14:0] m15_49;
   assign m15_49 =15'b0;

   // m15_50 = W*in
   wire signed [14:0] m15_50;
   assign m15_50 =15'b0;

   // m15_51 = W*in
   wire signed [14:0] m15_51;
   assign m15_51 =15'b0;

   // m15_52 = W*in
   wire signed [14:0] m15_52;
   assign m15_52 =15'b0;

   // m15_53 = W*in
   wire signed [14:0] m15_53;
   assign m15_53 =15'b0;

   // m15_54 = W*in
   wire signed [14:0] m15_54;
   assign m15_54 =15'b0;

   // m15_55 = W*in
   wire signed [14:0] m15_55;
   assign m15_55 ={ {4{in15[14]}} , in15[14:4] };

   // m15_56 = W*in
   wire signed [14:0] m15_56;
   assign m15_56 =15'b0;

   // m15_57 = W*in
   wire signed [14:0] m15_57;
   assign m15_57 ={ {3{in15[14]}} , in15[14:3] };

   // m15_58 = W*in
   wire signed [14:0] m15_58;
   assign m15_58 =15'b0;

   // m15_59 = W*in
   wire signed [14:0] m15_59;
   assign m15_59 =15'b0;

   // m15_60 = W*in
   wire signed [14:0] m15_60;
   assign m15_60 =15'b0;

   // m15_61 = W*in
   wire signed [14:0] m15_61;
   assign m15_61 =15'b0;

   // m15_62 = W*in
   wire signed [14:0] m15_62;
   assign m15_62 =15'b0;

   // m15_63 = W*in
   wire signed [14:0] m15_63;
   assign m15_63 =15'b0;

   // m15_64 = W*in
   wire signed [14:0] m15_64;
   assign m15_64 =15'b0;

   // m15_65 = W*in
   wire signed [14:0] m15_65;
   assign m15_65 =15'b0;

   // m15_66 = W*in
   wire signed [14:0] m15_66;
   assign m15_66 =15'b0;

   // m15_67 = W*in
   wire signed [14:0] m15_67;
   assign m15_67 =15'b0;

   // m15_68 = W*in
   wire signed [14:0] m15_68;
   assign m15_68 =15'b0;

   // m15_69 = W*in
   wire signed [14:0] m15_69;
   assign m15_69 =15'b0;

   // m15_70 = W*in
   wire signed [14:0] m15_70;
   assign m15_70 =15'b0;

   // m15_71 = W*in
   wire signed [14:0] m15_71;
   assign m15_71 =15'b0;

   // m15_72 = W*in
   wire signed [14:0] m15_72;
   assign m15_72 ={ {3{neg15[14]}} , neg15[14:3] };

   // m15_73 = W*in
   wire signed [14:0] m15_73;
   assign m15_73 =15'b0;

   // m15_74 = W*in
   wire signed [14:0] m15_74;
   assign m15_74 =15'b0;

   // m15_75 = W*in
   wire signed [14:0] m15_75;
   assign m15_75 =15'b0;

   // m15_76 = W*in
   wire signed [14:0] m15_76;
   assign m15_76 ={ {3{neg15[14]}} , neg15[14:3] };

   // m15_77 = W*in
   wire signed [14:0] m15_77;
   assign m15_77 =15'b0;

   // m15_78 = W*in
   wire signed [14:0] m15_78;
   assign m15_78 =15'b0;

   // m15_79 = W*in
   wire signed [14:0] m15_79;
   assign m15_79 =15'b0;

   // m15_80 = W*in
   wire signed [14:0] m15_80;
   assign m15_80 =15'b0;

   // m15_81 = W*in
   wire signed [14:0] m15_81;
   assign m15_81 ={ {3{in15[14]}} , in15[14:3] };

   // m15_82 = W*in
   wire signed [14:0] m15_82;
   assign m15_82 =15'b0;

   // m15_83 = W*in
   wire signed [14:0] m15_83;
   assign m15_83 =15'b0;

   // m15_84 = W*in
   wire signed [14:0] m15_84;
   assign m15_84 =15'b0;

   // m15_85 = W*in
   wire signed [14:0] m15_85;
   assign m15_85 =15'b0;

   // m15_86 = W*in
   wire signed [14:0] m15_86;
   assign m15_86 ={ {3{in15[14]}} , in15[14:3] };

   // m15_87 = W*in
   wire signed [14:0] m15_87;
   assign m15_87 =15'b0;

   // m15_88 = W*in
   wire signed [14:0] m15_88;
   assign m15_88 =15'b0;

   // m15_89 = W*in
   wire signed [14:0] m15_89;
   assign m15_89 =15'b0;

   // m15_90 = W*in
   wire signed [14:0] m15_90;
   assign m15_90 =15'b0;

   // m15_91 = W*in
   wire signed [14:0] m15_91;
   assign m15_91 =15'b0;

   // m15_92 = W*in
   wire signed [14:0] m15_92;
   assign m15_92 =15'b0;

   // m15_93 = W*in
   wire signed [14:0] m15_93;
   assign m15_93 ={ {2{in15[14]}} , in15[14:2] };

   // m15_94 = W*in
   wire signed [14:0] m15_94;
   assign m15_94 ={ {3{neg15[14]}} , neg15[14:3] };

   // m15_95 = W*in
   wire signed [14:0] m15_95;
   assign m15_95 =15'b0;

   // m15_96 = W*in
   wire signed [14:0] m15_96;
   assign m15_96 =15'b0;

   // m15_97 = W*in
   wire signed [14:0] m15_97;
   assign m15_97 =15'b0;

   // m15_98 = W*in
   wire signed [14:0] m15_98;
   assign m15_98 =15'b0;

   // m15_99 = W*in
   wire signed [14:0] m15_99;
   assign m15_99 =15'b0;

   // m15_100 = W*in
   wire signed [14:0] m15_100;
   assign m15_100 =15'b0;

   // m16_1 = W*in
   wire signed [14:0] m16_1;
   assign m16_1 =15'b0;

   // m16_2 = W*in
   wire signed [14:0] m16_2;
   assign m16_2 =15'b0;

   // m16_3 = W*in
   wire signed [14:0] m16_3;
   assign m16_3 =15'b0;

   // m16_4 = W*in
   wire signed [14:0] m16_4;
   assign m16_4 ={ {3{in16[14]}} , in16[14:3] };

   // m16_5 = W*in
   wire signed [14:0] m16_5;
   assign m16_5 =15'b0;

   // m16_6 = W*in
   wire signed [14:0] m16_6;
   assign m16_6 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_7 = W*in
   wire signed [14:0] m16_7;
   assign m16_7 =15'b0;

   // m16_8 = W*in
   wire signed [14:0] m16_8;
   assign m16_8 =15'b0;

   // m16_9 = W*in
   wire signed [14:0] m16_9;
   assign m16_9 =15'b0;

   // m16_10 = W*in
   wire signed [14:0] m16_10;
   assign m16_10 =15'b0;

   // m16_11 = W*in
   wire signed [14:0] m16_11;
   assign m16_11 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_12 = W*in
   wire signed [14:0] m16_12;
   assign m16_12 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_13 = W*in
   wire signed [14:0] m16_13;
   assign m16_13 =15'b0;

   // m16_14 = W*in
   wire signed [14:0] m16_14;
   assign m16_14 ={ {3{in16[14]}} , in16[14:3] };

   // m16_15 = W*in
   wire signed [14:0] m16_15;
   assign m16_15 =15'b0;

   // m16_16 = W*in
   wire signed [14:0] m16_16;
   assign m16_16 =15'b0;

   // m16_17 = W*in
   wire signed [14:0] m16_17;
   assign m16_17 =15'b0;

   // m16_18 = W*in
   wire signed [14:0] m16_18;
   assign m16_18 =15'b0;

   // m16_19 = W*in
   wire signed [14:0] m16_19;
   assign m16_19 =15'b0;

   // m16_20 = W*in
   wire signed [14:0] m16_20;
   assign m16_20 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_21 = W*in
   wire signed [14:0] m16_21;
   assign m16_21 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_22 = W*in
   wire signed [14:0] m16_22;
   assign m16_22 ={ {3{in16[14]}} , in16[14:3] };

   // m16_23 = W*in
   wire signed [14:0] m16_23;
   assign m16_23 =15'b0;

   // m16_24 = W*in
   wire signed [14:0] m16_24;
   assign m16_24 =15'b0;

   // m16_25 = W*in
   wire signed [14:0] m16_25;
   assign m16_25 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_26 = W*in
   wire signed [14:0] m16_26;
   assign m16_26 ={ {3{in16[14]}} , in16[14:3] };

   // m16_27 = W*in
   wire signed [14:0] m16_27;
   assign m16_27 =15'b0;

   // m16_28 = W*in
   wire signed [14:0] m16_28;
   assign m16_28 =15'b0;

   // m16_29 = W*in
   wire signed [14:0] m16_29;
   assign m16_29 =15'b0;

   // m16_30 = W*in
   wire signed [14:0] m16_30;
   assign m16_30 =15'b0;

   // m16_31 = W*in
   wire signed [14:0] m16_31;
   assign m16_31 =15'b0;

   // m16_32 = W*in
   wire signed [14:0] m16_32;
   assign m16_32 =15'b0;

   // m16_33 = W*in
   wire signed [14:0] m16_33;
   assign m16_33 =15'b0;

   // m16_34 = W*in
   wire signed [14:0] m16_34;
   assign m16_34 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_35 = W*in
   wire signed [14:0] m16_35;
   assign m16_35 =15'b0;

   // m16_36 = W*in
   wire signed [14:0] m16_36;
   assign m16_36 =15'b0;

   // m16_37 = W*in
   wire signed [14:0] m16_37;
   assign m16_37 =15'b0;

   // m16_38 = W*in
   wire signed [14:0] m16_38;
   assign m16_38 =15'b0;

   // m16_39 = W*in
   wire signed [14:0] m16_39;
   assign m16_39 =15'b0;

   // m16_40 = W*in
   wire signed [14:0] m16_40;
   assign m16_40 =15'b0;

   // m16_41 = W*in
   wire signed [14:0] m16_41;
   assign m16_41 =15'b0;

   // m16_42 = W*in
   wire signed [14:0] m16_42;
   assign m16_42 =15'b0;

   // m16_43 = W*in
   wire signed [14:0] m16_43;
   assign m16_43 =15'b0;

   // m16_44 = W*in
   wire signed [14:0] m16_44;
   assign m16_44 =15'b0;

   // m16_45 = W*in
   wire signed [14:0] m16_45;
   assign m16_45 =15'b0;

   // m16_46 = W*in
   wire signed [14:0] m16_46;
   assign m16_46 =15'b0;

   // m16_47 = W*in
   wire signed [14:0] m16_47;
   assign m16_47 =15'b0;

   // m16_48 = W*in
   wire signed [14:0] m16_48;
   assign m16_48 =15'b0;

   // m16_49 = W*in
   wire signed [14:0] m16_49;
   assign m16_49 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_50 = W*in
   wire signed [14:0] m16_50;
   assign m16_50 =15'b0;

   // m16_51 = W*in
   wire signed [14:0] m16_51;
   assign m16_51 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_52 = W*in
   wire signed [14:0] m16_52;
   assign m16_52 =15'b0;

   // m16_53 = W*in
   wire signed [14:0] m16_53;
   assign m16_53 =15'b0;

   // m16_54 = W*in
   wire signed [14:0] m16_54;
   assign m16_54 =15'b0;

   // m16_55 = W*in
   wire signed [14:0] m16_55;
   assign m16_55 =15'b0;

   // m16_56 = W*in
   wire signed [14:0] m16_56;
   assign m16_56 =15'b0;

   // m16_57 = W*in
   wire signed [14:0] m16_57;
   assign m16_57 ={ {3{in16[14]}} , in16[14:3] };

   // m16_58 = W*in
   wire signed [14:0] m16_58;
   assign m16_58 =15'b0;

   // m16_59 = W*in
   wire signed [14:0] m16_59;
   assign m16_59 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_60 = W*in
   wire signed [14:0] m16_60;
   assign m16_60 =15'b0;

   // m16_61 = W*in
   wire signed [14:0] m16_61;
   assign m16_61 ={ {3{in16[14]}} , in16[14:3] };

   // m16_62 = W*in
   wire signed [14:0] m16_62;
   assign m16_62 ={ {4{in16[14]}} , in16[14:4] };

   // m16_63 = W*in
   wire signed [14:0] m16_63;
   assign m16_63 ={ {3{in16[14]}} , in16[14:3] };

   // m16_64 = W*in
   wire signed [14:0] m16_64;
   assign m16_64 ={ {4{in16[14]}} , in16[14:4] };

   // m16_65 = W*in
   wire signed [14:0] m16_65;
   assign m16_65 =15'b0;

   // m16_66 = W*in
   wire signed [14:0] m16_66;
   assign m16_66 =15'b0;

   // m16_67 = W*in
   wire signed [14:0] m16_67;
   assign m16_67 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_68 = W*in
   wire signed [14:0] m16_68;
   assign m16_68 =15'b0;

   // m16_69 = W*in
   wire signed [14:0] m16_69;
   assign m16_69 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_70 = W*in
   wire signed [14:0] m16_70;
   assign m16_70 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_71 = W*in
   wire signed [14:0] m16_71;
   assign m16_71 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_72 = W*in
   wire signed [14:0] m16_72;
   assign m16_72 =15'b0;

   // m16_73 = W*in
   wire signed [14:0] m16_73;
   assign m16_73 =15'b0;

   // m16_74 = W*in
   wire signed [14:0] m16_74;
   assign m16_74 =15'b0;

   // m16_75 = W*in
   wire signed [14:0] m16_75;
   assign m16_75 ={ {4{neg16[14]}} , neg16[14:4] };

   // m16_76 = W*in
   wire signed [14:0] m16_76;
   assign m16_76 =15'b0;

   // m16_77 = W*in
   wire signed [14:0] m16_77;
   assign m16_77 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_78 = W*in
   wire signed [14:0] m16_78;
   assign m16_78 =15'b0;

   // m16_79 = W*in
   wire signed [14:0] m16_79;
   assign m16_79 =15'b0;

   // m16_80 = W*in
   wire signed [14:0] m16_80;
   assign m16_80 =15'b0;

   // m16_81 = W*in
   wire signed [14:0] m16_81;
   assign m16_81 =15'b0;

   // m16_82 = W*in
   wire signed [14:0] m16_82;
   assign m16_82 =15'b0;

   // m16_83 = W*in
   wire signed [14:0] m16_83;
   assign m16_83 =15'b0;

   // m16_84 = W*in
   wire signed [14:0] m16_84;
   assign m16_84 =15'b0;

   // m16_85 = W*in
   wire signed [14:0] m16_85;
   assign m16_85 =15'b0;

   // m16_86 = W*in
   wire signed [14:0] m16_86;
   assign m16_86 =15'b0;

   // m16_87 = W*in
   wire signed [14:0] m16_87;
   assign m16_87 =15'b0;

   // m16_88 = W*in
   wire signed [14:0] m16_88;
   assign m16_88 =15'b0;

   // m16_89 = W*in
   wire signed [14:0] m16_89;
   assign m16_89 =15'b0;

   // m16_90 = W*in
   wire signed [14:0] m16_90;
   assign m16_90 =15'b0;

   // m16_91 = W*in
   wire signed [14:0] m16_91;
   assign m16_91 =15'b0;

   // m16_92 = W*in
   wire signed [14:0] m16_92;
   assign m16_92 =15'b0;

   // m16_93 = W*in
   wire signed [14:0] m16_93;
   assign m16_93 =15'b0;

   // m16_94 = W*in
   wire signed [14:0] m16_94;
   assign m16_94 =15'b0;

   // m16_95 = W*in
   wire signed [14:0] m16_95;
   assign m16_95 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_96 = W*in
   wire signed [14:0] m16_96;
   assign m16_96 ={ {3{neg16[14]}} , neg16[14:3] };

   // m16_97 = W*in
   wire signed [14:0] m16_97;
   assign m16_97 ={ {3{in16[14]}} , in16[14:3] };

   // m16_98 = W*in
   wire signed [14:0] m16_98;
   assign m16_98 =15'b0;

   // m16_99 = W*in
   wire signed [14:0] m16_99;
   assign m16_99 =15'b0;

   // m16_100 = W*in
   wire signed [14:0] m16_100;
   assign m16_100 =15'b0;

   // m17_1 = W*in
   wire signed [14:0] m17_1;
   assign m17_1 =15'b0;

   // m17_2 = W*in
   wire signed [14:0] m17_2;
   assign m17_2 =15'b0;

   // m17_3 = W*in
   wire signed [14:0] m17_3;
   assign m17_3 =15'b0;

   // m17_4 = W*in
   wire signed [14:0] m17_4;
   assign m17_4 =15'b0;

   // m17_5 = W*in
   wire signed [14:0] m17_5;
   assign m17_5 =15'b0;

   // m17_6 = W*in
   wire signed [14:0] m17_6;
   assign m17_6 =15'b0;

   // m17_7 = W*in
   wire signed [14:0] m17_7;
   assign m17_7 ={ {3{in17[14]}} , in17[14:3] };

   // m17_8 = W*in
   wire signed [14:0] m17_8;
   assign m17_8 =15'b0;

   // m17_9 = W*in
   wire signed [14:0] m17_9;
   assign m17_9 =15'b0;

   // m17_10 = W*in
   wire signed [14:0] m17_10;
   assign m17_10 ={ {3{in17[14]}} , in17[14:3] };

   // m17_11 = W*in
   wire signed [14:0] m17_11;
   assign m17_11 =15'b0;

   // m17_12 = W*in
   wire signed [14:0] m17_12;
   assign m17_12 =15'b0;

   // m17_13 = W*in
   wire signed [14:0] m17_13;
   assign m17_13 =15'b0;

   // m17_14 = W*in
   wire signed [14:0] m17_14;
   assign m17_14 =15'b0;

   // m17_15 = W*in
   wire signed [14:0] m17_15;
   assign m17_15 =15'b0;

   // m17_16 = W*in
   wire signed [14:0] m17_16;
   assign m17_16 =15'b0;

   // m17_17 = W*in
   wire signed [14:0] m17_17;
   assign m17_17 =15'b0;

   // m17_18 = W*in
   wire signed [14:0] m17_18;
   assign m17_18 =15'b0;

   // m17_19 = W*in
   wire signed [14:0] m17_19;
   assign m17_19 =15'b0;

   // m17_20 = W*in
   wire signed [14:0] m17_20;
   assign m17_20 =15'b0;

   // m17_21 = W*in
   wire signed [14:0] m17_21;
   assign m17_21 =15'b0;

   // m17_22 = W*in
   wire signed [14:0] m17_22;
   assign m17_22 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_23 = W*in
   wire signed [14:0] m17_23;
   assign m17_23 =15'b0;

   // m17_24 = W*in
   wire signed [14:0] m17_24;
   assign m17_24 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_25 = W*in
   wire signed [14:0] m17_25;
   assign m17_25 ={ {4{in17[14]}} , in17[14:4] };

   // m17_26 = W*in
   wire signed [14:0] m17_26;
   assign m17_26 =15'b0;

   // m17_27 = W*in
   wire signed [14:0] m17_27;
   assign m17_27 =15'b0;

   // m17_28 = W*in
   wire signed [14:0] m17_28;
   assign m17_28 ={ {4{neg17[14]}} , neg17[14:4] };

   // m17_29 = W*in
   wire signed [14:0] m17_29;
   assign m17_29 =15'b0;

   // m17_30 = W*in
   wire signed [14:0] m17_30;
   assign m17_30 =15'b0;

   // m17_31 = W*in
   wire signed [14:0] m17_31;
   assign m17_31 =15'b0;

   // m17_32 = W*in
   wire signed [14:0] m17_32;
   assign m17_32 =15'b0;

   // m17_33 = W*in
   wire signed [14:0] m17_33;
   assign m17_33 =15'b0;

   // m17_34 = W*in
   wire signed [14:0] m17_34;
   assign m17_34 =15'b0;

   // m17_35 = W*in
   wire signed [14:0] m17_35;
   assign m17_35 =15'b0;

   // m17_36 = W*in
   wire signed [14:0] m17_36;
   assign m17_36 =15'b0;

   // m17_37 = W*in
   wire signed [14:0] m17_37;
   assign m17_37 =15'b0;

   // m17_38 = W*in
   wire signed [14:0] m17_38;
   assign m17_38 =15'b0;

   // m17_39 = W*in
   wire signed [14:0] m17_39;
   assign m17_39 =15'b0;

   // m17_40 = W*in
   wire signed [14:0] m17_40;
   assign m17_40 =15'b0;

   // m17_41 = W*in
   wire signed [14:0] m17_41;
   assign m17_41 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_42 = W*in
   wire signed [14:0] m17_42;
   assign m17_42 =15'b0;

   // m17_43 = W*in
   wire signed [14:0] m17_43;
   assign m17_43 =15'b0;

   // m17_44 = W*in
   wire signed [14:0] m17_44;
   assign m17_44 ={ {3{in17[14]}} , in17[14:3] };

   // m17_45 = W*in
   wire signed [14:0] m17_45;
   assign m17_45 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_46 = W*in
   wire signed [14:0] m17_46;
   assign m17_46 =15'b0;

   // m17_47 = W*in
   wire signed [14:0] m17_47;
   assign m17_47 =15'b0;

   // m17_48 = W*in
   wire signed [14:0] m17_48;
   assign m17_48 =15'b0;

   // m17_49 = W*in
   wire signed [14:0] m17_49;
   assign m17_49 =15'b0;

   // m17_50 = W*in
   wire signed [14:0] m17_50;
   assign m17_50 =15'b0;

   // m17_51 = W*in
   wire signed [14:0] m17_51;
   assign m17_51 =15'b0;

   // m17_52 = W*in
   wire signed [14:0] m17_52;
   assign m17_52 =15'b0;

   // m17_53 = W*in
   wire signed [14:0] m17_53;
   assign m17_53 =15'b0;

   // m17_54 = W*in
   wire signed [14:0] m17_54;
   assign m17_54 =15'b0;

   // m17_55 = W*in
   wire signed [14:0] m17_55;
   assign m17_55 =15'b0;

   // m17_56 = W*in
   wire signed [14:0] m17_56;
   assign m17_56 =15'b0;

   // m17_57 = W*in
   wire signed [14:0] m17_57;
   assign m17_57 =15'b0;

   // m17_58 = W*in
   wire signed [14:0] m17_58;
   assign m17_58 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_59 = W*in
   wire signed [14:0] m17_59;
   assign m17_59 =15'b0;

   // m17_60 = W*in
   wire signed [14:0] m17_60;
   assign m17_60 =15'b0;

   // m17_61 = W*in
   wire signed [14:0] m17_61;
   assign m17_61 ={ {4{neg17[14]}} , neg17[14:4] };

   // m17_62 = W*in
   wire signed [14:0] m17_62;
   assign m17_62 ={ {2{neg17[14]}} , neg17[14:2] };

   // m17_63 = W*in
   wire signed [14:0] m17_63;
   assign m17_63 =15'b0;

   // m17_64 = W*in
   wire signed [14:0] m17_64;
   assign m17_64 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_65 = W*in
   wire signed [14:0] m17_65;
   assign m17_65 =15'b0;

   // m17_66 = W*in
   wire signed [14:0] m17_66;
   assign m17_66 ={ {3{in17[14]}} , in17[14:3] };

   // m17_67 = W*in
   wire signed [14:0] m17_67;
   assign m17_67 ={ {4{neg17[14]}} , neg17[14:4] };

   // m17_68 = W*in
   wire signed [14:0] m17_68;
   assign m17_68 ={ {4{neg17[14]}} , neg17[14:4] };

   // m17_69 = W*in
   wire signed [14:0] m17_69;
   assign m17_69 =15'b0;

   // m17_70 = W*in
   wire signed [14:0] m17_70;
   assign m17_70 ={ {4{in17[14]}} , in17[14:4] };

   // m17_71 = W*in
   wire signed [14:0] m17_71;
   assign m17_71 =15'b0;

   // m17_72 = W*in
   wire signed [14:0] m17_72;
   assign m17_72 =15'b0;

   // m17_73 = W*in
   wire signed [14:0] m17_73;
   assign m17_73 =15'b0;

   // m17_74 = W*in
   wire signed [14:0] m17_74;
   assign m17_74 =15'b0;

   // m17_75 = W*in
   wire signed [14:0] m17_75;
   assign m17_75 ={ {3{neg17[14]}} , neg17[14:3] };

   // m17_76 = W*in
   wire signed [14:0] m17_76;
   assign m17_76 =15'b0;

   // m17_77 = W*in
   wire signed [14:0] m17_77;
   assign m17_77 =15'b0;

   // m17_78 = W*in
   wire signed [14:0] m17_78;
   assign m17_78 =15'b0;

   // m17_79 = W*in
   wire signed [14:0] m17_79;
   assign m17_79 ={ {4{in17[14]}} , in17[14:4] };

   // m17_80 = W*in
   wire signed [14:0] m17_80;
   assign m17_80 =15'b0;

   // m17_81 = W*in
   wire signed [14:0] m17_81;
   assign m17_81 ={ {2{neg17[14]}} , neg17[14:2] };

   // m17_82 = W*in
   wire signed [14:0] m17_82;
   assign m17_82 =15'b0;

   // m17_83 = W*in
   wire signed [14:0] m17_83;
   assign m17_83 =15'b0;

   // m17_84 = W*in
   wire signed [14:0] m17_84;
   assign m17_84 =15'b0;

   // m17_85 = W*in
   wire signed [14:0] m17_85;
   assign m17_85 ={ {2{neg17[14]}} , neg17[14:2] };

   // m17_86 = W*in
   wire signed [14:0] m17_86;
   assign m17_86 =15'b0;

   // m17_87 = W*in
   wire signed [14:0] m17_87;
   assign m17_87 ={ {2{neg17[14]}} , neg17[14:2] };

   // m17_88 = W*in
   wire signed [14:0] m17_88;
   assign m17_88 =15'b0;

   // m17_89 = W*in
   wire signed [14:0] m17_89;
   assign m17_89 =15'b0;

   // m17_90 = W*in
   wire signed [14:0] m17_90;
   assign m17_90 =15'b0;

   // m17_91 = W*in
   wire signed [14:0] m17_91;
   assign m17_91 =15'b0;

   // m17_92 = W*in
   wire signed [14:0] m17_92;
   assign m17_92 =15'b0;

   // m17_93 = W*in
   wire signed [14:0] m17_93;
   assign m17_93 =15'b0;

   // m17_94 = W*in
   wire signed [14:0] m17_94;
   assign m17_94 =15'b0;

   // m17_95 = W*in
   wire signed [14:0] m17_95;
   assign m17_95 =15'b0;

   // m17_96 = W*in
   wire signed [14:0] m17_96;
   assign m17_96 =15'b0;

   // m17_97 = W*in
   wire signed [14:0] m17_97;
   assign m17_97 =15'b0;

   // m17_98 = W*in
   wire signed [14:0] m17_98;
   assign m17_98 =15'b0;

   // m17_99 = W*in
   wire signed [14:0] m17_99;
   assign m17_99 =15'b0;

   // m17_100 = W*in
   wire signed [14:0] m17_100;
   assign m17_100 =15'b0;

   // m18_1 = W*in
   wire signed [14:0] m18_1;
   assign m18_1 =15'b0;

   // m18_2 = W*in
   wire signed [14:0] m18_2;
   assign m18_2 =15'b0;

   // m18_3 = W*in
   wire signed [14:0] m18_3;
   assign m18_3 =15'b0;

   // m18_4 = W*in
   wire signed [14:0] m18_4;
   assign m18_4 =15'b0;

   // m18_5 = W*in
   wire signed [14:0] m18_5;
   assign m18_5 ={ {3{in18[14]}} , in18[14:3] };

   // m18_6 = W*in
   wire signed [14:0] m18_6;
   assign m18_6 =15'b0;

   // m18_7 = W*in
   wire signed [14:0] m18_7;
   assign m18_7 =15'b0;

   // m18_8 = W*in
   wire signed [14:0] m18_8;
   assign m18_8 ={ {4{in18[14]}} , in18[14:4] };

   // m18_9 = W*in
   wire signed [14:0] m18_9;
   assign m18_9 =15'b0;

   // m18_10 = W*in
   wire signed [14:0] m18_10;
   assign m18_10 =15'b0;

   // m18_11 = W*in
   wire signed [14:0] m18_11;
   assign m18_11 ={ {2{neg18[14]}} , neg18[14:2] };

   // m18_12 = W*in
   wire signed [14:0] m18_12;
   assign m18_12 =15'b0;

   // m18_13 = W*in
   wire signed [14:0] m18_13;
   assign m18_13 =15'b0;

   // m18_14 = W*in
   wire signed [14:0] m18_14;
   assign m18_14 =15'b0;

   // m18_15 = W*in
   wire signed [14:0] m18_15;
   assign m18_15 =15'b0;

   // m18_16 = W*in
   wire signed [14:0] m18_16;
   assign m18_16 =15'b0;

   // m18_17 = W*in
   wire signed [14:0] m18_17;
   assign m18_17 =15'b0;

   // m18_18 = W*in
   wire signed [14:0] m18_18;
   assign m18_18 =15'b0;

   // m18_19 = W*in
   wire signed [14:0] m18_19;
   assign m18_19 =15'b0;

   // m18_20 = W*in
   wire signed [14:0] m18_20;
   assign m18_20 =15'b0;

   // m18_21 = W*in
   wire signed [14:0] m18_21;
   assign m18_21 =15'b0;

   // m18_22 = W*in
   wire signed [14:0] m18_22;
   assign m18_22 =15'b0;

   // m18_23 = W*in
   wire signed [14:0] m18_23;
   assign m18_23 =15'b0;

   // m18_24 = W*in
   wire signed [14:0] m18_24;
   assign m18_24 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_25 = W*in
   wire signed [14:0] m18_25;
   assign m18_25 =15'b0;

   // m18_26 = W*in
   wire signed [14:0] m18_26;
   assign m18_26 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_27 = W*in
   wire signed [14:0] m18_27;
   assign m18_27 =15'b0;

   // m18_28 = W*in
   wire signed [14:0] m18_28;
   assign m18_28 =15'b0;

   // m18_29 = W*in
   wire signed [14:0] m18_29;
   assign m18_29 =15'b0;

   // m18_30 = W*in
   wire signed [14:0] m18_30;
   assign m18_30 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_31 = W*in
   wire signed [14:0] m18_31;
   assign m18_31 ={ {4{in18[14]}} , in18[14:4] };

   // m18_32 = W*in
   wire signed [14:0] m18_32;
   assign m18_32 =15'b0;

   // m18_33 = W*in
   wire signed [14:0] m18_33;
   assign m18_33 =15'b0;

   // m18_34 = W*in
   wire signed [14:0] m18_34;
   assign m18_34 =15'b0;

   // m18_35 = W*in
   wire signed [14:0] m18_35;
   assign m18_35 =15'b0;

   // m18_36 = W*in
   wire signed [14:0] m18_36;
   assign m18_36 =15'b0;

   // m18_37 = W*in
   wire signed [14:0] m18_37;
   assign m18_37 =15'b0;

   // m18_38 = W*in
   wire signed [14:0] m18_38;
   assign m18_38 ={ {3{in18[14]}} , in18[14:3] };

   // m18_39 = W*in
   wire signed [14:0] m18_39;
   assign m18_39 =15'b0;

   // m18_40 = W*in
   wire signed [14:0] m18_40;
   assign m18_40 =15'b0;

   // m18_41 = W*in
   wire signed [14:0] m18_41;
   assign m18_41 =15'b0;

   // m18_42 = W*in
   wire signed [14:0] m18_42;
   assign m18_42 =15'b0;

   // m18_43 = W*in
   wire signed [14:0] m18_43;
   assign m18_43 =15'b0;

   // m18_44 = W*in
   wire signed [14:0] m18_44;
   assign m18_44 =15'b0;

   // m18_45 = W*in
   wire signed [14:0] m18_45;
   assign m18_45 =15'b0;

   // m18_46 = W*in
   wire signed [14:0] m18_46;
   assign m18_46 =15'b0;

   // m18_47 = W*in
   wire signed [14:0] m18_47;
   assign m18_47 =15'b0;

   // m18_48 = W*in
   wire signed [14:0] m18_48;
   assign m18_48 =15'b0;

   // m18_49 = W*in
   wire signed [14:0] m18_49;
   assign m18_49 =15'b0;

   // m18_50 = W*in
   wire signed [14:0] m18_50;
   assign m18_50 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_51 = W*in
   wire signed [14:0] m18_51;
   assign m18_51 =15'b0;

   // m18_52 = W*in
   wire signed [14:0] m18_52;
   assign m18_52 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_53 = W*in
   wire signed [14:0] m18_53;
   assign m18_53 =15'b0;

   // m18_54 = W*in
   wire signed [14:0] m18_54;
   assign m18_54 =15'b0;

   // m18_55 = W*in
   wire signed [14:0] m18_55;
   assign m18_55 =15'b0;

   // m18_56 = W*in
   wire signed [14:0] m18_56;
   assign m18_56 =15'b0;

   // m18_57 = W*in
   wire signed [14:0] m18_57;
   assign m18_57 ={ {3{in18[14]}} , in18[14:3] };

   // m18_58 = W*in
   wire signed [14:0] m18_58;
   assign m18_58 =15'b0;

   // m18_59 = W*in
   wire signed [14:0] m18_59;
   assign m18_59 =15'b0;

   // m18_60 = W*in
   wire signed [14:0] m18_60;
   assign m18_60 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_61 = W*in
   wire signed [14:0] m18_61;
   assign m18_61 =15'b0;

   // m18_62 = W*in
   wire signed [14:0] m18_62;
   assign m18_62 =15'b0;

   // m18_63 = W*in
   wire signed [14:0] m18_63;
   assign m18_63 =15'b0;

   // m18_64 = W*in
   wire signed [14:0] m18_64;
   assign m18_64 =15'b0;

   // m18_65 = W*in
   wire signed [14:0] m18_65;
   assign m18_65 =15'b0;

   // m18_66 = W*in
   wire signed [14:0] m18_66;
   assign m18_66 =15'b0;

   // m18_67 = W*in
   wire signed [14:0] m18_67;
   assign m18_67 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_68 = W*in
   wire signed [14:0] m18_68;
   assign m18_68 =15'b0;

   // m18_69 = W*in
   wire signed [14:0] m18_69;
   assign m18_69 =15'b0;

   // m18_70 = W*in
   wire signed [14:0] m18_70;
   assign m18_70 =15'b0;

   // m18_71 = W*in
   wire signed [14:0] m18_71;
   assign m18_71 =15'b0;

   // m18_72 = W*in
   wire signed [14:0] m18_72;
   assign m18_72 =15'b0;

   // m18_73 = W*in
   wire signed [14:0] m18_73;
   assign m18_73 ={ {4{neg18[14]}} , neg18[14:4] };

   // m18_74 = W*in
   wire signed [14:0] m18_74;
   assign m18_74 ={ {3{in18[14]}} , in18[14:3] };

   // m18_75 = W*in
   wire signed [14:0] m18_75;
   assign m18_75 =15'b0;

   // m18_76 = W*in
   wire signed [14:0] m18_76;
   assign m18_76 =15'b0;

   // m18_77 = W*in
   wire signed [14:0] m18_77;
   assign m18_77 =15'b0;

   // m18_78 = W*in
   wire signed [14:0] m18_78;
   assign m18_78 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_79 = W*in
   wire signed [14:0] m18_79;
   assign m18_79 =15'b0;

   // m18_80 = W*in
   wire signed [14:0] m18_80;
   assign m18_80 =15'b0;

   // m18_81 = W*in
   wire signed [14:0] m18_81;
   assign m18_81 =15'b0;

   // m18_82 = W*in
   wire signed [14:0] m18_82;
   assign m18_82 ={ {3{in18[14]}} , in18[14:3] };

   // m18_83 = W*in
   wire signed [14:0] m18_83;
   assign m18_83 ={ {2{in18[14]}} , in18[14:2] };

   // m18_84 = W*in
   wire signed [14:0] m18_84;
   assign m18_84 =15'b0;

   // m18_85 = W*in
   wire signed [14:0] m18_85;
   assign m18_85 =15'b0;

   // m18_86 = W*in
   wire signed [14:0] m18_86;
   assign m18_86 =15'b0;

   // m18_87 = W*in
   wire signed [14:0] m18_87;
   assign m18_87 =15'b0;

   // m18_88 = W*in
   wire signed [14:0] m18_88;
   assign m18_88 =15'b0;

   // m18_89 = W*in
   wire signed [14:0] m18_89;
   assign m18_89 ={ {3{in18[14]}} , in18[14:3] };

   // m18_90 = W*in
   wire signed [14:0] m18_90;
   assign m18_90 =15'b0;

   // m18_91 = W*in
   wire signed [14:0] m18_91;
   assign m18_91 =15'b0;

   // m18_92 = W*in
   wire signed [14:0] m18_92;
   assign m18_92 =15'b0;

   // m18_93 = W*in
   wire signed [14:0] m18_93;
   assign m18_93 =15'b0;

   // m18_94 = W*in
   wire signed [14:0] m18_94;
   assign m18_94 =15'b0;

   // m18_95 = W*in
   wire signed [14:0] m18_95;
   assign m18_95 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_96 = W*in
   wire signed [14:0] m18_96;
   assign m18_96 ={ {3{neg18[14]}} , neg18[14:3] };

   // m18_97 = W*in
   wire signed [14:0] m18_97;
   assign m18_97 =15'b0;

   // m18_98 = W*in
   wire signed [14:0] m18_98;
   assign m18_98 =15'b0;

   // m18_99 = W*in
   wire signed [14:0] m18_99;
   assign m18_99 =15'b0;

   // m18_100 = W*in
   wire signed [14:0] m18_100;
   assign m18_100 =15'b0;

   // m19_1 = W*in
   wire signed [14:0] m19_1;
   assign m19_1 =15'b0;

   // m19_2 = W*in
   wire signed [14:0] m19_2;
   assign m19_2 =15'b0;

   // m19_3 = W*in
   wire signed [14:0] m19_3;
   assign m19_3 =15'b0;

   // m19_4 = W*in
   wire signed [14:0] m19_4;
   assign m19_4 =15'b0;

   // m19_5 = W*in
   wire signed [14:0] m19_5;
   assign m19_5 =15'b0;

   // m19_6 = W*in
   wire signed [14:0] m19_6;
   assign m19_6 =15'b0;

   // m19_7 = W*in
   wire signed [14:0] m19_7;
   assign m19_7 =15'b0;

   // m19_8 = W*in
   wire signed [14:0] m19_8;
   assign m19_8 =15'b0;

   // m19_9 = W*in
   wire signed [14:0] m19_9;
   assign m19_9 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_10 = W*in
   wire signed [14:0] m19_10;
   assign m19_10 =15'b0;

   // m19_11 = W*in
   wire signed [14:0] m19_11;
   assign m19_11 =15'b0;

   // m19_12 = W*in
   wire signed [14:0] m19_12;
   assign m19_12 =15'b0;

   // m19_13 = W*in
   wire signed [14:0] m19_13;
   assign m19_13 ={ {3{in19[14]}} , in19[14:3] };

   // m19_14 = W*in
   wire signed [14:0] m19_14;
   assign m19_14 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_15 = W*in
   wire signed [14:0] m19_15;
   assign m19_15 =15'b0;

   // m19_16 = W*in
   wire signed [14:0] m19_16;
   assign m19_16 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_17 = W*in
   wire signed [14:0] m19_17;
   assign m19_17 =15'b0;

   // m19_18 = W*in
   wire signed [14:0] m19_18;
   assign m19_18 =15'b0;

   // m19_19 = W*in
   wire signed [14:0] m19_19;
   assign m19_19 =15'b0;

   // m19_20 = W*in
   wire signed [14:0] m19_20;
   assign m19_20 ={ {3{in19[14]}} , in19[14:3] };

   // m19_21 = W*in
   wire signed [14:0] m19_21;
   assign m19_21 =15'b0;

   // m19_22 = W*in
   wire signed [14:0] m19_22;
   assign m19_22 =15'b0;

   // m19_23 = W*in
   wire signed [14:0] m19_23;
   assign m19_23 =15'b0;

   // m19_24 = W*in
   wire signed [14:0] m19_24;
   assign m19_24 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_25 = W*in
   wire signed [14:0] m19_25;
   assign m19_25 =15'b0;

   // m19_26 = W*in
   wire signed [14:0] m19_26;
   assign m19_26 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_27 = W*in
   wire signed [14:0] m19_27;
   assign m19_27 =15'b0;

   // m19_28 = W*in
   wire signed [14:0] m19_28;
   assign m19_28 =15'b0;

   // m19_29 = W*in
   wire signed [14:0] m19_29;
   assign m19_29 ={ {4{neg19[14]}} , neg19[14:4] };

   // m19_30 = W*in
   wire signed [14:0] m19_30;
   assign m19_30 =15'b0;

   // m19_31 = W*in
   wire signed [14:0] m19_31;
   assign m19_31 =15'b0;

   // m19_32 = W*in
   wire signed [14:0] m19_32;
   assign m19_32 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_33 = W*in
   wire signed [14:0] m19_33;
   assign m19_33 =15'b0;

   // m19_34 = W*in
   wire signed [14:0] m19_34;
   assign m19_34 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_35 = W*in
   wire signed [14:0] m19_35;
   assign m19_35 =15'b0;

   // m19_36 = W*in
   wire signed [14:0] m19_36;
   assign m19_36 =15'b0;

   // m19_37 = W*in
   wire signed [14:0] m19_37;
   assign m19_37 =15'b0;

   // m19_38 = W*in
   wire signed [14:0] m19_38;
   assign m19_38 =15'b0;

   // m19_39 = W*in
   wire signed [14:0] m19_39;
   assign m19_39 =15'b0;

   // m19_40 = W*in
   wire signed [14:0] m19_40;
   assign m19_40 =15'b0;

   // m19_41 = W*in
   wire signed [14:0] m19_41;
   assign m19_41 =15'b0;

   // m19_42 = W*in
   wire signed [14:0] m19_42;
   assign m19_42 =15'b0;

   // m19_43 = W*in
   wire signed [14:0] m19_43;
   assign m19_43 =15'b0;

   // m19_44 = W*in
   wire signed [14:0] m19_44;
   assign m19_44 =15'b0;

   // m19_45 = W*in
   wire signed [14:0] m19_45;
   assign m19_45 =15'b0;

   // m19_46 = W*in
   wire signed [14:0] m19_46;
   assign m19_46 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_47 = W*in
   wire signed [14:0] m19_47;
   assign m19_47 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_48 = W*in
   wire signed [14:0] m19_48;
   assign m19_48 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_49 = W*in
   wire signed [14:0] m19_49;
   assign m19_49 =15'b0;

   // m19_50 = W*in
   wire signed [14:0] m19_50;
   assign m19_50 =15'b0;

   // m19_51 = W*in
   wire signed [14:0] m19_51;
   assign m19_51 =15'b0;

   // m19_52 = W*in
   wire signed [14:0] m19_52;
   assign m19_52 =15'b0;

   // m19_53 = W*in
   wire signed [14:0] m19_53;
   assign m19_53 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_54 = W*in
   wire signed [14:0] m19_54;
   assign m19_54 =15'b0;

   // m19_55 = W*in
   wire signed [14:0] m19_55;
   assign m19_55 =15'b0;

   // m19_56 = W*in
   wire signed [14:0] m19_56;
   assign m19_56 =15'b0;

   // m19_57 = W*in
   wire signed [14:0] m19_57;
   assign m19_57 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_58 = W*in
   wire signed [14:0] m19_58;
   assign m19_58 =15'b0;

   // m19_59 = W*in
   wire signed [14:0] m19_59;
   assign m19_59 ={ {4{neg19[14]}} , neg19[14:4] };

   // m19_60 = W*in
   wire signed [14:0] m19_60;
   assign m19_60 =15'b0;

   // m19_61 = W*in
   wire signed [14:0] m19_61;
   assign m19_61 =15'b0;

   // m19_62 = W*in
   wire signed [14:0] m19_62;
   assign m19_62 ={ {3{in19[14]}} , in19[14:3] };

   // m19_63 = W*in
   wire signed [14:0] m19_63;
   assign m19_63 =15'b0;

   // m19_64 = W*in
   wire signed [14:0] m19_64;
   assign m19_64 =15'b0;

   // m19_65 = W*in
   wire signed [14:0] m19_65;
   assign m19_65 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_66 = W*in
   wire signed [14:0] m19_66;
   assign m19_66 =15'b0;

   // m19_67 = W*in
   wire signed [14:0] m19_67;
   assign m19_67 =15'b0;

   // m19_68 = W*in
   wire signed [14:0] m19_68;
   assign m19_68 =15'b0;

   // m19_69 = W*in
   wire signed [14:0] m19_69;
   assign m19_69 =15'b0;

   // m19_70 = W*in
   wire signed [14:0] m19_70;
   assign m19_70 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_71 = W*in
   wire signed [14:0] m19_71;
   assign m19_71 =15'b0;

   // m19_72 = W*in
   wire signed [14:0] m19_72;
   assign m19_72 ={ {3{in19[14]}} , in19[14:3] };

   // m19_73 = W*in
   wire signed [14:0] m19_73;
   assign m19_73 =15'b0;

   // m19_74 = W*in
   wire signed [14:0] m19_74;
   assign m19_74 ={ {4{neg19[14]}} , neg19[14:4] };

   // m19_75 = W*in
   wire signed [14:0] m19_75;
   assign m19_75 =15'b0;

   // m19_76 = W*in
   wire signed [14:0] m19_76;
   assign m19_76 =15'b0;

   // m19_77 = W*in
   wire signed [14:0] m19_77;
   assign m19_77 =15'b0;

   // m19_78 = W*in
   wire signed [14:0] m19_78;
   assign m19_78 ={ {4{in19[14]}} , in19[14:4] };

   // m19_79 = W*in
   wire signed [14:0] m19_79;
   assign m19_79 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_80 = W*in
   wire signed [14:0] m19_80;
   assign m19_80 ={ {3{in19[14]}} , in19[14:3] };

   // m19_81 = W*in
   wire signed [14:0] m19_81;
   assign m19_81 =15'b0;

   // m19_82 = W*in
   wire signed [14:0] m19_82;
   assign m19_82 =15'b0;

   // m19_83 = W*in
   wire signed [14:0] m19_83;
   assign m19_83 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_84 = W*in
   wire signed [14:0] m19_84;
   assign m19_84 =15'b0;

   // m19_85 = W*in
   wire signed [14:0] m19_85;
   assign m19_85 =15'b0;

   // m19_86 = W*in
   wire signed [14:0] m19_86;
   assign m19_86 =15'b0;

   // m19_87 = W*in
   wire signed [14:0] m19_87;
   assign m19_87 =15'b0;

   // m19_88 = W*in
   wire signed [14:0] m19_88;
   assign m19_88 =15'b0;

   // m19_89 = W*in
   wire signed [14:0] m19_89;
   assign m19_89 =15'b0;

   // m19_90 = W*in
   wire signed [14:0] m19_90;
   assign m19_90 =15'b0;

   // m19_91 = W*in
   wire signed [14:0] m19_91;
   assign m19_91 =15'b0;

   // m19_92 = W*in
   wire signed [14:0] m19_92;
   assign m19_92 ={ {4{neg19[14]}} , neg19[14:4] };

   // m19_93 = W*in
   wire signed [14:0] m19_93;
   assign m19_93 =15'b0;

   // m19_94 = W*in
   wire signed [14:0] m19_94;
   assign m19_94 ={ {3{neg19[14]}} , neg19[14:3] };

   // m19_95 = W*in
   wire signed [14:0] m19_95;
   assign m19_95 =15'b0;

   // m19_96 = W*in
   wire signed [14:0] m19_96;
   assign m19_96 =15'b0;

   // m19_97 = W*in
   wire signed [14:0] m19_97;
   assign m19_97 =15'b0;

   // m19_98 = W*in
   wire signed [14:0] m19_98;
   assign m19_98 =15'b0;

   // m19_99 = W*in
   wire signed [14:0] m19_99;
   assign m19_99 =15'b0;

   // m19_100 = W*in
   wire signed [14:0] m19_100;
   assign m19_100 ={ {3{neg19[14]}} , neg19[14:3] };

   // m20_1 = W*in
   wire signed [14:0] m20_1;
   assign m20_1 =15'b0;

   // m20_2 = W*in
   wire signed [14:0] m20_2;
   assign m20_2 =15'b0;

   // m20_3 = W*in
   wire signed [14:0] m20_3;
   assign m20_3 =15'b0;

   // m20_4 = W*in
   wire signed [14:0] m20_4;
   assign m20_4 =15'b0;

   // m20_5 = W*in
   wire signed [14:0] m20_5;
   assign m20_5 =15'b0;

   // m20_6 = W*in
   wire signed [14:0] m20_6;
   assign m20_6 ={ {3{in20[14]}} , in20[14:3] };

   // m20_7 = W*in
   wire signed [14:0] m20_7;
   assign m20_7 =15'b0;

   // m20_8 = W*in
   wire signed [14:0] m20_8;
   assign m20_8 =15'b0;

   // m20_9 = W*in
   wire signed [14:0] m20_9;
   assign m20_9 =15'b0;

   // m20_10 = W*in
   wire signed [14:0] m20_10;
   assign m20_10 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_11 = W*in
   wire signed [14:0] m20_11;
   assign m20_11 =15'b0;

   // m20_12 = W*in
   wire signed [14:0] m20_12;
   assign m20_12 =15'b0;

   // m20_13 = W*in
   wire signed [14:0] m20_13;
   assign m20_13 =15'b0;

   // m20_14 = W*in
   wire signed [14:0] m20_14;
   assign m20_14 =15'b0;

   // m20_15 = W*in
   wire signed [14:0] m20_15;
   assign m20_15 =15'b0;

   // m20_16 = W*in
   wire signed [14:0] m20_16;
   assign m20_16 =15'b0;

   // m20_17 = W*in
   wire signed [14:0] m20_17;
   assign m20_17 =15'b0;

   // m20_18 = W*in
   wire signed [14:0] m20_18;
   assign m20_18 =15'b0;

   // m20_19 = W*in
   wire signed [14:0] m20_19;
   assign m20_19 ={ {4{neg20[14]}} , neg20[14:4] };

   // m20_20 = W*in
   wire signed [14:0] m20_20;
   assign m20_20 =15'b0;

   // m20_21 = W*in
   wire signed [14:0] m20_21;
   assign m20_21 =15'b0;

   // m20_22 = W*in
   wire signed [14:0] m20_22;
   assign m20_22 =15'b0;

   // m20_23 = W*in
   wire signed [14:0] m20_23;
   assign m20_23 =15'b0;

   // m20_24 = W*in
   wire signed [14:0] m20_24;
   assign m20_24 =15'b0;

   // m20_25 = W*in
   wire signed [14:0] m20_25;
   assign m20_25 =15'b0;

   // m20_26 = W*in
   wire signed [14:0] m20_26;
   assign m20_26 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_27 = W*in
   wire signed [14:0] m20_27;
   assign m20_27 ={ {4{neg20[14]}} , neg20[14:4] };

   // m20_28 = W*in
   wire signed [14:0] m20_28;
   assign m20_28 =15'b0;

   // m20_29 = W*in
   wire signed [14:0] m20_29;
   assign m20_29 =15'b0;

   // m20_30 = W*in
   wire signed [14:0] m20_30;
   assign m20_30 ={ {4{neg20[14]}} , neg20[14:4] };

   // m20_31 = W*in
   wire signed [14:0] m20_31;
   assign m20_31 =15'b0;

   // m20_32 = W*in
   wire signed [14:0] m20_32;
   assign m20_32 =15'b0;

   // m20_33 = W*in
   wire signed [14:0] m20_33;
   assign m20_33 =15'b0;

   // m20_34 = W*in
   wire signed [14:0] m20_34;
   assign m20_34 =15'b0;

   // m20_35 = W*in
   wire signed [14:0] m20_35;
   assign m20_35 =15'b0;

   // m20_36 = W*in
   wire signed [14:0] m20_36;
   assign m20_36 =15'b0;

   // m20_37 = W*in
   wire signed [14:0] m20_37;
   assign m20_37 =15'b0;

   // m20_38 = W*in
   wire signed [14:0] m20_38;
   assign m20_38 =15'b0;

   // m20_39 = W*in
   wire signed [14:0] m20_39;
   assign m20_39 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_40 = W*in
   wire signed [14:0] m20_40;
   assign m20_40 =15'b0;

   // m20_41 = W*in
   wire signed [14:0] m20_41;
   assign m20_41 ={ {3{in20[14]}} , in20[14:3] };

   // m20_42 = W*in
   wire signed [14:0] m20_42;
   assign m20_42 =15'b0;

   // m20_43 = W*in
   wire signed [14:0] m20_43;
   assign m20_43 =15'b0;

   // m20_44 = W*in
   wire signed [14:0] m20_44;
   assign m20_44 =15'b0;

   // m20_45 = W*in
   wire signed [14:0] m20_45;
   assign m20_45 =15'b0;

   // m20_46 = W*in
   wire signed [14:0] m20_46;
   assign m20_46 =15'b0;

   // m20_47 = W*in
   wire signed [14:0] m20_47;
   assign m20_47 =15'b0;

   // m20_48 = W*in
   wire signed [14:0] m20_48;
   assign m20_48 =15'b0;

   // m20_49 = W*in
   wire signed [14:0] m20_49;
   assign m20_49 =15'b0;

   // m20_50 = W*in
   wire signed [14:0] m20_50;
   assign m20_50 =15'b0;

   // m20_51 = W*in
   wire signed [14:0] m20_51;
   assign m20_51 =15'b0;

   // m20_52 = W*in
   wire signed [14:0] m20_52;
   assign m20_52 ={ {3{in20[14]}} , in20[14:3] };

   // m20_53 = W*in
   wire signed [14:0] m20_53;
   assign m20_53 =15'b0;

   // m20_54 = W*in
   wire signed [14:0] m20_54;
   assign m20_54 =15'b0;

   // m20_55 = W*in
   wire signed [14:0] m20_55;
   assign m20_55 =15'b0;

   // m20_56 = W*in
   wire signed [14:0] m20_56;
   assign m20_56 =15'b0;

   // m20_57 = W*in
   wire signed [14:0] m20_57;
   assign m20_57 =15'b0;

   // m20_58 = W*in
   wire signed [14:0] m20_58;
   assign m20_58 ={ {3{in20[14]}} , in20[14:3] };

   // m20_59 = W*in
   wire signed [14:0] m20_59;
   assign m20_59 =15'b0;

   // m20_60 = W*in
   wire signed [14:0] m20_60;
   assign m20_60 ={ {3{in20[14]}} , in20[14:3] };

   // m20_61 = W*in
   wire signed [14:0] m20_61;
   assign m20_61 =15'b0;

   // m20_62 = W*in
   wire signed [14:0] m20_62;
   assign m20_62 ={ {3{in20[14]}} , in20[14:3] };

   // m20_63 = W*in
   wire signed [14:0] m20_63;
   assign m20_63 =15'b0;

   // m20_64 = W*in
   wire signed [14:0] m20_64;
   assign m20_64 ={ {3{in20[14]}} , in20[14:3] };

   // m20_65 = W*in
   wire signed [14:0] m20_65;
   assign m20_65 =15'b0;

   // m20_66 = W*in
   wire signed [14:0] m20_66;
   assign m20_66 =15'b0;

   // m20_67 = W*in
   wire signed [14:0] m20_67;
   assign m20_67 =15'b0;

   // m20_68 = W*in
   wire signed [14:0] m20_68;
   assign m20_68 ={ {3{in20[14]}} , in20[14:3] };

   // m20_69 = W*in
   wire signed [14:0] m20_69;
   assign m20_69 =15'b0;

   // m20_70 = W*in
   wire signed [14:0] m20_70;
   assign m20_70 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_71 = W*in
   wire signed [14:0] m20_71;
   assign m20_71 =15'b0;

   // m20_72 = W*in
   wire signed [14:0] m20_72;
   assign m20_72 =15'b0;

   // m20_73 = W*in
   wire signed [14:0] m20_73;
   assign m20_73 =15'b0;

   // m20_74 = W*in
   wire signed [14:0] m20_74;
   assign m20_74 =15'b0;

   // m20_75 = W*in
   wire signed [14:0] m20_75;
   assign m20_75 =15'b0;

   // m20_76 = W*in
   wire signed [14:0] m20_76;
   assign m20_76 =15'b0;

   // m20_77 = W*in
   wire signed [14:0] m20_77;
   assign m20_77 =15'b0;

   // m20_78 = W*in
   wire signed [14:0] m20_78;
   assign m20_78 =15'b0;

   // m20_79 = W*in
   wire signed [14:0] m20_79;
   assign m20_79 =15'b0;

   // m20_80 = W*in
   wire signed [14:0] m20_80;
   assign m20_80 =15'b0;

   // m20_81 = W*in
   wire signed [14:0] m20_81;
   assign m20_81 =15'b0;

   // m20_82 = W*in
   wire signed [14:0] m20_82;
   assign m20_82 =15'b0;

   // m20_83 = W*in
   wire signed [14:0] m20_83;
   assign m20_83 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_84 = W*in
   wire signed [14:0] m20_84;
   assign m20_84 =15'b0;

   // m20_85 = W*in
   wire signed [14:0] m20_85;
   assign m20_85 =15'b0;

   // m20_86 = W*in
   wire signed [14:0] m20_86;
   assign m20_86 =15'b0;

   // m20_87 = W*in
   wire signed [14:0] m20_87;
   assign m20_87 ={ {3{in20[14]}} , in20[14:3] };

   // m20_88 = W*in
   wire signed [14:0] m20_88;
   assign m20_88 =15'b0;

   // m20_89 = W*in
   wire signed [14:0] m20_89;
   assign m20_89 =15'b0;

   // m20_90 = W*in
   wire signed [14:0] m20_90;
   assign m20_90 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_91 = W*in
   wire signed [14:0] m20_91;
   assign m20_91 =15'b0;

   // m20_92 = W*in
   wire signed [14:0] m20_92;
   assign m20_92 =15'b0;

   // m20_93 = W*in
   wire signed [14:0] m20_93;
   assign m20_93 =15'b0;

   // m20_94 = W*in
   wire signed [14:0] m20_94;
   assign m20_94 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_95 = W*in
   wire signed [14:0] m20_95;
   assign m20_95 ={ {3{neg20[14]}} , neg20[14:3] };

   // m20_96 = W*in
   wire signed [14:0] m20_96;
   assign m20_96 ={ {3{in20[14]}} , in20[14:3] };

   // m20_97 = W*in
   wire signed [14:0] m20_97;
   assign m20_97 =15'b0;

   // m20_98 = W*in
   wire signed [14:0] m20_98;
   assign m20_98 =15'b0;

   // m20_99 = W*in
   wire signed [14:0] m20_99;
   assign m20_99 =15'b0;

   // m20_100 = W*in
   wire signed [14:0] m20_100;
   assign m20_100 =15'b0;

   // m21_1 = W*in
   wire signed [14:0] m21_1;
   assign m21_1 =15'b0;

   // m21_2 = W*in
   wire signed [14:0] m21_2;
   assign m21_2 =15'b0;

   // m21_3 = W*in
   wire signed [14:0] m21_3;
   assign m21_3 =15'b0;

   // m21_4 = W*in
   wire signed [14:0] m21_4;
   assign m21_4 =15'b0;

   // m21_5 = W*in
   wire signed [14:0] m21_5;
   assign m21_5 =15'b0;

   // m21_6 = W*in
   wire signed [14:0] m21_6;
   assign m21_6 =15'b0;

   // m21_7 = W*in
   wire signed [14:0] m21_7;
   assign m21_7 =15'b0;

   // m21_8 = W*in
   wire signed [14:0] m21_8;
   assign m21_8 =15'b0;

   // m21_9 = W*in
   wire signed [14:0] m21_9;
   assign m21_9 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_10 = W*in
   wire signed [14:0] m21_10;
   assign m21_10 =15'b0;

   // m21_11 = W*in
   wire signed [14:0] m21_11;
   assign m21_11 =15'b0;

   // m21_12 = W*in
   wire signed [14:0] m21_12;
   assign m21_12 =15'b0;

   // m21_13 = W*in
   wire signed [14:0] m21_13;
   assign m21_13 =15'b0;

   // m21_14 = W*in
   wire signed [14:0] m21_14;
   assign m21_14 =15'b0;

   // m21_15 = W*in
   wire signed [14:0] m21_15;
   assign m21_15 =15'b0;

   // m21_16 = W*in
   wire signed [14:0] m21_16;
   assign m21_16 =15'b0;

   // m21_17 = W*in
   wire signed [14:0] m21_17;
   assign m21_17 ={ {3{in21[14]}} , in21[14:3] };

   // m21_18 = W*in
   wire signed [14:0] m21_18;
   assign m21_18 =15'b0;

   // m21_19 = W*in
   wire signed [14:0] m21_19;
   assign m21_19 =15'b0;

   // m21_20 = W*in
   wire signed [14:0] m21_20;
   assign m21_20 =15'b0;

   // m21_21 = W*in
   wire signed [14:0] m21_21;
   assign m21_21 =15'b0;

   // m21_22 = W*in
   wire signed [14:0] m21_22;
   assign m21_22 ={ {4{neg21[14]}} , neg21[14:4] };

   // m21_23 = W*in
   wire signed [14:0] m21_23;
   assign m21_23 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_24 = W*in
   wire signed [14:0] m21_24;
   assign m21_24 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_25 = W*in
   wire signed [14:0] m21_25;
   assign m21_25 =15'b0;

   // m21_26 = W*in
   wire signed [14:0] m21_26;
   assign m21_26 =15'b0;

   // m21_27 = W*in
   wire signed [14:0] m21_27;
   assign m21_27 =15'b0;

   // m21_28 = W*in
   wire signed [14:0] m21_28;
   assign m21_28 ={ {4{in21[14]}} , in21[14:4] };

   // m21_29 = W*in
   wire signed [14:0] m21_29;
   assign m21_29 =15'b0;

   // m21_30 = W*in
   wire signed [14:0] m21_30;
   assign m21_30 =15'b0;

   // m21_31 = W*in
   wire signed [14:0] m21_31;
   assign m21_31 =15'b0;

   // m21_32 = W*in
   wire signed [14:0] m21_32;
   assign m21_32 ={ {3{in21[14]}} , in21[14:3] };

   // m21_33 = W*in
   wire signed [14:0] m21_33;
   assign m21_33 =15'b0;

   // m21_34 = W*in
   wire signed [14:0] m21_34;
   assign m21_34 =15'b0;

   // m21_35 = W*in
   wire signed [14:0] m21_35;
   assign m21_35 =15'b0;

   // m21_36 = W*in
   wire signed [14:0] m21_36;
   assign m21_36 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_37 = W*in
   wire signed [14:0] m21_37;
   assign m21_37 =15'b0;

   // m21_38 = W*in
   wire signed [14:0] m21_38;
   assign m21_38 =15'b0;

   // m21_39 = W*in
   wire signed [14:0] m21_39;
   assign m21_39 =15'b0;

   // m21_40 = W*in
   wire signed [14:0] m21_40;
   assign m21_40 =15'b0;

   // m21_41 = W*in
   wire signed [14:0] m21_41;
   assign m21_41 =15'b0;

   // m21_42 = W*in
   wire signed [14:0] m21_42;
   assign m21_42 =15'b0;

   // m21_43 = W*in
   wire signed [14:0] m21_43;
   assign m21_43 =15'b0;

   // m21_44 = W*in
   wire signed [14:0] m21_44;
   assign m21_44 =15'b0;

   // m21_45 = W*in
   wire signed [14:0] m21_45;
   assign m21_45 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_46 = W*in
   wire signed [14:0] m21_46;
   assign m21_46 =15'b0;

   // m21_47 = W*in
   wire signed [14:0] m21_47;
   assign m21_47 =15'b0;

   // m21_48 = W*in
   wire signed [14:0] m21_48;
   assign m21_48 =15'b0;

   // m21_49 = W*in
   wire signed [14:0] m21_49;
   assign m21_49 =15'b0;

   // m21_50 = W*in
   wire signed [14:0] m21_50;
   assign m21_50 ={ {3{in21[14]}} , in21[14:3] };

   // m21_51 = W*in
   wire signed [14:0] m21_51;
   assign m21_51 ={ {4{in21[14]}} , in21[14:4] };

   // m21_52 = W*in
   wire signed [14:0] m21_52;
   assign m21_52 =15'b0;

   // m21_53 = W*in
   wire signed [14:0] m21_53;
   assign m21_53 ={ {3{in21[14]}} , in21[14:3] };

   // m21_54 = W*in
   wire signed [14:0] m21_54;
   assign m21_54 =15'b0;

   // m21_55 = W*in
   wire signed [14:0] m21_55;
   assign m21_55 ={ {2{in21[14]}} , in21[14:2] };

   // m21_56 = W*in
   wire signed [14:0] m21_56;
   assign m21_56 =15'b0;

   // m21_57 = W*in
   wire signed [14:0] m21_57;
   assign m21_57 =15'b0;

   // m21_58 = W*in
   wire signed [14:0] m21_58;
   assign m21_58 =15'b0;

   // m21_59 = W*in
   wire signed [14:0] m21_59;
   assign m21_59 =15'b0;

   // m21_60 = W*in
   wire signed [14:0] m21_60;
   assign m21_60 ={ {4{neg21[14]}} , neg21[14:4] };

   // m21_61 = W*in
   wire signed [14:0] m21_61;
   assign m21_61 =15'b0;

   // m21_62 = W*in
   wire signed [14:0] m21_62;
   assign m21_62 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_63 = W*in
   wire signed [14:0] m21_63;
   assign m21_63 ={ {2{in21[14]}} , in21[14:2] };

   // m21_64 = W*in
   wire signed [14:0] m21_64;
   assign m21_64 =15'b0;

   // m21_65 = W*in
   wire signed [14:0] m21_65;
   assign m21_65 =15'b0;

   // m21_66 = W*in
   wire signed [14:0] m21_66;
   assign m21_66 =15'b0;

   // m21_67 = W*in
   wire signed [14:0] m21_67;
   assign m21_67 =15'b0;

   // m21_68 = W*in
   wire signed [14:0] m21_68;
   assign m21_68 =15'b0;

   // m21_69 = W*in
   wire signed [14:0] m21_69;
   assign m21_69 =15'b0;

   // m21_70 = W*in
   wire signed [14:0] m21_70;
   assign m21_70 =15'b0;

   // m21_71 = W*in
   wire signed [14:0] m21_71;
   assign m21_71 =15'b0;

   // m21_72 = W*in
   wire signed [14:0] m21_72;
   assign m21_72 =15'b0;

   // m21_73 = W*in
   wire signed [14:0] m21_73;
   assign m21_73 =15'b0;

   // m21_74 = W*in
   wire signed [14:0] m21_74;
   assign m21_74 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_75 = W*in
   wire signed [14:0] m21_75;
   assign m21_75 ={ {4{neg21[14]}} , neg21[14:4] };

   // m21_76 = W*in
   wire signed [14:0] m21_76;
   assign m21_76 =15'b0;

   // m21_77 = W*in
   wire signed [14:0] m21_77;
   assign m21_77 ={ {4{in21[14]}} , in21[14:4] };

   // m21_78 = W*in
   wire signed [14:0] m21_78;
   assign m21_78 =15'b0;

   // m21_79 = W*in
   wire signed [14:0] m21_79;
   assign m21_79 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_80 = W*in
   wire signed [14:0] m21_80;
   assign m21_80 =15'b0;

   // m21_81 = W*in
   wire signed [14:0] m21_81;
   assign m21_81 =15'b0;

   // m21_82 = W*in
   wire signed [14:0] m21_82;
   assign m21_82 =15'b0;

   // m21_83 = W*in
   wire signed [14:0] m21_83;
   assign m21_83 =15'b0;

   // m21_84 = W*in
   wire signed [14:0] m21_84;
   assign m21_84 =15'b0;

   // m21_85 = W*in
   wire signed [14:0] m21_85;
   assign m21_85 =15'b0;

   // m21_86 = W*in
   wire signed [14:0] m21_86;
   assign m21_86 =15'b0;

   // m21_87 = W*in
   wire signed [14:0] m21_87;
   assign m21_87 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_88 = W*in
   wire signed [14:0] m21_88;
   assign m21_88 =15'b0;

   // m21_89 = W*in
   wire signed [14:0] m21_89;
   assign m21_89 =15'b0;

   // m21_90 = W*in
   wire signed [14:0] m21_90;
   assign m21_90 =15'b0;

   // m21_91 = W*in
   wire signed [14:0] m21_91;
   assign m21_91 =15'b0;

   // m21_92 = W*in
   wire signed [14:0] m21_92;
   assign m21_92 =15'b0;

   // m21_93 = W*in
   wire signed [14:0] m21_93;
   assign m21_93 ={ {3{neg21[14]}} , neg21[14:3] };

   // m21_94 = W*in
   wire signed [14:0] m21_94;
   assign m21_94 =15'b0;

   // m21_95 = W*in
   wire signed [14:0] m21_95;
   assign m21_95 =15'b0;

   // m21_96 = W*in
   wire signed [14:0] m21_96;
   assign m21_96 =15'b0;

   // m21_97 = W*in
   wire signed [14:0] m21_97;
   assign m21_97 =15'b0;

   // m21_98 = W*in
   wire signed [14:0] m21_98;
   assign m21_98 =15'b0;

   // m21_99 = W*in
   wire signed [14:0] m21_99;
   assign m21_99 =15'b0;

   // m21_100 = W*in
   wire signed [14:0] m21_100;
   assign m21_100 =15'b0;

   // m22_1 = W*in
   wire signed [14:0] m22_1;
   assign m22_1 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_2 = W*in
   wire signed [14:0] m22_2;
   assign m22_2 =15'b0;

   // m22_3 = W*in
   wire signed [14:0] m22_3;
   assign m22_3 =15'b0;

   // m22_4 = W*in
   wire signed [14:0] m22_4;
   assign m22_4 =15'b0;

   // m22_5 = W*in
   wire signed [14:0] m22_5;
   assign m22_5 =15'b0;

   // m22_6 = W*in
   wire signed [14:0] m22_6;
   assign m22_6 =15'b0;

   // m22_7 = W*in
   wire signed [14:0] m22_7;
   assign m22_7 =15'b0;

   // m22_8 = W*in
   wire signed [14:0] m22_8;
   assign m22_8 =15'b0;

   // m22_9 = W*in
   wire signed [14:0] m22_9;
   assign m22_9 =15'b0;

   // m22_10 = W*in
   wire signed [14:0] m22_10;
   assign m22_10 ={ {3{in22[14]}} , in22[14:3] };

   // m22_11 = W*in
   wire signed [14:0] m22_11;
   assign m22_11 =15'b0;

   // m22_12 = W*in
   wire signed [14:0] m22_12;
   assign m22_12 ={ {3{in22[14]}} , in22[14:3] };

   // m22_13 = W*in
   wire signed [14:0] m22_13;
   assign m22_13 =15'b0;

   // m22_14 = W*in
   wire signed [14:0] m22_14;
   assign m22_14 =15'b0;

   // m22_15 = W*in
   wire signed [14:0] m22_15;
   assign m22_15 =15'b0;

   // m22_16 = W*in
   wire signed [14:0] m22_16;
   assign m22_16 ={ {2{in22[14]}} , in22[14:2] };

   // m22_17 = W*in
   wire signed [14:0] m22_17;
   assign m22_17 =15'b0;

   // m22_18 = W*in
   wire signed [14:0] m22_18;
   assign m22_18 =15'b0;

   // m22_19 = W*in
   wire signed [14:0] m22_19;
   assign m22_19 =15'b0;

   // m22_20 = W*in
   wire signed [14:0] m22_20;
   assign m22_20 =15'b0;

   // m22_21 = W*in
   wire signed [14:0] m22_21;
   assign m22_21 =15'b0;

   // m22_22 = W*in
   wire signed [14:0] m22_22;
   assign m22_22 =15'b0;

   // m22_23 = W*in
   wire signed [14:0] m22_23;
   assign m22_23 =15'b0;

   // m22_24 = W*in
   wire signed [14:0] m22_24;
   assign m22_24 =15'b0;

   // m22_25 = W*in
   wire signed [14:0] m22_25;
   assign m22_25 ={ {4{neg22[14]}} , neg22[14:4] };

   // m22_26 = W*in
   wire signed [14:0] m22_26;
   assign m22_26 ={ {3{in22[14]}} , in22[14:3] };

   // m22_27 = W*in
   wire signed [14:0] m22_27;
   assign m22_27 =15'b0;

   // m22_28 = W*in
   wire signed [14:0] m22_28;
   assign m22_28 ={ {4{neg22[14]}} , neg22[14:4] };

   // m22_29 = W*in
   wire signed [14:0] m22_29;
   assign m22_29 ={ {3{in22[14]}} , in22[14:3] };

   // m22_30 = W*in
   wire signed [14:0] m22_30;
   assign m22_30 ={ {4{in22[14]}} , in22[14:4] };

   // m22_31 = W*in
   wire signed [14:0] m22_31;
   assign m22_31 =15'b0;

   // m22_32 = W*in
   wire signed [14:0] m22_32;
   assign m22_32 =15'b0;

   // m22_33 = W*in
   wire signed [14:0] m22_33;
   assign m22_33 =15'b0;

   // m22_34 = W*in
   wire signed [14:0] m22_34;
   assign m22_34 ={ {3{in22[14]}} , in22[14:3] };

   // m22_35 = W*in
   wire signed [14:0] m22_35;
   assign m22_35 =15'b0;

   // m22_36 = W*in
   wire signed [14:0] m22_36;
   assign m22_36 =15'b0;

   // m22_37 = W*in
   wire signed [14:0] m22_37;
   assign m22_37 =15'b0;

   // m22_38 = W*in
   wire signed [14:0] m22_38;
   assign m22_38 =15'b0;

   // m22_39 = W*in
   wire signed [14:0] m22_39;
   assign m22_39 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_40 = W*in
   wire signed [14:0] m22_40;
   assign m22_40 =15'b0;

   // m22_41 = W*in
   wire signed [14:0] m22_41;
   assign m22_41 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_42 = W*in
   wire signed [14:0] m22_42;
   assign m22_42 =15'b0;

   // m22_43 = W*in
   wire signed [14:0] m22_43;
   assign m22_43 =15'b0;

   // m22_44 = W*in
   wire signed [14:0] m22_44;
   assign m22_44 =15'b0;

   // m22_45 = W*in
   wire signed [14:0] m22_45;
   assign m22_45 =15'b0;

   // m22_46 = W*in
   wire signed [14:0] m22_46;
   assign m22_46 =15'b0;

   // m22_47 = W*in
   wire signed [14:0] m22_47;
   assign m22_47 ={ {4{neg22[14]}} , neg22[14:4] };

   // m22_48 = W*in
   wire signed [14:0] m22_48;
   assign m22_48 =15'b0;

   // m22_49 = W*in
   wire signed [14:0] m22_49;
   assign m22_49 =15'b0;

   // m22_50 = W*in
   wire signed [14:0] m22_50;
   assign m22_50 =15'b0;

   // m22_51 = W*in
   wire signed [14:0] m22_51;
   assign m22_51 =15'b0;

   // m22_52 = W*in
   wire signed [14:0] m22_52;
   assign m22_52 =15'b0;

   // m22_53 = W*in
   wire signed [14:0] m22_53;
   assign m22_53 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_54 = W*in
   wire signed [14:0] m22_54;
   assign m22_54 ={ {3{in22[14]}} , in22[14:3] };

   // m22_55 = W*in
   wire signed [14:0] m22_55;
   assign m22_55 =15'b0;

   // m22_56 = W*in
   wire signed [14:0] m22_56;
   assign m22_56 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_57 = W*in
   wire signed [14:0] m22_57;
   assign m22_57 =15'b0;

   // m22_58 = W*in
   wire signed [14:0] m22_58;
   assign m22_58 =15'b0;

   // m22_59 = W*in
   wire signed [14:0] m22_59;
   assign m22_59 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_60 = W*in
   wire signed [14:0] m22_60;
   assign m22_60 =15'b0;

   // m22_61 = W*in
   wire signed [14:0] m22_61;
   assign m22_61 =15'b0;

   // m22_62 = W*in
   wire signed [14:0] m22_62;
   assign m22_62 =15'b0;

   // m22_63 = W*in
   wire signed [14:0] m22_63;
   assign m22_63 ={ {3{in22[14]}} , in22[14:3] };

   // m22_64 = W*in
   wire signed [14:0] m22_64;
   assign m22_64 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_65 = W*in
   wire signed [14:0] m22_65;
   assign m22_65 ={ {3{in22[14]}} , in22[14:3] };

   // m22_66 = W*in
   wire signed [14:0] m22_66;
   assign m22_66 =15'b0;

   // m22_67 = W*in
   wire signed [14:0] m22_67;
   assign m22_67 ={ {4{neg22[14]}} , neg22[14:4] };

   // m22_68 = W*in
   wire signed [14:0] m22_68;
   assign m22_68 ={ {4{neg22[14]}} , neg22[14:4] };

   // m22_69 = W*in
   wire signed [14:0] m22_69;
   assign m22_69 =15'b0;

   // m22_70 = W*in
   wire signed [14:0] m22_70;
   assign m22_70 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_71 = W*in
   wire signed [14:0] m22_71;
   assign m22_71 =15'b0;

   // m22_72 = W*in
   wire signed [14:0] m22_72;
   assign m22_72 =15'b0;

   // m22_73 = W*in
   wire signed [14:0] m22_73;
   assign m22_73 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_74 = W*in
   wire signed [14:0] m22_74;
   assign m22_74 ={ {4{neg22[14]}} , neg22[14:4] };

   // m22_75 = W*in
   wire signed [14:0] m22_75;
   assign m22_75 =15'b0;

   // m22_76 = W*in
   wire signed [14:0] m22_76;
   assign m22_76 =15'b0;

   // m22_77 = W*in
   wire signed [14:0] m22_77;
   assign m22_77 =15'b0;

   // m22_78 = W*in
   wire signed [14:0] m22_78;
   assign m22_78 =15'b0;

   // m22_79 = W*in
   wire signed [14:0] m22_79;
   assign m22_79 =15'b0;

   // m22_80 = W*in
   wire signed [14:0] m22_80;
   assign m22_80 =15'b0;

   // m22_81 = W*in
   wire signed [14:0] m22_81;
   assign m22_81 =15'b0;

   // m22_82 = W*in
   wire signed [14:0] m22_82;
   assign m22_82 =15'b0;

   // m22_83 = W*in
   wire signed [14:0] m22_83;
   assign m22_83 =15'b0;

   // m22_84 = W*in
   wire signed [14:0] m22_84;
   assign m22_84 =15'b0;

   // m22_85 = W*in
   wire signed [14:0] m22_85;
   assign m22_85 =15'b0;

   // m22_86 = W*in
   wire signed [14:0] m22_86;
   assign m22_86 =15'b0;

   // m22_87 = W*in
   wire signed [14:0] m22_87;
   assign m22_87 =15'b0;

   // m22_88 = W*in
   wire signed [14:0] m22_88;
   assign m22_88 =15'b0;

   // m22_89 = W*in
   wire signed [14:0] m22_89;
   assign m22_89 =15'b0;

   // m22_90 = W*in
   wire signed [14:0] m22_90;
   assign m22_90 =15'b0;

   // m22_91 = W*in
   wire signed [14:0] m22_91;
   assign m22_91 =15'b0;

   // m22_92 = W*in
   wire signed [14:0] m22_92;
   assign m22_92 ={ {3{neg22[14]}} , neg22[14:3] };

   // m22_93 = W*in
   wire signed [14:0] m22_93;
   assign m22_93 =15'b0;

   // m22_94 = W*in
   wire signed [14:0] m22_94;
   assign m22_94 =15'b0;

   // m22_95 = W*in
   wire signed [14:0] m22_95;
   assign m22_95 =15'b0;

   // m22_96 = W*in
   wire signed [14:0] m22_96;
   assign m22_96 =15'b0;

   // m22_97 = W*in
   wire signed [14:0] m22_97;
   assign m22_97 ={ {3{in22[14]}} , in22[14:3] };

   // m22_98 = W*in
   wire signed [14:0] m22_98;
   assign m22_98 =15'b0;

   // m22_99 = W*in
   wire signed [14:0] m22_99;
   assign m22_99 =15'b0;

   // m22_100 = W*in
   wire signed [14:0] m22_100;
   assign m22_100 =15'b0;

   // m23_1 = W*in
   wire signed [14:0] m23_1;
   assign m23_1 =15'b0;

   // m23_2 = W*in
   wire signed [14:0] m23_2;
   assign m23_2 =15'b0;

   // m23_3 = W*in
   wire signed [14:0] m23_3;
   assign m23_3 =15'b0;

   // m23_4 = W*in
   wire signed [14:0] m23_4;
   assign m23_4 =15'b0;

   // m23_5 = W*in
   wire signed [14:0] m23_5;
   assign m23_5 =15'b0;

   // m23_6 = W*in
   wire signed [14:0] m23_6;
   assign m23_6 =15'b0;

   // m23_7 = W*in
   wire signed [14:0] m23_7;
   assign m23_7 ={ {3{neg23[14]}} , neg23[14:3] };

   // m23_8 = W*in
   wire signed [14:0] m23_8;
   assign m23_8 =15'b0;

   // m23_9 = W*in
   wire signed [14:0] m23_9;
   assign m23_9 ={ {3{in23[14]}} , in23[14:3] };

   // m23_10 = W*in
   wire signed [14:0] m23_10;
   assign m23_10 =15'b0;

   // m23_11 = W*in
   wire signed [14:0] m23_11;
   assign m23_11 =15'b0;

   // m23_12 = W*in
   wire signed [14:0] m23_12;
   assign m23_12 =15'b0;

   // m23_13 = W*in
   wire signed [14:0] m23_13;
   assign m23_13 =15'b0;

   // m23_14 = W*in
   wire signed [14:0] m23_14;
   assign m23_14 =15'b0;

   // m23_15 = W*in
   wire signed [14:0] m23_15;
   assign m23_15 ={ {3{neg23[14]}} , neg23[14:3] };

   // m23_16 = W*in
   wire signed [14:0] m23_16;
   assign m23_16 =15'b0;

   // m23_17 = W*in
   wire signed [14:0] m23_17;
   assign m23_17 =15'b0;

   // m23_18 = W*in
   wire signed [14:0] m23_18;
   assign m23_18 =15'b0;

   // m23_19 = W*in
   wire signed [14:0] m23_19;
   assign m23_19 =15'b0;

   // m23_20 = W*in
   wire signed [14:0] m23_20;
   assign m23_20 =15'b0;

   // m23_21 = W*in
   wire signed [14:0] m23_21;
   assign m23_21 ={ {3{in23[14]}} , in23[14:3] };

   // m23_22 = W*in
   wire signed [14:0] m23_22;
   assign m23_22 =15'b0;

   // m23_23 = W*in
   wire signed [14:0] m23_23;
   assign m23_23 =15'b0;

   // m23_24 = W*in
   wire signed [14:0] m23_24;
   assign m23_24 =15'b0;

   // m23_25 = W*in
   wire signed [14:0] m23_25;
   assign m23_25 ={ {4{in23[14]}} , in23[14:4] };

   // m23_26 = W*in
   wire signed [14:0] m23_26;
   assign m23_26 =15'b0;

   // m23_27 = W*in
   wire signed [14:0] m23_27;
   assign m23_27 =15'b0;

   // m23_28 = W*in
   wire signed [14:0] m23_28;
   assign m23_28 ={ {4{neg23[14]}} , neg23[14:4] };

   // m23_29 = W*in
   wire signed [14:0] m23_29;
   assign m23_29 =15'b0;

   // m23_30 = W*in
   wire signed [14:0] m23_30;
   assign m23_30 =15'b0;

   // m23_31 = W*in
   wire signed [14:0] m23_31;
   assign m23_31 =15'b0;

   // m23_32 = W*in
   wire signed [14:0] m23_32;
   assign m23_32 ={ {4{in23[14]}} , in23[14:4] };

   // m23_33 = W*in
   wire signed [14:0] m23_33;
   assign m23_33 ={ {4{neg23[14]}} , neg23[14:4] };

   // m23_34 = W*in
   wire signed [14:0] m23_34;
   assign m23_34 =15'b0;

   // m23_35 = W*in
   wire signed [14:0] m23_35;
   assign m23_35 =15'b0;

   // m23_36 = W*in
   wire signed [14:0] m23_36;
   assign m23_36 =15'b0;

   // m23_37 = W*in
   wire signed [14:0] m23_37;
   assign m23_37 =15'b0;

   // m23_38 = W*in
   wire signed [14:0] m23_38;
   assign m23_38 =15'b0;

   // m23_39 = W*in
   wire signed [14:0] m23_39;
   assign m23_39 =15'b0;

   // m23_40 = W*in
   wire signed [14:0] m23_40;
   assign m23_40 =15'b0;

   // m23_41 = W*in
   wire signed [14:0] m23_41;
   assign m23_41 =15'b0;

   // m23_42 = W*in
   wire signed [14:0] m23_42;
   assign m23_42 =15'b0;

   // m23_43 = W*in
   wire signed [14:0] m23_43;
   assign m23_43 =15'b0;

   // m23_44 = W*in
   wire signed [14:0] m23_44;
   assign m23_44 =15'b0;

   // m23_45 = W*in
   wire signed [14:0] m23_45;
   assign m23_45 =15'b0;

   // m23_46 = W*in
   wire signed [14:0] m23_46;
   assign m23_46 =15'b0;

   // m23_47 = W*in
   wire signed [14:0] m23_47;
   assign m23_47 =15'b0;

   // m23_48 = W*in
   wire signed [14:0] m23_48;
   assign m23_48 =15'b0;

   // m23_49 = W*in
   wire signed [14:0] m23_49;
   assign m23_49 =15'b0;

   // m23_50 = W*in
   wire signed [14:0] m23_50;
   assign m23_50 =15'b0;

   // m23_51 = W*in
   wire signed [14:0] m23_51;
   assign m23_51 =15'b0;

   // m23_52 = W*in
   wire signed [14:0] m23_52;
   assign m23_52 =15'b0;

   // m23_53 = W*in
   wire signed [14:0] m23_53;
   assign m23_53 =15'b0;

   // m23_54 = W*in
   wire signed [14:0] m23_54;
   assign m23_54 =15'b0;

   // m23_55 = W*in
   wire signed [14:0] m23_55;
   assign m23_55 =15'b0;

   // m23_56 = W*in
   wire signed [14:0] m23_56;
   assign m23_56 =15'b0;

   // m23_57 = W*in
   wire signed [14:0] m23_57;
   assign m23_57 =15'b0;

   // m23_58 = W*in
   wire signed [14:0] m23_58;
   assign m23_58 ={ {4{neg23[14]}} , neg23[14:4] };

   // m23_59 = W*in
   wire signed [14:0] m23_59;
   assign m23_59 ={ {4{in23[14]}} , in23[14:4] };

   // m23_60 = W*in
   wire signed [14:0] m23_60;
   assign m23_60 =15'b0;

   // m23_61 = W*in
   wire signed [14:0] m23_61;
   assign m23_61 ={ {4{neg23[14]}} , neg23[14:4] };

   // m23_62 = W*in
   wire signed [14:0] m23_62;
   assign m23_62 =15'b0;

   // m23_63 = W*in
   wire signed [14:0] m23_63;
   assign m23_63 =15'b0;

   // m23_64 = W*in
   wire signed [14:0] m23_64;
   assign m23_64 ={ {4{in23[14]}} , in23[14:4] };

   // m23_65 = W*in
   wire signed [14:0] m23_65;
   assign m23_65 =15'b0;

   // m23_66 = W*in
   wire signed [14:0] m23_66;
   assign m23_66 ={ {3{neg23[14]}} , neg23[14:3] };

   // m23_67 = W*in
   wire signed [14:0] m23_67;
   assign m23_67 =15'b0;

   // m23_68 = W*in
   wire signed [14:0] m23_68;
   assign m23_68 =15'b0;

   // m23_69 = W*in
   wire signed [14:0] m23_69;
   assign m23_69 ={ {4{in23[14]}} , in23[14:4] };

   // m23_70 = W*in
   wire signed [14:0] m23_70;
   assign m23_70 =15'b0;

   // m23_71 = W*in
   wire signed [14:0] m23_71;
   assign m23_71 =15'b0;

   // m23_72 = W*in
   wire signed [14:0] m23_72;
   assign m23_72 =15'b0;

   // m23_73 = W*in
   wire signed [14:0] m23_73;
   assign m23_73 ={ {3{in23[14]}} , in23[14:3] };

   // m23_74 = W*in
   wire signed [14:0] m23_74;
   assign m23_74 =15'b0;

   // m23_75 = W*in
   wire signed [14:0] m23_75;
   assign m23_75 =15'b0;

   // m23_76 = W*in
   wire signed [14:0] m23_76;
   assign m23_76 =15'b0;

   // m23_77 = W*in
   wire signed [14:0] m23_77;
   assign m23_77 =15'b0;

   // m23_78 = W*in
   wire signed [14:0] m23_78;
   assign m23_78 =15'b0;

   // m23_79 = W*in
   wire signed [14:0] m23_79;
   assign m23_79 =15'b0;

   // m23_80 = W*in
   wire signed [14:0] m23_80;
   assign m23_80 =15'b0;

   // m23_81 = W*in
   wire signed [14:0] m23_81;
   assign m23_81 =15'b0;

   // m23_82 = W*in
   wire signed [14:0] m23_82;
   assign m23_82 =15'b0;

   // m23_83 = W*in
   wire signed [14:0] m23_83;
   assign m23_83 ={ {3{neg23[14]}} , neg23[14:3] };

   // m23_84 = W*in
   wire signed [14:0] m23_84;
   assign m23_84 =15'b0;

   // m23_85 = W*in
   wire signed [14:0] m23_85;
   assign m23_85 =15'b0;

   // m23_86 = W*in
   wire signed [14:0] m23_86;
   assign m23_86 =15'b0;

   // m23_87 = W*in
   wire signed [14:0] m23_87;
   assign m23_87 =15'b0;

   // m23_88 = W*in
   wire signed [14:0] m23_88;
   assign m23_88 =15'b0;

   // m23_89 = W*in
   wire signed [14:0] m23_89;
   assign m23_89 =15'b0;

   // m23_90 = W*in
   wire signed [14:0] m23_90;
   assign m23_90 ={ {3{in23[14]}} , in23[14:3] };

   // m23_91 = W*in
   wire signed [14:0] m23_91;
   assign m23_91 =15'b0;

   // m23_92 = W*in
   wire signed [14:0] m23_92;
   assign m23_92 =15'b0;

   // m23_93 = W*in
   wire signed [14:0] m23_93;
   assign m23_93 =15'b0;

   // m23_94 = W*in
   wire signed [14:0] m23_94;
   assign m23_94 =15'b0;

   // m23_95 = W*in
   wire signed [14:0] m23_95;
   assign m23_95 =15'b0;

   // m23_96 = W*in
   wire signed [14:0] m23_96;
   assign m23_96 =15'b0;

   // m23_97 = W*in
   wire signed [14:0] m23_97;
   assign m23_97 =15'b0;

   // m23_98 = W*in
   wire signed [14:0] m23_98;
   assign m23_98 =15'b0;

   // m23_99 = W*in
   wire signed [14:0] m23_99;
   assign m23_99 =15'b0;

   // m23_100 = W*in
   wire signed [14:0] m23_100;
   assign m23_100 =15'b0;

   // m24_1 = W*in
   wire signed [14:0] m24_1;
   assign m24_1 =15'b0;

   // m24_2 = W*in
   wire signed [14:0] m24_2;
   assign m24_2 =15'b0;

   // m24_3 = W*in
   wire signed [14:0] m24_3;
   assign m24_3 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_4 = W*in
   wire signed [14:0] m24_4;
   assign m24_4 ={ {3{in24[14]}} , in24[14:3] };

   // m24_5 = W*in
   wire signed [14:0] m24_5;
   assign m24_5 =15'b0;

   // m24_6 = W*in
   wire signed [14:0] m24_6;
   assign m24_6 =15'b0;

   // m24_7 = W*in
   wire signed [14:0] m24_7;
   assign m24_7 =15'b0;

   // m24_8 = W*in
   wire signed [14:0] m24_8;
   assign m24_8 =15'b0;

   // m24_9 = W*in
   wire signed [14:0] m24_9;
   assign m24_9 ={ {3{in24[14]}} , in24[14:3] };

   // m24_10 = W*in
   wire signed [14:0] m24_10;
   assign m24_10 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_11 = W*in
   wire signed [14:0] m24_11;
   assign m24_11 =15'b0;

   // m24_12 = W*in
   wire signed [14:0] m24_12;
   assign m24_12 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_13 = W*in
   wire signed [14:0] m24_13;
   assign m24_13 =15'b0;

   // m24_14 = W*in
   wire signed [14:0] m24_14;
   assign m24_14 ={ {3{in24[14]}} , in24[14:3] };

   // m24_15 = W*in
   wire signed [14:0] m24_15;
   assign m24_15 =15'b0;

   // m24_16 = W*in
   wire signed [14:0] m24_16;
   assign m24_16 =15'b0;

   // m24_17 = W*in
   wire signed [14:0] m24_17;
   assign m24_17 =15'b0;

   // m24_18 = W*in
   wire signed [14:0] m24_18;
   assign m24_18 ={ {3{in24[14]}} , in24[14:3] };

   // m24_19 = W*in
   wire signed [14:0] m24_19;
   assign m24_19 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_20 = W*in
   wire signed [14:0] m24_20;
   assign m24_20 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_21 = W*in
   wire signed [14:0] m24_21;
   assign m24_21 =15'b0;

   // m24_22 = W*in
   wire signed [14:0] m24_22;
   assign m24_22 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_23 = W*in
   wire signed [14:0] m24_23;
   assign m24_23 =15'b0;

   // m24_24 = W*in
   wire signed [14:0] m24_24;
   assign m24_24 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_25 = W*in
   wire signed [14:0] m24_25;
   assign m24_25 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_26 = W*in
   wire signed [14:0] m24_26;
   assign m24_26 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_27 = W*in
   wire signed [14:0] m24_27;
   assign m24_27 =15'b0;

   // m24_28 = W*in
   wire signed [14:0] m24_28;
   assign m24_28 ={ {3{in24[14]}} , in24[14:3] };

   // m24_29 = W*in
   wire signed [14:0] m24_29;
   assign m24_29 =15'b0;

   // m24_30 = W*in
   wire signed [14:0] m24_30;
   assign m24_30 ={ {4{in24[14]}} , in24[14:4] };

   // m24_31 = W*in
   wire signed [14:0] m24_31;
   assign m24_31 =15'b0;

   // m24_32 = W*in
   wire signed [14:0] m24_32;
   assign m24_32 ={ {3{in24[14]}} , in24[14:3] };

   // m24_33 = W*in
   wire signed [14:0] m24_33;
   assign m24_33 ={ {3{in24[14]}} , in24[14:3] };

   // m24_34 = W*in
   wire signed [14:0] m24_34;
   assign m24_34 =15'b0;

   // m24_35 = W*in
   wire signed [14:0] m24_35;
   assign m24_35 =15'b0;

   // m24_36 = W*in
   wire signed [14:0] m24_36;
   assign m24_36 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_37 = W*in
   wire signed [14:0] m24_37;
   assign m24_37 =15'b0;

   // m24_38 = W*in
   wire signed [14:0] m24_38;
   assign m24_38 =15'b0;

   // m24_39 = W*in
   wire signed [14:0] m24_39;
   assign m24_39 =15'b0;

   // m24_40 = W*in
   wire signed [14:0] m24_40;
   assign m24_40 ={ {3{in24[14]}} , in24[14:3] };

   // m24_41 = W*in
   wire signed [14:0] m24_41;
   assign m24_41 =15'b0;

   // m24_42 = W*in
   wire signed [14:0] m24_42;
   assign m24_42 =15'b0;

   // m24_43 = W*in
   wire signed [14:0] m24_43;
   assign m24_43 =15'b0;

   // m24_44 = W*in
   wire signed [14:0] m24_44;
   assign m24_44 =15'b0;

   // m24_45 = W*in
   wire signed [14:0] m24_45;
   assign m24_45 =15'b0;

   // m24_46 = W*in
   wire signed [14:0] m24_46;
   assign m24_46 =15'b0;

   // m24_47 = W*in
   wire signed [14:0] m24_47;
   assign m24_47 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_48 = W*in
   wire signed [14:0] m24_48;
   assign m24_48 =15'b0;

   // m24_49 = W*in
   wire signed [14:0] m24_49;
   assign m24_49 =15'b0;

   // m24_50 = W*in
   wire signed [14:0] m24_50;
   assign m24_50 =15'b0;

   // m24_51 = W*in
   wire signed [14:0] m24_51;
   assign m24_51 =15'b0;

   // m24_52 = W*in
   wire signed [14:0] m24_52;
   assign m24_52 =15'b0;

   // m24_53 = W*in
   wire signed [14:0] m24_53;
   assign m24_53 =15'b0;

   // m24_54 = W*in
   wire signed [14:0] m24_54;
   assign m24_54 =15'b0;

   // m24_55 = W*in
   wire signed [14:0] m24_55;
   assign m24_55 ={ {3{in24[14]}} , in24[14:3] };

   // m24_56 = W*in
   wire signed [14:0] m24_56;
   assign m24_56 =15'b0;

   // m24_57 = W*in
   wire signed [14:0] m24_57;
   assign m24_57 =15'b0;

   // m24_58 = W*in
   wire signed [14:0] m24_58;
   assign m24_58 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_59 = W*in
   wire signed [14:0] m24_59;
   assign m24_59 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_60 = W*in
   wire signed [14:0] m24_60;
   assign m24_60 =15'b0;

   // m24_61 = W*in
   wire signed [14:0] m24_61;
   assign m24_61 =15'b0;

   // m24_62 = W*in
   wire signed [14:0] m24_62;
   assign m24_62 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_63 = W*in
   wire signed [14:0] m24_63;
   assign m24_63 =15'b0;

   // m24_64 = W*in
   wire signed [14:0] m24_64;
   assign m24_64 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_65 = W*in
   wire signed [14:0] m24_65;
   assign m24_65 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_66 = W*in
   wire signed [14:0] m24_66;
   assign m24_66 =15'b0;

   // m24_67 = W*in
   wire signed [14:0] m24_67;
   assign m24_67 =15'b0;

   // m24_68 = W*in
   wire signed [14:0] m24_68;
   assign m24_68 ={ {3{in24[14]}} , in24[14:3] };

   // m24_69 = W*in
   wire signed [14:0] m24_69;
   assign m24_69 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_70 = W*in
   wire signed [14:0] m24_70;
   assign m24_70 =15'b0;

   // m24_71 = W*in
   wire signed [14:0] m24_71;
   assign m24_71 =15'b0;

   // m24_72 = W*in
   wire signed [14:0] m24_72;
   assign m24_72 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_73 = W*in
   wire signed [14:0] m24_73;
   assign m24_73 =15'b0;

   // m24_74 = W*in
   wire signed [14:0] m24_74;
   assign m24_74 =15'b0;

   // m24_75 = W*in
   wire signed [14:0] m24_75;
   assign m24_75 =15'b0;

   // m24_76 = W*in
   wire signed [14:0] m24_76;
   assign m24_76 =15'b0;

   // m24_77 = W*in
   wire signed [14:0] m24_77;
   assign m24_77 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_78 = W*in
   wire signed [14:0] m24_78;
   assign m24_78 ={ {3{in24[14]}} , in24[14:3] };

   // m24_79 = W*in
   wire signed [14:0] m24_79;
   assign m24_79 ={ {4{neg24[14]}} , neg24[14:4] };

   // m24_80 = W*in
   wire signed [14:0] m24_80;
   assign m24_80 =15'b0;

   // m24_81 = W*in
   wire signed [14:0] m24_81;
   assign m24_81 =15'b0;

   // m24_82 = W*in
   wire signed [14:0] m24_82;
   assign m24_82 =15'b0;

   // m24_83 = W*in
   wire signed [14:0] m24_83;
   assign m24_83 =15'b0;

   // m24_84 = W*in
   wire signed [14:0] m24_84;
   assign m24_84 =15'b0;

   // m24_85 = W*in
   wire signed [14:0] m24_85;
   assign m24_85 =15'b0;

   // m24_86 = W*in
   wire signed [14:0] m24_86;
   assign m24_86 =15'b0;

   // m24_87 = W*in
   wire signed [14:0] m24_87;
   assign m24_87 =15'b0;

   // m24_88 = W*in
   wire signed [14:0] m24_88;
   assign m24_88 =15'b0;

   // m24_89 = W*in
   wire signed [14:0] m24_89;
   assign m24_89 =15'b0;

   // m24_90 = W*in
   wire signed [14:0] m24_90;
   assign m24_90 =15'b0;

   // m24_91 = W*in
   wire signed [14:0] m24_91;
   assign m24_91 =15'b0;

   // m24_92 = W*in
   wire signed [14:0] m24_92;
   assign m24_92 =15'b0;

   // m24_93 = W*in
   wire signed [14:0] m24_93;
   assign m24_93 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_94 = W*in
   wire signed [14:0] m24_94;
   assign m24_94 ={ {3{in24[14]}} , in24[14:3] };

   // m24_95 = W*in
   wire signed [14:0] m24_95;
   assign m24_95 =15'b0;

   // m24_96 = W*in
   wire signed [14:0] m24_96;
   assign m24_96 ={ {3{neg24[14]}} , neg24[14:3] };

   // m24_97 = W*in
   wire signed [14:0] m24_97;
   assign m24_97 =15'b0;

   // m24_98 = W*in
   wire signed [14:0] m24_98;
   assign m24_98 =15'b0;

   // m24_99 = W*in
   wire signed [14:0] m24_99;
   assign m24_99 =15'b0;

   // m24_100 = W*in
   wire signed [14:0] m24_100;
   assign m24_100 =15'b0;

   // m25_1 = W*in
   wire signed [14:0] m25_1;
   assign m25_1 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_2 = W*in
   wire signed [14:0] m25_2;
   assign m25_2 =15'b0;

   // m25_3 = W*in
   wire signed [14:0] m25_3;
   assign m25_3 =15'b0;

   // m25_4 = W*in
   wire signed [14:0] m25_4;
   assign m25_4 =15'b0;

   // m25_5 = W*in
   wire signed [14:0] m25_5;
   assign m25_5 =15'b0;

   // m25_6 = W*in
   wire signed [14:0] m25_6;
   assign m25_6 =15'b0;

   // m25_7 = W*in
   wire signed [14:0] m25_7;
   assign m25_7 =15'b0;

   // m25_8 = W*in
   wire signed [14:0] m25_8;
   assign m25_8 =15'b0;

   // m25_9 = W*in
   wire signed [14:0] m25_9;
   assign m25_9 =15'b0;

   // m25_10 = W*in
   wire signed [14:0] m25_10;
   assign m25_10 =15'b0;

   // m25_11 = W*in
   wire signed [14:0] m25_11;
   assign m25_11 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_12 = W*in
   wire signed [14:0] m25_12;
   assign m25_12 =15'b0;

   // m25_13 = W*in
   wire signed [14:0] m25_13;
   assign m25_13 =15'b0;

   // m25_14 = W*in
   wire signed [14:0] m25_14;
   assign m25_14 =15'b0;

   // m25_15 = W*in
   wire signed [14:0] m25_15;
   assign m25_15 =15'b0;

   // m25_16 = W*in
   wire signed [14:0] m25_16;
   assign m25_16 =15'b0;

   // m25_17 = W*in
   wire signed [14:0] m25_17;
   assign m25_17 =15'b0;

   // m25_18 = W*in
   wire signed [14:0] m25_18;
   assign m25_18 =15'b0;

   // m25_19 = W*in
   wire signed [14:0] m25_19;
   assign m25_19 =15'b0;

   // m25_20 = W*in
   wire signed [14:0] m25_20;
   assign m25_20 =15'b0;

   // m25_21 = W*in
   wire signed [14:0] m25_21;
   assign m25_21 =15'b0;

   // m25_22 = W*in
   wire signed [14:0] m25_22;
   assign m25_22 ={ {3{in25[14]}} , in25[14:3] };

   // m25_23 = W*in
   wire signed [14:0] m25_23;
   assign m25_23 =15'b0;

   // m25_24 = W*in
   wire signed [14:0] m25_24;
   assign m25_24 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_25 = W*in
   wire signed [14:0] m25_25;
   assign m25_25 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_26 = W*in
   wire signed [14:0] m25_26;
   assign m25_26 =15'b0;

   // m25_27 = W*in
   wire signed [14:0] m25_27;
   assign m25_27 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_28 = W*in
   wire signed [14:0] m25_28;
   assign m25_28 =15'b0;

   // m25_29 = W*in
   wire signed [14:0] m25_29;
   assign m25_29 =15'b0;

   // m25_30 = W*in
   wire signed [14:0] m25_30;
   assign m25_30 =15'b0;

   // m25_31 = W*in
   wire signed [14:0] m25_31;
   assign m25_31 =15'b0;

   // m25_32 = W*in
   wire signed [14:0] m25_32;
   assign m25_32 =15'b0;

   // m25_33 = W*in
   wire signed [14:0] m25_33;
   assign m25_33 =15'b0;

   // m25_34 = W*in
   wire signed [14:0] m25_34;
   assign m25_34 =15'b0;

   // m25_35 = W*in
   wire signed [14:0] m25_35;
   assign m25_35 =15'b0;

   // m25_36 = W*in
   wire signed [14:0] m25_36;
   assign m25_36 =15'b0;

   // m25_37 = W*in
   wire signed [14:0] m25_37;
   assign m25_37 ={ {3{in25[14]}} , in25[14:3] };

   // m25_38 = W*in
   wire signed [14:0] m25_38;
   assign m25_38 =15'b0;

   // m25_39 = W*in
   wire signed [14:0] m25_39;
   assign m25_39 =15'b0;

   // m25_40 = W*in
   wire signed [14:0] m25_40;
   assign m25_40 =15'b0;

   // m25_41 = W*in
   wire signed [14:0] m25_41;
   assign m25_41 ={ {4{neg25[14]}} , neg25[14:4] };

   // m25_42 = W*in
   wire signed [14:0] m25_42;
   assign m25_42 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_43 = W*in
   wire signed [14:0] m25_43;
   assign m25_43 =15'b0;

   // m25_44 = W*in
   wire signed [14:0] m25_44;
   assign m25_44 =15'b0;

   // m25_45 = W*in
   wire signed [14:0] m25_45;
   assign m25_45 =15'b0;

   // m25_46 = W*in
   wire signed [14:0] m25_46;
   assign m25_46 =15'b0;

   // m25_47 = W*in
   wire signed [14:0] m25_47;
   assign m25_47 =15'b0;

   // m25_48 = W*in
   wire signed [14:0] m25_48;
   assign m25_48 =15'b0;

   // m25_49 = W*in
   wire signed [14:0] m25_49;
   assign m25_49 =15'b0;

   // m25_50 = W*in
   wire signed [14:0] m25_50;
   assign m25_50 =15'b0;

   // m25_51 = W*in
   wire signed [14:0] m25_51;
   assign m25_51 =15'b0;

   // m25_52 = W*in
   wire signed [14:0] m25_52;
   assign m25_52 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_53 = W*in
   wire signed [14:0] m25_53;
   assign m25_53 =15'b0;

   // m25_54 = W*in
   wire signed [14:0] m25_54;
   assign m25_54 =15'b0;

   // m25_55 = W*in
   wire signed [14:0] m25_55;
   assign m25_55 =15'b0;

   // m25_56 = W*in
   wire signed [14:0] m25_56;
   assign m25_56 =15'b0;

   // m25_57 = W*in
   wire signed [14:0] m25_57;
   assign m25_57 =15'b0;

   // m25_58 = W*in
   wire signed [14:0] m25_58;
   assign m25_58 =15'b0;

   // m25_59 = W*in
   wire signed [14:0] m25_59;
   assign m25_59 =15'b0;

   // m25_60 = W*in
   wire signed [14:0] m25_60;
   assign m25_60 =15'b0;

   // m25_61 = W*in
   wire signed [14:0] m25_61;
   assign m25_61 ={ {3{in25[14]}} , in25[14:3] };

   // m25_62 = W*in
   wire signed [14:0] m25_62;
   assign m25_62 =15'b0;

   // m25_63 = W*in
   wire signed [14:0] m25_63;
   assign m25_63 ={ {3{in25[14]}} , in25[14:3] };

   // m25_64 = W*in
   wire signed [14:0] m25_64;
   assign m25_64 =15'b0;

   // m25_65 = W*in
   wire signed [14:0] m25_65;
   assign m25_65 =15'b0;

   // m25_66 = W*in
   wire signed [14:0] m25_66;
   assign m25_66 =15'b0;

   // m25_67 = W*in
   wire signed [14:0] m25_67;
   assign m25_67 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_68 = W*in
   wire signed [14:0] m25_68;
   assign m25_68 =15'b0;

   // m25_69 = W*in
   wire signed [14:0] m25_69;
   assign m25_69 =15'b0;

   // m25_70 = W*in
   wire signed [14:0] m25_70;
   assign m25_70 =15'b0;

   // m25_71 = W*in
   wire signed [14:0] m25_71;
   assign m25_71 =15'b0;

   // m25_72 = W*in
   wire signed [14:0] m25_72;
   assign m25_72 =15'b0;

   // m25_73 = W*in
   wire signed [14:0] m25_73;
   assign m25_73 =15'b0;

   // m25_74 = W*in
   wire signed [14:0] m25_74;
   assign m25_74 =15'b0;

   // m25_75 = W*in
   wire signed [14:0] m25_75;
   assign m25_75 =15'b0;

   // m25_76 = W*in
   wire signed [14:0] m25_76;
   assign m25_76 =15'b0;

   // m25_77 = W*in
   wire signed [14:0] m25_77;
   assign m25_77 =15'b0;

   // m25_78 = W*in
   wire signed [14:0] m25_78;
   assign m25_78 =15'b0;

   // m25_79 = W*in
   wire signed [14:0] m25_79;
   assign m25_79 =15'b0;

   // m25_80 = W*in
   wire signed [14:0] m25_80;
   assign m25_80 =15'b0;

   // m25_81 = W*in
   wire signed [14:0] m25_81;
   assign m25_81 =15'b0;

   // m25_82 = W*in
   wire signed [14:0] m25_82;
   assign m25_82 =15'b0;

   // m25_83 = W*in
   wire signed [14:0] m25_83;
   assign m25_83 =15'b0;

   // m25_84 = W*in
   wire signed [14:0] m25_84;
   assign m25_84 =15'b0;

   // m25_85 = W*in
   wire signed [14:0] m25_85;
   assign m25_85 =15'b0;

   // m25_86 = W*in
   wire signed [14:0] m25_86;
   assign m25_86 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_87 = W*in
   wire signed [14:0] m25_87;
   assign m25_87 =15'b0;

   // m25_88 = W*in
   wire signed [14:0] m25_88;
   assign m25_88 =15'b0;

   // m25_89 = W*in
   wire signed [14:0] m25_89;
   assign m25_89 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_90 = W*in
   wire signed [14:0] m25_90;
   assign m25_90 =15'b0;

   // m25_91 = W*in
   wire signed [14:0] m25_91;
   assign m25_91 ={ {4{in25[14]}} , in25[14:4] };

   // m25_92 = W*in
   wire signed [14:0] m25_92;
   assign m25_92 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_93 = W*in
   wire signed [14:0] m25_93;
   assign m25_93 ={ {4{in25[14]}} , in25[14:4] };

   // m25_94 = W*in
   wire signed [14:0] m25_94;
   assign m25_94 =15'b0;

   // m25_95 = W*in
   wire signed [14:0] m25_95;
   assign m25_95 ={ {3{neg25[14]}} , neg25[14:3] };

   // m25_96 = W*in
   wire signed [14:0] m25_96;
   assign m25_96 =15'b0;

   // m25_97 = W*in
   wire signed [14:0] m25_97;
   assign m25_97 =15'b0;

   // m25_98 = W*in
   wire signed [14:0] m25_98;
   assign m25_98 =15'b0;

   // m25_99 = W*in
   wire signed [14:0] m25_99;
   assign m25_99 =15'b0;

   // m25_100 = W*in
   wire signed [14:0] m25_100;
   assign m25_100 ={ {2{in25[14]}} , in25[14:2] };

   // m26_1 = W*in
   wire signed [14:0] m26_1;
   assign m26_1 =15'b0;

   // m26_2 = W*in
   wire signed [14:0] m26_2;
   assign m26_2 =15'b0;

   // m26_3 = W*in
   wire signed [14:0] m26_3;
   assign m26_3 =15'b0;

   // m26_4 = W*in
   wire signed [14:0] m26_4;
   assign m26_4 =15'b0;

   // m26_5 = W*in
   wire signed [14:0] m26_5;
   assign m26_5 =15'b0;

   // m26_6 = W*in
   wire signed [14:0] m26_6;
   assign m26_6 =15'b0;

   // m26_7 = W*in
   wire signed [14:0] m26_7;
   assign m26_7 =15'b0;

   // m26_8 = W*in
   wire signed [14:0] m26_8;
   assign m26_8 =15'b0;

   // m26_9 = W*in
   wire signed [14:0] m26_9;
   assign m26_9 =15'b0;

   // m26_10 = W*in
   wire signed [14:0] m26_10;
   assign m26_10 =15'b0;

   // m26_11 = W*in
   wire signed [14:0] m26_11;
   assign m26_11 =15'b0;

   // m26_12 = W*in
   wire signed [14:0] m26_12;
   assign m26_12 ={ {3{in26[14]}} , in26[14:3] };

   // m26_13 = W*in
   wire signed [14:0] m26_13;
   assign m26_13 =15'b0;

   // m26_14 = W*in
   wire signed [14:0] m26_14;
   assign m26_14 =15'b0;

   // m26_15 = W*in
   wire signed [14:0] m26_15;
   assign m26_15 =15'b0;

   // m26_16 = W*in
   wire signed [14:0] m26_16;
   assign m26_16 ={ {3{in26[14]}} , in26[14:3] };

   // m26_17 = W*in
   wire signed [14:0] m26_17;
   assign m26_17 =15'b0;

   // m26_18 = W*in
   wire signed [14:0] m26_18;
   assign m26_18 =15'b0;

   // m26_19 = W*in
   wire signed [14:0] m26_19;
   assign m26_19 =15'b0;

   // m26_20 = W*in
   wire signed [14:0] m26_20;
   assign m26_20 ={ {3{neg26[14]}} , neg26[14:3] };

   // m26_21 = W*in
   wire signed [14:0] m26_21;
   assign m26_21 =15'b0;

   // m26_22 = W*in
   wire signed [14:0] m26_22;
   assign m26_22 ={ {4{in26[14]}} , in26[14:4] };

   // m26_23 = W*in
   wire signed [14:0] m26_23;
   assign m26_23 =15'b0;

   // m26_24 = W*in
   wire signed [14:0] m26_24;
   assign m26_24 =15'b0;

   // m26_25 = W*in
   wire signed [14:0] m26_25;
   assign m26_25 =15'b0;

   // m26_26 = W*in
   wire signed [14:0] m26_26;
   assign m26_26 =15'b0;

   // m26_27 = W*in
   wire signed [14:0] m26_27;
   assign m26_27 =15'b0;

   // m26_28 = W*in
   wire signed [14:0] m26_28;
   assign m26_28 =15'b0;

   // m26_29 = W*in
   wire signed [14:0] m26_29;
   assign m26_29 =15'b0;

   // m26_30 = W*in
   wire signed [14:0] m26_30;
   assign m26_30 ={ {4{neg26[14]}} , neg26[14:4] };

   // m26_31 = W*in
   wire signed [14:0] m26_31;
   assign m26_31 =15'b0;

   // m26_32 = W*in
   wire signed [14:0] m26_32;
   assign m26_32 =15'b0;

   // m26_33 = W*in
   wire signed [14:0] m26_33;
   assign m26_33 =15'b0;

   // m26_34 = W*in
   wire signed [14:0] m26_34;
   assign m26_34 =15'b0;

   // m26_35 = W*in
   wire signed [14:0] m26_35;
   assign m26_35 =15'b0;

   // m26_36 = W*in
   wire signed [14:0] m26_36;
   assign m26_36 =15'b0;

   // m26_37 = W*in
   wire signed [14:0] m26_37;
   assign m26_37 =15'b0;

   // m26_38 = W*in
   wire signed [14:0] m26_38;
   assign m26_38 =15'b0;

   // m26_39 = W*in
   wire signed [14:0] m26_39;
   assign m26_39 =15'b0;

   // m26_40 = W*in
   wire signed [14:0] m26_40;
   assign m26_40 =15'b0;

   // m26_41 = W*in
   wire signed [14:0] m26_41;
   assign m26_41 =15'b0;

   // m26_42 = W*in
   wire signed [14:0] m26_42;
   assign m26_42 =15'b0;

   // m26_43 = W*in
   wire signed [14:0] m26_43;
   assign m26_43 =15'b0;

   // m26_44 = W*in
   wire signed [14:0] m26_44;
   assign m26_44 =15'b0;

   // m26_45 = W*in
   wire signed [14:0] m26_45;
   assign m26_45 =15'b0;

   // m26_46 = W*in
   wire signed [14:0] m26_46;
   assign m26_46 =15'b0;

   // m26_47 = W*in
   wire signed [14:0] m26_47;
   assign m26_47 =15'b0;

   // m26_48 = W*in
   wire signed [14:0] m26_48;
   assign m26_48 =15'b0;

   // m26_49 = W*in
   wire signed [14:0] m26_49;
   assign m26_49 =15'b0;

   // m26_50 = W*in
   wire signed [14:0] m26_50;
   assign m26_50 =15'b0;

   // m26_51 = W*in
   wire signed [14:0] m26_51;
   assign m26_51 =15'b0;

   // m26_52 = W*in
   wire signed [14:0] m26_52;
   assign m26_52 =15'b0;

   // m26_53 = W*in
   wire signed [14:0] m26_53;
   assign m26_53 =15'b0;

   // m26_54 = W*in
   wire signed [14:0] m26_54;
   assign m26_54 =15'b0;

   // m26_55 = W*in
   wire signed [14:0] m26_55;
   assign m26_55 =15'b0;

   // m26_56 = W*in
   wire signed [14:0] m26_56;
   assign m26_56 =15'b0;

   // m26_57 = W*in
   wire signed [14:0] m26_57;
   assign m26_57 =15'b0;

   // m26_58 = W*in
   wire signed [14:0] m26_58;
   assign m26_58 =15'b0;

   // m26_59 = W*in
   wire signed [14:0] m26_59;
   assign m26_59 =15'b0;

   // m26_60 = W*in
   wire signed [14:0] m26_60;
   assign m26_60 =15'b0;

   // m26_61 = W*in
   wire signed [14:0] m26_61;
   assign m26_61 =15'b0;

   // m26_62 = W*in
   wire signed [14:0] m26_62;
   assign m26_62 =15'b0;

   // m26_63 = W*in
   wire signed [14:0] m26_63;
   assign m26_63 =15'b0;

   // m26_64 = W*in
   wire signed [14:0] m26_64;
   assign m26_64 =15'b0;

   // m26_65 = W*in
   wire signed [14:0] m26_65;
   assign m26_65 =15'b0;

   // m26_66 = W*in
   wire signed [14:0] m26_66;
   assign m26_66 =15'b0;

   // m26_67 = W*in
   wire signed [14:0] m26_67;
   assign m26_67 =15'b0;

   // m26_68 = W*in
   wire signed [14:0] m26_68;
   assign m26_68 =15'b0;

   // m26_69 = W*in
   wire signed [14:0] m26_69;
   assign m26_69 =15'b0;

   // m26_70 = W*in
   wire signed [14:0] m26_70;
   assign m26_70 =15'b0;

   // m26_71 = W*in
   wire signed [14:0] m26_71;
   assign m26_71 =15'b0;

   // m26_72 = W*in
   wire signed [14:0] m26_72;
   assign m26_72 ={ {3{neg26[14]}} , neg26[14:3] };

   // m26_73 = W*in
   wire signed [14:0] m26_73;
   assign m26_73 =15'b0;

   // m26_74 = W*in
   wire signed [14:0] m26_74;
   assign m26_74 ={ {4{neg26[14]}} , neg26[14:4] };

   // m26_75 = W*in
   wire signed [14:0] m26_75;
   assign m26_75 =15'b0;

   // m26_76 = W*in
   wire signed [14:0] m26_76;
   assign m26_76 =15'b0;

   // m26_77 = W*in
   wire signed [14:0] m26_77;
   assign m26_77 =15'b0;

   // m26_78 = W*in
   wire signed [14:0] m26_78;
   assign m26_78 =15'b0;

   // m26_79 = W*in
   wire signed [14:0] m26_79;
   assign m26_79 ={ {2{in26[14]}} , in26[14:2] };

   // m26_80 = W*in
   wire signed [14:0] m26_80;
   assign m26_80 =15'b0;

   // m26_81 = W*in
   wire signed [14:0] m26_81;
   assign m26_81 =15'b0;

   // m26_82 = W*in
   wire signed [14:0] m26_82;
   assign m26_82 =15'b0;

   // m26_83 = W*in
   wire signed [14:0] m26_83;
   assign m26_83 ={ {4{in26[14]}} , in26[14:4] };

   // m26_84 = W*in
   wire signed [14:0] m26_84;
   assign m26_84 =15'b0;

   // m26_85 = W*in
   wire signed [14:0] m26_85;
   assign m26_85 =15'b0;

   // m26_86 = W*in
   wire signed [14:0] m26_86;
   assign m26_86 ={ {4{in26[14]}} , in26[14:4] };

   // m26_87 = W*in
   wire signed [14:0] m26_87;
   assign m26_87 =15'b0;

   // m26_88 = W*in
   wire signed [14:0] m26_88;
   assign m26_88 =15'b0;

   // m26_89 = W*in
   wire signed [14:0] m26_89;
   assign m26_89 =15'b0;

   // m26_90 = W*in
   wire signed [14:0] m26_90;
   assign m26_90 =15'b0;

   // m26_91 = W*in
   wire signed [14:0] m26_91;
   assign m26_91 =15'b0;

   // m26_92 = W*in
   wire signed [14:0] m26_92;
   assign m26_92 ={ {4{neg26[14]}} , neg26[14:4] };

   // m26_93 = W*in
   wire signed [14:0] m26_93;
   assign m26_93 =15'b0;

   // m26_94 = W*in
   wire signed [14:0] m26_94;
   assign m26_94 =15'b0;

   // m26_95 = W*in
   wire signed [14:0] m26_95;
   assign m26_95 ={ {4{neg26[14]}} , neg26[14:4] };

   // m26_96 = W*in
   wire signed [14:0] m26_96;
   assign m26_96 =15'b0;

   // m26_97 = W*in
   wire signed [14:0] m26_97;
   assign m26_97 ={ {4{neg26[14]}} , neg26[14:4] };

   // m26_98 = W*in
   wire signed [14:0] m26_98;
   assign m26_98 =15'b0;

   // m26_99 = W*in
   wire signed [14:0] m26_99;
   assign m26_99 ={ {3{neg26[14]}} , neg26[14:3] };

   // m26_100 = W*in
   wire signed [14:0] m26_100;
   assign m26_100 =15'b0;

   // m27_1 = W*in
   wire signed [14:0] m27_1;
   assign m27_1 =15'b0;

   // m27_2 = W*in
   wire signed [14:0] m27_2;
   assign m27_2 =15'b0;

   // m27_3 = W*in
   wire signed [14:0] m27_3;
   assign m27_3 =15'b0;

   // m27_4 = W*in
   wire signed [14:0] m27_4;
   assign m27_4 =15'b0;

   // m27_5 = W*in
   wire signed [14:0] m27_5;
   assign m27_5 =15'b0;

   // m27_6 = W*in
   wire signed [14:0] m27_6;
   assign m27_6 =15'b0;

   // m27_7 = W*in
   wire signed [14:0] m27_7;
   assign m27_7 =15'b0;

   // m27_8 = W*in
   wire signed [14:0] m27_8;
   assign m27_8 =15'b0;

   // m27_9 = W*in
   wire signed [14:0] m27_9;
   assign m27_9 =15'b0;

   // m27_10 = W*in
   wire signed [14:0] m27_10;
   assign m27_10 =15'b0;

   // m27_11 = W*in
   wire signed [14:0] m27_11;
   assign m27_11 ={ {3{neg27[14]}} , neg27[14:3] };

   // m27_12 = W*in
   wire signed [14:0] m27_12;
   assign m27_12 =15'b0;

   // m27_13 = W*in
   wire signed [14:0] m27_13;
   assign m27_13 =15'b0;

   // m27_14 = W*in
   wire signed [14:0] m27_14;
   assign m27_14 =15'b0;

   // m27_15 = W*in
   wire signed [14:0] m27_15;
   assign m27_15 =15'b0;

   // m27_16 = W*in
   wire signed [14:0] m27_16;
   assign m27_16 =15'b0;

   // m27_17 = W*in
   wire signed [14:0] m27_17;
   assign m27_17 =15'b0;

   // m27_18 = W*in
   wire signed [14:0] m27_18;
   assign m27_18 =15'b0;

   // m27_19 = W*in
   wire signed [14:0] m27_19;
   assign m27_19 =15'b0;

   // m27_20 = W*in
   wire signed [14:0] m27_20;
   assign m27_20 =15'b0;

   // m27_21 = W*in
   wire signed [14:0] m27_21;
   assign m27_21 ={ {4{in27[14]}} , in27[14:4] };

   // m27_22 = W*in
   wire signed [14:0] m27_22;
   assign m27_22 =15'b0;

   // m27_23 = W*in
   wire signed [14:0] m27_23;
   assign m27_23 =15'b0;

   // m27_24 = W*in
   wire signed [14:0] m27_24;
   assign m27_24 =15'b0;

   // m27_25 = W*in
   wire signed [14:0] m27_25;
   assign m27_25 =15'b0;

   // m27_26 = W*in
   wire signed [14:0] m27_26;
   assign m27_26 =15'b0;

   // m27_27 = W*in
   wire signed [14:0] m27_27;
   assign m27_27 =15'b0;

   // m27_28 = W*in
   wire signed [14:0] m27_28;
   assign m27_28 =15'b0;

   // m27_29 = W*in
   wire signed [14:0] m27_29;
   assign m27_29 =15'b0;

   // m27_30 = W*in
   wire signed [14:0] m27_30;
   assign m27_30 ={ {4{neg27[14]}} , neg27[14:4] };

   // m27_31 = W*in
   wire signed [14:0] m27_31;
   assign m27_31 =15'b0;

   // m27_32 = W*in
   wire signed [14:0] m27_32;
   assign m27_32 =15'b0;

   // m27_33 = W*in
   wire signed [14:0] m27_33;
   assign m27_33 =15'b0;

   // m27_34 = W*in
   wire signed [14:0] m27_34;
   assign m27_34 =15'b0;

   // m27_35 = W*in
   wire signed [14:0] m27_35;
   assign m27_35 =15'b0;

   // m27_36 = W*in
   wire signed [14:0] m27_36;
   assign m27_36 =15'b0;

   // m27_37 = W*in
   wire signed [14:0] m27_37;
   assign m27_37 =15'b0;

   // m27_38 = W*in
   wire signed [14:0] m27_38;
   assign m27_38 =15'b0;

   // m27_39 = W*in
   wire signed [14:0] m27_39;
   assign m27_39 =15'b0;

   // m27_40 = W*in
   wire signed [14:0] m27_40;
   assign m27_40 =15'b0;

   // m27_41 = W*in
   wire signed [14:0] m27_41;
   assign m27_41 =15'b0;

   // m27_42 = W*in
   wire signed [14:0] m27_42;
   assign m27_42 =15'b0;

   // m27_43 = W*in
   wire signed [14:0] m27_43;
   assign m27_43 =15'b0;

   // m27_44 = W*in
   wire signed [14:0] m27_44;
   assign m27_44 =15'b0;

   // m27_45 = W*in
   wire signed [14:0] m27_45;
   assign m27_45 =15'b0;

   // m27_46 = W*in
   wire signed [14:0] m27_46;
   assign m27_46 ={ {4{in27[14]}} , in27[14:4] };

   // m27_47 = W*in
   wire signed [14:0] m27_47;
   assign m27_47 =15'b0;

   // m27_48 = W*in
   wire signed [14:0] m27_48;
   assign m27_48 =15'b0;

   // m27_49 = W*in
   wire signed [14:0] m27_49;
   assign m27_49 =15'b0;

   // m27_50 = W*in
   wire signed [14:0] m27_50;
   assign m27_50 =15'b0;

   // m27_51 = W*in
   wire signed [14:0] m27_51;
   assign m27_51 =15'b0;

   // m27_52 = W*in
   wire signed [14:0] m27_52;
   assign m27_52 =15'b0;

   // m27_53 = W*in
   wire signed [14:0] m27_53;
   assign m27_53 =15'b0;

   // m27_54 = W*in
   wire signed [14:0] m27_54;
   assign m27_54 =15'b0;

   // m27_55 = W*in
   wire signed [14:0] m27_55;
   assign m27_55 =15'b0;

   // m27_56 = W*in
   wire signed [14:0] m27_56;
   assign m27_56 =15'b0;

   // m27_57 = W*in
   wire signed [14:0] m27_57;
   assign m27_57 =15'b0;

   // m27_58 = W*in
   wire signed [14:0] m27_58;
   assign m27_58 =15'b0;

   // m27_59 = W*in
   wire signed [14:0] m27_59;
   assign m27_59 =15'b0;

   // m27_60 = W*in
   wire signed [14:0] m27_60;
   assign m27_60 =15'b0;

   // m27_61 = W*in
   wire signed [14:0] m27_61;
   assign m27_61 =15'b0;

   // m27_62 = W*in
   wire signed [14:0] m27_62;
   assign m27_62 =15'b0;

   // m27_63 = W*in
   wire signed [14:0] m27_63;
   assign m27_63 =15'b0;

   // m27_64 = W*in
   wire signed [14:0] m27_64;
   assign m27_64 =15'b0;

   // m27_65 = W*in
   wire signed [14:0] m27_65;
   assign m27_65 =15'b0;

   // m27_66 = W*in
   wire signed [14:0] m27_66;
   assign m27_66 =15'b0;

   // m27_67 = W*in
   wire signed [14:0] m27_67;
   assign m27_67 =15'b0;

   // m27_68 = W*in
   wire signed [14:0] m27_68;
   assign m27_68 ={ {4{neg27[14]}} , neg27[14:4] };

   // m27_69 = W*in
   wire signed [14:0] m27_69;
   assign m27_69 =15'b0;

   // m27_70 = W*in
   wire signed [14:0] m27_70;
   assign m27_70 =15'b0;

   // m27_71 = W*in
   wire signed [14:0] m27_71;
   assign m27_71 =15'b0;

   // m27_72 = W*in
   wire signed [14:0] m27_72;
   assign m27_72 =15'b0;

   // m27_73 = W*in
   wire signed [14:0] m27_73;
   assign m27_73 =15'b0;

   // m27_74 = W*in
   wire signed [14:0] m27_74;
   assign m27_74 ={ {2{in27[14]}} , in27[14:2] };

   // m27_75 = W*in
   wire signed [14:0] m27_75;
   assign m27_75 =15'b0;

   // m27_76 = W*in
   wire signed [14:0] m27_76;
   assign m27_76 =15'b0;

   // m27_77 = W*in
   wire signed [14:0] m27_77;
   assign m27_77 =15'b0;

   // m27_78 = W*in
   wire signed [14:0] m27_78;
   assign m27_78 =15'b0;

   // m27_79 = W*in
   wire signed [14:0] m27_79;
   assign m27_79 =15'b0;

   // m27_80 = W*in
   wire signed [14:0] m27_80;
   assign m27_80 =15'b0;

   // m27_81 = W*in
   wire signed [14:0] m27_81;
   assign m27_81 ={ {3{in27[14]}} , in27[14:3] };

   // m27_82 = W*in
   wire signed [14:0] m27_82;
   assign m27_82 =15'b0;

   // m27_83 = W*in
   wire signed [14:0] m27_83;
   assign m27_83 =15'b0;

   // m27_84 = W*in
   wire signed [14:0] m27_84;
   assign m27_84 =15'b0;

   // m27_85 = W*in
   wire signed [14:0] m27_85;
   assign m27_85 =15'b0;

   // m27_86 = W*in
   wire signed [14:0] m27_86;
   assign m27_86 =15'b0;

   // m27_87 = W*in
   wire signed [14:0] m27_87;
   assign m27_87 =15'b0;

   // m27_88 = W*in
   wire signed [14:0] m27_88;
   assign m27_88 =15'b0;

   // m27_89 = W*in
   wire signed [14:0] m27_89;
   assign m27_89 =15'b0;

   // m27_90 = W*in
   wire signed [14:0] m27_90;
   assign m27_90 =15'b0;

   // m27_91 = W*in
   wire signed [14:0] m27_91;
   assign m27_91 =15'b0;

   // m27_92 = W*in
   wire signed [14:0] m27_92;
   assign m27_92 ={ {3{in27[14]}} , in27[14:3] };

   // m27_93 = W*in
   wire signed [14:0] m27_93;
   assign m27_93 =15'b0;

   // m27_94 = W*in
   wire signed [14:0] m27_94;
   assign m27_94 =15'b0;

   // m27_95 = W*in
   wire signed [14:0] m27_95;
   assign m27_95 =15'b0;

   // m27_96 = W*in
   wire signed [14:0] m27_96;
   assign m27_96 =15'b0;

   // m27_97 = W*in
   wire signed [14:0] m27_97;
   assign m27_97 =15'b0;

   // m27_98 = W*in
   wire signed [14:0] m27_98;
   assign m27_98 =15'b0;

   // m27_99 = W*in
   wire signed [14:0] m27_99;
   assign m27_99 =15'b0;

   // m27_100 = W*in
   wire signed [14:0] m27_100;
   assign m27_100 =15'b0;

   // m28_1 = W*in
   wire signed [14:0] m28_1;
   assign m28_1 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_2 = W*in
   wire signed [14:0] m28_2;
   assign m28_2 =15'b0;

   // m28_3 = W*in
   wire signed [14:0] m28_3;
   assign m28_3 =15'b0;

   // m28_4 = W*in
   wire signed [14:0] m28_4;
   assign m28_4 =15'b0;

   // m28_5 = W*in
   wire signed [14:0] m28_5;
   assign m28_5 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_6 = W*in
   wire signed [14:0] m28_6;
   assign m28_6 =15'b0;

   // m28_7 = W*in
   wire signed [14:0] m28_7;
   assign m28_7 =15'b0;

   // m28_8 = W*in
   wire signed [14:0] m28_8;
   assign m28_8 =15'b0;

   // m28_9 = W*in
   wire signed [14:0] m28_9;
   assign m28_9 ={ {3{in28[14]}} , in28[14:3] };

   // m28_10 = W*in
   wire signed [14:0] m28_10;
   assign m28_10 =15'b0;

   // m28_11 = W*in
   wire signed [14:0] m28_11;
   assign m28_11 =15'b0;

   // m28_12 = W*in
   wire signed [14:0] m28_12;
   assign m28_12 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_13 = W*in
   wire signed [14:0] m28_13;
   assign m28_13 =15'b0;

   // m28_14 = W*in
   wire signed [14:0] m28_14;
   assign m28_14 =15'b0;

   // m28_15 = W*in
   wire signed [14:0] m28_15;
   assign m28_15 =15'b0;

   // m28_16 = W*in
   wire signed [14:0] m28_16;
   assign m28_16 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_17 = W*in
   wire signed [14:0] m28_17;
   assign m28_17 ={ {3{in28[14]}} , in28[14:3] };

   // m28_18 = W*in
   wire signed [14:0] m28_18;
   assign m28_18 ={ {4{in28[14]}} , in28[14:4] };

   // m28_19 = W*in
   wire signed [14:0] m28_19;
   assign m28_19 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_20 = W*in
   wire signed [14:0] m28_20;
   assign m28_20 =15'b0;

   // m28_21 = W*in
   wire signed [14:0] m28_21;
   assign m28_21 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_22 = W*in
   wire signed [14:0] m28_22;
   assign m28_22 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_23 = W*in
   wire signed [14:0] m28_23;
   assign m28_23 =15'b0;

   // m28_24 = W*in
   wire signed [14:0] m28_24;
   assign m28_24 =15'b0;

   // m28_25 = W*in
   wire signed [14:0] m28_25;
   assign m28_25 =15'b0;

   // m28_26 = W*in
   wire signed [14:0] m28_26;
   assign m28_26 =15'b0;

   // m28_27 = W*in
   wire signed [14:0] m28_27;
   assign m28_27 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_28 = W*in
   wire signed [14:0] m28_28;
   assign m28_28 =15'b0;

   // m28_29 = W*in
   wire signed [14:0] m28_29;
   assign m28_29 =15'b0;

   // m28_30 = W*in
   wire signed [14:0] m28_30;
   assign m28_30 =15'b0;

   // m28_31 = W*in
   wire signed [14:0] m28_31;
   assign m28_31 =15'b0;

   // m28_32 = W*in
   wire signed [14:0] m28_32;
   assign m28_32 =15'b0;

   // m28_33 = W*in
   wire signed [14:0] m28_33;
   assign m28_33 ={ {3{in28[14]}} , in28[14:3] };

   // m28_34 = W*in
   wire signed [14:0] m28_34;
   assign m28_34 =15'b0;

   // m28_35 = W*in
   wire signed [14:0] m28_35;
   assign m28_35 =15'b0;

   // m28_36 = W*in
   wire signed [14:0] m28_36;
   assign m28_36 =15'b0;

   // m28_37 = W*in
   wire signed [14:0] m28_37;
   assign m28_37 =15'b0;

   // m28_38 = W*in
   wire signed [14:0] m28_38;
   assign m28_38 =15'b0;

   // m28_39 = W*in
   wire signed [14:0] m28_39;
   assign m28_39 =15'b0;

   // m28_40 = W*in
   wire signed [14:0] m28_40;
   assign m28_40 =15'b0;

   // m28_41 = W*in
   wire signed [14:0] m28_41;
   assign m28_41 =15'b0;

   // m28_42 = W*in
   wire signed [14:0] m28_42;
   assign m28_42 =15'b0;

   // m28_43 = W*in
   wire signed [14:0] m28_43;
   assign m28_43 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_44 = W*in
   wire signed [14:0] m28_44;
   assign m28_44 =15'b0;

   // m28_45 = W*in
   wire signed [14:0] m28_45;
   assign m28_45 =15'b0;

   // m28_46 = W*in
   wire signed [14:0] m28_46;
   assign m28_46 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_47 = W*in
   wire signed [14:0] m28_47;
   assign m28_47 =15'b0;

   // m28_48 = W*in
   wire signed [14:0] m28_48;
   assign m28_48 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_49 = W*in
   wire signed [14:0] m28_49;
   assign m28_49 =15'b0;

   // m28_50 = W*in
   wire signed [14:0] m28_50;
   assign m28_50 =15'b0;

   // m28_51 = W*in
   wire signed [14:0] m28_51;
   assign m28_51 =15'b0;

   // m28_52 = W*in
   wire signed [14:0] m28_52;
   assign m28_52 =15'b0;

   // m28_53 = W*in
   wire signed [14:0] m28_53;
   assign m28_53 =15'b0;

   // m28_54 = W*in
   wire signed [14:0] m28_54;
   assign m28_54 =15'b0;

   // m28_55 = W*in
   wire signed [14:0] m28_55;
   assign m28_55 =15'b0;

   // m28_56 = W*in
   wire signed [14:0] m28_56;
   assign m28_56 =15'b0;

   // m28_57 = W*in
   wire signed [14:0] m28_57;
   assign m28_57 ={ {3{in28[14]}} , in28[14:3] };

   // m28_58 = W*in
   wire signed [14:0] m28_58;
   assign m28_58 =15'b0;

   // m28_59 = W*in
   wire signed [14:0] m28_59;
   assign m28_59 =15'b0;

   // m28_60 = W*in
   wire signed [14:0] m28_60;
   assign m28_60 =15'b0;

   // m28_61 = W*in
   wire signed [14:0] m28_61;
   assign m28_61 ={ {4{neg28[14]}} , neg28[14:4] };

   // m28_62 = W*in
   wire signed [14:0] m28_62;
   assign m28_62 =15'b0;

   // m28_63 = W*in
   wire signed [14:0] m28_63;
   assign m28_63 =15'b0;

   // m28_64 = W*in
   wire signed [14:0] m28_64;
   assign m28_64 =15'b0;

   // m28_65 = W*in
   wire signed [14:0] m28_65;
   assign m28_65 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_66 = W*in
   wire signed [14:0] m28_66;
   assign m28_66 =15'b0;

   // m28_67 = W*in
   wire signed [14:0] m28_67;
   assign m28_67 =15'b0;

   // m28_68 = W*in
   wire signed [14:0] m28_68;
   assign m28_68 =15'b0;

   // m28_69 = W*in
   wire signed [14:0] m28_69;
   assign m28_69 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_70 = W*in
   wire signed [14:0] m28_70;
   assign m28_70 ={ {2{in28[14]}} , in28[14:2] };

   // m28_71 = W*in
   wire signed [14:0] m28_71;
   assign m28_71 =15'b0;

   // m28_72 = W*in
   wire signed [14:0] m28_72;
   assign m28_72 =15'b0;

   // m28_73 = W*in
   wire signed [14:0] m28_73;
   assign m28_73 =15'b0;

   // m28_74 = W*in
   wire signed [14:0] m28_74;
   assign m28_74 =15'b0;

   // m28_75 = W*in
   wire signed [14:0] m28_75;
   assign m28_75 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_76 = W*in
   wire signed [14:0] m28_76;
   assign m28_76 =15'b0;

   // m28_77 = W*in
   wire signed [14:0] m28_77;
   assign m28_77 =15'b0;

   // m28_78 = W*in
   wire signed [14:0] m28_78;
   assign m28_78 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_79 = W*in
   wire signed [14:0] m28_79;
   assign m28_79 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_80 = W*in
   wire signed [14:0] m28_80;
   assign m28_80 =15'b0;

   // m28_81 = W*in
   wire signed [14:0] m28_81;
   assign m28_81 ={ {3{in28[14]}} , in28[14:3] };

   // m28_82 = W*in
   wire signed [14:0] m28_82;
   assign m28_82 =15'b0;

   // m28_83 = W*in
   wire signed [14:0] m28_83;
   assign m28_83 =15'b0;

   // m28_84 = W*in
   wire signed [14:0] m28_84;
   assign m28_84 =15'b0;

   // m28_85 = W*in
   wire signed [14:0] m28_85;
   assign m28_85 =15'b0;

   // m28_86 = W*in
   wire signed [14:0] m28_86;
   assign m28_86 ={ {3{in28[14]}} , in28[14:3] };

   // m28_87 = W*in
   wire signed [14:0] m28_87;
   assign m28_87 =15'b0;

   // m28_88 = W*in
   wire signed [14:0] m28_88;
   assign m28_88 =15'b0;

   // m28_89 = W*in
   wire signed [14:0] m28_89;
   assign m28_89 =15'b0;

   // m28_90 = W*in
   wire signed [14:0] m28_90;
   assign m28_90 =15'b0;

   // m28_91 = W*in
   wire signed [14:0] m28_91;
   assign m28_91 =15'b0;

   // m28_92 = W*in
   wire signed [14:0] m28_92;
   assign m28_92 =15'b0;

   // m28_93 = W*in
   wire signed [14:0] m28_93;
   assign m28_93 =15'b0;

   // m28_94 = W*in
   wire signed [14:0] m28_94;
   assign m28_94 =15'b0;

   // m28_95 = W*in
   wire signed [14:0] m28_95;
   assign m28_95 =15'b0;

   // m28_96 = W*in
   wire signed [14:0] m28_96;
   assign m28_96 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_97 = W*in
   wire signed [14:0] m28_97;
   assign m28_97 ={ {3{neg28[14]}} , neg28[14:3] };

   // m28_98 = W*in
   wire signed [14:0] m28_98;
   assign m28_98 =15'b0;

   // m28_99 = W*in
   wire signed [14:0] m28_99;
   assign m28_99 =15'b0;

   // m28_100 = W*in
   wire signed [14:0] m28_100;
   assign m28_100 =15'b0;

   // m29_1 = W*in
   wire signed [14:0] m29_1;
   assign m29_1 =15'b0;

   // m29_2 = W*in
   wire signed [14:0] m29_2;
   assign m29_2 =15'b0;

   // m29_3 = W*in
   wire signed [14:0] m29_3;
   assign m29_3 =15'b0;

   // m29_4 = W*in
   wire signed [14:0] m29_4;
   assign m29_4 =15'b0;

   // m29_5 = W*in
   wire signed [14:0] m29_5;
   assign m29_5 =15'b0;

   // m29_6 = W*in
   wire signed [14:0] m29_6;
   assign m29_6 =15'b0;

   // m29_7 = W*in
   wire signed [14:0] m29_7;
   assign m29_7 =15'b0;

   // m29_8 = W*in
   wire signed [14:0] m29_8;
   assign m29_8 =15'b0;

   // m29_9 = W*in
   wire signed [14:0] m29_9;
   assign m29_9 =15'b0;

   // m29_10 = W*in
   wire signed [14:0] m29_10;
   assign m29_10 =15'b0;

   // m29_11 = W*in
   wire signed [14:0] m29_11;
   assign m29_11 =15'b0;

   // m29_12 = W*in
   wire signed [14:0] m29_12;
   assign m29_12 =15'b0;

   // m29_13 = W*in
   wire signed [14:0] m29_13;
   assign m29_13 ={ {4{in29[14]}} , in29[14:4] };

   // m29_14 = W*in
   wire signed [14:0] m29_14;
   assign m29_14 =15'b0;

   // m29_15 = W*in
   wire signed [14:0] m29_15;
   assign m29_15 =15'b0;

   // m29_16 = W*in
   wire signed [14:0] m29_16;
   assign m29_16 =15'b0;

   // m29_17 = W*in
   wire signed [14:0] m29_17;
   assign m29_17 =15'b0;

   // m29_18 = W*in
   wire signed [14:0] m29_18;
   assign m29_18 =15'b0;

   // m29_19 = W*in
   wire signed [14:0] m29_19;
   assign m29_19 =15'b0;

   // m29_20 = W*in
   wire signed [14:0] m29_20;
   assign m29_20 =15'b0;

   // m29_21 = W*in
   wire signed [14:0] m29_21;
   assign m29_21 =15'b0;

   // m29_22 = W*in
   wire signed [14:0] m29_22;
   assign m29_22 =15'b0;

   // m29_23 = W*in
   wire signed [14:0] m29_23;
   assign m29_23 =15'b0;

   // m29_24 = W*in
   wire signed [14:0] m29_24;
   assign m29_24 =15'b0;

   // m29_25 = W*in
   wire signed [14:0] m29_25;
   assign m29_25 =15'b0;

   // m29_26 = W*in
   wire signed [14:0] m29_26;
   assign m29_26 =15'b0;

   // m29_27 = W*in
   wire signed [14:0] m29_27;
   assign m29_27 =15'b0;

   // m29_28 = W*in
   wire signed [14:0] m29_28;
   assign m29_28 =15'b0;

   // m29_29 = W*in
   wire signed [14:0] m29_29;
   assign m29_29 =15'b0;

   // m29_30 = W*in
   wire signed [14:0] m29_30;
   assign m29_30 =15'b0;

   // m29_31 = W*in
   wire signed [14:0] m29_31;
   assign m29_31 =15'b0;

   // m29_32 = W*in
   wire signed [14:0] m29_32;
   assign m29_32 =15'b0;

   // m29_33 = W*in
   wire signed [14:0] m29_33;
   assign m29_33 =15'b0;

   // m29_34 = W*in
   wire signed [14:0] m29_34;
   assign m29_34 =15'b0;

   // m29_35 = W*in
   wire signed [14:0] m29_35;
   assign m29_35 =15'b0;

   // m29_36 = W*in
   wire signed [14:0] m29_36;
   assign m29_36 =15'b0;

   // m29_37 = W*in
   wire signed [14:0] m29_37;
   assign m29_37 =15'b0;

   // m29_38 = W*in
   wire signed [14:0] m29_38;
   assign m29_38 =15'b0;

   // m29_39 = W*in
   wire signed [14:0] m29_39;
   assign m29_39 =15'b0;

   // m29_40 = W*in
   wire signed [14:0] m29_40;
   assign m29_40 =15'b0;

   // m29_41 = W*in
   wire signed [14:0] m29_41;
   assign m29_41 ={ {4{in29[14]}} , in29[14:4] };

   // m29_42 = W*in
   wire signed [14:0] m29_42;
   assign m29_42 =15'b0;

   // m29_43 = W*in
   wire signed [14:0] m29_43;
   assign m29_43 =15'b0;

   // m29_44 = W*in
   wire signed [14:0] m29_44;
   assign m29_44 =15'b0;

   // m29_45 = W*in
   wire signed [14:0] m29_45;
   assign m29_45 =15'b0;

   // m29_46 = W*in
   wire signed [14:0] m29_46;
   assign m29_46 =15'b0;

   // m29_47 = W*in
   wire signed [14:0] m29_47;
   assign m29_47 =15'b0;

   // m29_48 = W*in
   wire signed [14:0] m29_48;
   assign m29_48 =15'b0;

   // m29_49 = W*in
   wire signed [14:0] m29_49;
   assign m29_49 =15'b0;

   // m29_50 = W*in
   wire signed [14:0] m29_50;
   assign m29_50 ={ {4{neg29[14]}} , neg29[14:4] };

   // m29_51 = W*in
   wire signed [14:0] m29_51;
   assign m29_51 =15'b0;

   // m29_52 = W*in
   wire signed [14:0] m29_52;
   assign m29_52 =15'b0;

   // m29_53 = W*in
   wire signed [14:0] m29_53;
   assign m29_53 =15'b0;

   // m29_54 = W*in
   wire signed [14:0] m29_54;
   assign m29_54 =15'b0;

   // m29_55 = W*in
   wire signed [14:0] m29_55;
   assign m29_55 ={ {4{in29[14]}} , in29[14:4] };

   // m29_56 = W*in
   wire signed [14:0] m29_56;
   assign m29_56 =15'b0;

   // m29_57 = W*in
   wire signed [14:0] m29_57;
   assign m29_57 =15'b0;

   // m29_58 = W*in
   wire signed [14:0] m29_58;
   assign m29_58 =15'b0;

   // m29_59 = W*in
   wire signed [14:0] m29_59;
   assign m29_59 =15'b0;

   // m29_60 = W*in
   wire signed [14:0] m29_60;
   assign m29_60 =15'b0;

   // m29_61 = W*in
   wire signed [14:0] m29_61;
   assign m29_61 =15'b0;

   // m29_62 = W*in
   wire signed [14:0] m29_62;
   assign m29_62 =15'b0;

   // m29_63 = W*in
   wire signed [14:0] m29_63;
   assign m29_63 =15'b0;

   // m29_64 = W*in
   wire signed [14:0] m29_64;
   assign m29_64 =15'b0;

   // m29_65 = W*in
   wire signed [14:0] m29_65;
   assign m29_65 =15'b0;

   // m29_66 = W*in
   wire signed [14:0] m29_66;
   assign m29_66 ={ {4{neg29[14]}} , neg29[14:4] };

   // m29_67 = W*in
   wire signed [14:0] m29_67;
   assign m29_67 =15'b0;

   // m29_68 = W*in
   wire signed [14:0] m29_68;
   assign m29_68 =15'b0;

   // m29_69 = W*in
   wire signed [14:0] m29_69;
   assign m29_69 =15'b0;

   // m29_70 = W*in
   wire signed [14:0] m29_70;
   assign m29_70 =15'b0;

   // m29_71 = W*in
   wire signed [14:0] m29_71;
   assign m29_71 =15'b0;

   // m29_72 = W*in
   wire signed [14:0] m29_72;
   assign m29_72 =15'b0;

   // m29_73 = W*in
   wire signed [14:0] m29_73;
   assign m29_73 =15'b0;

   // m29_74 = W*in
   wire signed [14:0] m29_74;
   assign m29_74 ={ {4{neg29[14]}} , neg29[14:4] };

   // m29_75 = W*in
   wire signed [14:0] m29_75;
   assign m29_75 =15'b0;

   // m29_76 = W*in
   wire signed [14:0] m29_76;
   assign m29_76 ={ {3{neg29[14]}} , neg29[14:3] };

   // m29_77 = W*in
   wire signed [14:0] m29_77;
   assign m29_77 =15'b0;

   // m29_78 = W*in
   wire signed [14:0] m29_78;
   assign m29_78 =15'b0;

   // m29_79 = W*in
   wire signed [14:0] m29_79;
   assign m29_79 =15'b0;

   // m29_80 = W*in
   wire signed [14:0] m29_80;
   assign m29_80 =15'b0;

   // m29_81 = W*in
   wire signed [14:0] m29_81;
   assign m29_81 ={ {4{in29[14]}} , in29[14:4] };

   // m29_82 = W*in
   wire signed [14:0] m29_82;
   assign m29_82 =15'b0;

   // m29_83 = W*in
   wire signed [14:0] m29_83;
   assign m29_83 =15'b0;

   // m29_84 = W*in
   wire signed [14:0] m29_84;
   assign m29_84 =15'b0;

   // m29_85 = W*in
   wire signed [14:0] m29_85;
   assign m29_85 =15'b0;

   // m29_86 = W*in
   wire signed [14:0] m29_86;
   assign m29_86 =15'b0;

   // m29_87 = W*in
   wire signed [14:0] m29_87;
   assign m29_87 =15'b0;

   // m29_88 = W*in
   wire signed [14:0] m29_88;
   assign m29_88 =15'b0;

   // m29_89 = W*in
   wire signed [14:0] m29_89;
   assign m29_89 =15'b0;

   // m29_90 = W*in
   wire signed [14:0] m29_90;
   assign m29_90 =15'b0;

   // m29_91 = W*in
   wire signed [14:0] m29_91;
   assign m29_91 =15'b0;

   // m29_92 = W*in
   wire signed [14:0] m29_92;
   assign m29_92 =15'b0;

   // m29_93 = W*in
   wire signed [14:0] m29_93;
   assign m29_93 ={ {3{neg29[14]}} , neg29[14:3] };

   // m29_94 = W*in
   wire signed [14:0] m29_94;
   assign m29_94 ={ {4{neg29[14]}} , neg29[14:4] };

   // m29_95 = W*in
   wire signed [14:0] m29_95;
   assign m29_95 =15'b0;

   // m29_96 = W*in
   wire signed [14:0] m29_96;
   assign m29_96 =15'b0;

   // m29_97 = W*in
   wire signed [14:0] m29_97;
   assign m29_97 =15'b0;

   // m29_98 = W*in
   wire signed [14:0] m29_98;
   assign m29_98 ={ {4{neg29[14]}} , neg29[14:4] };

   // m29_99 = W*in
   wire signed [14:0] m29_99;
   assign m29_99 =15'b0;

   // m29_100 = W*in
   wire signed [14:0] m29_100;
   assign m29_100 =15'b0;

   // m30_1 = W*in
   wire signed [14:0] m30_1;
   assign m30_1 =15'b0;

   // m30_2 = W*in
   wire signed [14:0] m30_2;
   assign m30_2 =15'b0;

   // m30_3 = W*in
   wire signed [14:0] m30_3;
   assign m30_3 ={ {3{in30[14]}} , in30[14:3] };

   // m30_4 = W*in
   wire signed [14:0] m30_4;
   assign m30_4 =15'b0;

   // m30_5 = W*in
   wire signed [14:0] m30_5;
   assign m30_5 =15'b0;

   // m30_6 = W*in
   wire signed [14:0] m30_6;
   assign m30_6 =15'b0;

   // m30_7 = W*in
   wire signed [14:0] m30_7;
   assign m30_7 =15'b0;

   // m30_8 = W*in
   wire signed [14:0] m30_8;
   assign m30_8 ={ {3{in30[14]}} , in30[14:3] };

   // m30_9 = W*in
   wire signed [14:0] m30_9;
   assign m30_9 =15'b0;

   // m30_10 = W*in
   wire signed [14:0] m30_10;
   assign m30_10 =15'b0;

   // m30_11 = W*in
   wire signed [14:0] m30_11;
   assign m30_11 =15'b0;

   // m30_12 = W*in
   wire signed [14:0] m30_12;
   assign m30_12 =15'b0;

   // m30_13 = W*in
   wire signed [14:0] m30_13;
   assign m30_13 =15'b0;

   // m30_14 = W*in
   wire signed [14:0] m30_14;
   assign m30_14 =15'b0;

   // m30_15 = W*in
   wire signed [14:0] m30_15;
   assign m30_15 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_16 = W*in
   wire signed [14:0] m30_16;
   assign m30_16 =15'b0;

   // m30_17 = W*in
   wire signed [14:0] m30_17;
   assign m30_17 ={ {3{in30[14]}} , in30[14:3] };

   // m30_18 = W*in
   wire signed [14:0] m30_18;
   assign m30_18 =15'b0;

   // m30_19 = W*in
   wire signed [14:0] m30_19;
   assign m30_19 =15'b0;

   // m30_20 = W*in
   wire signed [14:0] m30_20;
   assign m30_20 =15'b0;

   // m30_21 = W*in
   wire signed [14:0] m30_21;
   assign m30_21 =15'b0;

   // m30_22 = W*in
   wire signed [14:0] m30_22;
   assign m30_22 =15'b0;

   // m30_23 = W*in
   wire signed [14:0] m30_23;
   assign m30_23 =15'b0;

   // m30_24 = W*in
   wire signed [14:0] m30_24;
   assign m30_24 =15'b0;

   // m30_25 = W*in
   wire signed [14:0] m30_25;
   assign m30_25 =15'b0;

   // m30_26 = W*in
   wire signed [14:0] m30_26;
   assign m30_26 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_27 = W*in
   wire signed [14:0] m30_27;
   assign m30_27 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_28 = W*in
   wire signed [14:0] m30_28;
   assign m30_28 =15'b0;

   // m30_29 = W*in
   wire signed [14:0] m30_29;
   assign m30_29 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_30 = W*in
   wire signed [14:0] m30_30;
   assign m30_30 =15'b0;

   // m30_31 = W*in
   wire signed [14:0] m30_31;
   assign m30_31 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_32 = W*in
   wire signed [14:0] m30_32;
   assign m30_32 =15'b0;

   // m30_33 = W*in
   wire signed [14:0] m30_33;
   assign m30_33 =15'b0;

   // m30_34 = W*in
   wire signed [14:0] m30_34;
   assign m30_34 =15'b0;

   // m30_35 = W*in
   wire signed [14:0] m30_35;
   assign m30_35 =15'b0;

   // m30_36 = W*in
   wire signed [14:0] m30_36;
   assign m30_36 =15'b0;

   // m30_37 = W*in
   wire signed [14:0] m30_37;
   assign m30_37 =15'b0;

   // m30_38 = W*in
   wire signed [14:0] m30_38;
   assign m30_38 =15'b0;

   // m30_39 = W*in
   wire signed [14:0] m30_39;
   assign m30_39 =15'b0;

   // m30_40 = W*in
   wire signed [14:0] m30_40;
   assign m30_40 =15'b0;

   // m30_41 = W*in
   wire signed [14:0] m30_41;
   assign m30_41 =15'b0;

   // m30_42 = W*in
   wire signed [14:0] m30_42;
   assign m30_42 =15'b0;

   // m30_43 = W*in
   wire signed [14:0] m30_43;
   assign m30_43 =15'b0;

   // m30_44 = W*in
   wire signed [14:0] m30_44;
   assign m30_44 ={ {3{in30[14]}} , in30[14:3] };

   // m30_45 = W*in
   wire signed [14:0] m30_45;
   assign m30_45 =15'b0;

   // m30_46 = W*in
   wire signed [14:0] m30_46;
   assign m30_46 =15'b0;

   // m30_47 = W*in
   wire signed [14:0] m30_47;
   assign m30_47 =15'b0;

   // m30_48 = W*in
   wire signed [14:0] m30_48;
   assign m30_48 =15'b0;

   // m30_49 = W*in
   wire signed [14:0] m30_49;
   assign m30_49 =15'b0;

   // m30_50 = W*in
   wire signed [14:0] m30_50;
   assign m30_50 =15'b0;

   // m30_51 = W*in
   wire signed [14:0] m30_51;
   assign m30_51 =15'b0;

   // m30_52 = W*in
   wire signed [14:0] m30_52;
   assign m30_52 =15'b0;

   // m30_53 = W*in
   wire signed [14:0] m30_53;
   assign m30_53 =15'b0;

   // m30_54 = W*in
   wire signed [14:0] m30_54;
   assign m30_54 =15'b0;

   // m30_55 = W*in
   wire signed [14:0] m30_55;
   assign m30_55 =15'b0;

   // m30_56 = W*in
   wire signed [14:0] m30_56;
   assign m30_56 =15'b0;

   // m30_57 = W*in
   wire signed [14:0] m30_57;
   assign m30_57 =15'b0;

   // m30_58 = W*in
   wire signed [14:0] m30_58;
   assign m30_58 =15'b0;

   // m30_59 = W*in
   wire signed [14:0] m30_59;
   assign m30_59 =15'b0;

   // m30_60 = W*in
   wire signed [14:0] m30_60;
   assign m30_60 ={ {4{neg30[14]}} , neg30[14:4] };

   // m30_61 = W*in
   wire signed [14:0] m30_61;
   assign m30_61 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_62 = W*in
   wire signed [14:0] m30_62;
   assign m30_62 =15'b0;

   // m30_63 = W*in
   wire signed [14:0] m30_63;
   assign m30_63 =15'b0;

   // m30_64 = W*in
   wire signed [14:0] m30_64;
   assign m30_64 =15'b0;

   // m30_65 = W*in
   wire signed [14:0] m30_65;
   assign m30_65 =15'b0;

   // m30_66 = W*in
   wire signed [14:0] m30_66;
   assign m30_66 =15'b0;

   // m30_67 = W*in
   wire signed [14:0] m30_67;
   assign m30_67 =15'b0;

   // m30_68 = W*in
   wire signed [14:0] m30_68;
   assign m30_68 =15'b0;

   // m30_69 = W*in
   wire signed [14:0] m30_69;
   assign m30_69 ={ {3{in30[14]}} , in30[14:3] };

   // m30_70 = W*in
   wire signed [14:0] m30_70;
   assign m30_70 ={ {3{in30[14]}} , in30[14:3] };

   // m30_71 = W*in
   wire signed [14:0] m30_71;
   assign m30_71 =15'b0;

   // m30_72 = W*in
   wire signed [14:0] m30_72;
   assign m30_72 =15'b0;

   // m30_73 = W*in
   wire signed [14:0] m30_73;
   assign m30_73 =15'b0;

   // m30_74 = W*in
   wire signed [14:0] m30_74;
   assign m30_74 ={ {3{in30[14]}} , in30[14:3] };

   // m30_75 = W*in
   wire signed [14:0] m30_75;
   assign m30_75 =15'b0;

   // m30_76 = W*in
   wire signed [14:0] m30_76;
   assign m30_76 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_77 = W*in
   wire signed [14:0] m30_77;
   assign m30_77 =15'b0;

   // m30_78 = W*in
   wire signed [14:0] m30_78;
   assign m30_78 ={ {4{neg30[14]}} , neg30[14:4] };

   // m30_79 = W*in
   wire signed [14:0] m30_79;
   assign m30_79 =15'b0;

   // m30_80 = W*in
   wire signed [14:0] m30_80;
   assign m30_80 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_81 = W*in
   wire signed [14:0] m30_81;
   assign m30_81 =15'b0;

   // m30_82 = W*in
   wire signed [14:0] m30_82;
   assign m30_82 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_83 = W*in
   wire signed [14:0] m30_83;
   assign m30_83 =15'b0;

   // m30_84 = W*in
   wire signed [14:0] m30_84;
   assign m30_84 =15'b0;

   // m30_85 = W*in
   wire signed [14:0] m30_85;
   assign m30_85 =15'b0;

   // m30_86 = W*in
   wire signed [14:0] m30_86;
   assign m30_86 ={ {3{neg30[14]}} , neg30[14:3] };

   // m30_87 = W*in
   wire signed [14:0] m30_87;
   assign m30_87 =15'b0;

   // m30_88 = W*in
   wire signed [14:0] m30_88;
   assign m30_88 =15'b0;

   // m30_89 = W*in
   wire signed [14:0] m30_89;
   assign m30_89 =15'b0;

   // m30_90 = W*in
   wire signed [14:0] m30_90;
   assign m30_90 =15'b0;

   // m30_91 = W*in
   wire signed [14:0] m30_91;
   assign m30_91 =15'b0;

   // m30_92 = W*in
   wire signed [14:0] m30_92;
   assign m30_92 =15'b0;

   // m30_93 = W*in
   wire signed [14:0] m30_93;
   assign m30_93 =15'b0;

   // m30_94 = W*in
   wire signed [14:0] m30_94;
   assign m30_94 =15'b0;

   // m30_95 = W*in
   wire signed [14:0] m30_95;
   assign m30_95 =15'b0;

   // m30_96 = W*in
   wire signed [14:0] m30_96;
   assign m30_96 =15'b0;

   // m30_97 = W*in
   wire signed [14:0] m30_97;
   assign m30_97 =15'b0;

   // m30_98 = W*in
   wire signed [14:0] m30_98;
   assign m30_98 =15'b0;

   // m30_99 = W*in
   wire signed [14:0] m30_99;
   assign m30_99 ={ {3{in30[14]}} , in30[14:3] };

   // m30_100 = W*in
   wire signed [14:0] m30_100;
   assign m30_100 =15'b0;

   // m31_1 = W*in
   wire signed [14:0] m31_1;
   assign m31_1 ={ {3{in31[14]}} , in31[14:3] };

   // m31_2 = W*in
   wire signed [14:0] m31_2;
   assign m31_2 =15'b0;

   // m31_3 = W*in
   wire signed [14:0] m31_3;
   assign m31_3 =15'b0;

   // m31_4 = W*in
   wire signed [14:0] m31_4;
   assign m31_4 =15'b0;

   // m31_5 = W*in
   wire signed [14:0] m31_5;
   assign m31_5 =15'b0;

   // m31_6 = W*in
   wire signed [14:0] m31_6;
   assign m31_6 =15'b0;

   // m31_7 = W*in
   wire signed [14:0] m31_7;
   assign m31_7 =15'b0;

   // m31_8 = W*in
   wire signed [14:0] m31_8;
   assign m31_8 =15'b0;

   // m31_9 = W*in
   wire signed [14:0] m31_9;
   assign m31_9 ={ {4{neg31[14]}} , neg31[14:4] };

   // m31_10 = W*in
   wire signed [14:0] m31_10;
   assign m31_10 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_11 = W*in
   wire signed [14:0] m31_11;
   assign m31_11 =15'b0;

   // m31_12 = W*in
   wire signed [14:0] m31_12;
   assign m31_12 =15'b0;

   // m31_13 = W*in
   wire signed [14:0] m31_13;
   assign m31_13 =15'b0;

   // m31_14 = W*in
   wire signed [14:0] m31_14;
   assign m31_14 =15'b0;

   // m31_15 = W*in
   wire signed [14:0] m31_15;
   assign m31_15 =15'b0;

   // m31_16 = W*in
   wire signed [14:0] m31_16;
   assign m31_16 =15'b0;

   // m31_17 = W*in
   wire signed [14:0] m31_17;
   assign m31_17 =15'b0;

   // m31_18 = W*in
   wire signed [14:0] m31_18;
   assign m31_18 =15'b0;

   // m31_19 = W*in
   wire signed [14:0] m31_19;
   assign m31_19 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_20 = W*in
   wire signed [14:0] m31_20;
   assign m31_20 =15'b0;

   // m31_21 = W*in
   wire signed [14:0] m31_21;
   assign m31_21 =15'b0;

   // m31_22 = W*in
   wire signed [14:0] m31_22;
   assign m31_22 =15'b0;

   // m31_23 = W*in
   wire signed [14:0] m31_23;
   assign m31_23 ={ {3{in31[14]}} , in31[14:3] };

   // m31_24 = W*in
   wire signed [14:0] m31_24;
   assign m31_24 =15'b0;

   // m31_25 = W*in
   wire signed [14:0] m31_25;
   assign m31_25 =15'b0;

   // m31_26 = W*in
   wire signed [14:0] m31_26;
   assign m31_26 =15'b0;

   // m31_27 = W*in
   wire signed [14:0] m31_27;
   assign m31_27 =15'b0;

   // m31_28 = W*in
   wire signed [14:0] m31_28;
   assign m31_28 =15'b0;

   // m31_29 = W*in
   wire signed [14:0] m31_29;
   assign m31_29 =15'b0;

   // m31_30 = W*in
   wire signed [14:0] m31_30;
   assign m31_30 ={ {3{in31[14]}} , in31[14:3] };

   // m31_31 = W*in
   wire signed [14:0] m31_31;
   assign m31_31 =15'b0;

   // m31_32 = W*in
   wire signed [14:0] m31_32;
   assign m31_32 =15'b0;

   // m31_33 = W*in
   wire signed [14:0] m31_33;
   assign m31_33 =15'b0;

   // m31_34 = W*in
   wire signed [14:0] m31_34;
   assign m31_34 =15'b0;

   // m31_35 = W*in
   wire signed [14:0] m31_35;
   assign m31_35 =15'b0;

   // m31_36 = W*in
   wire signed [14:0] m31_36;
   assign m31_36 =15'b0;

   // m31_37 = W*in
   wire signed [14:0] m31_37;
   assign m31_37 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_38 = W*in
   wire signed [14:0] m31_38;
   assign m31_38 =15'b0;

   // m31_39 = W*in
   wire signed [14:0] m31_39;
   assign m31_39 =15'b0;

   // m31_40 = W*in
   wire signed [14:0] m31_40;
   assign m31_40 =15'b0;

   // m31_41 = W*in
   wire signed [14:0] m31_41;
   assign m31_41 ={ {3{in31[14]}} , in31[14:3] };

   // m31_42 = W*in
   wire signed [14:0] m31_42;
   assign m31_42 =15'b0;

   // m31_43 = W*in
   wire signed [14:0] m31_43;
   assign m31_43 =15'b0;

   // m31_44 = W*in
   wire signed [14:0] m31_44;
   assign m31_44 =15'b0;

   // m31_45 = W*in
   wire signed [14:0] m31_45;
   assign m31_45 =15'b0;

   // m31_46 = W*in
   wire signed [14:0] m31_46;
   assign m31_46 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_47 = W*in
   wire signed [14:0] m31_47;
   assign m31_47 =15'b0;

   // m31_48 = W*in
   wire signed [14:0] m31_48;
   assign m31_48 =15'b0;

   // m31_49 = W*in
   wire signed [14:0] m31_49;
   assign m31_49 =15'b0;

   // m31_50 = W*in
   wire signed [14:0] m31_50;
   assign m31_50 =15'b0;

   // m31_51 = W*in
   wire signed [14:0] m31_51;
   assign m31_51 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_52 = W*in
   wire signed [14:0] m31_52;
   assign m31_52 =15'b0;

   // m31_53 = W*in
   wire signed [14:0] m31_53;
   assign m31_53 =15'b0;

   // m31_54 = W*in
   wire signed [14:0] m31_54;
   assign m31_54 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_55 = W*in
   wire signed [14:0] m31_55;
   assign m31_55 =15'b0;

   // m31_56 = W*in
   wire signed [14:0] m31_56;
   assign m31_56 =15'b0;

   // m31_57 = W*in
   wire signed [14:0] m31_57;
   assign m31_57 =15'b0;

   // m31_58 = W*in
   wire signed [14:0] m31_58;
   assign m31_58 ={ {4{neg31[14]}} , neg31[14:4] };

   // m31_59 = W*in
   wire signed [14:0] m31_59;
   assign m31_59 =15'b0;

   // m31_60 = W*in
   wire signed [14:0] m31_60;
   assign m31_60 =15'b0;

   // m31_61 = W*in
   wire signed [14:0] m31_61;
   assign m31_61 =15'b0;

   // m31_62 = W*in
   wire signed [14:0] m31_62;
   assign m31_62 =15'b0;

   // m31_63 = W*in
   wire signed [14:0] m31_63;
   assign m31_63 =15'b0;

   // m31_64 = W*in
   wire signed [14:0] m31_64;
   assign m31_64 ={ {4{in31[14]}} , in31[14:4] };

   // m31_65 = W*in
   wire signed [14:0] m31_65;
   assign m31_65 =15'b0;

   // m31_66 = W*in
   wire signed [14:0] m31_66;
   assign m31_66 =15'b0;

   // m31_67 = W*in
   wire signed [14:0] m31_67;
   assign m31_67 =15'b0;

   // m31_68 = W*in
   wire signed [14:0] m31_68;
   assign m31_68 =15'b0;

   // m31_69 = W*in
   wire signed [14:0] m31_69;
   assign m31_69 =15'b0;

   // m31_70 = W*in
   wire signed [14:0] m31_70;
   assign m31_70 =15'b0;

   // m31_71 = W*in
   wire signed [14:0] m31_71;
   assign m31_71 ={ {3{neg31[14]}} , neg31[14:3] };

   // m31_72 = W*in
   wire signed [14:0] m31_72;
   assign m31_72 =15'b0;

   // m31_73 = W*in
   wire signed [14:0] m31_73;
   assign m31_73 =15'b0;

   // m31_74 = W*in
   wire signed [14:0] m31_74;
   assign m31_74 =15'b0;

   // m31_75 = W*in
   wire signed [14:0] m31_75;
   assign m31_75 =15'b0;

   // m31_76 = W*in
   wire signed [14:0] m31_76;
   assign m31_76 =15'b0;

   // m31_77 = W*in
   wire signed [14:0] m31_77;
   assign m31_77 =15'b0;

   // m31_78 = W*in
   wire signed [14:0] m31_78;
   assign m31_78 =15'b0;

   // m31_79 = W*in
   wire signed [14:0] m31_79;
   assign m31_79 =15'b0;

   // m31_80 = W*in
   wire signed [14:0] m31_80;
   assign m31_80 =15'b0;

   // m31_81 = W*in
   wire signed [14:0] m31_81;
   assign m31_81 =15'b0;

   // m31_82 = W*in
   wire signed [14:0] m31_82;
   assign m31_82 =15'b0;

   // m31_83 = W*in
   wire signed [14:0] m31_83;
   assign m31_83 =15'b0;

   // m31_84 = W*in
   wire signed [14:0] m31_84;
   assign m31_84 =15'b0;

   // m31_85 = W*in
   wire signed [14:0] m31_85;
   assign m31_85 =15'b0;

   // m31_86 = W*in
   wire signed [14:0] m31_86;
   assign m31_86 =15'b0;

   // m31_87 = W*in
   wire signed [14:0] m31_87;
   assign m31_87 ={ {3{in31[14]}} , in31[14:3] };

   // m31_88 = W*in
   wire signed [14:0] m31_88;
   assign m31_88 =15'b0;

   // m31_89 = W*in
   wire signed [14:0] m31_89;
   assign m31_89 =15'b0;

   // m31_90 = W*in
   wire signed [14:0] m31_90;
   assign m31_90 =15'b0;

   // m31_91 = W*in
   wire signed [14:0] m31_91;
   assign m31_91 =15'b0;

   // m31_92 = W*in
   wire signed [14:0] m31_92;
   assign m31_92 =15'b0;

   // m31_93 = W*in
   wire signed [14:0] m31_93;
   assign m31_93 =15'b0;

   // m31_94 = W*in
   wire signed [14:0] m31_94;
   assign m31_94 =15'b0;

   // m31_95 = W*in
   wire signed [14:0] m31_95;
   assign m31_95 =15'b0;

   // m31_96 = W*in
   wire signed [14:0] m31_96;
   assign m31_96 ={ {3{in31[14]}} , in31[14:3] };

   // m31_97 = W*in
   wire signed [14:0] m31_97;
   assign m31_97 =15'b0;

   // m31_98 = W*in
   wire signed [14:0] m31_98;
   assign m31_98 =15'b0;

   // m31_99 = W*in
   wire signed [14:0] m31_99;
   assign m31_99 =15'b0;

   // m31_100 = W*in
   wire signed [14:0] m31_100;
   assign m31_100 =15'b0;

   // m32_1 = W*in
   wire signed [14:0] m32_1;
   assign m32_1 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_2 = W*in
   wire signed [14:0] m32_2;
   assign m32_2 =15'b0;

   // m32_3 = W*in
   wire signed [14:0] m32_3;
   assign m32_3 =15'b0;

   // m32_4 = W*in
   wire signed [14:0] m32_4;
   assign m32_4 =15'b0;

   // m32_5 = W*in
   wire signed [14:0] m32_5;
   assign m32_5 =15'b0;

   // m32_6 = W*in
   wire signed [14:0] m32_6;
   assign m32_6 =15'b0;

   // m32_7 = W*in
   wire signed [14:0] m32_7;
   assign m32_7 =15'b0;

   // m32_8 = W*in
   wire signed [14:0] m32_8;
   assign m32_8 =15'b0;

   // m32_9 = W*in
   wire signed [14:0] m32_9;
   assign m32_9 =15'b0;

   // m32_10 = W*in
   wire signed [14:0] m32_10;
   assign m32_10 =15'b0;

   // m32_11 = W*in
   wire signed [14:0] m32_11;
   assign m32_11 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_12 = W*in
   wire signed [14:0] m32_12;
   assign m32_12 =15'b0;

   // m32_13 = W*in
   wire signed [14:0] m32_13;
   assign m32_13 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_14 = W*in
   wire signed [14:0] m32_14;
   assign m32_14 =15'b0;

   // m32_15 = W*in
   wire signed [14:0] m32_15;
   assign m32_15 =15'b0;

   // m32_16 = W*in
   wire signed [14:0] m32_16;
   assign m32_16 =15'b0;

   // m32_17 = W*in
   wire signed [14:0] m32_17;
   assign m32_17 =15'b0;

   // m32_18 = W*in
   wire signed [14:0] m32_18;
   assign m32_18 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_19 = W*in
   wire signed [14:0] m32_19;
   assign m32_19 ={ {3{in32[14]}} , in32[14:3] };

   // m32_20 = W*in
   wire signed [14:0] m32_20;
   assign m32_20 ={ {4{neg32[14]}} , neg32[14:4] };

   // m32_21 = W*in
   wire signed [14:0] m32_21;
   assign m32_21 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_22 = W*in
   wire signed [14:0] m32_22;
   assign m32_22 =15'b0;

   // m32_23 = W*in
   wire signed [14:0] m32_23;
   assign m32_23 =15'b0;

   // m32_24 = W*in
   wire signed [14:0] m32_24;
   assign m32_24 ={ {3{in32[14]}} , in32[14:3] };

   // m32_25 = W*in
   wire signed [14:0] m32_25;
   assign m32_25 =15'b0;

   // m32_26 = W*in
   wire signed [14:0] m32_26;
   assign m32_26 ={ {3{in32[14]}} , in32[14:3] };

   // m32_27 = W*in
   wire signed [14:0] m32_27;
   assign m32_27 =15'b0;

   // m32_28 = W*in
   wire signed [14:0] m32_28;
   assign m32_28 =15'b0;

   // m32_29 = W*in
   wire signed [14:0] m32_29;
   assign m32_29 =15'b0;

   // m32_30 = W*in
   wire signed [14:0] m32_30;
   assign m32_30 =15'b0;

   // m32_31 = W*in
   wire signed [14:0] m32_31;
   assign m32_31 =15'b0;

   // m32_32 = W*in
   wire signed [14:0] m32_32;
   assign m32_32 ={ {3{in32[14]}} , in32[14:3] };

   // m32_33 = W*in
   wire signed [14:0] m32_33;
   assign m32_33 =15'b0;

   // m32_34 = W*in
   wire signed [14:0] m32_34;
   assign m32_34 =15'b0;

   // m32_35 = W*in
   wire signed [14:0] m32_35;
   assign m32_35 ={ {3{in32[14]}} , in32[14:3] };

   // m32_36 = W*in
   wire signed [14:0] m32_36;
   assign m32_36 =15'b0;

   // m32_37 = W*in
   wire signed [14:0] m32_37;
   assign m32_37 =15'b0;

   // m32_38 = W*in
   wire signed [14:0] m32_38;
   assign m32_38 =15'b0;

   // m32_39 = W*in
   wire signed [14:0] m32_39;
   assign m32_39 =15'b0;

   // m32_40 = W*in
   wire signed [14:0] m32_40;
   assign m32_40 ={ {3{in32[14]}} , in32[14:3] };

   // m32_41 = W*in
   wire signed [14:0] m32_41;
   assign m32_41 =15'b0;

   // m32_42 = W*in
   wire signed [14:0] m32_42;
   assign m32_42 ={ {2{in32[14]}} , in32[14:2] };

   // m32_43 = W*in
   wire signed [14:0] m32_43;
   assign m32_43 =15'b0;

   // m32_44 = W*in
   wire signed [14:0] m32_44;
   assign m32_44 =15'b0;

   // m32_45 = W*in
   wire signed [14:0] m32_45;
   assign m32_45 =15'b0;

   // m32_46 = W*in
   wire signed [14:0] m32_46;
   assign m32_46 =15'b0;

   // m32_47 = W*in
   wire signed [14:0] m32_47;
   assign m32_47 =15'b0;

   // m32_48 = W*in
   wire signed [14:0] m32_48;
   assign m32_48 =15'b0;

   // m32_49 = W*in
   wire signed [14:0] m32_49;
   assign m32_49 =15'b0;

   // m32_50 = W*in
   wire signed [14:0] m32_50;
   assign m32_50 =15'b0;

   // m32_51 = W*in
   wire signed [14:0] m32_51;
   assign m32_51 =15'b0;

   // m32_52 = W*in
   wire signed [14:0] m32_52;
   assign m32_52 =15'b0;

   // m32_53 = W*in
   wire signed [14:0] m32_53;
   assign m32_53 =15'b0;

   // m32_54 = W*in
   wire signed [14:0] m32_54;
   assign m32_54 =15'b0;

   // m32_55 = W*in
   wire signed [14:0] m32_55;
   assign m32_55 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_56 = W*in
   wire signed [14:0] m32_56;
   assign m32_56 =15'b0;

   // m32_57 = W*in
   wire signed [14:0] m32_57;
   assign m32_57 ={ {3{in32[14]}} , in32[14:3] };

   // m32_58 = W*in
   wire signed [14:0] m32_58;
   assign m32_58 =15'b0;

   // m32_59 = W*in
   wire signed [14:0] m32_59;
   assign m32_59 ={ {3{in32[14]}} , in32[14:3] };

   // m32_60 = W*in
   wire signed [14:0] m32_60;
   assign m32_60 =15'b0;

   // m32_61 = W*in
   wire signed [14:0] m32_61;
   assign m32_61 =15'b0;

   // m32_62 = W*in
   wire signed [14:0] m32_62;
   assign m32_62 =15'b0;

   // m32_63 = W*in
   wire signed [14:0] m32_63;
   assign m32_63 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_64 = W*in
   wire signed [14:0] m32_64;
   assign m32_64 ={ {4{neg32[14]}} , neg32[14:4] };

   // m32_65 = W*in
   wire signed [14:0] m32_65;
   assign m32_65 ={ {4{neg32[14]}} , neg32[14:4] };

   // m32_66 = W*in
   wire signed [14:0] m32_66;
   assign m32_66 ={ {3{in32[14]}} , in32[14:3] };

   // m32_67 = W*in
   wire signed [14:0] m32_67;
   assign m32_67 =15'b0;

   // m32_68 = W*in
   wire signed [14:0] m32_68;
   assign m32_68 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_69 = W*in
   wire signed [14:0] m32_69;
   assign m32_69 ={ {4{neg32[14]}} , neg32[14:4] };

   // m32_70 = W*in
   wire signed [14:0] m32_70;
   assign m32_70 ={ {3{in32[14]}} , in32[14:3] };

   // m32_71 = W*in
   wire signed [14:0] m32_71;
   assign m32_71 =15'b0;

   // m32_72 = W*in
   wire signed [14:0] m32_72;
   assign m32_72 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_73 = W*in
   wire signed [14:0] m32_73;
   assign m32_73 =15'b0;

   // m32_74 = W*in
   wire signed [14:0] m32_74;
   assign m32_74 =15'b0;

   // m32_75 = W*in
   wire signed [14:0] m32_75;
   assign m32_75 =15'b0;

   // m32_76 = W*in
   wire signed [14:0] m32_76;
   assign m32_76 =15'b0;

   // m32_77 = W*in
   wire signed [14:0] m32_77;
   assign m32_77 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_78 = W*in
   wire signed [14:0] m32_78;
   assign m32_78 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_79 = W*in
   wire signed [14:0] m32_79;
   assign m32_79 ={ {3{in32[14]}} , in32[14:3] };

   // m32_80 = W*in
   wire signed [14:0] m32_80;
   assign m32_80 =15'b0;

   // m32_81 = W*in
   wire signed [14:0] m32_81;
   assign m32_81 =15'b0;

   // m32_82 = W*in
   wire signed [14:0] m32_82;
   assign m32_82 =15'b0;

   // m32_83 = W*in
   wire signed [14:0] m32_83;
   assign m32_83 =15'b0;

   // m32_84 = W*in
   wire signed [14:0] m32_84;
   assign m32_84 =15'b0;

   // m32_85 = W*in
   wire signed [14:0] m32_85;
   assign m32_85 =15'b0;

   // m32_86 = W*in
   wire signed [14:0] m32_86;
   assign m32_86 =15'b0;

   // m32_87 = W*in
   wire signed [14:0] m32_87;
   assign m32_87 =15'b0;

   // m32_88 = W*in
   wire signed [14:0] m32_88;
   assign m32_88 =15'b0;

   // m32_89 = W*in
   wire signed [14:0] m32_89;
   assign m32_89 =15'b0;

   // m32_90 = W*in
   wire signed [14:0] m32_90;
   assign m32_90 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_91 = W*in
   wire signed [14:0] m32_91;
   assign m32_91 =15'b0;

   // m32_92 = W*in
   wire signed [14:0] m32_92;
   assign m32_92 =15'b0;

   // m32_93 = W*in
   wire signed [14:0] m32_93;
   assign m32_93 =15'b0;

   // m32_94 = W*in
   wire signed [14:0] m32_94;
   assign m32_94 =15'b0;

   // m32_95 = W*in
   wire signed [14:0] m32_95;
   assign m32_95 ={ {4{neg32[14]}} , neg32[14:4] };

   // m32_96 = W*in
   wire signed [14:0] m32_96;
   assign m32_96 =15'b0;

   // m32_97 = W*in
   wire signed [14:0] m32_97;
   assign m32_97 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_98 = W*in
   wire signed [14:0] m32_98;
   assign m32_98 =15'b0;

   // m32_99 = W*in
   wire signed [14:0] m32_99;
   assign m32_99 ={ {3{neg32[14]}} , neg32[14:3] };

   // m32_100 = W*in
   wire signed [14:0] m32_100;
   assign m32_100 =15'b0;

   // m33_1 = W*in
   wire signed [14:0] m33_1;
   assign m33_1 =15'b0;

   // m33_2 = W*in
   wire signed [14:0] m33_2;
   assign m33_2 =15'b0;

   // m33_3 = W*in
   wire signed [14:0] m33_3;
   assign m33_3 =15'b0;

   // m33_4 = W*in
   wire signed [14:0] m33_4;
   assign m33_4 =15'b0;

   // m33_5 = W*in
   wire signed [14:0] m33_5;
   assign m33_5 =15'b0;

   // m33_6 = W*in
   wire signed [14:0] m33_6;
   assign m33_6 =15'b0;

   // m33_7 = W*in
   wire signed [14:0] m33_7;
   assign m33_7 =15'b0;

   // m33_8 = W*in
   wire signed [14:0] m33_8;
   assign m33_8 =15'b0;

   // m33_9 = W*in
   wire signed [14:0] m33_9;
   assign m33_9 ={ {3{neg33[14]}} , neg33[14:3] };

   // m33_10 = W*in
   wire signed [14:0] m33_10;
   assign m33_10 ={ {4{neg33[14]}} , neg33[14:4] };

   // m33_11 = W*in
   wire signed [14:0] m33_11;
   assign m33_11 =15'b0;

   // m33_12 = W*in
   wire signed [14:0] m33_12;
   assign m33_12 =15'b0;

   // m33_13 = W*in
   wire signed [14:0] m33_13;
   assign m33_13 =15'b0;

   // m33_14 = W*in
   wire signed [14:0] m33_14;
   assign m33_14 =15'b0;

   // m33_15 = W*in
   wire signed [14:0] m33_15;
   assign m33_15 =15'b0;

   // m33_16 = W*in
   wire signed [14:0] m33_16;
   assign m33_16 =15'b0;

   // m33_17 = W*in
   wire signed [14:0] m33_17;
   assign m33_17 =15'b0;

   // m33_18 = W*in
   wire signed [14:0] m33_18;
   assign m33_18 ={ {3{in33[14]}} , in33[14:3] };

   // m33_19 = W*in
   wire signed [14:0] m33_19;
   assign m33_19 ={ {4{neg33[14]}} , neg33[14:4] };

   // m33_20 = W*in
   wire signed [14:0] m33_20;
   assign m33_20 =15'b0;

   // m33_21 = W*in
   wire signed [14:0] m33_21;
   assign m33_21 =15'b0;

   // m33_22 = W*in
   wire signed [14:0] m33_22;
   assign m33_22 =15'b0;

   // m33_23 = W*in
   wire signed [14:0] m33_23;
   assign m33_23 =15'b0;

   // m33_24 = W*in
   wire signed [14:0] m33_24;
   assign m33_24 =15'b0;

   // m33_25 = W*in
   wire signed [14:0] m33_25;
   assign m33_25 =15'b0;

   // m33_26 = W*in
   wire signed [14:0] m33_26;
   assign m33_26 =15'b0;

   // m33_27 = W*in
   wire signed [14:0] m33_27;
   assign m33_27 =15'b0;

   // m33_28 = W*in
   wire signed [14:0] m33_28;
   assign m33_28 =15'b0;

   // m33_29 = W*in
   wire signed [14:0] m33_29;
   assign m33_29 =15'b0;

   // m33_30 = W*in
   wire signed [14:0] m33_30;
   assign m33_30 =15'b0;

   // m33_31 = W*in
   wire signed [14:0] m33_31;
   assign m33_31 =15'b0;

   // m33_32 = W*in
   wire signed [14:0] m33_32;
   assign m33_32 =15'b0;

   // m33_33 = W*in
   wire signed [14:0] m33_33;
   assign m33_33 =15'b0;

   // m33_34 = W*in
   wire signed [14:0] m33_34;
   assign m33_34 =15'b0;

   // m33_35 = W*in
   wire signed [14:0] m33_35;
   assign m33_35 =15'b0;

   // m33_36 = W*in
   wire signed [14:0] m33_36;
   assign m33_36 =15'b0;

   // m33_37 = W*in
   wire signed [14:0] m33_37;
   assign m33_37 =15'b0;

   // m33_38 = W*in
   wire signed [14:0] m33_38;
   assign m33_38 ={ {3{in33[14]}} , in33[14:3] };

   // m33_39 = W*in
   wire signed [14:0] m33_39;
   assign m33_39 =15'b0;

   // m33_40 = W*in
   wire signed [14:0] m33_40;
   assign m33_40 =15'b0;

   // m33_41 = W*in
   wire signed [14:0] m33_41;
   assign m33_41 =15'b0;

   // m33_42 = W*in
   wire signed [14:0] m33_42;
   assign m33_42 =15'b0;

   // m33_43 = W*in
   wire signed [14:0] m33_43;
   assign m33_43 ={ {4{neg33[14]}} , neg33[14:4] };

   // m33_44 = W*in
   wire signed [14:0] m33_44;
   assign m33_44 =15'b0;

   // m33_45 = W*in
   wire signed [14:0] m33_45;
   assign m33_45 =15'b0;

   // m33_46 = W*in
   wire signed [14:0] m33_46;
   assign m33_46 =15'b0;

   // m33_47 = W*in
   wire signed [14:0] m33_47;
   assign m33_47 =15'b0;

   // m33_48 = W*in
   wire signed [14:0] m33_48;
   assign m33_48 =15'b0;

   // m33_49 = W*in
   wire signed [14:0] m33_49;
   assign m33_49 =15'b0;

   // m33_50 = W*in
   wire signed [14:0] m33_50;
   assign m33_50 =15'b0;

   // m33_51 = W*in
   wire signed [14:0] m33_51;
   assign m33_51 =15'b0;

   // m33_52 = W*in
   wire signed [14:0] m33_52;
   assign m33_52 =15'b0;

   // m33_53 = W*in
   wire signed [14:0] m33_53;
   assign m33_53 =15'b0;

   // m33_54 = W*in
   wire signed [14:0] m33_54;
   assign m33_54 =15'b0;

   // m33_55 = W*in
   wire signed [14:0] m33_55;
   assign m33_55 =15'b0;

   // m33_56 = W*in
   wire signed [14:0] m33_56;
   assign m33_56 =15'b0;

   // m33_57 = W*in
   wire signed [14:0] m33_57;
   assign m33_57 =15'b0;

   // m33_58 = W*in
   wire signed [14:0] m33_58;
   assign m33_58 =15'b0;

   // m33_59 = W*in
   wire signed [14:0] m33_59;
   assign m33_59 =15'b0;

   // m33_60 = W*in
   wire signed [14:0] m33_60;
   assign m33_60 =15'b0;

   // m33_61 = W*in
   wire signed [14:0] m33_61;
   assign m33_61 =15'b0;

   // m33_62 = W*in
   wire signed [14:0] m33_62;
   assign m33_62 =15'b0;

   // m33_63 = W*in
   wire signed [14:0] m33_63;
   assign m33_63 =15'b0;

   // m33_64 = W*in
   wire signed [14:0] m33_64;
   assign m33_64 ={ {4{in33[14]}} , in33[14:4] };

   // m33_65 = W*in
   wire signed [14:0] m33_65;
   assign m33_65 =15'b0;

   // m33_66 = W*in
   wire signed [14:0] m33_66;
   assign m33_66 =15'b0;

   // m33_67 = W*in
   wire signed [14:0] m33_67;
   assign m33_67 =15'b0;

   // m33_68 = W*in
   wire signed [14:0] m33_68;
   assign m33_68 ={ {3{neg33[14]}} , neg33[14:3] };

   // m33_69 = W*in
   wire signed [14:0] m33_69;
   assign m33_69 =15'b0;

   // m33_70 = W*in
   wire signed [14:0] m33_70;
   assign m33_70 =15'b0;

   // m33_71 = W*in
   wire signed [14:0] m33_71;
   assign m33_71 =15'b0;

   // m33_72 = W*in
   wire signed [14:0] m33_72;
   assign m33_72 =15'b0;

   // m33_73 = W*in
   wire signed [14:0] m33_73;
   assign m33_73 =15'b0;

   // m33_74 = W*in
   wire signed [14:0] m33_74;
   assign m33_74 =15'b0;

   // m33_75 = W*in
   wire signed [14:0] m33_75;
   assign m33_75 ={ {4{in33[14]}} , in33[14:4] };

   // m33_76 = W*in
   wire signed [14:0] m33_76;
   assign m33_76 =15'b0;

   // m33_77 = W*in
   wire signed [14:0] m33_77;
   assign m33_77 ={ {4{neg33[14]}} , neg33[14:4] };

   // m33_78 = W*in
   wire signed [14:0] m33_78;
   assign m33_78 =15'b0;

   // m33_79 = W*in
   wire signed [14:0] m33_79;
   assign m33_79 ={ {3{neg33[14]}} , neg33[14:3] };

   // m33_80 = W*in
   wire signed [14:0] m33_80;
   assign m33_80 =15'b0;

   // m33_81 = W*in
   wire signed [14:0] m33_81;
   assign m33_81 =15'b0;

   // m33_82 = W*in
   wire signed [14:0] m33_82;
   assign m33_82 =15'b0;

   // m33_83 = W*in
   wire signed [14:0] m33_83;
   assign m33_83 =15'b0;

   // m33_84 = W*in
   wire signed [14:0] m33_84;
   assign m33_84 =15'b0;

   // m33_85 = W*in
   wire signed [14:0] m33_85;
   assign m33_85 =15'b0;

   // m33_86 = W*in
   wire signed [14:0] m33_86;
   assign m33_86 ={ {3{in33[14]}} , in33[14:3] };

   // m33_87 = W*in
   wire signed [14:0] m33_87;
   assign m33_87 =15'b0;

   // m33_88 = W*in
   wire signed [14:0] m33_88;
   assign m33_88 =15'b0;

   // m33_89 = W*in
   wire signed [14:0] m33_89;
   assign m33_89 =15'b0;

   // m33_90 = W*in
   wire signed [14:0] m33_90;
   assign m33_90 =15'b0;

   // m33_91 = W*in
   wire signed [14:0] m33_91;
   assign m33_91 =15'b0;

   // m33_92 = W*in
   wire signed [14:0] m33_92;
   assign m33_92 =15'b0;

   // m33_93 = W*in
   wire signed [14:0] m33_93;
   assign m33_93 =15'b0;

   // m33_94 = W*in
   wire signed [14:0] m33_94;
   assign m33_94 =15'b0;

   // m33_95 = W*in
   wire signed [14:0] m33_95;
   assign m33_95 =15'b0;

   // m33_96 = W*in
   wire signed [14:0] m33_96;
   assign m33_96 ={ {4{in33[14]}} , in33[14:4] };

   // m33_97 = W*in
   wire signed [14:0] m33_97;
   assign m33_97 =15'b0;

   // m33_98 = W*in
   wire signed [14:0] m33_98;
   assign m33_98 =15'b0;

   // m33_99 = W*in
   wire signed [14:0] m33_99;
   assign m33_99 =15'b0;

   // m33_100 = W*in
   wire signed [14:0] m33_100;
   assign m33_100 =15'b0;

   // m34_1 = W*in
   wire signed [14:0] m34_1;
   assign m34_1 =15'b0;

   // m34_2 = W*in
   wire signed [14:0] m34_2;
   assign m34_2 =15'b0;

   // m34_3 = W*in
   wire signed [14:0] m34_3;
   assign m34_3 =15'b0;

   // m34_4 = W*in
   wire signed [14:0] m34_4;
   assign m34_4 =15'b0;

   // m34_5 = W*in
   wire signed [14:0] m34_5;
   assign m34_5 =15'b0;

   // m34_6 = W*in
   wire signed [14:0] m34_6;
   assign m34_6 =15'b0;

   // m34_7 = W*in
   wire signed [14:0] m34_7;
   assign m34_7 =15'b0;

   // m34_8 = W*in
   wire signed [14:0] m34_8;
   assign m34_8 =15'b0;

   // m34_9 = W*in
   wire signed [14:0] m34_9;
   assign m34_9 =15'b0;

   // m34_10 = W*in
   wire signed [14:0] m34_10;
   assign m34_10 =15'b0;

   // m34_11 = W*in
   wire signed [14:0] m34_11;
   assign m34_11 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_12 = W*in
   wire signed [14:0] m34_12;
   assign m34_12 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_13 = W*in
   wire signed [14:0] m34_13;
   assign m34_13 =15'b0;

   // m34_14 = W*in
   wire signed [14:0] m34_14;
   assign m34_14 =15'b0;

   // m34_15 = W*in
   wire signed [14:0] m34_15;
   assign m34_15 =15'b0;

   // m34_16 = W*in
   wire signed [14:0] m34_16;
   assign m34_16 =15'b0;

   // m34_17 = W*in
   wire signed [14:0] m34_17;
   assign m34_17 =15'b0;

   // m34_18 = W*in
   wire signed [14:0] m34_18;
   assign m34_18 =15'b0;

   // m34_19 = W*in
   wire signed [14:0] m34_19;
   assign m34_19 =15'b0;

   // m34_20 = W*in
   wire signed [14:0] m34_20;
   assign m34_20 =15'b0;

   // m34_21 = W*in
   wire signed [14:0] m34_21;
   assign m34_21 =15'b0;

   // m34_22 = W*in
   wire signed [14:0] m34_22;
   assign m34_22 =15'b0;

   // m34_23 = W*in
   wire signed [14:0] m34_23;
   assign m34_23 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_24 = W*in
   wire signed [14:0] m34_24;
   assign m34_24 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_25 = W*in
   wire signed [14:0] m34_25;
   assign m34_25 =15'b0;

   // m34_26 = W*in
   wire signed [14:0] m34_26;
   assign m34_26 =15'b0;

   // m34_27 = W*in
   wire signed [14:0] m34_27;
   assign m34_27 ={ {3{in34[14]}} , in34[14:3] };

   // m34_28 = W*in
   wire signed [14:0] m34_28;
   assign m34_28 =15'b0;

   // m34_29 = W*in
   wire signed [14:0] m34_29;
   assign m34_29 =15'b0;

   // m34_30 = W*in
   wire signed [14:0] m34_30;
   assign m34_30 =15'b0;

   // m34_31 = W*in
   wire signed [14:0] m34_31;
   assign m34_31 =15'b0;

   // m34_32 = W*in
   wire signed [14:0] m34_32;
   assign m34_32 =15'b0;

   // m34_33 = W*in
   wire signed [14:0] m34_33;
   assign m34_33 ={ {4{in34[14]}} , in34[14:4] };

   // m34_34 = W*in
   wire signed [14:0] m34_34;
   assign m34_34 =15'b0;

   // m34_35 = W*in
   wire signed [14:0] m34_35;
   assign m34_35 =15'b0;

   // m34_36 = W*in
   wire signed [14:0] m34_36;
   assign m34_36 =15'b0;

   // m34_37 = W*in
   wire signed [14:0] m34_37;
   assign m34_37 =15'b0;

   // m34_38 = W*in
   wire signed [14:0] m34_38;
   assign m34_38 =15'b0;

   // m34_39 = W*in
   wire signed [14:0] m34_39;
   assign m34_39 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_40 = W*in
   wire signed [14:0] m34_40;
   assign m34_40 =15'b0;

   // m34_41 = W*in
   wire signed [14:0] m34_41;
   assign m34_41 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_42 = W*in
   wire signed [14:0] m34_42;
   assign m34_42 ={ {3{in34[14]}} , in34[14:3] };

   // m34_43 = W*in
   wire signed [14:0] m34_43;
   assign m34_43 =15'b0;

   // m34_44 = W*in
   wire signed [14:0] m34_44;
   assign m34_44 =15'b0;

   // m34_45 = W*in
   wire signed [14:0] m34_45;
   assign m34_45 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_46 = W*in
   wire signed [14:0] m34_46;
   assign m34_46 =15'b0;

   // m34_47 = W*in
   wire signed [14:0] m34_47;
   assign m34_47 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_48 = W*in
   wire signed [14:0] m34_48;
   assign m34_48 =15'b0;

   // m34_49 = W*in
   wire signed [14:0] m34_49;
   assign m34_49 =15'b0;

   // m34_50 = W*in
   wire signed [14:0] m34_50;
   assign m34_50 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_51 = W*in
   wire signed [14:0] m34_51;
   assign m34_51 =15'b0;

   // m34_52 = W*in
   wire signed [14:0] m34_52;
   assign m34_52 =15'b0;

   // m34_53 = W*in
   wire signed [14:0] m34_53;
   assign m34_53 =15'b0;

   // m34_54 = W*in
   wire signed [14:0] m34_54;
   assign m34_54 =15'b0;

   // m34_55 = W*in
   wire signed [14:0] m34_55;
   assign m34_55 ={ {3{in34[14]}} , in34[14:3] };

   // m34_56 = W*in
   wire signed [14:0] m34_56;
   assign m34_56 =15'b0;

   // m34_57 = W*in
   wire signed [14:0] m34_57;
   assign m34_57 ={ {3{in34[14]}} , in34[14:3] };

   // m34_58 = W*in
   wire signed [14:0] m34_58;
   assign m34_58 =15'b0;

   // m34_59 = W*in
   wire signed [14:0] m34_59;
   assign m34_59 =15'b0;

   // m34_60 = W*in
   wire signed [14:0] m34_60;
   assign m34_60 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_61 = W*in
   wire signed [14:0] m34_61;
   assign m34_61 ={ {3{in34[14]}} , in34[14:3] };

   // m34_62 = W*in
   wire signed [14:0] m34_62;
   assign m34_62 =15'b0;

   // m34_63 = W*in
   wire signed [14:0] m34_63;
   assign m34_63 =15'b0;

   // m34_64 = W*in
   wire signed [14:0] m34_64;
   assign m34_64 ={ {4{neg34[14]}} , neg34[14:4] };

   // m34_65 = W*in
   wire signed [14:0] m34_65;
   assign m34_65 =15'b0;

   // m34_66 = W*in
   wire signed [14:0] m34_66;
   assign m34_66 =15'b0;

   // m34_67 = W*in
   wire signed [14:0] m34_67;
   assign m34_67 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_68 = W*in
   wire signed [14:0] m34_68;
   assign m34_68 ={ {3{in34[14]}} , in34[14:3] };

   // m34_69 = W*in
   wire signed [14:0] m34_69;
   assign m34_69 =15'b0;

   // m34_70 = W*in
   wire signed [14:0] m34_70;
   assign m34_70 =15'b0;

   // m34_71 = W*in
   wire signed [14:0] m34_71;
   assign m34_71 =15'b0;

   // m34_72 = W*in
   wire signed [14:0] m34_72;
   assign m34_72 =15'b0;

   // m34_73 = W*in
   wire signed [14:0] m34_73;
   assign m34_73 =15'b0;

   // m34_74 = W*in
   wire signed [14:0] m34_74;
   assign m34_74 =15'b0;

   // m34_75 = W*in
   wire signed [14:0] m34_75;
   assign m34_75 ={ {4{neg34[14]}} , neg34[14:4] };

   // m34_76 = W*in
   wire signed [14:0] m34_76;
   assign m34_76 =15'b0;

   // m34_77 = W*in
   wire signed [14:0] m34_77;
   assign m34_77 =15'b0;

   // m34_78 = W*in
   wire signed [14:0] m34_78;
   assign m34_78 =15'b0;

   // m34_79 = W*in
   wire signed [14:0] m34_79;
   assign m34_79 =15'b0;

   // m34_80 = W*in
   wire signed [14:0] m34_80;
   assign m34_80 =15'b0;

   // m34_81 = W*in
   wire signed [14:0] m34_81;
   assign m34_81 =15'b0;

   // m34_82 = W*in
   wire signed [14:0] m34_82;
   assign m34_82 =15'b0;

   // m34_83 = W*in
   wire signed [14:0] m34_83;
   assign m34_83 ={ {3{in34[14]}} , in34[14:3] };

   // m34_84 = W*in
   wire signed [14:0] m34_84;
   assign m34_84 =15'b0;

   // m34_85 = W*in
   wire signed [14:0] m34_85;
   assign m34_85 =15'b0;

   // m34_86 = W*in
   wire signed [14:0] m34_86;
   assign m34_86 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_87 = W*in
   wire signed [14:0] m34_87;
   assign m34_87 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_88 = W*in
   wire signed [14:0] m34_88;
   assign m34_88 =15'b0;

   // m34_89 = W*in
   wire signed [14:0] m34_89;
   assign m34_89 =15'b0;

   // m34_90 = W*in
   wire signed [14:0] m34_90;
   assign m34_90 =15'b0;

   // m34_91 = W*in
   wire signed [14:0] m34_91;
   assign m34_91 =15'b0;

   // m34_92 = W*in
   wire signed [14:0] m34_92;
   assign m34_92 ={ {3{in34[14]}} , in34[14:3] };

   // m34_93 = W*in
   wire signed [14:0] m34_93;
   assign m34_93 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_94 = W*in
   wire signed [14:0] m34_94;
   assign m34_94 =15'b0;

   // m34_95 = W*in
   wire signed [14:0] m34_95;
   assign m34_95 ={ {3{neg34[14]}} , neg34[14:3] };

   // m34_96 = W*in
   wire signed [14:0] m34_96;
   assign m34_96 =15'b0;

   // m34_97 = W*in
   wire signed [14:0] m34_97;
   assign m34_97 ={ {3{in34[14]}} , in34[14:3] };

   // m34_98 = W*in
   wire signed [14:0] m34_98;
   assign m34_98 =15'b0;

   // m34_99 = W*in
   wire signed [14:0] m34_99;
   assign m34_99 =15'b0;

   // m34_100 = W*in
   wire signed [14:0] m34_100;
   assign m34_100 =15'b0;

   // m35_1 = W*in
   wire signed [14:0] m35_1;
   assign m35_1 =15'b0;

   // m35_2 = W*in
   wire signed [14:0] m35_2;
   assign m35_2 =15'b0;

   // m35_3 = W*in
   wire signed [14:0] m35_3;
   assign m35_3 =15'b0;

   // m35_4 = W*in
   wire signed [14:0] m35_4;
   assign m35_4 =15'b0;

   // m35_5 = W*in
   wire signed [14:0] m35_5;
   assign m35_5 ={ {3{neg35[14]}} , neg35[14:3] };

   // m35_6 = W*in
   wire signed [14:0] m35_6;
   assign m35_6 =15'b0;

   // m35_7 = W*in
   wire signed [14:0] m35_7;
   assign m35_7 =15'b0;

   // m35_8 = W*in
   wire signed [14:0] m35_8;
   assign m35_8 =15'b0;

   // m35_9 = W*in
   wire signed [14:0] m35_9;
   assign m35_9 =15'b0;

   // m35_10 = W*in
   wire signed [14:0] m35_10;
   assign m35_10 =15'b0;

   // m35_11 = W*in
   wire signed [14:0] m35_11;
   assign m35_11 =15'b0;

   // m35_12 = W*in
   wire signed [14:0] m35_12;
   assign m35_12 =15'b0;

   // m35_13 = W*in
   wire signed [14:0] m35_13;
   assign m35_13 =15'b0;

   // m35_14 = W*in
   wire signed [14:0] m35_14;
   assign m35_14 =15'b0;

   // m35_15 = W*in
   wire signed [14:0] m35_15;
   assign m35_15 =15'b0;

   // m35_16 = W*in
   wire signed [14:0] m35_16;
   assign m35_16 =15'b0;

   // m35_17 = W*in
   wire signed [14:0] m35_17;
   assign m35_17 =15'b0;

   // m35_18 = W*in
   wire signed [14:0] m35_18;
   assign m35_18 =15'b0;

   // m35_19 = W*in
   wire signed [14:0] m35_19;
   assign m35_19 =15'b0;

   // m35_20 = W*in
   wire signed [14:0] m35_20;
   assign m35_20 =15'b0;

   // m35_21 = W*in
   wire signed [14:0] m35_21;
   assign m35_21 =15'b0;

   // m35_22 = W*in
   wire signed [14:0] m35_22;
   assign m35_22 =15'b0;

   // m35_23 = W*in
   wire signed [14:0] m35_23;
   assign m35_23 =15'b0;

   // m35_24 = W*in
   wire signed [14:0] m35_24;
   assign m35_24 =15'b0;

   // m35_25 = W*in
   wire signed [14:0] m35_25;
   assign m35_25 =15'b0;

   // m35_26 = W*in
   wire signed [14:0] m35_26;
   assign m35_26 =15'b0;

   // m35_27 = W*in
   wire signed [14:0] m35_27;
   assign m35_27 =15'b0;

   // m35_28 = W*in
   wire signed [14:0] m35_28;
   assign m35_28 ={ {4{in35[14]}} , in35[14:4] };

   // m35_29 = W*in
   wire signed [14:0] m35_29;
   assign m35_29 ={ {3{in35[14]}} , in35[14:3] };

   // m35_30 = W*in
   wire signed [14:0] m35_30;
   assign m35_30 =15'b0;

   // m35_31 = W*in
   wire signed [14:0] m35_31;
   assign m35_31 =15'b0;

   // m35_32 = W*in
   wire signed [14:0] m35_32;
   assign m35_32 =15'b0;

   // m35_33 = W*in
   wire signed [14:0] m35_33;
   assign m35_33 =15'b0;

   // m35_34 = W*in
   wire signed [14:0] m35_34;
   assign m35_34 =15'b0;

   // m35_35 = W*in
   wire signed [14:0] m35_35;
   assign m35_35 =15'b0;

   // m35_36 = W*in
   wire signed [14:0] m35_36;
   assign m35_36 ={ {3{neg35[14]}} , neg35[14:3] };

   // m35_37 = W*in
   wire signed [14:0] m35_37;
   assign m35_37 =15'b0;

   // m35_38 = W*in
   wire signed [14:0] m35_38;
   assign m35_38 =15'b0;

   // m35_39 = W*in
   wire signed [14:0] m35_39;
   assign m35_39 =15'b0;

   // m35_40 = W*in
   wire signed [14:0] m35_40;
   assign m35_40 =15'b0;

   // m35_41 = W*in
   wire signed [14:0] m35_41;
   assign m35_41 ={ {3{in35[14]}} , in35[14:3] };

   // m35_42 = W*in
   wire signed [14:0] m35_42;
   assign m35_42 =15'b0;

   // m35_43 = W*in
   wire signed [14:0] m35_43;
   assign m35_43 =15'b0;

   // m35_44 = W*in
   wire signed [14:0] m35_44;
   assign m35_44 =15'b0;

   // m35_45 = W*in
   wire signed [14:0] m35_45;
   assign m35_45 =15'b0;

   // m35_46 = W*in
   wire signed [14:0] m35_46;
   assign m35_46 =15'b0;

   // m35_47 = W*in
   wire signed [14:0] m35_47;
   assign m35_47 =15'b0;

   // m35_48 = W*in
   wire signed [14:0] m35_48;
   assign m35_48 =15'b0;

   // m35_49 = W*in
   wire signed [14:0] m35_49;
   assign m35_49 =15'b0;

   // m35_50 = W*in
   wire signed [14:0] m35_50;
   assign m35_50 =15'b0;

   // m35_51 = W*in
   wire signed [14:0] m35_51;
   assign m35_51 =15'b0;

   // m35_52 = W*in
   wire signed [14:0] m35_52;
   assign m35_52 =15'b0;

   // m35_53 = W*in
   wire signed [14:0] m35_53;
   assign m35_53 ={ {3{neg35[14]}} , neg35[14:3] };

   // m35_54 = W*in
   wire signed [14:0] m35_54;
   assign m35_54 =15'b0;

   // m35_55 = W*in
   wire signed [14:0] m35_55;
   assign m35_55 ={ {4{in35[14]}} , in35[14:4] };

   // m35_56 = W*in
   wire signed [14:0] m35_56;
   assign m35_56 ={ {4{in35[14]}} , in35[14:4] };

   // m35_57 = W*in
   wire signed [14:0] m35_57;
   assign m35_57 =15'b0;

   // m35_58 = W*in
   wire signed [14:0] m35_58;
   assign m35_58 =15'b0;

   // m35_59 = W*in
   wire signed [14:0] m35_59;
   assign m35_59 ={ {4{neg35[14]}} , neg35[14:4] };

   // m35_60 = W*in
   wire signed [14:0] m35_60;
   assign m35_60 ={ {3{in35[14]}} , in35[14:3] };

   // m35_61 = W*in
   wire signed [14:0] m35_61;
   assign m35_61 =15'b0;

   // m35_62 = W*in
   wire signed [14:0] m35_62;
   assign m35_62 =15'b0;

   // m35_63 = W*in
   wire signed [14:0] m35_63;
   assign m35_63 =15'b0;

   // m35_64 = W*in
   wire signed [14:0] m35_64;
   assign m35_64 =15'b0;

   // m35_65 = W*in
   wire signed [14:0] m35_65;
   assign m35_65 =15'b0;

   // m35_66 = W*in
   wire signed [14:0] m35_66;
   assign m35_66 =15'b0;

   // m35_67 = W*in
   wire signed [14:0] m35_67;
   assign m35_67 ={ {4{in35[14]}} , in35[14:4] };

   // m35_68 = W*in
   wire signed [14:0] m35_68;
   assign m35_68 ={ {3{neg35[14]}} , neg35[14:3] };

   // m35_69 = W*in
   wire signed [14:0] m35_69;
   assign m35_69 ={ {3{in35[14]}} , in35[14:3] };

   // m35_70 = W*in
   wire signed [14:0] m35_70;
   assign m35_70 =15'b0;

   // m35_71 = W*in
   wire signed [14:0] m35_71;
   assign m35_71 =15'b0;

   // m35_72 = W*in
   wire signed [14:0] m35_72;
   assign m35_72 =15'b0;

   // m35_73 = W*in
   wire signed [14:0] m35_73;
   assign m35_73 =15'b0;

   // m35_74 = W*in
   wire signed [14:0] m35_74;
   assign m35_74 ={ {4{neg35[14]}} , neg35[14:4] };

   // m35_75 = W*in
   wire signed [14:0] m35_75;
   assign m35_75 =15'b0;

   // m35_76 = W*in
   wire signed [14:0] m35_76;
   assign m35_76 =15'b0;

   // m35_77 = W*in
   wire signed [14:0] m35_77;
   assign m35_77 =15'b0;

   // m35_78 = W*in
   wire signed [14:0] m35_78;
   assign m35_78 =15'b0;

   // m35_79 = W*in
   wire signed [14:0] m35_79;
   assign m35_79 =15'b0;

   // m35_80 = W*in
   wire signed [14:0] m35_80;
   assign m35_80 ={ {4{in35[14]}} , in35[14:4] };

   // m35_81 = W*in
   wire signed [14:0] m35_81;
   assign m35_81 =15'b0;

   // m35_82 = W*in
   wire signed [14:0] m35_82;
   assign m35_82 =15'b0;

   // m35_83 = W*in
   wire signed [14:0] m35_83;
   assign m35_83 =15'b0;

   // m35_84 = W*in
   wire signed [14:0] m35_84;
   assign m35_84 =15'b0;

   // m35_85 = W*in
   wire signed [14:0] m35_85;
   assign m35_85 =15'b0;

   // m35_86 = W*in
   wire signed [14:0] m35_86;
   assign m35_86 =15'b0;

   // m35_87 = W*in
   wire signed [14:0] m35_87;
   assign m35_87 =15'b0;

   // m35_88 = W*in
   wire signed [14:0] m35_88;
   assign m35_88 =15'b0;

   // m35_89 = W*in
   wire signed [14:0] m35_89;
   assign m35_89 =15'b0;

   // m35_90 = W*in
   wire signed [14:0] m35_90;
   assign m35_90 =15'b0;

   // m35_91 = W*in
   wire signed [14:0] m35_91;
   assign m35_91 =15'b0;

   // m35_92 = W*in
   wire signed [14:0] m35_92;
   assign m35_92 =15'b0;

   // m35_93 = W*in
   wire signed [14:0] m35_93;
   assign m35_93 ={ {3{in35[14]}} , in35[14:3] };

   // m35_94 = W*in
   wire signed [14:0] m35_94;
   assign m35_94 =15'b0;

   // m35_95 = W*in
   wire signed [14:0] m35_95;
   assign m35_95 ={ {4{in35[14]}} , in35[14:4] };

   // m35_96 = W*in
   wire signed [14:0] m35_96;
   assign m35_96 =15'b0;

   // m35_97 = W*in
   wire signed [14:0] m35_97;
   assign m35_97 =15'b0;

   // m35_98 = W*in
   wire signed [14:0] m35_98;
   assign m35_98 ={ {4{in35[14]}} , in35[14:4] };

   // m35_99 = W*in
   wire signed [14:0] m35_99;
   assign m35_99 =15'b0;

   // m35_100 = W*in
   wire signed [14:0] m35_100;
   assign m35_100 =15'b0;

   // m36_1 = W*in
   wire signed [14:0] m36_1;
   assign m36_1 =15'b0;

   // m36_2 = W*in
   wire signed [14:0] m36_2;
   assign m36_2 =15'b0;

   // m36_3 = W*in
   wire signed [14:0] m36_3;
   assign m36_3 =15'b0;

   // m36_4 = W*in
   wire signed [14:0] m36_4;
   assign m36_4 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_5 = W*in
   wire signed [14:0] m36_5;
   assign m36_5 =15'b0;

   // m36_6 = W*in
   wire signed [14:0] m36_6;
   assign m36_6 =15'b0;

   // m36_7 = W*in
   wire signed [14:0] m36_7;
   assign m36_7 =15'b0;

   // m36_8 = W*in
   wire signed [14:0] m36_8;
   assign m36_8 ={ {3{in36[14]}} , in36[14:3] };

   // m36_9 = W*in
   wire signed [14:0] m36_9;
   assign m36_9 =15'b0;

   // m36_10 = W*in
   wire signed [14:0] m36_10;
   assign m36_10 =15'b0;

   // m36_11 = W*in
   wire signed [14:0] m36_11;
   assign m36_11 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_12 = W*in
   wire signed [14:0] m36_12;
   assign m36_12 =15'b0;

   // m36_13 = W*in
   wire signed [14:0] m36_13;
   assign m36_13 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_14 = W*in
   wire signed [14:0] m36_14;
   assign m36_14 =15'b0;

   // m36_15 = W*in
   wire signed [14:0] m36_15;
   assign m36_15 =15'b0;

   // m36_16 = W*in
   wire signed [14:0] m36_16;
   assign m36_16 =15'b0;

   // m36_17 = W*in
   wire signed [14:0] m36_17;
   assign m36_17 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_18 = W*in
   wire signed [14:0] m36_18;
   assign m36_18 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_19 = W*in
   wire signed [14:0] m36_19;
   assign m36_19 =15'b0;

   // m36_20 = W*in
   wire signed [14:0] m36_20;
   assign m36_20 ={ {4{neg36[14]}} , neg36[14:4] };

   // m36_21 = W*in
   wire signed [14:0] m36_21;
   assign m36_21 ={ {4{neg36[14]}} , neg36[14:4] };

   // m36_22 = W*in
   wire signed [14:0] m36_22;
   assign m36_22 =15'b0;

   // m36_23 = W*in
   wire signed [14:0] m36_23;
   assign m36_23 =15'b0;

   // m36_24 = W*in
   wire signed [14:0] m36_24;
   assign m36_24 =15'b0;

   // m36_25 = W*in
   wire signed [14:0] m36_25;
   assign m36_25 =15'b0;

   // m36_26 = W*in
   wire signed [14:0] m36_26;
   assign m36_26 ={ {3{in36[14]}} , in36[14:3] };

   // m36_27 = W*in
   wire signed [14:0] m36_27;
   assign m36_27 =15'b0;

   // m36_28 = W*in
   wire signed [14:0] m36_28;
   assign m36_28 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_29 = W*in
   wire signed [14:0] m36_29;
   assign m36_29 =15'b0;

   // m36_30 = W*in
   wire signed [14:0] m36_30;
   assign m36_30 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_31 = W*in
   wire signed [14:0] m36_31;
   assign m36_31 =15'b0;

   // m36_32 = W*in
   wire signed [14:0] m36_32;
   assign m36_32 ={ {4{neg36[14]}} , neg36[14:4] };

   // m36_33 = W*in
   wire signed [14:0] m36_33;
   assign m36_33 =15'b0;

   // m36_34 = W*in
   wire signed [14:0] m36_34;
   assign m36_34 =15'b0;

   // m36_35 = W*in
   wire signed [14:0] m36_35;
   assign m36_35 ={ {3{in36[14]}} , in36[14:3] };

   // m36_36 = W*in
   wire signed [14:0] m36_36;
   assign m36_36 =15'b0;

   // m36_37 = W*in
   wire signed [14:0] m36_37;
   assign m36_37 =15'b0;

   // m36_38 = W*in
   wire signed [14:0] m36_38;
   assign m36_38 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_39 = W*in
   wire signed [14:0] m36_39;
   assign m36_39 =15'b0;

   // m36_40 = W*in
   wire signed [14:0] m36_40;
   assign m36_40 =15'b0;

   // m36_41 = W*in
   wire signed [14:0] m36_41;
   assign m36_41 =15'b0;

   // m36_42 = W*in
   wire signed [14:0] m36_42;
   assign m36_42 ={ {3{in36[14]}} , in36[14:3] };

   // m36_43 = W*in
   wire signed [14:0] m36_43;
   assign m36_43 =15'b0;

   // m36_44 = W*in
   wire signed [14:0] m36_44;
   assign m36_44 =15'b0;

   // m36_45 = W*in
   wire signed [14:0] m36_45;
   assign m36_45 =15'b0;

   // m36_46 = W*in
   wire signed [14:0] m36_46;
   assign m36_46 =15'b0;

   // m36_47 = W*in
   wire signed [14:0] m36_47;
   assign m36_47 ={ {3{in36[14]}} , in36[14:3] };

   // m36_48 = W*in
   wire signed [14:0] m36_48;
   assign m36_48 =15'b0;

   // m36_49 = W*in
   wire signed [14:0] m36_49;
   assign m36_49 =15'b0;

   // m36_50 = W*in
   wire signed [14:0] m36_50;
   assign m36_50 =15'b0;

   // m36_51 = W*in
   wire signed [14:0] m36_51;
   assign m36_51 =15'b0;

   // m36_52 = W*in
   wire signed [14:0] m36_52;
   assign m36_52 =15'b0;

   // m36_53 = W*in
   wire signed [14:0] m36_53;
   assign m36_53 =15'b0;

   // m36_54 = W*in
   wire signed [14:0] m36_54;
   assign m36_54 =15'b0;

   // m36_55 = W*in
   wire signed [14:0] m36_55;
   assign m36_55 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_56 = W*in
   wire signed [14:0] m36_56;
   assign m36_56 =15'b0;

   // m36_57 = W*in
   wire signed [14:0] m36_57;
   assign m36_57 ={ {4{in36[14]}} , in36[14:4] };

   // m36_58 = W*in
   wire signed [14:0] m36_58;
   assign m36_58 =15'b0;

   // m36_59 = W*in
   wire signed [14:0] m36_59;
   assign m36_59 =15'b0;

   // m36_60 = W*in
   wire signed [14:0] m36_60;
   assign m36_60 =15'b0;

   // m36_61 = W*in
   wire signed [14:0] m36_61;
   assign m36_61 =15'b0;

   // m36_62 = W*in
   wire signed [14:0] m36_62;
   assign m36_62 =15'b0;

   // m36_63 = W*in
   wire signed [14:0] m36_63;
   assign m36_63 =15'b0;

   // m36_64 = W*in
   wire signed [14:0] m36_64;
   assign m36_64 =15'b0;

   // m36_65 = W*in
   wire signed [14:0] m36_65;
   assign m36_65 =15'b0;

   // m36_66 = W*in
   wire signed [14:0] m36_66;
   assign m36_66 =15'b0;

   // m36_67 = W*in
   wire signed [14:0] m36_67;
   assign m36_67 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_68 = W*in
   wire signed [14:0] m36_68;
   assign m36_68 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_69 = W*in
   wire signed [14:0] m36_69;
   assign m36_69 =15'b0;

   // m36_70 = W*in
   wire signed [14:0] m36_70;
   assign m36_70 =15'b0;

   // m36_71 = W*in
   wire signed [14:0] m36_71;
   assign m36_71 =15'b0;

   // m36_72 = W*in
   wire signed [14:0] m36_72;
   assign m36_72 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_73 = W*in
   wire signed [14:0] m36_73;
   assign m36_73 =15'b0;

   // m36_74 = W*in
   wire signed [14:0] m36_74;
   assign m36_74 =15'b0;

   // m36_75 = W*in
   wire signed [14:0] m36_75;
   assign m36_75 =15'b0;

   // m36_76 = W*in
   wire signed [14:0] m36_76;
   assign m36_76 =15'b0;

   // m36_77 = W*in
   wire signed [14:0] m36_77;
   assign m36_77 =15'b0;

   // m36_78 = W*in
   wire signed [14:0] m36_78;
   assign m36_78 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_79 = W*in
   wire signed [14:0] m36_79;
   assign m36_79 ={ {3{in36[14]}} , in36[14:3] };

   // m36_80 = W*in
   wire signed [14:0] m36_80;
   assign m36_80 =15'b0;

   // m36_81 = W*in
   wire signed [14:0] m36_81;
   assign m36_81 =15'b0;

   // m36_82 = W*in
   wire signed [14:0] m36_82;
   assign m36_82 =15'b0;

   // m36_83 = W*in
   wire signed [14:0] m36_83;
   assign m36_83 =15'b0;

   // m36_84 = W*in
   wire signed [14:0] m36_84;
   assign m36_84 =15'b0;

   // m36_85 = W*in
   wire signed [14:0] m36_85;
   assign m36_85 =15'b0;

   // m36_86 = W*in
   wire signed [14:0] m36_86;
   assign m36_86 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_87 = W*in
   wire signed [14:0] m36_87;
   assign m36_87 =15'b0;

   // m36_88 = W*in
   wire signed [14:0] m36_88;
   assign m36_88 =15'b0;

   // m36_89 = W*in
   wire signed [14:0] m36_89;
   assign m36_89 =15'b0;

   // m36_90 = W*in
   wire signed [14:0] m36_90;
   assign m36_90 =15'b0;

   // m36_91 = W*in
   wire signed [14:0] m36_91;
   assign m36_91 =15'b0;

   // m36_92 = W*in
   wire signed [14:0] m36_92;
   assign m36_92 =15'b0;

   // m36_93 = W*in
   wire signed [14:0] m36_93;
   assign m36_93 =15'b0;

   // m36_94 = W*in
   wire signed [14:0] m36_94;
   assign m36_94 =15'b0;

   // m36_95 = W*in
   wire signed [14:0] m36_95;
   assign m36_95 ={ {3{neg36[14]}} , neg36[14:3] };

   // m36_96 = W*in
   wire signed [14:0] m36_96;
   assign m36_96 =15'b0;

   // m36_97 = W*in
   wire signed [14:0] m36_97;
   assign m36_97 ={ {4{neg36[14]}} , neg36[14:4] };

   // m36_98 = W*in
   wire signed [14:0] m36_98;
   assign m36_98 =15'b0;

   // m36_99 = W*in
   wire signed [14:0] m36_99;
   assign m36_99 =15'b0;

   // m36_100 = W*in
   wire signed [14:0] m36_100;
   assign m36_100 ={ {3{in36[14]}} , in36[14:3] };

   // m37_1 = W*in
   wire signed [14:0] m37_1;
   assign m37_1 ={ {3{in37[14]}} , in37[14:3] };

   // m37_2 = W*in
   wire signed [14:0] m37_2;
   assign m37_2 =15'b0;

   // m37_3 = W*in
   wire signed [14:0] m37_3;
   assign m37_3 =15'b0;

   // m37_4 = W*in
   wire signed [14:0] m37_4;
   assign m37_4 =15'b0;

   // m37_5 = W*in
   wire signed [14:0] m37_5;
   assign m37_5 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_6 = W*in
   wire signed [14:0] m37_6;
   assign m37_6 =15'b0;

   // m37_7 = W*in
   wire signed [14:0] m37_7;
   assign m37_7 =15'b0;

   // m37_8 = W*in
   wire signed [14:0] m37_8;
   assign m37_8 ={ {3{in37[14]}} , in37[14:3] };

   // m37_9 = W*in
   wire signed [14:0] m37_9;
   assign m37_9 =15'b0;

   // m37_10 = W*in
   wire signed [14:0] m37_10;
   assign m37_10 =15'b0;

   // m37_11 = W*in
   wire signed [14:0] m37_11;
   assign m37_11 ={ {3{in37[14]}} , in37[14:3] };

   // m37_12 = W*in
   wire signed [14:0] m37_12;
   assign m37_12 =15'b0;

   // m37_13 = W*in
   wire signed [14:0] m37_13;
   assign m37_13 =15'b0;

   // m37_14 = W*in
   wire signed [14:0] m37_14;
   assign m37_14 =15'b0;

   // m37_15 = W*in
   wire signed [14:0] m37_15;
   assign m37_15 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_16 = W*in
   wire signed [14:0] m37_16;
   assign m37_16 =15'b0;

   // m37_17 = W*in
   wire signed [14:0] m37_17;
   assign m37_17 =15'b0;

   // m37_18 = W*in
   wire signed [14:0] m37_18;
   assign m37_18 =15'b0;

   // m37_19 = W*in
   wire signed [14:0] m37_19;
   assign m37_19 =15'b0;

   // m37_20 = W*in
   wire signed [14:0] m37_20;
   assign m37_20 =15'b0;

   // m37_21 = W*in
   wire signed [14:0] m37_21;
   assign m37_21 ={ {3{in37[14]}} , in37[14:3] };

   // m37_22 = W*in
   wire signed [14:0] m37_22;
   assign m37_22 =15'b0;

   // m37_23 = W*in
   wire signed [14:0] m37_23;
   assign m37_23 =15'b0;

   // m37_24 = W*in
   wire signed [14:0] m37_24;
   assign m37_24 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_25 = W*in
   wire signed [14:0] m37_25;
   assign m37_25 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_26 = W*in
   wire signed [14:0] m37_26;
   assign m37_26 =15'b0;

   // m37_27 = W*in
   wire signed [14:0] m37_27;
   assign m37_27 =15'b0;

   // m37_28 = W*in
   wire signed [14:0] m37_28;
   assign m37_28 =15'b0;

   // m37_29 = W*in
   wire signed [14:0] m37_29;
   assign m37_29 =15'b0;

   // m37_30 = W*in
   wire signed [14:0] m37_30;
   assign m37_30 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_31 = W*in
   wire signed [14:0] m37_31;
   assign m37_31 =15'b0;

   // m37_32 = W*in
   wire signed [14:0] m37_32;
   assign m37_32 =15'b0;

   // m37_33 = W*in
   wire signed [14:0] m37_33;
   assign m37_33 =15'b0;

   // m37_34 = W*in
   wire signed [14:0] m37_34;
   assign m37_34 =15'b0;

   // m37_35 = W*in
   wire signed [14:0] m37_35;
   assign m37_35 =15'b0;

   // m37_36 = W*in
   wire signed [14:0] m37_36;
   assign m37_36 =15'b0;

   // m37_37 = W*in
   wire signed [14:0] m37_37;
   assign m37_37 =15'b0;

   // m37_38 = W*in
   wire signed [14:0] m37_38;
   assign m37_38 =15'b0;

   // m37_39 = W*in
   wire signed [14:0] m37_39;
   assign m37_39 =15'b0;

   // m37_40 = W*in
   wire signed [14:0] m37_40;
   assign m37_40 =15'b0;

   // m37_41 = W*in
   wire signed [14:0] m37_41;
   assign m37_41 =15'b0;

   // m37_42 = W*in
   wire signed [14:0] m37_42;
   assign m37_42 =15'b0;

   // m37_43 = W*in
   wire signed [14:0] m37_43;
   assign m37_43 =15'b0;

   // m37_44 = W*in
   wire signed [14:0] m37_44;
   assign m37_44 =15'b0;

   // m37_45 = W*in
   wire signed [14:0] m37_45;
   assign m37_45 =15'b0;

   // m37_46 = W*in
   wire signed [14:0] m37_46;
   assign m37_46 =15'b0;

   // m37_47 = W*in
   wire signed [14:0] m37_47;
   assign m37_47 =15'b0;

   // m37_48 = W*in
   wire signed [14:0] m37_48;
   assign m37_48 =15'b0;

   // m37_49 = W*in
   wire signed [14:0] m37_49;
   assign m37_49 =15'b0;

   // m37_50 = W*in
   wire signed [14:0] m37_50;
   assign m37_50 =15'b0;

   // m37_51 = W*in
   wire signed [14:0] m37_51;
   assign m37_51 =15'b0;

   // m37_52 = W*in
   wire signed [14:0] m37_52;
   assign m37_52 ={ {3{in37[14]}} , in37[14:3] };

   // m37_53 = W*in
   wire signed [14:0] m37_53;
   assign m37_53 =15'b0;

   // m37_54 = W*in
   wire signed [14:0] m37_54;
   assign m37_54 =15'b0;

   // m37_55 = W*in
   wire signed [14:0] m37_55;
   assign m37_55 =15'b0;

   // m37_56 = W*in
   wire signed [14:0] m37_56;
   assign m37_56 =15'b0;

   // m37_57 = W*in
   wire signed [14:0] m37_57;
   assign m37_57 =15'b0;

   // m37_58 = W*in
   wire signed [14:0] m37_58;
   assign m37_58 =15'b0;

   // m37_59 = W*in
   wire signed [14:0] m37_59;
   assign m37_59 =15'b0;

   // m37_60 = W*in
   wire signed [14:0] m37_60;
   assign m37_60 ={ {3{in37[14]}} , in37[14:3] };

   // m37_61 = W*in
   wire signed [14:0] m37_61;
   assign m37_61 ={ {4{neg37[14]}} , neg37[14:4] };

   // m37_62 = W*in
   wire signed [14:0] m37_62;
   assign m37_62 =15'b0;

   // m37_63 = W*in
   wire signed [14:0] m37_63;
   assign m37_63 =15'b0;

   // m37_64 = W*in
   wire signed [14:0] m37_64;
   assign m37_64 =15'b0;

   // m37_65 = W*in
   wire signed [14:0] m37_65;
   assign m37_65 =15'b0;

   // m37_66 = W*in
   wire signed [14:0] m37_66;
   assign m37_66 =15'b0;

   // m37_67 = W*in
   wire signed [14:0] m37_67;
   assign m37_67 =15'b0;

   // m37_68 = W*in
   wire signed [14:0] m37_68;
   assign m37_68 =15'b0;

   // m37_69 = W*in
   wire signed [14:0] m37_69;
   assign m37_69 =15'b0;

   // m37_70 = W*in
   wire signed [14:0] m37_70;
   assign m37_70 =15'b0;

   // m37_71 = W*in
   wire signed [14:0] m37_71;
   assign m37_71 =15'b0;

   // m37_72 = W*in
   wire signed [14:0] m37_72;
   assign m37_72 =15'b0;

   // m37_73 = W*in
   wire signed [14:0] m37_73;
   assign m37_73 ={ {3{in37[14]}} , in37[14:3] };

   // m37_74 = W*in
   wire signed [14:0] m37_74;
   assign m37_74 =15'b0;

   // m37_75 = W*in
   wire signed [14:0] m37_75;
   assign m37_75 =15'b0;

   // m37_76 = W*in
   wire signed [14:0] m37_76;
   assign m37_76 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_77 = W*in
   wire signed [14:0] m37_77;
   assign m37_77 =15'b0;

   // m37_78 = W*in
   wire signed [14:0] m37_78;
   assign m37_78 =15'b0;

   // m37_79 = W*in
   wire signed [14:0] m37_79;
   assign m37_79 =15'b0;

   // m37_80 = W*in
   wire signed [14:0] m37_80;
   assign m37_80 =15'b0;

   // m37_81 = W*in
   wire signed [14:0] m37_81;
   assign m37_81 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_82 = W*in
   wire signed [14:0] m37_82;
   assign m37_82 =15'b0;

   // m37_83 = W*in
   wire signed [14:0] m37_83;
   assign m37_83 =15'b0;

   // m37_84 = W*in
   wire signed [14:0] m37_84;
   assign m37_84 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_85 = W*in
   wire signed [14:0] m37_85;
   assign m37_85 =15'b0;

   // m37_86 = W*in
   wire signed [14:0] m37_86;
   assign m37_86 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_87 = W*in
   wire signed [14:0] m37_87;
   assign m37_87 =15'b0;

   // m37_88 = W*in
   wire signed [14:0] m37_88;
   assign m37_88 ={ {3{in37[14]}} , in37[14:3] };

   // m37_89 = W*in
   wire signed [14:0] m37_89;
   assign m37_89 =15'b0;

   // m37_90 = W*in
   wire signed [14:0] m37_90;
   assign m37_90 =15'b0;

   // m37_91 = W*in
   wire signed [14:0] m37_91;
   assign m37_91 =15'b0;

   // m37_92 = W*in
   wire signed [14:0] m37_92;
   assign m37_92 =15'b0;

   // m37_93 = W*in
   wire signed [14:0] m37_93;
   assign m37_93 =15'b0;

   // m37_94 = W*in
   wire signed [14:0] m37_94;
   assign m37_94 =15'b0;

   // m37_95 = W*in
   wire signed [14:0] m37_95;
   assign m37_95 =15'b0;

   // m37_96 = W*in
   wire signed [14:0] m37_96;
   assign m37_96 =15'b0;

   // m37_97 = W*in
   wire signed [14:0] m37_97;
   assign m37_97 =15'b0;

   // m37_98 = W*in
   wire signed [14:0] m37_98;
   assign m37_98 ={ {3{neg37[14]}} , neg37[14:3] };

   // m37_99 = W*in
   wire signed [14:0] m37_99;
   assign m37_99 =15'b0;

   // m37_100 = W*in
   wire signed [14:0] m37_100;
   assign m37_100 =15'b0;

   // m38_1 = W*in
   wire signed [14:0] m38_1;
   assign m38_1 =15'b0;

   // m38_2 = W*in
   wire signed [14:0] m38_2;
   assign m38_2 =15'b0;

   // m38_3 = W*in
   wire signed [14:0] m38_3;
   assign m38_3 =15'b0;

   // m38_4 = W*in
   wire signed [14:0] m38_4;
   assign m38_4 =15'b0;

   // m38_5 = W*in
   wire signed [14:0] m38_5;
   assign m38_5 =15'b0;

   // m38_6 = W*in
   wire signed [14:0] m38_6;
   assign m38_6 =15'b0;

   // m38_7 = W*in
   wire signed [14:0] m38_7;
   assign m38_7 =15'b0;

   // m38_8 = W*in
   wire signed [14:0] m38_8;
   assign m38_8 ={ {3{in38[14]}} , in38[14:3] };

   // m38_9 = W*in
   wire signed [14:0] m38_9;
   assign m38_9 ={ {3{neg38[14]}} , neg38[14:3] };

   // m38_10 = W*in
   wire signed [14:0] m38_10;
   assign m38_10 =15'b0;

   // m38_11 = W*in
   wire signed [14:0] m38_11;
   assign m38_11 =15'b0;

   // m38_12 = W*in
   wire signed [14:0] m38_12;
   assign m38_12 =15'b0;

   // m38_13 = W*in
   wire signed [14:0] m38_13;
   assign m38_13 =15'b0;

   // m38_14 = W*in
   wire signed [14:0] m38_14;
   assign m38_14 =15'b0;

   // m38_15 = W*in
   wire signed [14:0] m38_15;
   assign m38_15 =15'b0;

   // m38_16 = W*in
   wire signed [14:0] m38_16;
   assign m38_16 =15'b0;

   // m38_17 = W*in
   wire signed [14:0] m38_17;
   assign m38_17 =15'b0;

   // m38_18 = W*in
   wire signed [14:0] m38_18;
   assign m38_18 =15'b0;

   // m38_19 = W*in
   wire signed [14:0] m38_19;
   assign m38_19 =15'b0;

   // m38_20 = W*in
   wire signed [14:0] m38_20;
   assign m38_20 =15'b0;

   // m38_21 = W*in
   wire signed [14:0] m38_21;
   assign m38_21 ={ {4{neg38[14]}} , neg38[14:4] };

   // m38_22 = W*in
   wire signed [14:0] m38_22;
   assign m38_22 =15'b0;

   // m38_23 = W*in
   wire signed [14:0] m38_23;
   assign m38_23 ={ {3{neg38[14]}} , neg38[14:3] };

   // m38_24 = W*in
   wire signed [14:0] m38_24;
   assign m38_24 =15'b0;

   // m38_25 = W*in
   wire signed [14:0] m38_25;
   assign m38_25 =15'b0;

   // m38_26 = W*in
   wire signed [14:0] m38_26;
   assign m38_26 =15'b0;

   // m38_27 = W*in
   wire signed [14:0] m38_27;
   assign m38_27 =15'b0;

   // m38_28 = W*in
   wire signed [14:0] m38_28;
   assign m38_28 ={ {3{in38[14]}} , in38[14:3] };

   // m38_29 = W*in
   wire signed [14:0] m38_29;
   assign m38_29 =15'b0;

   // m38_30 = W*in
   wire signed [14:0] m38_30;
   assign m38_30 =15'b0;

   // m38_31 = W*in
   wire signed [14:0] m38_31;
   assign m38_31 =15'b0;

   // m38_32 = W*in
   wire signed [14:0] m38_32;
   assign m38_32 =15'b0;

   // m38_33 = W*in
   wire signed [14:0] m38_33;
   assign m38_33 ={ {3{in38[14]}} , in38[14:3] };

   // m38_34 = W*in
   wire signed [14:0] m38_34;
   assign m38_34 ={ {3{neg38[14]}} , neg38[14:3] };

   // m38_35 = W*in
   wire signed [14:0] m38_35;
   assign m38_35 =15'b0;

   // m38_36 = W*in
   wire signed [14:0] m38_36;
   assign m38_36 ={ {3{neg38[14]}} , neg38[14:3] };

   // m38_37 = W*in
   wire signed [14:0] m38_37;
   assign m38_37 =15'b0;

   // m38_38 = W*in
   wire signed [14:0] m38_38;
   assign m38_38 =15'b0;

   // m38_39 = W*in
   wire signed [14:0] m38_39;
   assign m38_39 =15'b0;

   // m38_40 = W*in
   wire signed [14:0] m38_40;
   assign m38_40 =15'b0;

   // m38_41 = W*in
   wire signed [14:0] m38_41;
   assign m38_41 =15'b0;

   // m38_42 = W*in
   wire signed [14:0] m38_42;
   assign m38_42 =15'b0;

   // m38_43 = W*in
   wire signed [14:0] m38_43;
   assign m38_43 =15'b0;

   // m38_44 = W*in
   wire signed [14:0] m38_44;
   assign m38_44 =15'b0;

   // m38_45 = W*in
   wire signed [14:0] m38_45;
   assign m38_45 =15'b0;

   // m38_46 = W*in
   wire signed [14:0] m38_46;
   assign m38_46 =15'b0;

   // m38_47 = W*in
   wire signed [14:0] m38_47;
   assign m38_47 =15'b0;

   // m38_48 = W*in
   wire signed [14:0] m38_48;
   assign m38_48 =15'b0;

   // m38_49 = W*in
   wire signed [14:0] m38_49;
   assign m38_49 =15'b0;

   // m38_50 = W*in
   wire signed [14:0] m38_50;
   assign m38_50 =15'b0;

   // m38_51 = W*in
   wire signed [14:0] m38_51;
   assign m38_51 =15'b0;

   // m38_52 = W*in
   wire signed [14:0] m38_52;
   assign m38_52 =15'b0;

   // m38_53 = W*in
   wire signed [14:0] m38_53;
   assign m38_53 ={ {3{in38[14]}} , in38[14:3] };

   // m38_54 = W*in
   wire signed [14:0] m38_54;
   assign m38_54 =15'b0;

   // m38_55 = W*in
   wire signed [14:0] m38_55;
   assign m38_55 =15'b0;

   // m38_56 = W*in
   wire signed [14:0] m38_56;
   assign m38_56 =15'b0;

   // m38_57 = W*in
   wire signed [14:0] m38_57;
   assign m38_57 =15'b0;

   // m38_58 = W*in
   wire signed [14:0] m38_58;
   assign m38_58 ={ {3{neg38[14]}} , neg38[14:3] };

   // m38_59 = W*in
   wire signed [14:0] m38_59;
   assign m38_59 =15'b0;

   // m38_60 = W*in
   wire signed [14:0] m38_60;
   assign m38_60 =15'b0;

   // m38_61 = W*in
   wire signed [14:0] m38_61;
   assign m38_61 =15'b0;

   // m38_62 = W*in
   wire signed [14:0] m38_62;
   assign m38_62 =15'b0;

   // m38_63 = W*in
   wire signed [14:0] m38_63;
   assign m38_63 =15'b0;

   // m38_64 = W*in
   wire signed [14:0] m38_64;
   assign m38_64 =15'b0;

   // m38_65 = W*in
   wire signed [14:0] m38_65;
   assign m38_65 =15'b0;

   // m38_66 = W*in
   wire signed [14:0] m38_66;
   assign m38_66 =15'b0;

   // m38_67 = W*in
   wire signed [14:0] m38_67;
   assign m38_67 =15'b0;

   // m38_68 = W*in
   wire signed [14:0] m38_68;
   assign m38_68 ={ {3{in38[14]}} , in38[14:3] };

   // m38_69 = W*in
   wire signed [14:0] m38_69;
   assign m38_69 =15'b0;

   // m38_70 = W*in
   wire signed [14:0] m38_70;
   assign m38_70 =15'b0;

   // m38_71 = W*in
   wire signed [14:0] m38_71;
   assign m38_71 =15'b0;

   // m38_72 = W*in
   wire signed [14:0] m38_72;
   assign m38_72 =15'b0;

   // m38_73 = W*in
   wire signed [14:0] m38_73;
   assign m38_73 =15'b0;

   // m38_74 = W*in
   wire signed [14:0] m38_74;
   assign m38_74 =15'b0;

   // m38_75 = W*in
   wire signed [14:0] m38_75;
   assign m38_75 =15'b0;

   // m38_76 = W*in
   wire signed [14:0] m38_76;
   assign m38_76 =15'b0;

   // m38_77 = W*in
   wire signed [14:0] m38_77;
   assign m38_77 =15'b0;

   // m38_78 = W*in
   wire signed [14:0] m38_78;
   assign m38_78 =15'b0;

   // m38_79 = W*in
   wire signed [14:0] m38_79;
   assign m38_79 =15'b0;

   // m38_80 = W*in
   wire signed [14:0] m38_80;
   assign m38_80 =15'b0;

   // m38_81 = W*in
   wire signed [14:0] m38_81;
   assign m38_81 =15'b0;

   // m38_82 = W*in
   wire signed [14:0] m38_82;
   assign m38_82 =15'b0;

   // m38_83 = W*in
   wire signed [14:0] m38_83;
   assign m38_83 =15'b0;

   // m38_84 = W*in
   wire signed [14:0] m38_84;
   assign m38_84 =15'b0;

   // m38_85 = W*in
   wire signed [14:0] m38_85;
   assign m38_85 =15'b0;

   // m38_86 = W*in
   wire signed [14:0] m38_86;
   assign m38_86 =15'b0;

   // m38_87 = W*in
   wire signed [14:0] m38_87;
   assign m38_87 =15'b0;

   // m38_88 = W*in
   wire signed [14:0] m38_88;
   assign m38_88 =15'b0;

   // m38_89 = W*in
   wire signed [14:0] m38_89;
   assign m38_89 =15'b0;

   // m38_90 = W*in
   wire signed [14:0] m38_90;
   assign m38_90 =15'b0;

   // m38_91 = W*in
   wire signed [14:0] m38_91;
   assign m38_91 =15'b0;

   // m38_92 = W*in
   wire signed [14:0] m38_92;
   assign m38_92 =15'b0;

   // m38_93 = W*in
   wire signed [14:0] m38_93;
   assign m38_93 ={ {3{neg38[14]}} , neg38[14:3] };

   // m38_94 = W*in
   wire signed [14:0] m38_94;
   assign m38_94 ={ {4{neg38[14]}} , neg38[14:4] };

   // m38_95 = W*in
   wire signed [14:0] m38_95;
   assign m38_95 =15'b0;

   // m38_96 = W*in
   wire signed [14:0] m38_96;
   assign m38_96 =15'b0;

   // m38_97 = W*in
   wire signed [14:0] m38_97;
   assign m38_97 =15'b0;

   // m38_98 = W*in
   wire signed [14:0] m38_98;
   assign m38_98 ={ {4{neg38[14]}} , neg38[14:4] };

   // m38_99 = W*in
   wire signed [14:0] m38_99;
   assign m38_99 =15'b0;

   // m38_100 = W*in
   wire signed [14:0] m38_100;
   assign m38_100 =15'b0;

   // m39_1 = W*in
   wire signed [14:0] m39_1;
   assign m39_1 =15'b0;

   // m39_2 = W*in
   wire signed [14:0] m39_2;
   assign m39_2 =15'b0;

   // m39_3 = W*in
   wire signed [14:0] m39_3;
   assign m39_3 =15'b0;

   // m39_4 = W*in
   wire signed [14:0] m39_4;
   assign m39_4 =15'b0;

   // m39_5 = W*in
   wire signed [14:0] m39_5;
   assign m39_5 =15'b0;

   // m39_6 = W*in
   wire signed [14:0] m39_6;
   assign m39_6 =15'b0;

   // m39_7 = W*in
   wire signed [14:0] m39_7;
   assign m39_7 =15'b0;

   // m39_8 = W*in
   wire signed [14:0] m39_8;
   assign m39_8 =15'b0;

   // m39_9 = W*in
   wire signed [14:0] m39_9;
   assign m39_9 =15'b0;

   // m39_10 = W*in
   wire signed [14:0] m39_10;
   assign m39_10 =15'b0;

   // m39_11 = W*in
   wire signed [14:0] m39_11;
   assign m39_11 ={ {3{in39[14]}} , in39[14:3] };

   // m39_12 = W*in
   wire signed [14:0] m39_12;
   assign m39_12 =15'b0;

   // m39_13 = W*in
   wire signed [14:0] m39_13;
   assign m39_13 =15'b0;

   // m39_14 = W*in
   wire signed [14:0] m39_14;
   assign m39_14 =15'b0;

   // m39_15 = W*in
   wire signed [14:0] m39_15;
   assign m39_15 =15'b0;

   // m39_16 = W*in
   wire signed [14:0] m39_16;
   assign m39_16 =15'b0;

   // m39_17 = W*in
   wire signed [14:0] m39_17;
   assign m39_17 ={ {3{in39[14]}} , in39[14:3] };

   // m39_18 = W*in
   wire signed [14:0] m39_18;
   assign m39_18 =15'b0;

   // m39_19 = W*in
   wire signed [14:0] m39_19;
   assign m39_19 =15'b0;

   // m39_20 = W*in
   wire signed [14:0] m39_20;
   assign m39_20 =15'b0;

   // m39_21 = W*in
   wire signed [14:0] m39_21;
   assign m39_21 =15'b0;

   // m39_22 = W*in
   wire signed [14:0] m39_22;
   assign m39_22 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_23 = W*in
   wire signed [14:0] m39_23;
   assign m39_23 =15'b0;

   // m39_24 = W*in
   wire signed [14:0] m39_24;
   assign m39_24 =15'b0;

   // m39_25 = W*in
   wire signed [14:0] m39_25;
   assign m39_25 =15'b0;

   // m39_26 = W*in
   wire signed [14:0] m39_26;
   assign m39_26 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_27 = W*in
   wire signed [14:0] m39_27;
   assign m39_27 =15'b0;

   // m39_28 = W*in
   wire signed [14:0] m39_28;
   assign m39_28 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_29 = W*in
   wire signed [14:0] m39_29;
   assign m39_29 =15'b0;

   // m39_30 = W*in
   wire signed [14:0] m39_30;
   assign m39_30 ={ {4{in39[14]}} , in39[14:4] };

   // m39_31 = W*in
   wire signed [14:0] m39_31;
   assign m39_31 =15'b0;

   // m39_32 = W*in
   wire signed [14:0] m39_32;
   assign m39_32 =15'b0;

   // m39_33 = W*in
   wire signed [14:0] m39_33;
   assign m39_33 =15'b0;

   // m39_34 = W*in
   wire signed [14:0] m39_34;
   assign m39_34 =15'b0;

   // m39_35 = W*in
   wire signed [14:0] m39_35;
   assign m39_35 =15'b0;

   // m39_36 = W*in
   wire signed [14:0] m39_36;
   assign m39_36 =15'b0;

   // m39_37 = W*in
   wire signed [14:0] m39_37;
   assign m39_37 =15'b0;

   // m39_38 = W*in
   wire signed [14:0] m39_38;
   assign m39_38 =15'b0;

   // m39_39 = W*in
   wire signed [14:0] m39_39;
   assign m39_39 =15'b0;

   // m39_40 = W*in
   wire signed [14:0] m39_40;
   assign m39_40 =15'b0;

   // m39_41 = W*in
   wire signed [14:0] m39_41;
   assign m39_41 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_42 = W*in
   wire signed [14:0] m39_42;
   assign m39_42 =15'b0;

   // m39_43 = W*in
   wire signed [14:0] m39_43;
   assign m39_43 =15'b0;

   // m39_44 = W*in
   wire signed [14:0] m39_44;
   assign m39_44 =15'b0;

   // m39_45 = W*in
   wire signed [14:0] m39_45;
   assign m39_45 =15'b0;

   // m39_46 = W*in
   wire signed [14:0] m39_46;
   assign m39_46 ={ {3{neg39[14]}} , neg39[14:3] };

   // m39_47 = W*in
   wire signed [14:0] m39_47;
   assign m39_47 =15'b0;

   // m39_48 = W*in
   wire signed [14:0] m39_48;
   assign m39_48 =15'b0;

   // m39_49 = W*in
   wire signed [14:0] m39_49;
   assign m39_49 =15'b0;

   // m39_50 = W*in
   wire signed [14:0] m39_50;
   assign m39_50 =15'b0;

   // m39_51 = W*in
   wire signed [14:0] m39_51;
   assign m39_51 =15'b0;

   // m39_52 = W*in
   wire signed [14:0] m39_52;
   assign m39_52 =15'b0;

   // m39_53 = W*in
   wire signed [14:0] m39_53;
   assign m39_53 =15'b0;

   // m39_54 = W*in
   wire signed [14:0] m39_54;
   assign m39_54 =15'b0;

   // m39_55 = W*in
   wire signed [14:0] m39_55;
   assign m39_55 =15'b0;

   // m39_56 = W*in
   wire signed [14:0] m39_56;
   assign m39_56 ={ {3{in39[14]}} , in39[14:3] };

   // m39_57 = W*in
   wire signed [14:0] m39_57;
   assign m39_57 =15'b0;

   // m39_58 = W*in
   wire signed [14:0] m39_58;
   assign m39_58 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_59 = W*in
   wire signed [14:0] m39_59;
   assign m39_59 =15'b0;

   // m39_60 = W*in
   wire signed [14:0] m39_60;
   assign m39_60 =15'b0;

   // m39_61 = W*in
   wire signed [14:0] m39_61;
   assign m39_61 =15'b0;

   // m39_62 = W*in
   wire signed [14:0] m39_62;
   assign m39_62 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_63 = W*in
   wire signed [14:0] m39_63;
   assign m39_63 ={ {3{neg39[14]}} , neg39[14:3] };

   // m39_64 = W*in
   wire signed [14:0] m39_64;
   assign m39_64 =15'b0;

   // m39_65 = W*in
   wire signed [14:0] m39_65;
   assign m39_65 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_66 = W*in
   wire signed [14:0] m39_66;
   assign m39_66 =15'b0;

   // m39_67 = W*in
   wire signed [14:0] m39_67;
   assign m39_67 ={ {3{in39[14]}} , in39[14:3] };

   // m39_68 = W*in
   wire signed [14:0] m39_68;
   assign m39_68 =15'b0;

   // m39_69 = W*in
   wire signed [14:0] m39_69;
   assign m39_69 =15'b0;

   // m39_70 = W*in
   wire signed [14:0] m39_70;
   assign m39_70 =15'b0;

   // m39_71 = W*in
   wire signed [14:0] m39_71;
   assign m39_71 ={ {4{neg39[14]}} , neg39[14:4] };

   // m39_72 = W*in
   wire signed [14:0] m39_72;
   assign m39_72 =15'b0;

   // m39_73 = W*in
   wire signed [14:0] m39_73;
   assign m39_73 =15'b0;

   // m39_74 = W*in
   wire signed [14:0] m39_74;
   assign m39_74 =15'b0;

   // m39_75 = W*in
   wire signed [14:0] m39_75;
   assign m39_75 =15'b0;

   // m39_76 = W*in
   wire signed [14:0] m39_76;
   assign m39_76 =15'b0;

   // m39_77 = W*in
   wire signed [14:0] m39_77;
   assign m39_77 =15'b0;

   // m39_78 = W*in
   wire signed [14:0] m39_78;
   assign m39_78 =15'b0;

   // m39_79 = W*in
   wire signed [14:0] m39_79;
   assign m39_79 =15'b0;

   // m39_80 = W*in
   wire signed [14:0] m39_80;
   assign m39_80 =15'b0;

   // m39_81 = W*in
   wire signed [14:0] m39_81;
   assign m39_81 =15'b0;

   // m39_82 = W*in
   wire signed [14:0] m39_82;
   assign m39_82 =15'b0;

   // m39_83 = W*in
   wire signed [14:0] m39_83;
   assign m39_83 =15'b0;

   // m39_84 = W*in
   wire signed [14:0] m39_84;
   assign m39_84 =15'b0;

   // m39_85 = W*in
   wire signed [14:0] m39_85;
   assign m39_85 =15'b0;

   // m39_86 = W*in
   wire signed [14:0] m39_86;
   assign m39_86 ={ {3{in39[14]}} , in39[14:3] };

   // m39_87 = W*in
   wire signed [14:0] m39_87;
   assign m39_87 =15'b0;

   // m39_88 = W*in
   wire signed [14:0] m39_88;
   assign m39_88 =15'b0;

   // m39_89 = W*in
   wire signed [14:0] m39_89;
   assign m39_89 =15'b0;

   // m39_90 = W*in
   wire signed [14:0] m39_90;
   assign m39_90 =15'b0;

   // m39_91 = W*in
   wire signed [14:0] m39_91;
   assign m39_91 =15'b0;

   // m39_92 = W*in
   wire signed [14:0] m39_92;
   assign m39_92 =15'b0;

   // m39_93 = W*in
   wire signed [14:0] m39_93;
   assign m39_93 =15'b0;

   // m39_94 = W*in
   wire signed [14:0] m39_94;
   assign m39_94 ={ {4{in39[14]}} , in39[14:4] };

   // m39_95 = W*in
   wire signed [14:0] m39_95;
   assign m39_95 ={ {3{in39[14]}} , in39[14:3] };

   // m39_96 = W*in
   wire signed [14:0] m39_96;
   assign m39_96 =15'b0;

   // m39_97 = W*in
   wire signed [14:0] m39_97;
   assign m39_97 =15'b0;

   // m39_98 = W*in
   wire signed [14:0] m39_98;
   assign m39_98 ={ {3{in39[14]}} , in39[14:3] };

   // m39_99 = W*in
   wire signed [14:0] m39_99;
   assign m39_99 =15'b0;

   // m39_100 = W*in
   wire signed [14:0] m39_100;
   assign m39_100 =15'b0;

   // m40_1 = W*in
   wire signed [14:0] m40_1;
   assign m40_1 =15'b0;

   // m40_2 = W*in
   wire signed [14:0] m40_2;
   assign m40_2 =15'b0;

   // m40_3 = W*in
   wire signed [14:0] m40_3;
   assign m40_3 =15'b0;

   // m40_4 = W*in
   wire signed [14:0] m40_4;
   assign m40_4 =15'b0;

   // m40_5 = W*in
   wire signed [14:0] m40_5;
   assign m40_5 ={ {3{in40[14]}} , in40[14:3] };

   // m40_6 = W*in
   wire signed [14:0] m40_6;
   assign m40_6 =15'b0;

   // m40_7 = W*in
   wire signed [14:0] m40_7;
   assign m40_7 =15'b0;

   // m40_8 = W*in
   wire signed [14:0] m40_8;
   assign m40_8 =15'b0;

   // m40_9 = W*in
   wire signed [14:0] m40_9;
   assign m40_9 =15'b0;

   // m40_10 = W*in
   wire signed [14:0] m40_10;
   assign m40_10 ={ {3{in40[14]}} , in40[14:3] };

   // m40_11 = W*in
   wire signed [14:0] m40_11;
   assign m40_11 ={ {3{neg40[14]}} , neg40[14:3] };

   // m40_12 = W*in
   wire signed [14:0] m40_12;
   assign m40_12 =15'b0;

   // m40_13 = W*in
   wire signed [14:0] m40_13;
   assign m40_13 =15'b0;

   // m40_14 = W*in
   wire signed [14:0] m40_14;
   assign m40_14 =15'b0;

   // m40_15 = W*in
   wire signed [14:0] m40_15;
   assign m40_15 =15'b0;

   // m40_16 = W*in
   wire signed [14:0] m40_16;
   assign m40_16 =15'b0;

   // m40_17 = W*in
   wire signed [14:0] m40_17;
   assign m40_17 ={ {3{neg40[14]}} , neg40[14:3] };

   // m40_18 = W*in
   wire signed [14:0] m40_18;
   assign m40_18 =15'b0;

   // m40_19 = W*in
   wire signed [14:0] m40_19;
   assign m40_19 ={ {4{in40[14]}} , in40[14:4] };

   // m40_20 = W*in
   wire signed [14:0] m40_20;
   assign m40_20 =15'b0;

   // m40_21 = W*in
   wire signed [14:0] m40_21;
   assign m40_21 =15'b0;

   // m40_22 = W*in
   wire signed [14:0] m40_22;
   assign m40_22 =15'b0;

   // m40_23 = W*in
   wire signed [14:0] m40_23;
   assign m40_23 =15'b0;

   // m40_24 = W*in
   wire signed [14:0] m40_24;
   assign m40_24 =15'b0;

   // m40_25 = W*in
   wire signed [14:0] m40_25;
   assign m40_25 =15'b0;

   // m40_26 = W*in
   wire signed [14:0] m40_26;
   assign m40_26 =15'b0;

   // m40_27 = W*in
   wire signed [14:0] m40_27;
   assign m40_27 ={ {3{in40[14]}} , in40[14:3] };

   // m40_28 = W*in
   wire signed [14:0] m40_28;
   assign m40_28 =15'b0;

   // m40_29 = W*in
   wire signed [14:0] m40_29;
   assign m40_29 =15'b0;

   // m40_30 = W*in
   wire signed [14:0] m40_30;
   assign m40_30 =15'b0;

   // m40_31 = W*in
   wire signed [14:0] m40_31;
   assign m40_31 =15'b0;

   // m40_32 = W*in
   wire signed [14:0] m40_32;
   assign m40_32 =15'b0;

   // m40_33 = W*in
   wire signed [14:0] m40_33;
   assign m40_33 =15'b0;

   // m40_34 = W*in
   wire signed [14:0] m40_34;
   assign m40_34 =15'b0;

   // m40_35 = W*in
   wire signed [14:0] m40_35;
   assign m40_35 =15'b0;

   // m40_36 = W*in
   wire signed [14:0] m40_36;
   assign m40_36 =15'b0;

   // m40_37 = W*in
   wire signed [14:0] m40_37;
   assign m40_37 =15'b0;

   // m40_38 = W*in
   wire signed [14:0] m40_38;
   assign m40_38 =15'b0;

   // m40_39 = W*in
   wire signed [14:0] m40_39;
   assign m40_39 =15'b0;

   // m40_40 = W*in
   wire signed [14:0] m40_40;
   assign m40_40 =15'b0;

   // m40_41 = W*in
   wire signed [14:0] m40_41;
   assign m40_41 ={ {3{neg40[14]}} , neg40[14:3] };

   // m40_42 = W*in
   wire signed [14:0] m40_42;
   assign m40_42 =15'b0;

   // m40_43 = W*in
   wire signed [14:0] m40_43;
   assign m40_43 ={ {3{in40[14]}} , in40[14:3] };

   // m40_44 = W*in
   wire signed [14:0] m40_44;
   assign m40_44 =15'b0;

   // m40_45 = W*in
   wire signed [14:0] m40_45;
   assign m40_45 =15'b0;

   // m40_46 = W*in
   wire signed [14:0] m40_46;
   assign m40_46 ={ {3{in40[14]}} , in40[14:3] };

   // m40_47 = W*in
   wire signed [14:0] m40_47;
   assign m40_47 =15'b0;

   // m40_48 = W*in
   wire signed [14:0] m40_48;
   assign m40_48 =15'b0;

   // m40_49 = W*in
   wire signed [14:0] m40_49;
   assign m40_49 =15'b0;

   // m40_50 = W*in
   wire signed [14:0] m40_50;
   assign m40_50 ={ {3{neg40[14]}} , neg40[14:3] };

   // m40_51 = W*in
   wire signed [14:0] m40_51;
   assign m40_51 =15'b0;

   // m40_52 = W*in
   wire signed [14:0] m40_52;
   assign m40_52 =15'b0;

   // m40_53 = W*in
   wire signed [14:0] m40_53;
   assign m40_53 =15'b0;

   // m40_54 = W*in
   wire signed [14:0] m40_54;
   assign m40_54 =15'b0;

   // m40_55 = W*in
   wire signed [14:0] m40_55;
   assign m40_55 =15'b0;

   // m40_56 = W*in
   wire signed [14:0] m40_56;
   assign m40_56 =15'b0;

   // m40_57 = W*in
   wire signed [14:0] m40_57;
   assign m40_57 =15'b0;

   // m40_58 = W*in
   wire signed [14:0] m40_58;
   assign m40_58 =15'b0;

   // m40_59 = W*in
   wire signed [14:0] m40_59;
   assign m40_59 ={ {4{in40[14]}} , in40[14:4] };

   // m40_60 = W*in
   wire signed [14:0] m40_60;
   assign m40_60 ={ {3{neg40[14]}} , neg40[14:3] };

   // m40_61 = W*in
   wire signed [14:0] m40_61;
   assign m40_61 =15'b0;

   // m40_62 = W*in
   wire signed [14:0] m40_62;
   assign m40_62 =15'b0;

   // m40_63 = W*in
   wire signed [14:0] m40_63;
   assign m40_63 ={ {3{in40[14]}} , in40[14:3] };

   // m40_64 = W*in
   wire signed [14:0] m40_64;
   assign m40_64 =15'b0;

   // m40_65 = W*in
   wire signed [14:0] m40_65;
   assign m40_65 ={ {3{in40[14]}} , in40[14:3] };

   // m40_66 = W*in
   wire signed [14:0] m40_66;
   assign m40_66 ={ {4{in40[14]}} , in40[14:4] };

   // m40_67 = W*in
   wire signed [14:0] m40_67;
   assign m40_67 =15'b0;

   // m40_68 = W*in
   wire signed [14:0] m40_68;
   assign m40_68 =15'b0;

   // m40_69 = W*in
   wire signed [14:0] m40_69;
   assign m40_69 =15'b0;

   // m40_70 = W*in
   wire signed [14:0] m40_70;
   assign m40_70 ={ {4{neg40[14]}} , neg40[14:4] };

   // m40_71 = W*in
   wire signed [14:0] m40_71;
   assign m40_71 =15'b0;

   // m40_72 = W*in
   wire signed [14:0] m40_72;
   assign m40_72 =15'b0;

   // m40_73 = W*in
   wire signed [14:0] m40_73;
   assign m40_73 =15'b0;

   // m40_74 = W*in
   wire signed [14:0] m40_74;
   assign m40_74 =15'b0;

   // m40_75 = W*in
   wire signed [14:0] m40_75;
   assign m40_75 =15'b0;

   // m40_76 = W*in
   wire signed [14:0] m40_76;
   assign m40_76 ={ {3{in40[14]}} , in40[14:3] };

   // m40_77 = W*in
   wire signed [14:0] m40_77;
   assign m40_77 =15'b0;

   // m40_78 = W*in
   wire signed [14:0] m40_78;
   assign m40_78 =15'b0;

   // m40_79 = W*in
   wire signed [14:0] m40_79;
   assign m40_79 ={ {4{in40[14]}} , in40[14:4] };

   // m40_80 = W*in
   wire signed [14:0] m40_80;
   assign m40_80 =15'b0;

   // m40_81 = W*in
   wire signed [14:0] m40_81;
   assign m40_81 =15'b0;

   // m40_82 = W*in
   wire signed [14:0] m40_82;
   assign m40_82 ={ {3{in40[14]}} , in40[14:3] };

   // m40_83 = W*in
   wire signed [14:0] m40_83;
   assign m40_83 =15'b0;

   // m40_84 = W*in
   wire signed [14:0] m40_84;
   assign m40_84 =15'b0;

   // m40_85 = W*in
   wire signed [14:0] m40_85;
   assign m40_85 =15'b0;

   // m40_86 = W*in
   wire signed [14:0] m40_86;
   assign m40_86 =15'b0;

   // m40_87 = W*in
   wire signed [14:0] m40_87;
   assign m40_87 =15'b0;

   // m40_88 = W*in
   wire signed [14:0] m40_88;
   assign m40_88 =15'b0;

   // m40_89 = W*in
   wire signed [14:0] m40_89;
   assign m40_89 =15'b0;

   // m40_90 = W*in
   wire signed [14:0] m40_90;
   assign m40_90 =15'b0;

   // m40_91 = W*in
   wire signed [14:0] m40_91;
   assign m40_91 =15'b0;

   // m40_92 = W*in
   wire signed [14:0] m40_92;
   assign m40_92 =15'b0;

   // m40_93 = W*in
   wire signed [14:0] m40_93;
   assign m40_93 =15'b0;

   // m40_94 = W*in
   wire signed [14:0] m40_94;
   assign m40_94 =15'b0;

   // m40_95 = W*in
   wire signed [14:0] m40_95;
   assign m40_95 =15'b0;

   // m40_96 = W*in
   wire signed [14:0] m40_96;
   assign m40_96 =15'b0;

   // m40_97 = W*in
   wire signed [14:0] m40_97;
   assign m40_97 ={ {3{in40[14]}} , in40[14:3] };

   // m40_98 = W*in
   wire signed [14:0] m40_98;
   assign m40_98 =15'b0;

   // m40_99 = W*in
   wire signed [14:0] m40_99;
   assign m40_99 =15'b0;

   // m40_100 = W*in
   wire signed [14:0] m40_100;
   assign m40_100 =15'b0;

   // m41_1 = W*in
   wire signed [14:0] m41_1;
   assign m41_1 =15'b0;

   // m41_2 = W*in
   wire signed [14:0] m41_2;
   assign m41_2 =15'b0;

   // m41_3 = W*in
   wire signed [14:0] m41_3;
   assign m41_3 =15'b0;

   // m41_4 = W*in
   wire signed [14:0] m41_4;
   assign m41_4 =15'b0;

   // m41_5 = W*in
   wire signed [14:0] m41_5;
   assign m41_5 =15'b0;

   // m41_6 = W*in
   wire signed [14:0] m41_6;
   assign m41_6 =15'b0;

   // m41_7 = W*in
   wire signed [14:0] m41_7;
   assign m41_7 ={ {3{in41[14]}} , in41[14:3] };

   // m41_8 = W*in
   wire signed [14:0] m41_8;
   assign m41_8 =15'b0;

   // m41_9 = W*in
   wire signed [14:0] m41_9;
   assign m41_9 =15'b0;

   // m41_10 = W*in
   wire signed [14:0] m41_10;
   assign m41_10 =15'b0;

   // m41_11 = W*in
   wire signed [14:0] m41_11;
   assign m41_11 =15'b0;

   // m41_12 = W*in
   wire signed [14:0] m41_12;
   assign m41_12 =15'b0;

   // m41_13 = W*in
   wire signed [14:0] m41_13;
   assign m41_13 =15'b0;

   // m41_14 = W*in
   wire signed [14:0] m41_14;
   assign m41_14 ={ {3{in41[14]}} , in41[14:3] };

   // m41_15 = W*in
   wire signed [14:0] m41_15;
   assign m41_15 =15'b0;

   // m41_16 = W*in
   wire signed [14:0] m41_16;
   assign m41_16 =15'b0;

   // m41_17 = W*in
   wire signed [14:0] m41_17;
   assign m41_17 ={ {3{in41[14]}} , in41[14:3] };

   // m41_18 = W*in
   wire signed [14:0] m41_18;
   assign m41_18 =15'b0;

   // m41_19 = W*in
   wire signed [14:0] m41_19;
   assign m41_19 =15'b0;

   // m41_20 = W*in
   wire signed [14:0] m41_20;
   assign m41_20 ={ {4{neg41[14]}} , neg41[14:4] };

   // m41_21 = W*in
   wire signed [14:0] m41_21;
   assign m41_21 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_22 = W*in
   wire signed [14:0] m41_22;
   assign m41_22 =15'b0;

   // m41_23 = W*in
   wire signed [14:0] m41_23;
   assign m41_23 =15'b0;

   // m41_24 = W*in
   wire signed [14:0] m41_24;
   assign m41_24 =15'b0;

   // m41_25 = W*in
   wire signed [14:0] m41_25;
   assign m41_25 =15'b0;

   // m41_26 = W*in
   wire signed [14:0] m41_26;
   assign m41_26 =15'b0;

   // m41_27 = W*in
   wire signed [14:0] m41_27;
   assign m41_27 =15'b0;

   // m41_28 = W*in
   wire signed [14:0] m41_28;
   assign m41_28 =15'b0;

   // m41_29 = W*in
   wire signed [14:0] m41_29;
   assign m41_29 =15'b0;

   // m41_30 = W*in
   wire signed [14:0] m41_30;
   assign m41_30 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_31 = W*in
   wire signed [14:0] m41_31;
   assign m41_31 =15'b0;

   // m41_32 = W*in
   wire signed [14:0] m41_32;
   assign m41_32 ={ {3{in41[14]}} , in41[14:3] };

   // m41_33 = W*in
   wire signed [14:0] m41_33;
   assign m41_33 ={ {3{in41[14]}} , in41[14:3] };

   // m41_34 = W*in
   wire signed [14:0] m41_34;
   assign m41_34 =15'b0;

   // m41_35 = W*in
   wire signed [14:0] m41_35;
   assign m41_35 ={ {3{in41[14]}} , in41[14:3] };

   // m41_36 = W*in
   wire signed [14:0] m41_36;
   assign m41_36 =15'b0;

   // m41_37 = W*in
   wire signed [14:0] m41_37;
   assign m41_37 =15'b0;

   // m41_38 = W*in
   wire signed [14:0] m41_38;
   assign m41_38 =15'b0;

   // m41_39 = W*in
   wire signed [14:0] m41_39;
   assign m41_39 ={ {3{in41[14]}} , in41[14:3] };

   // m41_40 = W*in
   wire signed [14:0] m41_40;
   assign m41_40 ={ {3{in41[14]}} , in41[14:3] };

   // m41_41 = W*in
   wire signed [14:0] m41_41;
   assign m41_41 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_42 = W*in
   wire signed [14:0] m41_42;
   assign m41_42 ={ {3{in41[14]}} , in41[14:3] };

   // m41_43 = W*in
   wire signed [14:0] m41_43;
   assign m41_43 =15'b0;

   // m41_44 = W*in
   wire signed [14:0] m41_44;
   assign m41_44 ={ {3{in41[14]}} , in41[14:3] };

   // m41_45 = W*in
   wire signed [14:0] m41_45;
   assign m41_45 =15'b0;

   // m41_46 = W*in
   wire signed [14:0] m41_46;
   assign m41_46 =15'b0;

   // m41_47 = W*in
   wire signed [14:0] m41_47;
   assign m41_47 =15'b0;

   // m41_48 = W*in
   wire signed [14:0] m41_48;
   assign m41_48 =15'b0;

   // m41_49 = W*in
   wire signed [14:0] m41_49;
   assign m41_49 =15'b0;

   // m41_50 = W*in
   wire signed [14:0] m41_50;
   assign m41_50 =15'b0;

   // m41_51 = W*in
   wire signed [14:0] m41_51;
   assign m41_51 =15'b0;

   // m41_52 = W*in
   wire signed [14:0] m41_52;
   assign m41_52 =15'b0;

   // m41_53 = W*in
   wire signed [14:0] m41_53;
   assign m41_53 =15'b0;

   // m41_54 = W*in
   wire signed [14:0] m41_54;
   assign m41_54 ={ {3{in41[14]}} , in41[14:3] };

   // m41_55 = W*in
   wire signed [14:0] m41_55;
   assign m41_55 =15'b0;

   // m41_56 = W*in
   wire signed [14:0] m41_56;
   assign m41_56 =15'b0;

   // m41_57 = W*in
   wire signed [14:0] m41_57;
   assign m41_57 ={ {3{in41[14]}} , in41[14:3] };

   // m41_58 = W*in
   wire signed [14:0] m41_58;
   assign m41_58 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_59 = W*in
   wire signed [14:0] m41_59;
   assign m41_59 =15'b0;

   // m41_60 = W*in
   wire signed [14:0] m41_60;
   assign m41_60 =15'b0;

   // m41_61 = W*in
   wire signed [14:0] m41_61;
   assign m41_61 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_62 = W*in
   wire signed [14:0] m41_62;
   assign m41_62 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_63 = W*in
   wire signed [14:0] m41_63;
   assign m41_63 =15'b0;

   // m41_64 = W*in
   wire signed [14:0] m41_64;
   assign m41_64 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_65 = W*in
   wire signed [14:0] m41_65;
   assign m41_65 =15'b0;

   // m41_66 = W*in
   wire signed [14:0] m41_66;
   assign m41_66 ={ {3{in41[14]}} , in41[14:3] };

   // m41_67 = W*in
   wire signed [14:0] m41_67;
   assign m41_67 =15'b0;

   // m41_68 = W*in
   wire signed [14:0] m41_68;
   assign m41_68 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_69 = W*in
   wire signed [14:0] m41_69;
   assign m41_69 =15'b0;

   // m41_70 = W*in
   wire signed [14:0] m41_70;
   assign m41_70 ={ {4{in41[14]}} , in41[14:4] };

   // m41_71 = W*in
   wire signed [14:0] m41_71;
   assign m41_71 =15'b0;

   // m41_72 = W*in
   wire signed [14:0] m41_72;
   assign m41_72 =15'b0;

   // m41_73 = W*in
   wire signed [14:0] m41_73;
   assign m41_73 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_74 = W*in
   wire signed [14:0] m41_74;
   assign m41_74 =15'b0;

   // m41_75 = W*in
   wire signed [14:0] m41_75;
   assign m41_75 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_76 = W*in
   wire signed [14:0] m41_76;
   assign m41_76 =15'b0;

   // m41_77 = W*in
   wire signed [14:0] m41_77;
   assign m41_77 =15'b0;

   // m41_78 = W*in
   wire signed [14:0] m41_78;
   assign m41_78 =15'b0;

   // m41_79 = W*in
   wire signed [14:0] m41_79;
   assign m41_79 =15'b0;

   // m41_80 = W*in
   wire signed [14:0] m41_80;
   assign m41_80 =15'b0;

   // m41_81 = W*in
   wire signed [14:0] m41_81;
   assign m41_81 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_82 = W*in
   wire signed [14:0] m41_82;
   assign m41_82 =15'b0;

   // m41_83 = W*in
   wire signed [14:0] m41_83;
   assign m41_83 =15'b0;

   // m41_84 = W*in
   wire signed [14:0] m41_84;
   assign m41_84 =15'b0;

   // m41_85 = W*in
   wire signed [14:0] m41_85;
   assign m41_85 =15'b0;

   // m41_86 = W*in
   wire signed [14:0] m41_86;
   assign m41_86 =15'b0;

   // m41_87 = W*in
   wire signed [14:0] m41_87;
   assign m41_87 =15'b0;

   // m41_88 = W*in
   wire signed [14:0] m41_88;
   assign m41_88 =15'b0;

   // m41_89 = W*in
   wire signed [14:0] m41_89;
   assign m41_89 =15'b0;

   // m41_90 = W*in
   wire signed [14:0] m41_90;
   assign m41_90 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_91 = W*in
   wire signed [14:0] m41_91;
   assign m41_91 =15'b0;

   // m41_92 = W*in
   wire signed [14:0] m41_92;
   assign m41_92 ={ {3{neg41[14]}} , neg41[14:3] };

   // m41_93 = W*in
   wire signed [14:0] m41_93;
   assign m41_93 =15'b0;

   // m41_94 = W*in
   wire signed [14:0] m41_94;
   assign m41_94 ={ {3{in41[14]}} , in41[14:3] };

   // m41_95 = W*in
   wire signed [14:0] m41_95;
   assign m41_95 =15'b0;

   // m41_96 = W*in
   wire signed [14:0] m41_96;
   assign m41_96 =15'b0;

   // m41_97 = W*in
   wire signed [14:0] m41_97;
   assign m41_97 =15'b0;

   // m41_98 = W*in
   wire signed [14:0] m41_98;
   assign m41_98 =15'b0;

   // m41_99 = W*in
   wire signed [14:0] m41_99;
   assign m41_99 =15'b0;

   // m41_100 = W*in
   wire signed [14:0] m41_100;
   assign m41_100 ={ {3{in41[14]}} , in41[14:3] };

   // m42_1 = W*in
   wire signed [14:0] m42_1;
   assign m42_1 =15'b0;

   // m42_2 = W*in
   wire signed [14:0] m42_2;
   assign m42_2 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_3 = W*in
   wire signed [14:0] m42_3;
   assign m42_3 =15'b0;

   // m42_4 = W*in
   wire signed [14:0] m42_4;
   assign m42_4 =15'b0;

   // m42_5 = W*in
   wire signed [14:0] m42_5;
   assign m42_5 =15'b0;

   // m42_6 = W*in
   wire signed [14:0] m42_6;
   assign m42_6 =15'b0;

   // m42_7 = W*in
   wire signed [14:0] m42_7;
   assign m42_7 =15'b0;

   // m42_8 = W*in
   wire signed [14:0] m42_8;
   assign m42_8 ={ {3{in42[14]}} , in42[14:3] };

   // m42_9 = W*in
   wire signed [14:0] m42_9;
   assign m42_9 =15'b0;

   // m42_10 = W*in
   wire signed [14:0] m42_10;
   assign m42_10 =15'b0;

   // m42_11 = W*in
   wire signed [14:0] m42_11;
   assign m42_11 ={ {3{in42[14]}} , in42[14:3] };

   // m42_12 = W*in
   wire signed [14:0] m42_12;
   assign m42_12 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_13 = W*in
   wire signed [14:0] m42_13;
   assign m42_13 =15'b0;

   // m42_14 = W*in
   wire signed [14:0] m42_14;
   assign m42_14 =15'b0;

   // m42_15 = W*in
   wire signed [14:0] m42_15;
   assign m42_15 =15'b0;

   // m42_16 = W*in
   wire signed [14:0] m42_16;
   assign m42_16 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_17 = W*in
   wire signed [14:0] m42_17;
   assign m42_17 =15'b0;

   // m42_18 = W*in
   wire signed [14:0] m42_18;
   assign m42_18 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_19 = W*in
   wire signed [14:0] m42_19;
   assign m42_19 ={ {4{in42[14]}} , in42[14:4] };

   // m42_20 = W*in
   wire signed [14:0] m42_20;
   assign m42_20 ={ {4{neg42[14]}} , neg42[14:4] };

   // m42_21 = W*in
   wire signed [14:0] m42_21;
   assign m42_21 ={ {4{in42[14]}} , in42[14:4] };

   // m42_22 = W*in
   wire signed [14:0] m42_22;
   assign m42_22 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_23 = W*in
   wire signed [14:0] m42_23;
   assign m42_23 =15'b0;

   // m42_24 = W*in
   wire signed [14:0] m42_24;
   assign m42_24 =15'b0;

   // m42_25 = W*in
   wire signed [14:0] m42_25;
   assign m42_25 ={ {3{in42[14]}} , in42[14:3] };

   // m42_26 = W*in
   wire signed [14:0] m42_26;
   assign m42_26 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_27 = W*in
   wire signed [14:0] m42_27;
   assign m42_27 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_28 = W*in
   wire signed [14:0] m42_28;
   assign m42_28 =15'b0;

   // m42_29 = W*in
   wire signed [14:0] m42_29;
   assign m42_29 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_30 = W*in
   wire signed [14:0] m42_30;
   assign m42_30 =15'b0;

   // m42_31 = W*in
   wire signed [14:0] m42_31;
   assign m42_31 =15'b0;

   // m42_32 = W*in
   wire signed [14:0] m42_32;
   assign m42_32 =15'b0;

   // m42_33 = W*in
   wire signed [14:0] m42_33;
   assign m42_33 ={ {4{neg42[14]}} , neg42[14:4] };

   // m42_34 = W*in
   wire signed [14:0] m42_34;
   assign m42_34 =15'b0;

   // m42_35 = W*in
   wire signed [14:0] m42_35;
   assign m42_35 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_36 = W*in
   wire signed [14:0] m42_36;
   assign m42_36 =15'b0;

   // m42_37 = W*in
   wire signed [14:0] m42_37;
   assign m42_37 ={ {3{in42[14]}} , in42[14:3] };

   // m42_38 = W*in
   wire signed [14:0] m42_38;
   assign m42_38 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_39 = W*in
   wire signed [14:0] m42_39;
   assign m42_39 =15'b0;

   // m42_40 = W*in
   wire signed [14:0] m42_40;
   assign m42_40 =15'b0;

   // m42_41 = W*in
   wire signed [14:0] m42_41;
   assign m42_41 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_42 = W*in
   wire signed [14:0] m42_42;
   assign m42_42 =15'b0;

   // m42_43 = W*in
   wire signed [14:0] m42_43;
   assign m42_43 =15'b0;

   // m42_44 = W*in
   wire signed [14:0] m42_44;
   assign m42_44 =15'b0;

   // m42_45 = W*in
   wire signed [14:0] m42_45;
   assign m42_45 =15'b0;

   // m42_46 = W*in
   wire signed [14:0] m42_46;
   assign m42_46 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_47 = W*in
   wire signed [14:0] m42_47;
   assign m42_47 ={ {3{in42[14]}} , in42[14:3] };

   // m42_48 = W*in
   wire signed [14:0] m42_48;
   assign m42_48 ={ {4{in42[14]}} , in42[14:4] };

   // m42_49 = W*in
   wire signed [14:0] m42_49;
   assign m42_49 ={ {3{in42[14]}} , in42[14:3] };

   // m42_50 = W*in
   wire signed [14:0] m42_50;
   assign m42_50 =15'b0;

   // m42_51 = W*in
   wire signed [14:0] m42_51;
   assign m42_51 ={ {3{in42[14]}} , in42[14:3] };

   // m42_52 = W*in
   wire signed [14:0] m42_52;
   assign m42_52 =15'b0;

   // m42_53 = W*in
   wire signed [14:0] m42_53;
   assign m42_53 ={ {3{in42[14]}} , in42[14:3] };

   // m42_54 = W*in
   wire signed [14:0] m42_54;
   assign m42_54 ={ {3{in42[14]}} , in42[14:3] };

   // m42_55 = W*in
   wire signed [14:0] m42_55;
   assign m42_55 =15'b0;

   // m42_56 = W*in
   wire signed [14:0] m42_56;
   assign m42_56 =15'b0;

   // m42_57 = W*in
   wire signed [14:0] m42_57;
   assign m42_57 =15'b0;

   // m42_58 = W*in
   wire signed [14:0] m42_58;
   assign m42_58 =15'b0;

   // m42_59 = W*in
   wire signed [14:0] m42_59;
   assign m42_59 ={ {3{in42[14]}} , in42[14:3] };

   // m42_60 = W*in
   wire signed [14:0] m42_60;
   assign m42_60 ={ {4{in42[14]}} , in42[14:4] };

   // m42_61 = W*in
   wire signed [14:0] m42_61;
   assign m42_61 =15'b0;

   // m42_62 = W*in
   wire signed [14:0] m42_62;
   assign m42_62 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_63 = W*in
   wire signed [14:0] m42_63;
   assign m42_63 =15'b0;

   // m42_64 = W*in
   wire signed [14:0] m42_64;
   assign m42_64 ={ {4{neg42[14]}} , neg42[14:4] };

   // m42_65 = W*in
   wire signed [14:0] m42_65;
   assign m42_65 ={ {4{neg42[14]}} , neg42[14:4] };

   // m42_66 = W*in
   wire signed [14:0] m42_66;
   assign m42_66 ={ {4{neg42[14]}} , neg42[14:4] };

   // m42_67 = W*in
   wire signed [14:0] m42_67;
   assign m42_67 ={ {4{in42[14]}} , in42[14:4] };

   // m42_68 = W*in
   wire signed [14:0] m42_68;
   assign m42_68 =15'b0;

   // m42_69 = W*in
   wire signed [14:0] m42_69;
   assign m42_69 ={ {3{in42[14]}} , in42[14:3] };

   // m42_70 = W*in
   wire signed [14:0] m42_70;
   assign m42_70 ={ {4{in42[14]}} , in42[14:4] };

   // m42_71 = W*in
   wire signed [14:0] m42_71;
   assign m42_71 ={ {3{in42[14]}} , in42[14:3] };

   // m42_72 = W*in
   wire signed [14:0] m42_72;
   assign m42_72 ={ {3{in42[14]}} , in42[14:3] };

   // m42_73 = W*in
   wire signed [14:0] m42_73;
   assign m42_73 =15'b0;

   // m42_74 = W*in
   wire signed [14:0] m42_74;
   assign m42_74 ={ {4{neg42[14]}} , neg42[14:4] };

   // m42_75 = W*in
   wire signed [14:0] m42_75;
   assign m42_75 =15'b0;

   // m42_76 = W*in
   wire signed [14:0] m42_76;
   assign m42_76 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_77 = W*in
   wire signed [14:0] m42_77;
   assign m42_77 ={ {3{in42[14]}} , in42[14:3] };

   // m42_78 = W*in
   wire signed [14:0] m42_78;
   assign m42_78 =15'b0;

   // m42_79 = W*in
   wire signed [14:0] m42_79;
   assign m42_79 ={ {3{in42[14]}} , in42[14:3] };

   // m42_80 = W*in
   wire signed [14:0] m42_80;
   assign m42_80 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_81 = W*in
   wire signed [14:0] m42_81;
   assign m42_81 =15'b0;

   // m42_82 = W*in
   wire signed [14:0] m42_82;
   assign m42_82 =15'b0;

   // m42_83 = W*in
   wire signed [14:0] m42_83;
   assign m42_83 =15'b0;

   // m42_84 = W*in
   wire signed [14:0] m42_84;
   assign m42_84 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_85 = W*in
   wire signed [14:0] m42_85;
   assign m42_85 =15'b0;

   // m42_86 = W*in
   wire signed [14:0] m42_86;
   assign m42_86 =15'b0;

   // m42_87 = W*in
   wire signed [14:0] m42_87;
   assign m42_87 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_88 = W*in
   wire signed [14:0] m42_88;
   assign m42_88 =15'b0;

   // m42_89 = W*in
   wire signed [14:0] m42_89;
   assign m42_89 ={ {3{in42[14]}} , in42[14:3] };

   // m42_90 = W*in
   wire signed [14:0] m42_90;
   assign m42_90 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_91 = W*in
   wire signed [14:0] m42_91;
   assign m42_91 ={ {3{in42[14]}} , in42[14:3] };

   // m42_92 = W*in
   wire signed [14:0] m42_92;
   assign m42_92 ={ {3{in42[14]}} , in42[14:3] };

   // m42_93 = W*in
   wire signed [14:0] m42_93;
   assign m42_93 =15'b0;

   // m42_94 = W*in
   wire signed [14:0] m42_94;
   assign m42_94 =15'b0;

   // m42_95 = W*in
   wire signed [14:0] m42_95;
   assign m42_95 ={ {3{in42[14]}} , in42[14:3] };

   // m42_96 = W*in
   wire signed [14:0] m42_96;
   assign m42_96 =15'b0;

   // m42_97 = W*in
   wire signed [14:0] m42_97;
   assign m42_97 ={ {3{neg42[14]}} , neg42[14:3] };

   // m42_98 = W*in
   wire signed [14:0] m42_98;
   assign m42_98 ={ {3{in42[14]}} , in42[14:3] };

   // m42_99 = W*in
   wire signed [14:0] m42_99;
   assign m42_99 =15'b0;

   // m42_100 = W*in
   wire signed [14:0] m42_100;
   assign m42_100 =15'b0;

   // m43_1 = W*in
   wire signed [14:0] m43_1;
   assign m43_1 ={ {3{in43[14]}} , in43[14:3] };

   // m43_2 = W*in
   wire signed [14:0] m43_2;
   assign m43_2 =15'b0;

   // m43_3 = W*in
   wire signed [14:0] m43_3;
   assign m43_3 =15'b0;

   // m43_4 = W*in
   wire signed [14:0] m43_4;
   assign m43_4 =15'b0;

   // m43_5 = W*in
   wire signed [14:0] m43_5;
   assign m43_5 =15'b0;

   // m43_6 = W*in
   wire signed [14:0] m43_6;
   assign m43_6 =15'b0;

   // m43_7 = W*in
   wire signed [14:0] m43_7;
   assign m43_7 =15'b0;

   // m43_8 = W*in
   wire signed [14:0] m43_8;
   assign m43_8 =15'b0;

   // m43_9 = W*in
   wire signed [14:0] m43_9;
   assign m43_9 =15'b0;

   // m43_10 = W*in
   wire signed [14:0] m43_10;
   assign m43_10 =15'b0;

   // m43_11 = W*in
   wire signed [14:0] m43_11;
   assign m43_11 =15'b0;

   // m43_12 = W*in
   wire signed [14:0] m43_12;
   assign m43_12 =15'b0;

   // m43_13 = W*in
   wire signed [14:0] m43_13;
   assign m43_13 ={ {4{in43[14]}} , in43[14:4] };

   // m43_14 = W*in
   wire signed [14:0] m43_14;
   assign m43_14 =15'b0;

   // m43_15 = W*in
   wire signed [14:0] m43_15;
   assign m43_15 =15'b0;

   // m43_16 = W*in
   wire signed [14:0] m43_16;
   assign m43_16 =15'b0;

   // m43_17 = W*in
   wire signed [14:0] m43_17;
   assign m43_17 =15'b0;

   // m43_18 = W*in
   wire signed [14:0] m43_18;
   assign m43_18 =15'b0;

   // m43_19 = W*in
   wire signed [14:0] m43_19;
   assign m43_19 =15'b0;

   // m43_20 = W*in
   wire signed [14:0] m43_20;
   assign m43_20 =15'b0;

   // m43_21 = W*in
   wire signed [14:0] m43_21;
   assign m43_21 =15'b0;

   // m43_22 = W*in
   wire signed [14:0] m43_22;
   assign m43_22 =15'b0;

   // m43_23 = W*in
   wire signed [14:0] m43_23;
   assign m43_23 =15'b0;

   // m43_24 = W*in
   wire signed [14:0] m43_24;
   assign m43_24 =15'b0;

   // m43_25 = W*in
   wire signed [14:0] m43_25;
   assign m43_25 =15'b0;

   // m43_26 = W*in
   wire signed [14:0] m43_26;
   assign m43_26 =15'b0;

   // m43_27 = W*in
   wire signed [14:0] m43_27;
   assign m43_27 =15'b0;

   // m43_28 = W*in
   wire signed [14:0] m43_28;
   assign m43_28 =15'b0;

   // m43_29 = W*in
   wire signed [14:0] m43_29;
   assign m43_29 ={ {4{neg43[14]}} , neg43[14:4] };

   // m43_30 = W*in
   wire signed [14:0] m43_30;
   assign m43_30 =15'b0;

   // m43_31 = W*in
   wire signed [14:0] m43_31;
   assign m43_31 =15'b0;

   // m43_32 = W*in
   wire signed [14:0] m43_32;
   assign m43_32 =15'b0;

   // m43_33 = W*in
   wire signed [14:0] m43_33;
   assign m43_33 =15'b0;

   // m43_34 = W*in
   wire signed [14:0] m43_34;
   assign m43_34 =15'b0;

   // m43_35 = W*in
   wire signed [14:0] m43_35;
   assign m43_35 =15'b0;

   // m43_36 = W*in
   wire signed [14:0] m43_36;
   assign m43_36 =15'b0;

   // m43_37 = W*in
   wire signed [14:0] m43_37;
   assign m43_37 =15'b0;

   // m43_38 = W*in
   wire signed [14:0] m43_38;
   assign m43_38 =15'b0;

   // m43_39 = W*in
   wire signed [14:0] m43_39;
   assign m43_39 ={ {3{neg43[14]}} , neg43[14:3] };

   // m43_40 = W*in
   wire signed [14:0] m43_40;
   assign m43_40 =15'b0;

   // m43_41 = W*in
   wire signed [14:0] m43_41;
   assign m43_41 =15'b0;

   // m43_42 = W*in
   wire signed [14:0] m43_42;
   assign m43_42 =15'b0;

   // m43_43 = W*in
   wire signed [14:0] m43_43;
   assign m43_43 =15'b0;

   // m43_44 = W*in
   wire signed [14:0] m43_44;
   assign m43_44 =15'b0;

   // m43_45 = W*in
   wire signed [14:0] m43_45;
   assign m43_45 =15'b0;

   // m43_46 = W*in
   wire signed [14:0] m43_46;
   assign m43_46 =15'b0;

   // m43_47 = W*in
   wire signed [14:0] m43_47;
   assign m43_47 =15'b0;

   // m43_48 = W*in
   wire signed [14:0] m43_48;
   assign m43_48 =15'b0;

   // m43_49 = W*in
   wire signed [14:0] m43_49;
   assign m43_49 =15'b0;

   // m43_50 = W*in
   wire signed [14:0] m43_50;
   assign m43_50 ={ {3{in43[14]}} , in43[14:3] };

   // m43_51 = W*in
   wire signed [14:0] m43_51;
   assign m43_51 =15'b0;

   // m43_52 = W*in
   wire signed [14:0] m43_52;
   assign m43_52 =15'b0;

   // m43_53 = W*in
   wire signed [14:0] m43_53;
   assign m43_53 =15'b0;

   // m43_54 = W*in
   wire signed [14:0] m43_54;
   assign m43_54 =15'b0;

   // m43_55 = W*in
   wire signed [14:0] m43_55;
   assign m43_55 =15'b0;

   // m43_56 = W*in
   wire signed [14:0] m43_56;
   assign m43_56 =15'b0;

   // m43_57 = W*in
   wire signed [14:0] m43_57;
   assign m43_57 =15'b0;

   // m43_58 = W*in
   wire signed [14:0] m43_58;
   assign m43_58 =15'b0;

   // m43_59 = W*in
   wire signed [14:0] m43_59;
   assign m43_59 =15'b0;

   // m43_60 = W*in
   wire signed [14:0] m43_60;
   assign m43_60 ={ {3{neg43[14]}} , neg43[14:3] };

   // m43_61 = W*in
   wire signed [14:0] m43_61;
   assign m43_61 =15'b0;

   // m43_62 = W*in
   wire signed [14:0] m43_62;
   assign m43_62 ={ {3{in43[14]}} , in43[14:3] };

   // m43_63 = W*in
   wire signed [14:0] m43_63;
   assign m43_63 =15'b0;

   // m43_64 = W*in
   wire signed [14:0] m43_64;
   assign m43_64 =15'b0;

   // m43_65 = W*in
   wire signed [14:0] m43_65;
   assign m43_65 =15'b0;

   // m43_66 = W*in
   wire signed [14:0] m43_66;
   assign m43_66 =15'b0;

   // m43_67 = W*in
   wire signed [14:0] m43_67;
   assign m43_67 =15'b0;

   // m43_68 = W*in
   wire signed [14:0] m43_68;
   assign m43_68 =15'b0;

   // m43_69 = W*in
   wire signed [14:0] m43_69;
   assign m43_69 =15'b0;

   // m43_70 = W*in
   wire signed [14:0] m43_70;
   assign m43_70 =15'b0;

   // m43_71 = W*in
   wire signed [14:0] m43_71;
   assign m43_71 =15'b0;

   // m43_72 = W*in
   wire signed [14:0] m43_72;
   assign m43_72 =15'b0;

   // m43_73 = W*in
   wire signed [14:0] m43_73;
   assign m43_73 ={ {3{in43[14]}} , in43[14:3] };

   // m43_74 = W*in
   wire signed [14:0] m43_74;
   assign m43_74 =15'b0;

   // m43_75 = W*in
   wire signed [14:0] m43_75;
   assign m43_75 ={ {3{in43[14]}} , in43[14:3] };

   // m43_76 = W*in
   wire signed [14:0] m43_76;
   assign m43_76 =15'b0;

   // m43_77 = W*in
   wire signed [14:0] m43_77;
   assign m43_77 =15'b0;

   // m43_78 = W*in
   wire signed [14:0] m43_78;
   assign m43_78 =15'b0;

   // m43_79 = W*in
   wire signed [14:0] m43_79;
   assign m43_79 =15'b0;

   // m43_80 = W*in
   wire signed [14:0] m43_80;
   assign m43_80 =15'b0;

   // m43_81 = W*in
   wire signed [14:0] m43_81;
   assign m43_81 =15'b0;

   // m43_82 = W*in
   wire signed [14:0] m43_82;
   assign m43_82 =15'b0;

   // m43_83 = W*in
   wire signed [14:0] m43_83;
   assign m43_83 =15'b0;

   // m43_84 = W*in
   wire signed [14:0] m43_84;
   assign m43_84 =15'b0;

   // m43_85 = W*in
   wire signed [14:0] m43_85;
   assign m43_85 =15'b0;

   // m43_86 = W*in
   wire signed [14:0] m43_86;
   assign m43_86 =15'b0;

   // m43_87 = W*in
   wire signed [14:0] m43_87;
   assign m43_87 =15'b0;

   // m43_88 = W*in
   wire signed [14:0] m43_88;
   assign m43_88 =15'b0;

   // m43_89 = W*in
   wire signed [14:0] m43_89;
   assign m43_89 =15'b0;

   // m43_90 = W*in
   wire signed [14:0] m43_90;
   assign m43_90 =15'b0;

   // m43_91 = W*in
   wire signed [14:0] m43_91;
   assign m43_91 =15'b0;

   // m43_92 = W*in
   wire signed [14:0] m43_92;
   assign m43_92 ={ {3{in43[14]}} , in43[14:3] };

   // m43_93 = W*in
   wire signed [14:0] m43_93;
   assign m43_93 =15'b0;

   // m43_94 = W*in
   wire signed [14:0] m43_94;
   assign m43_94 =15'b0;

   // m43_95 = W*in
   wire signed [14:0] m43_95;
   assign m43_95 =15'b0;

   // m43_96 = W*in
   wire signed [14:0] m43_96;
   assign m43_96 =15'b0;

   // m43_97 = W*in
   wire signed [14:0] m43_97;
   assign m43_97 =15'b0;

   // m43_98 = W*in
   wire signed [14:0] m43_98;
   assign m43_98 =15'b0;

   // m43_99 = W*in
   wire signed [14:0] m43_99;
   assign m43_99 =15'b0;

   // m43_100 = W*in
   wire signed [14:0] m43_100;
   assign m43_100 =15'b0;

   // m44_1 = W*in
   wire signed [14:0] m44_1;
   assign m44_1 =15'b0;

   // m44_2 = W*in
   wire signed [14:0] m44_2;
   assign m44_2 =15'b0;

   // m44_3 = W*in
   wire signed [14:0] m44_3;
   assign m44_3 ={ {3{neg44[14]}} , neg44[14:3] };

   // m44_4 = W*in
   wire signed [14:0] m44_4;
   assign m44_4 =15'b0;

   // m44_5 = W*in
   wire signed [14:0] m44_5;
   assign m44_5 =15'b0;

   // m44_6 = W*in
   wire signed [14:0] m44_6;
   assign m44_6 =15'b0;

   // m44_7 = W*in
   wire signed [14:0] m44_7;
   assign m44_7 =15'b0;

   // m44_8 = W*in
   wire signed [14:0] m44_8;
   assign m44_8 =15'b0;

   // m44_9 = W*in
   wire signed [14:0] m44_9;
   assign m44_9 =15'b0;

   // m44_10 = W*in
   wire signed [14:0] m44_10;
   assign m44_10 =15'b0;

   // m44_11 = W*in
   wire signed [14:0] m44_11;
   assign m44_11 =15'b0;

   // m44_12 = W*in
   wire signed [14:0] m44_12;
   assign m44_12 =15'b0;

   // m44_13 = W*in
   wire signed [14:0] m44_13;
   assign m44_13 =15'b0;

   // m44_14 = W*in
   wire signed [14:0] m44_14;
   assign m44_14 =15'b0;

   // m44_15 = W*in
   wire signed [14:0] m44_15;
   assign m44_15 =15'b0;

   // m44_16 = W*in
   wire signed [14:0] m44_16;
   assign m44_16 =15'b0;

   // m44_17 = W*in
   wire signed [14:0] m44_17;
   assign m44_17 =15'b0;

   // m44_18 = W*in
   wire signed [14:0] m44_18;
   assign m44_18 =15'b0;

   // m44_19 = W*in
   wire signed [14:0] m44_19;
   assign m44_19 =15'b0;

   // m44_20 = W*in
   wire signed [14:0] m44_20;
   assign m44_20 =15'b0;

   // m44_21 = W*in
   wire signed [14:0] m44_21;
   assign m44_21 ={ {3{in44[14]}} , in44[14:3] };

   // m44_22 = W*in
   wire signed [14:0] m44_22;
   assign m44_22 =15'b0;

   // m44_23 = W*in
   wire signed [14:0] m44_23;
   assign m44_23 =15'b0;

   // m44_24 = W*in
   wire signed [14:0] m44_24;
   assign m44_24 =15'b0;

   // m44_25 = W*in
   wire signed [14:0] m44_25;
   assign m44_25 =15'b0;

   // m44_26 = W*in
   wire signed [14:0] m44_26;
   assign m44_26 =15'b0;

   // m44_27 = W*in
   wire signed [14:0] m44_27;
   assign m44_27 =15'b0;

   // m44_28 = W*in
   wire signed [14:0] m44_28;
   assign m44_28 =15'b0;

   // m44_29 = W*in
   wire signed [14:0] m44_29;
   assign m44_29 =15'b0;

   // m44_30 = W*in
   wire signed [14:0] m44_30;
   assign m44_30 =15'b0;

   // m44_31 = W*in
   wire signed [14:0] m44_31;
   assign m44_31 =15'b0;

   // m44_32 = W*in
   wire signed [14:0] m44_32;
   assign m44_32 ={ {4{in44[14]}} , in44[14:4] };

   // m44_33 = W*in
   wire signed [14:0] m44_33;
   assign m44_33 ={ {4{neg44[14]}} , neg44[14:4] };

   // m44_34 = W*in
   wire signed [14:0] m44_34;
   assign m44_34 =15'b0;

   // m44_35 = W*in
   wire signed [14:0] m44_35;
   assign m44_35 =15'b0;

   // m44_36 = W*in
   wire signed [14:0] m44_36;
   assign m44_36 =15'b0;

   // m44_37 = W*in
   wire signed [14:0] m44_37;
   assign m44_37 =15'b0;

   // m44_38 = W*in
   wire signed [14:0] m44_38;
   assign m44_38 ={ {3{neg44[14]}} , neg44[14:3] };

   // m44_39 = W*in
   wire signed [14:0] m44_39;
   assign m44_39 =15'b0;

   // m44_40 = W*in
   wire signed [14:0] m44_40;
   assign m44_40 =15'b0;

   // m44_41 = W*in
   wire signed [14:0] m44_41;
   assign m44_41 =15'b0;

   // m44_42 = W*in
   wire signed [14:0] m44_42;
   assign m44_42 =15'b0;

   // m44_43 = W*in
   wire signed [14:0] m44_43;
   assign m44_43 =15'b0;

   // m44_44 = W*in
   wire signed [14:0] m44_44;
   assign m44_44 =15'b0;

   // m44_45 = W*in
   wire signed [14:0] m44_45;
   assign m44_45 =15'b0;

   // m44_46 = W*in
   wire signed [14:0] m44_46;
   assign m44_46 =15'b0;

   // m44_47 = W*in
   wire signed [14:0] m44_47;
   assign m44_47 =15'b0;

   // m44_48 = W*in
   wire signed [14:0] m44_48;
   assign m44_48 =15'b0;

   // m44_49 = W*in
   wire signed [14:0] m44_49;
   assign m44_49 =15'b0;

   // m44_50 = W*in
   wire signed [14:0] m44_50;
   assign m44_50 =15'b0;

   // m44_51 = W*in
   wire signed [14:0] m44_51;
   assign m44_51 =15'b0;

   // m44_52 = W*in
   wire signed [14:0] m44_52;
   assign m44_52 =15'b0;

   // m44_53 = W*in
   wire signed [14:0] m44_53;
   assign m44_53 =15'b0;

   // m44_54 = W*in
   wire signed [14:0] m44_54;
   assign m44_54 =15'b0;

   // m44_55 = W*in
   wire signed [14:0] m44_55;
   assign m44_55 =15'b0;

   // m44_56 = W*in
   wire signed [14:0] m44_56;
   assign m44_56 =15'b0;

   // m44_57 = W*in
   wire signed [14:0] m44_57;
   assign m44_57 =15'b0;

   // m44_58 = W*in
   wire signed [14:0] m44_58;
   assign m44_58 =15'b0;

   // m44_59 = W*in
   wire signed [14:0] m44_59;
   assign m44_59 =15'b0;

   // m44_60 = W*in
   wire signed [14:0] m44_60;
   assign m44_60 =15'b0;

   // m44_61 = W*in
   wire signed [14:0] m44_61;
   assign m44_61 =15'b0;

   // m44_62 = W*in
   wire signed [14:0] m44_62;
   assign m44_62 =15'b0;

   // m44_63 = W*in
   wire signed [14:0] m44_63;
   assign m44_63 ={ {3{neg44[14]}} , neg44[14:3] };

   // m44_64 = W*in
   wire signed [14:0] m44_64;
   assign m44_64 ={ {3{in44[14]}} , in44[14:3] };

   // m44_65 = W*in
   wire signed [14:0] m44_65;
   assign m44_65 =15'b0;

   // m44_66 = W*in
   wire signed [14:0] m44_66;
   assign m44_66 =15'b0;

   // m44_67 = W*in
   wire signed [14:0] m44_67;
   assign m44_67 =15'b0;

   // m44_68 = W*in
   wire signed [14:0] m44_68;
   assign m44_68 =15'b0;

   // m44_69 = W*in
   wire signed [14:0] m44_69;
   assign m44_69 ={ {3{in44[14]}} , in44[14:3] };

   // m44_70 = W*in
   wire signed [14:0] m44_70;
   assign m44_70 =15'b0;

   // m44_71 = W*in
   wire signed [14:0] m44_71;
   assign m44_71 =15'b0;

   // m44_72 = W*in
   wire signed [14:0] m44_72;
   assign m44_72 ={ {3{neg44[14]}} , neg44[14:3] };

   // m44_73 = W*in
   wire signed [14:0] m44_73;
   assign m44_73 =15'b0;

   // m44_74 = W*in
   wire signed [14:0] m44_74;
   assign m44_74 =15'b0;

   // m44_75 = W*in
   wire signed [14:0] m44_75;
   assign m44_75 =15'b0;

   // m44_76 = W*in
   wire signed [14:0] m44_76;
   assign m44_76 ={ {3{neg44[14]}} , neg44[14:3] };

   // m44_77 = W*in
   wire signed [14:0] m44_77;
   assign m44_77 =15'b0;

   // m44_78 = W*in
   wire signed [14:0] m44_78;
   assign m44_78 =15'b0;

   // m44_79 = W*in
   wire signed [14:0] m44_79;
   assign m44_79 =15'b0;

   // m44_80 = W*in
   wire signed [14:0] m44_80;
   assign m44_80 =15'b0;

   // m44_81 = W*in
   wire signed [14:0] m44_81;
   assign m44_81 =15'b0;

   // m44_82 = W*in
   wire signed [14:0] m44_82;
   assign m44_82 =15'b0;

   // m44_83 = W*in
   wire signed [14:0] m44_83;
   assign m44_83 ={ {3{neg44[14]}} , neg44[14:3] };

   // m44_84 = W*in
   wire signed [14:0] m44_84;
   assign m44_84 =15'b0;

   // m44_85 = W*in
   wire signed [14:0] m44_85;
   assign m44_85 =15'b0;

   // m44_86 = W*in
   wire signed [14:0] m44_86;
   assign m44_86 ={ {3{in44[14]}} , in44[14:3] };

   // m44_87 = W*in
   wire signed [14:0] m44_87;
   assign m44_87 =15'b0;

   // m44_88 = W*in
   wire signed [14:0] m44_88;
   assign m44_88 ={ {3{in44[14]}} , in44[14:3] };

   // m44_89 = W*in
   wire signed [14:0] m44_89;
   assign m44_89 =15'b0;

   // m44_90 = W*in
   wire signed [14:0] m44_90;
   assign m44_90 =15'b0;

   // m44_91 = W*in
   wire signed [14:0] m44_91;
   assign m44_91 =15'b0;

   // m44_92 = W*in
   wire signed [14:0] m44_92;
   assign m44_92 =15'b0;

   // m44_93 = W*in
   wire signed [14:0] m44_93;
   assign m44_93 =15'b0;

   // m44_94 = W*in
   wire signed [14:0] m44_94;
   assign m44_94 ={ {4{neg44[14]}} , neg44[14:4] };

   // m44_95 = W*in
   wire signed [14:0] m44_95;
   assign m44_95 ={ {3{in44[14]}} , in44[14:3] };

   // m44_96 = W*in
   wire signed [14:0] m44_96;
   assign m44_96 =15'b0;

   // m44_97 = W*in
   wire signed [14:0] m44_97;
   assign m44_97 =15'b0;

   // m44_98 = W*in
   wire signed [14:0] m44_98;
   assign m44_98 ={ {3{in44[14]}} , in44[14:3] };

   // m44_99 = W*in
   wire signed [14:0] m44_99;
   assign m44_99 =15'b0;

   // m44_100 = W*in
   wire signed [14:0] m44_100;
   assign m44_100 ={ {3{neg44[14]}} , neg44[14:3] };

   // m45_1 = W*in
   wire signed [14:0] m45_1;
   assign m45_1 =15'b0;

   // m45_2 = W*in
   wire signed [14:0] m45_2;
   assign m45_2 =15'b0;

   // m45_3 = W*in
   wire signed [14:0] m45_3;
   assign m45_3 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_4 = W*in
   wire signed [14:0] m45_4;
   assign m45_4 =15'b0;

   // m45_5 = W*in
   wire signed [14:0] m45_5;
   assign m45_5 =15'b0;

   // m45_6 = W*in
   wire signed [14:0] m45_6;
   assign m45_6 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_7 = W*in
   wire signed [14:0] m45_7;
   assign m45_7 ={ {4{in45[14]}} , in45[14:4] };

   // m45_8 = W*in
   wire signed [14:0] m45_8;
   assign m45_8 =15'b0;

   // m45_9 = W*in
   wire signed [14:0] m45_9;
   assign m45_9 =15'b0;

   // m45_10 = W*in
   wire signed [14:0] m45_10;
   assign m45_10 ={ {3{in45[14]}} , in45[14:3] };

   // m45_11 = W*in
   wire signed [14:0] m45_11;
   assign m45_11 ={ {4{in45[14]}} , in45[14:4] };

   // m45_12 = W*in
   wire signed [14:0] m45_12;
   assign m45_12 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_13 = W*in
   wire signed [14:0] m45_13;
   assign m45_13 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_14 = W*in
   wire signed [14:0] m45_14;
   assign m45_14 =15'b0;

   // m45_15 = W*in
   wire signed [14:0] m45_15;
   assign m45_15 =15'b0;

   // m45_16 = W*in
   wire signed [14:0] m45_16;
   assign m45_16 =15'b0;

   // m45_17 = W*in
   wire signed [14:0] m45_17;
   assign m45_17 =15'b0;

   // m45_18 = W*in
   wire signed [14:0] m45_18;
   assign m45_18 =15'b0;

   // m45_19 = W*in
   wire signed [14:0] m45_19;
   assign m45_19 ={ {3{in45[14]}} , in45[14:3] };

   // m45_20 = W*in
   wire signed [14:0] m45_20;
   assign m45_20 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_21 = W*in
   wire signed [14:0] m45_21;
   assign m45_21 =15'b0;

   // m45_22 = W*in
   wire signed [14:0] m45_22;
   assign m45_22 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_23 = W*in
   wire signed [14:0] m45_23;
   assign m45_23 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_24 = W*in
   wire signed [14:0] m45_24;
   assign m45_24 =15'b0;

   // m45_25 = W*in
   wire signed [14:0] m45_25;
   assign m45_25 =15'b0;

   // m45_26 = W*in
   wire signed [14:0] m45_26;
   assign m45_26 =15'b0;

   // m45_27 = W*in
   wire signed [14:0] m45_27;
   assign m45_27 =15'b0;

   // m45_28 = W*in
   wire signed [14:0] m45_28;
   assign m45_28 ={ {4{in45[14]}} , in45[14:4] };

   // m45_29 = W*in
   wire signed [14:0] m45_29;
   assign m45_29 =15'b0;

   // m45_30 = W*in
   wire signed [14:0] m45_30;
   assign m45_30 ={ {3{in45[14]}} , in45[14:3] };

   // m45_31 = W*in
   wire signed [14:0] m45_31;
   assign m45_31 ={ {3{in45[14]}} , in45[14:3] };

   // m45_32 = W*in
   wire signed [14:0] m45_32;
   assign m45_32 ={ {3{in45[14]}} , in45[14:3] };

   // m45_33 = W*in
   wire signed [14:0] m45_33;
   assign m45_33 ={ {3{in45[14]}} , in45[14:3] };

   // m45_34 = W*in
   wire signed [14:0] m45_34;
   assign m45_34 =15'b0;

   // m45_35 = W*in
   wire signed [14:0] m45_35;
   assign m45_35 =15'b0;

   // m45_36 = W*in
   wire signed [14:0] m45_36;
   assign m45_36 =15'b0;

   // m45_37 = W*in
   wire signed [14:0] m45_37;
   assign m45_37 =15'b0;

   // m45_38 = W*in
   wire signed [14:0] m45_38;
   assign m45_38 =15'b0;

   // m45_39 = W*in
   wire signed [14:0] m45_39;
   assign m45_39 =15'b0;

   // m45_40 = W*in
   wire signed [14:0] m45_40;
   assign m45_40 =15'b0;

   // m45_41 = W*in
   wire signed [14:0] m45_41;
   assign m45_41 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_42 = W*in
   wire signed [14:0] m45_42;
   assign m45_42 =15'b0;

   // m45_43 = W*in
   wire signed [14:0] m45_43;
   assign m45_43 =15'b0;

   // m45_44 = W*in
   wire signed [14:0] m45_44;
   assign m45_44 ={ {3{in45[14]}} , in45[14:3] };

   // m45_45 = W*in
   wire signed [14:0] m45_45;
   assign m45_45 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_46 = W*in
   wire signed [14:0] m45_46;
   assign m45_46 =15'b0;

   // m45_47 = W*in
   wire signed [14:0] m45_47;
   assign m45_47 =15'b0;

   // m45_48 = W*in
   wire signed [14:0] m45_48;
   assign m45_48 =15'b0;

   // m45_49 = W*in
   wire signed [14:0] m45_49;
   assign m45_49 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_50 = W*in
   wire signed [14:0] m45_50;
   assign m45_50 =15'b0;

   // m45_51 = W*in
   wire signed [14:0] m45_51;
   assign m45_51 =15'b0;

   // m45_52 = W*in
   wire signed [14:0] m45_52;
   assign m45_52 =15'b0;

   // m45_53 = W*in
   wire signed [14:0] m45_53;
   assign m45_53 =15'b0;

   // m45_54 = W*in
   wire signed [14:0] m45_54;
   assign m45_54 ={ {3{in45[14]}} , in45[14:3] };

   // m45_55 = W*in
   wire signed [14:0] m45_55;
   assign m45_55 =15'b0;

   // m45_56 = W*in
   wire signed [14:0] m45_56;
   assign m45_56 =15'b0;

   // m45_57 = W*in
   wire signed [14:0] m45_57;
   assign m45_57 =15'b0;

   // m45_58 = W*in
   wire signed [14:0] m45_58;
   assign m45_58 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_59 = W*in
   wire signed [14:0] m45_59;
   assign m45_59 ={ {4{neg45[14]}} , neg45[14:4] };

   // m45_60 = W*in
   wire signed [14:0] m45_60;
   assign m45_60 =15'b0;

   // m45_61 = W*in
   wire signed [14:0] m45_61;
   assign m45_61 ={ {4{neg45[14]}} , neg45[14:4] };

   // m45_62 = W*in
   wire signed [14:0] m45_62;
   assign m45_62 ={ {2{neg45[14]}} , neg45[14:2] };

   // m45_63 = W*in
   wire signed [14:0] m45_63;
   assign m45_63 ={ {3{in45[14]}} , in45[14:3] };

   // m45_64 = W*in
   wire signed [14:0] m45_64;
   assign m45_64 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_65 = W*in
   wire signed [14:0] m45_65;
   assign m45_65 ={ {3{in45[14]}} , in45[14:3] };

   // m45_66 = W*in
   wire signed [14:0] m45_66;
   assign m45_66 =15'b0;

   // m45_67 = W*in
   wire signed [14:0] m45_67;
   assign m45_67 =15'b0;

   // m45_68 = W*in
   wire signed [14:0] m45_68;
   assign m45_68 =15'b0;

   // m45_69 = W*in
   wire signed [14:0] m45_69;
   assign m45_69 ={ {3{in45[14]}} , in45[14:3] };

   // m45_70 = W*in
   wire signed [14:0] m45_70;
   assign m45_70 ={ {4{in45[14]}} , in45[14:4] };

   // m45_71 = W*in
   wire signed [14:0] m45_71;
   assign m45_71 ={ {4{in45[14]}} , in45[14:4] };

   // m45_72 = W*in
   wire signed [14:0] m45_72;
   assign m45_72 =15'b0;

   // m45_73 = W*in
   wire signed [14:0] m45_73;
   assign m45_73 =15'b0;

   // m45_74 = W*in
   wire signed [14:0] m45_74;
   assign m45_74 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_75 = W*in
   wire signed [14:0] m45_75;
   assign m45_75 ={ {2{neg45[14]}} , neg45[14:2] };

   // m45_76 = W*in
   wire signed [14:0] m45_76;
   assign m45_76 =15'b0;

   // m45_77 = W*in
   wire signed [14:0] m45_77;
   assign m45_77 =15'b0;

   // m45_78 = W*in
   wire signed [14:0] m45_78;
   assign m45_78 =15'b0;

   // m45_79 = W*in
   wire signed [14:0] m45_79;
   assign m45_79 ={ {3{in45[14]}} , in45[14:3] };

   // m45_80 = W*in
   wire signed [14:0] m45_80;
   assign m45_80 ={ {3{in45[14]}} , in45[14:3] };

   // m45_81 = W*in
   wire signed [14:0] m45_81;
   assign m45_81 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_82 = W*in
   wire signed [14:0] m45_82;
   assign m45_82 =15'b0;

   // m45_83 = W*in
   wire signed [14:0] m45_83;
   assign m45_83 =15'b0;

   // m45_84 = W*in
   wire signed [14:0] m45_84;
   assign m45_84 =15'b0;

   // m45_85 = W*in
   wire signed [14:0] m45_85;
   assign m45_85 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_86 = W*in
   wire signed [14:0] m45_86;
   assign m45_86 =15'b0;

   // m45_87 = W*in
   wire signed [14:0] m45_87;
   assign m45_87 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_88 = W*in
   wire signed [14:0] m45_88;
   assign m45_88 =15'b0;

   // m45_89 = W*in
   wire signed [14:0] m45_89;
   assign m45_89 =15'b0;

   // m45_90 = W*in
   wire signed [14:0] m45_90;
   assign m45_90 =15'b0;

   // m45_91 = W*in
   wire signed [14:0] m45_91;
   assign m45_91 =15'b0;

   // m45_92 = W*in
   wire signed [14:0] m45_92;
   assign m45_92 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_93 = W*in
   wire signed [14:0] m45_93;
   assign m45_93 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_94 = W*in
   wire signed [14:0] m45_94;
   assign m45_94 ={ {3{in45[14]}} , in45[14:3] };

   // m45_95 = W*in
   wire signed [14:0] m45_95;
   assign m45_95 =15'b0;

   // m45_96 = W*in
   wire signed [14:0] m45_96;
   assign m45_96 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_97 = W*in
   wire signed [14:0] m45_97;
   assign m45_97 ={ {3{neg45[14]}} , neg45[14:3] };

   // m45_98 = W*in
   wire signed [14:0] m45_98;
   assign m45_98 ={ {3{in45[14]}} , in45[14:3] };

   // m45_99 = W*in
   wire signed [14:0] m45_99;
   assign m45_99 =15'b0;

   // m45_100 = W*in
   wire signed [14:0] m45_100;
   assign m45_100 =15'b0;

   // m46_1 = W*in
   wire signed [14:0] m46_1;
   assign m46_1 =15'b0;

   // m46_2 = W*in
   wire signed [14:0] m46_2;
   assign m46_2 =15'b0;

   // m46_3 = W*in
   wire signed [14:0] m46_3;
   assign m46_3 =15'b0;

   // m46_4 = W*in
   wire signed [14:0] m46_4;
   assign m46_4 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_5 = W*in
   wire signed [14:0] m46_5;
   assign m46_5 =15'b0;

   // m46_6 = W*in
   wire signed [14:0] m46_6;
   assign m46_6 =15'b0;

   // m46_7 = W*in
   wire signed [14:0] m46_7;
   assign m46_7 ={ {4{neg46[14]}} , neg46[14:4] };

   // m46_8 = W*in
   wire signed [14:0] m46_8;
   assign m46_8 =15'b0;

   // m46_9 = W*in
   wire signed [14:0] m46_9;
   assign m46_9 =15'b0;

   // m46_10 = W*in
   wire signed [14:0] m46_10;
   assign m46_10 =15'b0;

   // m46_11 = W*in
   wire signed [14:0] m46_11;
   assign m46_11 =15'b0;

   // m46_12 = W*in
   wire signed [14:0] m46_12;
   assign m46_12 ={ {3{in46[14]}} , in46[14:3] };

   // m46_13 = W*in
   wire signed [14:0] m46_13;
   assign m46_13 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_14 = W*in
   wire signed [14:0] m46_14;
   assign m46_14 =15'b0;

   // m46_15 = W*in
   wire signed [14:0] m46_15;
   assign m46_15 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_16 = W*in
   wire signed [14:0] m46_16;
   assign m46_16 =15'b0;

   // m46_17 = W*in
   wire signed [14:0] m46_17;
   assign m46_17 =15'b0;

   // m46_18 = W*in
   wire signed [14:0] m46_18;
   assign m46_18 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_19 = W*in
   wire signed [14:0] m46_19;
   assign m46_19 ={ {3{in46[14]}} , in46[14:3] };

   // m46_20 = W*in
   wire signed [14:0] m46_20;
   assign m46_20 ={ {4{neg46[14]}} , neg46[14:4] };

   // m46_21 = W*in
   wire signed [14:0] m46_21;
   assign m46_21 =15'b0;

   // m46_22 = W*in
   wire signed [14:0] m46_22;
   assign m46_22 =15'b0;

   // m46_23 = W*in
   wire signed [14:0] m46_23;
   assign m46_23 =15'b0;

   // m46_24 = W*in
   wire signed [14:0] m46_24;
   assign m46_24 =15'b0;

   // m46_25 = W*in
   wire signed [14:0] m46_25;
   assign m46_25 =15'b0;

   // m46_26 = W*in
   wire signed [14:0] m46_26;
   assign m46_26 ={ {3{in46[14]}} , in46[14:3] };

   // m46_27 = W*in
   wire signed [14:0] m46_27;
   assign m46_27 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_28 = W*in
   wire signed [14:0] m46_28;
   assign m46_28 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_29 = W*in
   wire signed [14:0] m46_29;
   assign m46_29 =15'b0;

   // m46_30 = W*in
   wire signed [14:0] m46_30;
   assign m46_30 ={ {4{neg46[14]}} , neg46[14:4] };

   // m46_31 = W*in
   wire signed [14:0] m46_31;
   assign m46_31 =15'b0;

   // m46_32 = W*in
   wire signed [14:0] m46_32;
   assign m46_32 =15'b0;

   // m46_33 = W*in
   wire signed [14:0] m46_33;
   assign m46_33 ={ {4{neg46[14]}} , neg46[14:4] };

   // m46_34 = W*in
   wire signed [14:0] m46_34;
   assign m46_34 =15'b0;

   // m46_35 = W*in
   wire signed [14:0] m46_35;
   assign m46_35 =15'b0;

   // m46_36 = W*in
   wire signed [14:0] m46_36;
   assign m46_36 =15'b0;

   // m46_37 = W*in
   wire signed [14:0] m46_37;
   assign m46_37 =15'b0;

   // m46_38 = W*in
   wire signed [14:0] m46_38;
   assign m46_38 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_39 = W*in
   wire signed [14:0] m46_39;
   assign m46_39 ={ {3{in46[14]}} , in46[14:3] };

   // m46_40 = W*in
   wire signed [14:0] m46_40;
   assign m46_40 =15'b0;

   // m46_41 = W*in
   wire signed [14:0] m46_41;
   assign m46_41 =15'b0;

   // m46_42 = W*in
   wire signed [14:0] m46_42;
   assign m46_42 =15'b0;

   // m46_43 = W*in
   wire signed [14:0] m46_43;
   assign m46_43 =15'b0;

   // m46_44 = W*in
   wire signed [14:0] m46_44;
   assign m46_44 =15'b0;

   // m46_45 = W*in
   wire signed [14:0] m46_45;
   assign m46_45 =15'b0;

   // m46_46 = W*in
   wire signed [14:0] m46_46;
   assign m46_46 =15'b0;

   // m46_47 = W*in
   wire signed [14:0] m46_47;
   assign m46_47 ={ {2{in46[14]}} , in46[14:2] };

   // m46_48 = W*in
   wire signed [14:0] m46_48;
   assign m46_48 =15'b0;

   // m46_49 = W*in
   wire signed [14:0] m46_49;
   assign m46_49 =15'b0;

   // m46_50 = W*in
   wire signed [14:0] m46_50;
   assign m46_50 =15'b0;

   // m46_51 = W*in
   wire signed [14:0] m46_51;
   assign m46_51 =15'b0;

   // m46_52 = W*in
   wire signed [14:0] m46_52;
   assign m46_52 =15'b0;

   // m46_53 = W*in
   wire signed [14:0] m46_53;
   assign m46_53 =15'b0;

   // m46_54 = W*in
   wire signed [14:0] m46_54;
   assign m46_54 =15'b0;

   // m46_55 = W*in
   wire signed [14:0] m46_55;
   assign m46_55 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_56 = W*in
   wire signed [14:0] m46_56;
   assign m46_56 =15'b0;

   // m46_57 = W*in
   wire signed [14:0] m46_57;
   assign m46_57 =15'b0;

   // m46_58 = W*in
   wire signed [14:0] m46_58;
   assign m46_58 =15'b0;

   // m46_59 = W*in
   wire signed [14:0] m46_59;
   assign m46_59 ={ {3{in46[14]}} , in46[14:3] };

   // m46_60 = W*in
   wire signed [14:0] m46_60;
   assign m46_60 =15'b0;

   // m46_61 = W*in
   wire signed [14:0] m46_61;
   assign m46_61 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_62 = W*in
   wire signed [14:0] m46_62;
   assign m46_62 =15'b0;

   // m46_63 = W*in
   wire signed [14:0] m46_63;
   assign m46_63 =15'b0;

   // m46_64 = W*in
   wire signed [14:0] m46_64;
   assign m46_64 =15'b0;

   // m46_65 = W*in
   wire signed [14:0] m46_65;
   assign m46_65 =15'b0;

   // m46_66 = W*in
   wire signed [14:0] m46_66;
   assign m46_66 =15'b0;

   // m46_67 = W*in
   wire signed [14:0] m46_67;
   assign m46_67 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_68 = W*in
   wire signed [14:0] m46_68;
   assign m46_68 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_69 = W*in
   wire signed [14:0] m46_69;
   assign m46_69 =15'b0;

   // m46_70 = W*in
   wire signed [14:0] m46_70;
   assign m46_70 =15'b0;

   // m46_71 = W*in
   wire signed [14:0] m46_71;
   assign m46_71 =15'b0;

   // m46_72 = W*in
   wire signed [14:0] m46_72;
   assign m46_72 =15'b0;

   // m46_73 = W*in
   wire signed [14:0] m46_73;
   assign m46_73 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_74 = W*in
   wire signed [14:0] m46_74;
   assign m46_74 =15'b0;

   // m46_75 = W*in
   wire signed [14:0] m46_75;
   assign m46_75 ={ {3{in46[14]}} , in46[14:3] };

   // m46_76 = W*in
   wire signed [14:0] m46_76;
   assign m46_76 =15'b0;

   // m46_77 = W*in
   wire signed [14:0] m46_77;
   assign m46_77 =15'b0;

   // m46_78 = W*in
   wire signed [14:0] m46_78;
   assign m46_78 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_79 = W*in
   wire signed [14:0] m46_79;
   assign m46_79 ={ {2{in46[14]}} , in46[14:2] };

   // m46_80 = W*in
   wire signed [14:0] m46_80;
   assign m46_80 =15'b0;

   // m46_81 = W*in
   wire signed [14:0] m46_81;
   assign m46_81 =15'b0;

   // m46_82 = W*in
   wire signed [14:0] m46_82;
   assign m46_82 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_83 = W*in
   wire signed [14:0] m46_83;
   assign m46_83 =15'b0;

   // m46_84 = W*in
   wire signed [14:0] m46_84;
   assign m46_84 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_85 = W*in
   wire signed [14:0] m46_85;
   assign m46_85 =15'b0;

   // m46_86 = W*in
   wire signed [14:0] m46_86;
   assign m46_86 =15'b0;

   // m46_87 = W*in
   wire signed [14:0] m46_87;
   assign m46_87 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_88 = W*in
   wire signed [14:0] m46_88;
   assign m46_88 =15'b0;

   // m46_89 = W*in
   wire signed [14:0] m46_89;
   assign m46_89 =15'b0;

   // m46_90 = W*in
   wire signed [14:0] m46_90;
   assign m46_90 =15'b0;

   // m46_91 = W*in
   wire signed [14:0] m46_91;
   assign m46_91 =15'b0;

   // m46_92 = W*in
   wire signed [14:0] m46_92;
   assign m46_92 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_93 = W*in
   wire signed [14:0] m46_93;
   assign m46_93 ={ {4{in46[14]}} , in46[14:4] };

   // m46_94 = W*in
   wire signed [14:0] m46_94;
   assign m46_94 =15'b0;

   // m46_95 = W*in
   wire signed [14:0] m46_95;
   assign m46_95 =15'b0;

   // m46_96 = W*in
   wire signed [14:0] m46_96;
   assign m46_96 =15'b0;

   // m46_97 = W*in
   wire signed [14:0] m46_97;
   assign m46_97 ={ {3{neg46[14]}} , neg46[14:3] };

   // m46_98 = W*in
   wire signed [14:0] m46_98;
   assign m46_98 =15'b0;

   // m46_99 = W*in
   wire signed [14:0] m46_99;
   assign m46_99 =15'b0;

   // m46_100 = W*in
   wire signed [14:0] m46_100;
   assign m46_100 =15'b0;

   // m47_1 = W*in
   wire signed [14:0] m47_1;
   assign m47_1 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_2 = W*in
   wire signed [14:0] m47_2;
   assign m47_2 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_3 = W*in
   wire signed [14:0] m47_3;
   assign m47_3 =15'b0;

   // m47_4 = W*in
   wire signed [14:0] m47_4;
   assign m47_4 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_5 = W*in
   wire signed [14:0] m47_5;
   assign m47_5 =15'b0;

   // m47_6 = W*in
   wire signed [14:0] m47_6;
   assign m47_6 =15'b0;

   // m47_7 = W*in
   wire signed [14:0] m47_7;
   assign m47_7 =15'b0;

   // m47_8 = W*in
   wire signed [14:0] m47_8;
   assign m47_8 =15'b0;

   // m47_9 = W*in
   wire signed [14:0] m47_9;
   assign m47_9 =15'b0;

   // m47_10 = W*in
   wire signed [14:0] m47_10;
   assign m47_10 =15'b0;

   // m47_11 = W*in
   wire signed [14:0] m47_11;
   assign m47_11 =15'b0;

   // m47_12 = W*in
   wire signed [14:0] m47_12;
   assign m47_12 =15'b0;

   // m47_13 = W*in
   wire signed [14:0] m47_13;
   assign m47_13 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_14 = W*in
   wire signed [14:0] m47_14;
   assign m47_14 =15'b0;

   // m47_15 = W*in
   wire signed [14:0] m47_15;
   assign m47_15 =15'b0;

   // m47_16 = W*in
   wire signed [14:0] m47_16;
   assign m47_16 =15'b0;

   // m47_17 = W*in
   wire signed [14:0] m47_17;
   assign m47_17 =15'b0;

   // m47_18 = W*in
   wire signed [14:0] m47_18;
   assign m47_18 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_19 = W*in
   wire signed [14:0] m47_19;
   assign m47_19 ={ {3{in47[14]}} , in47[14:3] };

   // m47_20 = W*in
   wire signed [14:0] m47_20;
   assign m47_20 ={ {4{neg47[14]}} , neg47[14:4] };

   // m47_21 = W*in
   wire signed [14:0] m47_21;
   assign m47_21 ={ {4{neg47[14]}} , neg47[14:4] };

   // m47_22 = W*in
   wire signed [14:0] m47_22;
   assign m47_22 =15'b0;

   // m47_23 = W*in
   wire signed [14:0] m47_23;
   assign m47_23 =15'b0;

   // m47_24 = W*in
   wire signed [14:0] m47_24;
   assign m47_24 =15'b0;

   // m47_25 = W*in
   wire signed [14:0] m47_25;
   assign m47_25 =15'b0;

   // m47_26 = W*in
   wire signed [14:0] m47_26;
   assign m47_26 =15'b0;

   // m47_27 = W*in
   wire signed [14:0] m47_27;
   assign m47_27 =15'b0;

   // m47_28 = W*in
   wire signed [14:0] m47_28;
   assign m47_28 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_29 = W*in
   wire signed [14:0] m47_29;
   assign m47_29 =15'b0;

   // m47_30 = W*in
   wire signed [14:0] m47_30;
   assign m47_30 ={ {4{neg47[14]}} , neg47[14:4] };

   // m47_31 = W*in
   wire signed [14:0] m47_31;
   assign m47_31 =15'b0;

   // m47_32 = W*in
   wire signed [14:0] m47_32;
   assign m47_32 =15'b0;

   // m47_33 = W*in
   wire signed [14:0] m47_33;
   assign m47_33 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_34 = W*in
   wire signed [14:0] m47_34;
   assign m47_34 =15'b0;

   // m47_35 = W*in
   wire signed [14:0] m47_35;
   assign m47_35 =15'b0;

   // m47_36 = W*in
   wire signed [14:0] m47_36;
   assign m47_36 =15'b0;

   // m47_37 = W*in
   wire signed [14:0] m47_37;
   assign m47_37 =15'b0;

   // m47_38 = W*in
   wire signed [14:0] m47_38;
   assign m47_38 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_39 = W*in
   wire signed [14:0] m47_39;
   assign m47_39 ={ {3{in47[14]}} , in47[14:3] };

   // m47_40 = W*in
   wire signed [14:0] m47_40;
   assign m47_40 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_41 = W*in
   wire signed [14:0] m47_41;
   assign m47_41 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_42 = W*in
   wire signed [14:0] m47_42;
   assign m47_42 =15'b0;

   // m47_43 = W*in
   wire signed [14:0] m47_43;
   assign m47_43 =15'b0;

   // m47_44 = W*in
   wire signed [14:0] m47_44;
   assign m47_44 =15'b0;

   // m47_45 = W*in
   wire signed [14:0] m47_45;
   assign m47_45 =15'b0;

   // m47_46 = W*in
   wire signed [14:0] m47_46;
   assign m47_46 =15'b0;

   // m47_47 = W*in
   wire signed [14:0] m47_47;
   assign m47_47 ={ {3{in47[14]}} , in47[14:3] };

   // m47_48 = W*in
   wire signed [14:0] m47_48;
   assign m47_48 =15'b0;

   // m47_49 = W*in
   wire signed [14:0] m47_49;
   assign m47_49 =15'b0;

   // m47_50 = W*in
   wire signed [14:0] m47_50;
   assign m47_50 =15'b0;

   // m47_51 = W*in
   wire signed [14:0] m47_51;
   assign m47_51 =15'b0;

   // m47_52 = W*in
   wire signed [14:0] m47_52;
   assign m47_52 =15'b0;

   // m47_53 = W*in
   wire signed [14:0] m47_53;
   assign m47_53 =15'b0;

   // m47_54 = W*in
   wire signed [14:0] m47_54;
   assign m47_54 =15'b0;

   // m47_55 = W*in
   wire signed [14:0] m47_55;
   assign m47_55 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_56 = W*in
   wire signed [14:0] m47_56;
   assign m47_56 =15'b0;

   // m47_57 = W*in
   wire signed [14:0] m47_57;
   assign m47_57 =15'b0;

   // m47_58 = W*in
   wire signed [14:0] m47_58;
   assign m47_58 =15'b0;

   // m47_59 = W*in
   wire signed [14:0] m47_59;
   assign m47_59 =15'b0;

   // m47_60 = W*in
   wire signed [14:0] m47_60;
   assign m47_60 =15'b0;

   // m47_61 = W*in
   wire signed [14:0] m47_61;
   assign m47_61 =15'b0;

   // m47_62 = W*in
   wire signed [14:0] m47_62;
   assign m47_62 =15'b0;

   // m47_63 = W*in
   wire signed [14:0] m47_63;
   assign m47_63 ={ {3{in47[14]}} , in47[14:3] };

   // m47_64 = W*in
   wire signed [14:0] m47_64;
   assign m47_64 =15'b0;

   // m47_65 = W*in
   wire signed [14:0] m47_65;
   assign m47_65 =15'b0;

   // m47_66 = W*in
   wire signed [14:0] m47_66;
   assign m47_66 =15'b0;

   // m47_67 = W*in
   wire signed [14:0] m47_67;
   assign m47_67 ={ {4{neg47[14]}} , neg47[14:4] };

   // m47_68 = W*in
   wire signed [14:0] m47_68;
   assign m47_68 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_69 = W*in
   wire signed [14:0] m47_69;
   assign m47_69 =15'b0;

   // m47_70 = W*in
   wire signed [14:0] m47_70;
   assign m47_70 =15'b0;

   // m47_71 = W*in
   wire signed [14:0] m47_71;
   assign m47_71 =15'b0;

   // m47_72 = W*in
   wire signed [14:0] m47_72;
   assign m47_72 =15'b0;

   // m47_73 = W*in
   wire signed [14:0] m47_73;
   assign m47_73 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_74 = W*in
   wire signed [14:0] m47_74;
   assign m47_74 =15'b0;

   // m47_75 = W*in
   wire signed [14:0] m47_75;
   assign m47_75 =15'b0;

   // m47_76 = W*in
   wire signed [14:0] m47_76;
   assign m47_76 =15'b0;

   // m47_77 = W*in
   wire signed [14:0] m47_77;
   assign m47_77 =15'b0;

   // m47_78 = W*in
   wire signed [14:0] m47_78;
   assign m47_78 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_79 = W*in
   wire signed [14:0] m47_79;
   assign m47_79 ={ {3{in47[14]}} , in47[14:3] };

   // m47_80 = W*in
   wire signed [14:0] m47_80;
   assign m47_80 =15'b0;

   // m47_81 = W*in
   wire signed [14:0] m47_81;
   assign m47_81 =15'b0;

   // m47_82 = W*in
   wire signed [14:0] m47_82;
   assign m47_82 =15'b0;

   // m47_83 = W*in
   wire signed [14:0] m47_83;
   assign m47_83 =15'b0;

   // m47_84 = W*in
   wire signed [14:0] m47_84;
   assign m47_84 =15'b0;

   // m47_85 = W*in
   wire signed [14:0] m47_85;
   assign m47_85 =15'b0;

   // m47_86 = W*in
   wire signed [14:0] m47_86;
   assign m47_86 =15'b0;

   // m47_87 = W*in
   wire signed [14:0] m47_87;
   assign m47_87 =15'b0;

   // m47_88 = W*in
   wire signed [14:0] m47_88;
   assign m47_88 =15'b0;

   // m47_89 = W*in
   wire signed [14:0] m47_89;
   assign m47_89 =15'b0;

   // m47_90 = W*in
   wire signed [14:0] m47_90;
   assign m47_90 =15'b0;

   // m47_91 = W*in
   wire signed [14:0] m47_91;
   assign m47_91 ={ {3{in47[14]}} , in47[14:3] };

   // m47_92 = W*in
   wire signed [14:0] m47_92;
   assign m47_92 =15'b0;

   // m47_93 = W*in
   wire signed [14:0] m47_93;
   assign m47_93 =15'b0;

   // m47_94 = W*in
   wire signed [14:0] m47_94;
   assign m47_94 ={ {4{in47[14]}} , in47[14:4] };

   // m47_95 = W*in
   wire signed [14:0] m47_95;
   assign m47_95 =15'b0;

   // m47_96 = W*in
   wire signed [14:0] m47_96;
   assign m47_96 =15'b0;

   // m47_97 = W*in
   wire signed [14:0] m47_97;
   assign m47_97 ={ {3{neg47[14]}} , neg47[14:3] };

   // m47_98 = W*in
   wire signed [14:0] m47_98;
   assign m47_98 =15'b0;

   // m47_99 = W*in
   wire signed [14:0] m47_99;
   assign m47_99 =15'b0;

   // m47_100 = W*in
   wire signed [14:0] m47_100;
   assign m47_100 ={ {3{in47[14]}} , in47[14:3] };

   // m48_1 = W*in
   wire signed [14:0] m48_1;
   assign m48_1 =15'b0;

   // m48_2 = W*in
   wire signed [14:0] m48_2;
   assign m48_2 =15'b0;

   // m48_3 = W*in
   wire signed [14:0] m48_3;
   assign m48_3 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_4 = W*in
   wire signed [14:0] m48_4;
   assign m48_4 =15'b0;

   // m48_5 = W*in
   wire signed [14:0] m48_5;
   assign m48_5 =15'b0;

   // m48_6 = W*in
   wire signed [14:0] m48_6;
   assign m48_6 =15'b0;

   // m48_7 = W*in
   wire signed [14:0] m48_7;
   assign m48_7 ={ {3{in48[14]}} , in48[14:3] };

   // m48_8 = W*in
   wire signed [14:0] m48_8;
   assign m48_8 =15'b0;

   // m48_9 = W*in
   wire signed [14:0] m48_9;
   assign m48_9 =15'b0;

   // m48_10 = W*in
   wire signed [14:0] m48_10;
   assign m48_10 ={ {3{in48[14]}} , in48[14:3] };

   // m48_11 = W*in
   wire signed [14:0] m48_11;
   assign m48_11 ={ {3{in48[14]}} , in48[14:3] };

   // m48_12 = W*in
   wire signed [14:0] m48_12;
   assign m48_12 =15'b0;

   // m48_13 = W*in
   wire signed [14:0] m48_13;
   assign m48_13 =15'b0;

   // m48_14 = W*in
   wire signed [14:0] m48_14;
   assign m48_14 =15'b0;

   // m48_15 = W*in
   wire signed [14:0] m48_15;
   assign m48_15 =15'b0;

   // m48_16 = W*in
   wire signed [14:0] m48_16;
   assign m48_16 =15'b0;

   // m48_17 = W*in
   wire signed [14:0] m48_17;
   assign m48_17 =15'b0;

   // m48_18 = W*in
   wire signed [14:0] m48_18;
   assign m48_18 =15'b0;

   // m48_19 = W*in
   wire signed [14:0] m48_19;
   assign m48_19 ={ {4{in48[14]}} , in48[14:4] };

   // m48_20 = W*in
   wire signed [14:0] m48_20;
   assign m48_20 ={ {4{neg48[14]}} , neg48[14:4] };

   // m48_21 = W*in
   wire signed [14:0] m48_21;
   assign m48_21 =15'b0;

   // m48_22 = W*in
   wire signed [14:0] m48_22;
   assign m48_22 ={ {2{neg48[14]}} , neg48[14:2] };

   // m48_23 = W*in
   wire signed [14:0] m48_23;
   assign m48_23 =15'b0;

   // m48_24 = W*in
   wire signed [14:0] m48_24;
   assign m48_24 =15'b0;

   // m48_25 = W*in
   wire signed [14:0] m48_25;
   assign m48_25 =15'b0;

   // m48_26 = W*in
   wire signed [14:0] m48_26;
   assign m48_26 =15'b0;

   // m48_27 = W*in
   wire signed [14:0] m48_27;
   assign m48_27 =15'b0;

   // m48_28 = W*in
   wire signed [14:0] m48_28;
   assign m48_28 ={ {4{neg48[14]}} , neg48[14:4] };

   // m48_29 = W*in
   wire signed [14:0] m48_29;
   assign m48_29 =15'b0;

   // m48_30 = W*in
   wire signed [14:0] m48_30;
   assign m48_30 ={ {4{in48[14]}} , in48[14:4] };

   // m48_31 = W*in
   wire signed [14:0] m48_31;
   assign m48_31 =15'b0;

   // m48_32 = W*in
   wire signed [14:0] m48_32;
   assign m48_32 ={ {3{in48[14]}} , in48[14:3] };

   // m48_33 = W*in
   wire signed [14:0] m48_33;
   assign m48_33 =15'b0;

   // m48_34 = W*in
   wire signed [14:0] m48_34;
   assign m48_34 =15'b0;

   // m48_35 = W*in
   wire signed [14:0] m48_35;
   assign m48_35 =15'b0;

   // m48_36 = W*in
   wire signed [14:0] m48_36;
   assign m48_36 =15'b0;

   // m48_37 = W*in
   wire signed [14:0] m48_37;
   assign m48_37 =15'b0;

   // m48_38 = W*in
   wire signed [14:0] m48_38;
   assign m48_38 =15'b0;

   // m48_39 = W*in
   wire signed [14:0] m48_39;
   assign m48_39 =15'b0;

   // m48_40 = W*in
   wire signed [14:0] m48_40;
   assign m48_40 =15'b0;

   // m48_41 = W*in
   wire signed [14:0] m48_41;
   assign m48_41 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_42 = W*in
   wire signed [14:0] m48_42;
   assign m48_42 =15'b0;

   // m48_43 = W*in
   wire signed [14:0] m48_43;
   assign m48_43 =15'b0;

   // m48_44 = W*in
   wire signed [14:0] m48_44;
   assign m48_44 =15'b0;

   // m48_45 = W*in
   wire signed [14:0] m48_45;
   assign m48_45 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_46 = W*in
   wire signed [14:0] m48_46;
   assign m48_46 =15'b0;

   // m48_47 = W*in
   wire signed [14:0] m48_47;
   assign m48_47 ={ {4{in48[14]}} , in48[14:4] };

   // m48_48 = W*in
   wire signed [14:0] m48_48;
   assign m48_48 =15'b0;

   // m48_49 = W*in
   wire signed [14:0] m48_49;
   assign m48_49 =15'b0;

   // m48_50 = W*in
   wire signed [14:0] m48_50;
   assign m48_50 =15'b0;

   // m48_51 = W*in
   wire signed [14:0] m48_51;
   assign m48_51 ={ {3{in48[14]}} , in48[14:3] };

   // m48_52 = W*in
   wire signed [14:0] m48_52;
   assign m48_52 =15'b0;

   // m48_53 = W*in
   wire signed [14:0] m48_53;
   assign m48_53 =15'b0;

   // m48_54 = W*in
   wire signed [14:0] m48_54;
   assign m48_54 =15'b0;

   // m48_55 = W*in
   wire signed [14:0] m48_55;
   assign m48_55 =15'b0;

   // m48_56 = W*in
   wire signed [14:0] m48_56;
   assign m48_56 =15'b0;

   // m48_57 = W*in
   wire signed [14:0] m48_57;
   assign m48_57 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_58 = W*in
   wire signed [14:0] m48_58;
   assign m48_58 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_59 = W*in
   wire signed [14:0] m48_59;
   assign m48_59 =15'b0;

   // m48_60 = W*in
   wire signed [14:0] m48_60;
   assign m48_60 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_61 = W*in
   wire signed [14:0] m48_61;
   assign m48_61 ={ {4{neg48[14]}} , neg48[14:4] };

   // m48_62 = W*in
   wire signed [14:0] m48_62;
   assign m48_62 ={ {2{neg48[14]}} , neg48[14:2] };

   // m48_63 = W*in
   wire signed [14:0] m48_63;
   assign m48_63 =15'b0;

   // m48_64 = W*in
   wire signed [14:0] m48_64;
   assign m48_64 ={ {4{neg48[14]}} , neg48[14:4] };

   // m48_65 = W*in
   wire signed [14:0] m48_65;
   assign m48_65 =15'b0;

   // m48_66 = W*in
   wire signed [14:0] m48_66;
   assign m48_66 ={ {3{in48[14]}} , in48[14:3] };

   // m48_67 = W*in
   wire signed [14:0] m48_67;
   assign m48_67 =15'b0;

   // m48_68 = W*in
   wire signed [14:0] m48_68;
   assign m48_68 =15'b0;

   // m48_69 = W*in
   wire signed [14:0] m48_69;
   assign m48_69 ={ {4{in48[14]}} , in48[14:4] };

   // m48_70 = W*in
   wire signed [14:0] m48_70;
   assign m48_70 =15'b0;

   // m48_71 = W*in
   wire signed [14:0] m48_71;
   assign m48_71 ={ {4{in48[14]}} , in48[14:4] };

   // m48_72 = W*in
   wire signed [14:0] m48_72;
   assign m48_72 =15'b0;

   // m48_73 = W*in
   wire signed [14:0] m48_73;
   assign m48_73 =15'b0;

   // m48_74 = W*in
   wire signed [14:0] m48_74;
   assign m48_74 ={ {4{neg48[14]}} , neg48[14:4] };

   // m48_75 = W*in
   wire signed [14:0] m48_75;
   assign m48_75 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_76 = W*in
   wire signed [14:0] m48_76;
   assign m48_76 =15'b0;

   // m48_77 = W*in
   wire signed [14:0] m48_77;
   assign m48_77 =15'b0;

   // m48_78 = W*in
   wire signed [14:0] m48_78;
   assign m48_78 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_79 = W*in
   wire signed [14:0] m48_79;
   assign m48_79 ={ {3{in48[14]}} , in48[14:3] };

   // m48_80 = W*in
   wire signed [14:0] m48_80;
   assign m48_80 =15'b0;

   // m48_81 = W*in
   wire signed [14:0] m48_81;
   assign m48_81 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_82 = W*in
   wire signed [14:0] m48_82;
   assign m48_82 =15'b0;

   // m48_83 = W*in
   wire signed [14:0] m48_83;
   assign m48_83 =15'b0;

   // m48_84 = W*in
   wire signed [14:0] m48_84;
   assign m48_84 =15'b0;

   // m48_85 = W*in
   wire signed [14:0] m48_85;
   assign m48_85 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_86 = W*in
   wire signed [14:0] m48_86;
   assign m48_86 =15'b0;

   // m48_87 = W*in
   wire signed [14:0] m48_87;
   assign m48_87 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_88 = W*in
   wire signed [14:0] m48_88;
   assign m48_88 =15'b0;

   // m48_89 = W*in
   wire signed [14:0] m48_89;
   assign m48_89 =15'b0;

   // m48_90 = W*in
   wire signed [14:0] m48_90;
   assign m48_90 =15'b0;

   // m48_91 = W*in
   wire signed [14:0] m48_91;
   assign m48_91 =15'b0;

   // m48_92 = W*in
   wire signed [14:0] m48_92;
   assign m48_92 =15'b0;

   // m48_93 = W*in
   wire signed [14:0] m48_93;
   assign m48_93 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_94 = W*in
   wire signed [14:0] m48_94;
   assign m48_94 =15'b0;

   // m48_95 = W*in
   wire signed [14:0] m48_95;
   assign m48_95 ={ {3{in48[14]}} , in48[14:3] };

   // m48_96 = W*in
   wire signed [14:0] m48_96;
   assign m48_96 ={ {3{neg48[14]}} , neg48[14:3] };

   // m48_97 = W*in
   wire signed [14:0] m48_97;
   assign m48_97 =15'b0;

   // m48_98 = W*in
   wire signed [14:0] m48_98;
   assign m48_98 =15'b0;

   // m48_99 = W*in
   wire signed [14:0] m48_99;
   assign m48_99 =15'b0;

   // m48_100 = W*in
   wire signed [14:0] m48_100;
   assign m48_100 =15'b0;

   // m49_1 = W*in
   wire signed [14:0] m49_1;
   assign m49_1 =15'b0;

   // m49_2 = W*in
   wire signed [14:0] m49_2;
   assign m49_2 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_3 = W*in
   wire signed [14:0] m49_3;
   assign m49_3 =15'b0;

   // m49_4 = W*in
   wire signed [14:0] m49_4;
   assign m49_4 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_5 = W*in
   wire signed [14:0] m49_5;
   assign m49_5 =15'b0;

   // m49_6 = W*in
   wire signed [14:0] m49_6;
   assign m49_6 =15'b0;

   // m49_7 = W*in
   wire signed [14:0] m49_7;
   assign m49_7 =15'b0;

   // m49_8 = W*in
   wire signed [14:0] m49_8;
   assign m49_8 =15'b0;

   // m49_9 = W*in
   wire signed [14:0] m49_9;
   assign m49_9 =15'b0;

   // m49_10 = W*in
   wire signed [14:0] m49_10;
   assign m49_10 =15'b0;

   // m49_11 = W*in
   wire signed [14:0] m49_11;
   assign m49_11 =15'b0;

   // m49_12 = W*in
   wire signed [14:0] m49_12;
   assign m49_12 =15'b0;

   // m49_13 = W*in
   wire signed [14:0] m49_13;
   assign m49_13 ={ {2{neg49[14]}} , neg49[14:2] };

   // m49_14 = W*in
   wire signed [14:0] m49_14;
   assign m49_14 ={ {3{in49[14]}} , in49[14:3] };

   // m49_15 = W*in
   wire signed [14:0] m49_15;
   assign m49_15 =15'b0;

   // m49_16 = W*in
   wire signed [14:0] m49_16;
   assign m49_16 =15'b0;

   // m49_17 = W*in
   wire signed [14:0] m49_17;
   assign m49_17 =15'b0;

   // m49_18 = W*in
   wire signed [14:0] m49_18;
   assign m49_18 =15'b0;

   // m49_19 = W*in
   wire signed [14:0] m49_19;
   assign m49_19 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_20 = W*in
   wire signed [14:0] m49_20;
   assign m49_20 =15'b0;

   // m49_21 = W*in
   wire signed [14:0] m49_21;
   assign m49_21 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_22 = W*in
   wire signed [14:0] m49_22;
   assign m49_22 =15'b0;

   // m49_23 = W*in
   wire signed [14:0] m49_23;
   assign m49_23 =15'b0;

   // m49_24 = W*in
   wire signed [14:0] m49_24;
   assign m49_24 =15'b0;

   // m49_25 = W*in
   wire signed [14:0] m49_25;
   assign m49_25 =15'b0;

   // m49_26 = W*in
   wire signed [14:0] m49_26;
   assign m49_26 =15'b0;

   // m49_27 = W*in
   wire signed [14:0] m49_27;
   assign m49_27 =15'b0;

   // m49_28 = W*in
   wire signed [14:0] m49_28;
   assign m49_28 =15'b0;

   // m49_29 = W*in
   wire signed [14:0] m49_29;
   assign m49_29 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_30 = W*in
   wire signed [14:0] m49_30;
   assign m49_30 =15'b0;

   // m49_31 = W*in
   wire signed [14:0] m49_31;
   assign m49_31 ={ {3{in49[14]}} , in49[14:3] };

   // m49_32 = W*in
   wire signed [14:0] m49_32;
   assign m49_32 =15'b0;

   // m49_33 = W*in
   wire signed [14:0] m49_33;
   assign m49_33 =15'b0;

   // m49_34 = W*in
   wire signed [14:0] m49_34;
   assign m49_34 =15'b0;

   // m49_35 = W*in
   wire signed [14:0] m49_35;
   assign m49_35 =15'b0;

   // m49_36 = W*in
   wire signed [14:0] m49_36;
   assign m49_36 =15'b0;

   // m49_37 = W*in
   wire signed [14:0] m49_37;
   assign m49_37 =15'b0;

   // m49_38 = W*in
   wire signed [14:0] m49_38;
   assign m49_38 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_39 = W*in
   wire signed [14:0] m49_39;
   assign m49_39 =15'b0;

   // m49_40 = W*in
   wire signed [14:0] m49_40;
   assign m49_40 =15'b0;

   // m49_41 = W*in
   wire signed [14:0] m49_41;
   assign m49_41 =15'b0;

   // m49_42 = W*in
   wire signed [14:0] m49_42;
   assign m49_42 =15'b0;

   // m49_43 = W*in
   wire signed [14:0] m49_43;
   assign m49_43 ={ {3{in49[14]}} , in49[14:3] };

   // m49_44 = W*in
   wire signed [14:0] m49_44;
   assign m49_44 =15'b0;

   // m49_45 = W*in
   wire signed [14:0] m49_45;
   assign m49_45 =15'b0;

   // m49_46 = W*in
   wire signed [14:0] m49_46;
   assign m49_46 =15'b0;

   // m49_47 = W*in
   wire signed [14:0] m49_47;
   assign m49_47 ={ {2{in49[14]}} , in49[14:2] };

   // m49_48 = W*in
   wire signed [14:0] m49_48;
   assign m49_48 =15'b0;

   // m49_49 = W*in
   wire signed [14:0] m49_49;
   assign m49_49 =15'b0;

   // m49_50 = W*in
   wire signed [14:0] m49_50;
   assign m49_50 =15'b0;

   // m49_51 = W*in
   wire signed [14:0] m49_51;
   assign m49_51 =15'b0;

   // m49_52 = W*in
   wire signed [14:0] m49_52;
   assign m49_52 =15'b0;

   // m49_53 = W*in
   wire signed [14:0] m49_53;
   assign m49_53 ={ {3{in49[14]}} , in49[14:3] };

   // m49_54 = W*in
   wire signed [14:0] m49_54;
   assign m49_54 =15'b0;

   // m49_55 = W*in
   wire signed [14:0] m49_55;
   assign m49_55 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_56 = W*in
   wire signed [14:0] m49_56;
   assign m49_56 ={ {3{in49[14]}} , in49[14:3] };

   // m49_57 = W*in
   wire signed [14:0] m49_57;
   assign m49_57 =15'b0;

   // m49_58 = W*in
   wire signed [14:0] m49_58;
   assign m49_58 =15'b0;

   // m49_59 = W*in
   wire signed [14:0] m49_59;
   assign m49_59 ={ {3{in49[14]}} , in49[14:3] };

   // m49_60 = W*in
   wire signed [14:0] m49_60;
   assign m49_60 ={ {4{neg49[14]}} , neg49[14:4] };

   // m49_61 = W*in
   wire signed [14:0] m49_61;
   assign m49_61 =15'b0;

   // m49_62 = W*in
   wire signed [14:0] m49_62;
   assign m49_62 =15'b0;

   // m49_63 = W*in
   wire signed [14:0] m49_63;
   assign m49_63 =15'b0;

   // m49_64 = W*in
   wire signed [14:0] m49_64;
   assign m49_64 =15'b0;

   // m49_65 = W*in
   wire signed [14:0] m49_65;
   assign m49_65 =15'b0;

   // m49_66 = W*in
   wire signed [14:0] m49_66;
   assign m49_66 =15'b0;

   // m49_67 = W*in
   wire signed [14:0] m49_67;
   assign m49_67 =15'b0;

   // m49_68 = W*in
   wire signed [14:0] m49_68;
   assign m49_68 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_69 = W*in
   wire signed [14:0] m49_69;
   assign m49_69 =15'b0;

   // m49_70 = W*in
   wire signed [14:0] m49_70;
   assign m49_70 =15'b0;

   // m49_71 = W*in
   wire signed [14:0] m49_71;
   assign m49_71 =15'b0;

   // m49_72 = W*in
   wire signed [14:0] m49_72;
   assign m49_72 =15'b0;

   // m49_73 = W*in
   wire signed [14:0] m49_73;
   assign m49_73 =15'b0;

   // m49_74 = W*in
   wire signed [14:0] m49_74;
   assign m49_74 =15'b0;

   // m49_75 = W*in
   wire signed [14:0] m49_75;
   assign m49_75 =15'b0;

   // m49_76 = W*in
   wire signed [14:0] m49_76;
   assign m49_76 =15'b0;

   // m49_77 = W*in
   wire signed [14:0] m49_77;
   assign m49_77 =15'b0;

   // m49_78 = W*in
   wire signed [14:0] m49_78;
   assign m49_78 =15'b0;

   // m49_79 = W*in
   wire signed [14:0] m49_79;
   assign m49_79 ={ {3{in49[14]}} , in49[14:3] };

   // m49_80 = W*in
   wire signed [14:0] m49_80;
   assign m49_80 =15'b0;

   // m49_81 = W*in
   wire signed [14:0] m49_81;
   assign m49_81 =15'b0;

   // m49_82 = W*in
   wire signed [14:0] m49_82;
   assign m49_82 =15'b0;

   // m49_83 = W*in
   wire signed [14:0] m49_83;
   assign m49_83 =15'b0;

   // m49_84 = W*in
   wire signed [14:0] m49_84;
   assign m49_84 ={ {3{neg49[14]}} , neg49[14:3] };

   // m49_85 = W*in
   wire signed [14:0] m49_85;
   assign m49_85 =15'b0;

   // m49_86 = W*in
   wire signed [14:0] m49_86;
   assign m49_86 =15'b0;

   // m49_87 = W*in
   wire signed [14:0] m49_87;
   assign m49_87 =15'b0;

   // m49_88 = W*in
   wire signed [14:0] m49_88;
   assign m49_88 =15'b0;

   // m49_89 = W*in
   wire signed [14:0] m49_89;
   assign m49_89 =15'b0;

   // m49_90 = W*in
   wire signed [14:0] m49_90;
   assign m49_90 =15'b0;

   // m49_91 = W*in
   wire signed [14:0] m49_91;
   assign m49_91 ={ {3{in49[14]}} , in49[14:3] };

   // m49_92 = W*in
   wire signed [14:0] m49_92;
   assign m49_92 =15'b0;

   // m49_93 = W*in
   wire signed [14:0] m49_93;
   assign m49_93 ={ {3{in49[14]}} , in49[14:3] };

   // m49_94 = W*in
   wire signed [14:0] m49_94;
   assign m49_94 ={ {3{in49[14]}} , in49[14:3] };

   // m49_95 = W*in
   wire signed [14:0] m49_95;
   assign m49_95 =15'b0;

   // m49_96 = W*in
   wire signed [14:0] m49_96;
   assign m49_96 =15'b0;

   // m49_97 = W*in
   wire signed [14:0] m49_97;
   assign m49_97 =15'b0;

   // m49_98 = W*in
   wire signed [14:0] m49_98;
   assign m49_98 =15'b0;

   // m49_99 = W*in
   wire signed [14:0] m49_99;
   assign m49_99 =15'b0;

   // m49_100 = W*in
   wire signed [14:0] m49_100;
   assign m49_100 =15'b0;

   // m50_1 = W*in
   wire signed [14:0] m50_1;
   assign m50_1 =15'b0;

   // m50_2 = W*in
   wire signed [14:0] m50_2;
   assign m50_2 =15'b0;

   // m50_3 = W*in
   wire signed [14:0] m50_3;
   assign m50_3 =15'b0;

   // m50_4 = W*in
   wire signed [14:0] m50_4;
   assign m50_4 =15'b0;

   // m50_5 = W*in
   wire signed [14:0] m50_5;
   assign m50_5 =15'b0;

   // m50_6 = W*in
   wire signed [14:0] m50_6;
   assign m50_6 =15'b0;

   // m50_7 = W*in
   wire signed [14:0] m50_7;
   assign m50_7 =15'b0;

   // m50_8 = W*in
   wire signed [14:0] m50_8;
   assign m50_8 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_9 = W*in
   wire signed [14:0] m50_9;
   assign m50_9 =15'b0;

   // m50_10 = W*in
   wire signed [14:0] m50_10;
   assign m50_10 =15'b0;

   // m50_11 = W*in
   wire signed [14:0] m50_11;
   assign m50_11 ={ {3{in50[14]}} , in50[14:3] };

   // m50_12 = W*in
   wire signed [14:0] m50_12;
   assign m50_12 ={ {3{in50[14]}} , in50[14:3] };

   // m50_13 = W*in
   wire signed [14:0] m50_13;
   assign m50_13 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_14 = W*in
   wire signed [14:0] m50_14;
   assign m50_14 =15'b0;

   // m50_15 = W*in
   wire signed [14:0] m50_15;
   assign m50_15 =15'b0;

   // m50_16 = W*in
   wire signed [14:0] m50_16;
   assign m50_16 ={ {3{in50[14]}} , in50[14:3] };

   // m50_17 = W*in
   wire signed [14:0] m50_17;
   assign m50_17 =15'b0;

   // m50_18 = W*in
   wire signed [14:0] m50_18;
   assign m50_18 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_19 = W*in
   wire signed [14:0] m50_19;
   assign m50_19 ={ {3{in50[14]}} , in50[14:3] };

   // m50_20 = W*in
   wire signed [14:0] m50_20;
   assign m50_20 ={ {4{neg50[14]}} , neg50[14:4] };

   // m50_21 = W*in
   wire signed [14:0] m50_21;
   assign m50_21 =15'b0;

   // m50_22 = W*in
   wire signed [14:0] m50_22;
   assign m50_22 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_23 = W*in
   wire signed [14:0] m50_23;
   assign m50_23 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_24 = W*in
   wire signed [14:0] m50_24;
   assign m50_24 =15'b0;

   // m50_25 = W*in
   wire signed [14:0] m50_25;
   assign m50_25 =15'b0;

   // m50_26 = W*in
   wire signed [14:0] m50_26;
   assign m50_26 =15'b0;

   // m50_27 = W*in
   wire signed [14:0] m50_27;
   assign m50_27 =15'b0;

   // m50_28 = W*in
   wire signed [14:0] m50_28;
   assign m50_28 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_29 = W*in
   wire signed [14:0] m50_29;
   assign m50_29 =15'b0;

   // m50_30 = W*in
   wire signed [14:0] m50_30;
   assign m50_30 ={ {3{in50[14]}} , in50[14:3] };

   // m50_31 = W*in
   wire signed [14:0] m50_31;
   assign m50_31 =15'b0;

   // m50_32 = W*in
   wire signed [14:0] m50_32;
   assign m50_32 =15'b0;

   // m50_33 = W*in
   wire signed [14:0] m50_33;
   assign m50_33 =15'b0;

   // m50_34 = W*in
   wire signed [14:0] m50_34;
   assign m50_34 =15'b0;

   // m50_35 = W*in
   wire signed [14:0] m50_35;
   assign m50_35 =15'b0;

   // m50_36 = W*in
   wire signed [14:0] m50_36;
   assign m50_36 =15'b0;

   // m50_37 = W*in
   wire signed [14:0] m50_37;
   assign m50_37 =15'b0;

   // m50_38 = W*in
   wire signed [14:0] m50_38;
   assign m50_38 =15'b0;

   // m50_39 = W*in
   wire signed [14:0] m50_39;
   assign m50_39 =15'b0;

   // m50_40 = W*in
   wire signed [14:0] m50_40;
   assign m50_40 =15'b0;

   // m50_41 = W*in
   wire signed [14:0] m50_41;
   assign m50_41 =15'b0;

   // m50_42 = W*in
   wire signed [14:0] m50_42;
   assign m50_42 =15'b0;

   // m50_43 = W*in
   wire signed [14:0] m50_43;
   assign m50_43 =15'b0;

   // m50_44 = W*in
   wire signed [14:0] m50_44;
   assign m50_44 =15'b0;

   // m50_45 = W*in
   wire signed [14:0] m50_45;
   assign m50_45 =15'b0;

   // m50_46 = W*in
   wire signed [14:0] m50_46;
   assign m50_46 ={ {3{in50[14]}} , in50[14:3] };

   // m50_47 = W*in
   wire signed [14:0] m50_47;
   assign m50_47 ={ {3{in50[14]}} , in50[14:3] };

   // m50_48 = W*in
   wire signed [14:0] m50_48;
   assign m50_48 =15'b0;

   // m50_49 = W*in
   wire signed [14:0] m50_49;
   assign m50_49 =15'b0;

   // m50_50 = W*in
   wire signed [14:0] m50_50;
   assign m50_50 =15'b0;

   // m50_51 = W*in
   wire signed [14:0] m50_51;
   assign m50_51 =15'b0;

   // m50_52 = W*in
   wire signed [14:0] m50_52;
   assign m50_52 =15'b0;

   // m50_53 = W*in
   wire signed [14:0] m50_53;
   assign m50_53 =15'b0;

   // m50_54 = W*in
   wire signed [14:0] m50_54;
   assign m50_54 =15'b0;

   // m50_55 = W*in
   wire signed [14:0] m50_55;
   assign m50_55 =15'b0;

   // m50_56 = W*in
   wire signed [14:0] m50_56;
   assign m50_56 =15'b0;

   // m50_57 = W*in
   wire signed [14:0] m50_57;
   assign m50_57 =15'b0;

   // m50_58 = W*in
   wire signed [14:0] m50_58;
   assign m50_58 =15'b0;

   // m50_59 = W*in
   wire signed [14:0] m50_59;
   assign m50_59 ={ {3{in50[14]}} , in50[14:3] };

   // m50_60 = W*in
   wire signed [14:0] m50_60;
   assign m50_60 ={ {4{neg50[14]}} , neg50[14:4] };

   // m50_61 = W*in
   wire signed [14:0] m50_61;
   assign m50_61 =15'b0;

   // m50_62 = W*in
   wire signed [14:0] m50_62;
   assign m50_62 =15'b0;

   // m50_63 = W*in
   wire signed [14:0] m50_63;
   assign m50_63 =15'b0;

   // m50_64 = W*in
   wire signed [14:0] m50_64;
   assign m50_64 =15'b0;

   // m50_65 = W*in
   wire signed [14:0] m50_65;
   assign m50_65 ={ {3{in50[14]}} , in50[14:3] };

   // m50_66 = W*in
   wire signed [14:0] m50_66;
   assign m50_66 =15'b0;

   // m50_67 = W*in
   wire signed [14:0] m50_67;
   assign m50_67 =15'b0;

   // m50_68 = W*in
   wire signed [14:0] m50_68;
   assign m50_68 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_69 = W*in
   wire signed [14:0] m50_69;
   assign m50_69 ={ {3{in50[14]}} , in50[14:3] };

   // m50_70 = W*in
   wire signed [14:0] m50_70;
   assign m50_70 =15'b0;

   // m50_71 = W*in
   wire signed [14:0] m50_71;
   assign m50_71 =15'b0;

   // m50_72 = W*in
   wire signed [14:0] m50_72;
   assign m50_72 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_73 = W*in
   wire signed [14:0] m50_73;
   assign m50_73 =15'b0;

   // m50_74 = W*in
   wire signed [14:0] m50_74;
   assign m50_74 ={ {4{neg50[14]}} , neg50[14:4] };

   // m50_75 = W*in
   wire signed [14:0] m50_75;
   assign m50_75 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_76 = W*in
   wire signed [14:0] m50_76;
   assign m50_76 =15'b0;

   // m50_77 = W*in
   wire signed [14:0] m50_77;
   assign m50_77 ={ {3{in50[14]}} , in50[14:3] };

   // m50_78 = W*in
   wire signed [14:0] m50_78;
   assign m50_78 ={ {3{neg50[14]}} , neg50[14:3] };

   // m50_79 = W*in
   wire signed [14:0] m50_79;
   assign m50_79 ={ {3{in50[14]}} , in50[14:3] };

   // m50_80 = W*in
   wire signed [14:0] m50_80;
   assign m50_80 =15'b0;

   // m50_81 = W*in
   wire signed [14:0] m50_81;
   assign m50_81 =15'b0;

   // m50_82 = W*in
   wire signed [14:0] m50_82;
   assign m50_82 =15'b0;

   // m50_83 = W*in
   wire signed [14:0] m50_83;
   assign m50_83 =15'b0;

   // m50_84 = W*in
   wire signed [14:0] m50_84;
   assign m50_84 =15'b0;

   // m50_85 = W*in
   wire signed [14:0] m50_85;
   assign m50_85 =15'b0;

   // m50_86 = W*in
   wire signed [14:0] m50_86;
   assign m50_86 ={ {3{in50[14]}} , in50[14:3] };

   // m50_87 = W*in
   wire signed [14:0] m50_87;
   assign m50_87 =15'b0;

   // m50_88 = W*in
   wire signed [14:0] m50_88;
   assign m50_88 =15'b0;

   // m50_89 = W*in
   wire signed [14:0] m50_89;
   assign m50_89 =15'b0;

   // m50_90 = W*in
   wire signed [14:0] m50_90;
   assign m50_90 =15'b0;

   // m50_91 = W*in
   wire signed [14:0] m50_91;
   assign m50_91 =15'b0;

   // m50_92 = W*in
   wire signed [14:0] m50_92;
   assign m50_92 ={ {3{in50[14]}} , in50[14:3] };

   // m50_93 = W*in
   wire signed [14:0] m50_93;
   assign m50_93 =15'b0;

   // m50_94 = W*in
   wire signed [14:0] m50_94;
   assign m50_94 ={ {3{in50[14]}} , in50[14:3] };

   // m50_95 = W*in
   wire signed [14:0] m50_95;
   assign m50_95 ={ {3{in50[14]}} , in50[14:3] };

   // m50_96 = W*in
   wire signed [14:0] m50_96;
   assign m50_96 =15'b0;

   // m50_97 = W*in
   wire signed [14:0] m50_97;
   assign m50_97 =15'b0;

   // m50_98 = W*in
   wire signed [14:0] m50_98;
   assign m50_98 =15'b0;

   // m50_99 = W*in
   wire signed [14:0] m50_99;
   assign m50_99 =15'b0;

   // m50_100 = W*in
   wire signed [14:0] m50_100;
   assign m50_100 =15'b0;

   // m51_1 = W*in
   wire signed [14:0] m51_1;
   assign m51_1 =15'b0;

   // m51_2 = W*in
   wire signed [14:0] m51_2;
   assign m51_2 =15'b0;

   // m51_3 = W*in
   wire signed [14:0] m51_3;
   assign m51_3 =15'b0;

   // m51_4 = W*in
   wire signed [14:0] m51_4;
   assign m51_4 =15'b0;

   // m51_5 = W*in
   wire signed [14:0] m51_5;
   assign m51_5 =15'b0;

   // m51_6 = W*in
   wire signed [14:0] m51_6;
   assign m51_6 =15'b0;

   // m51_7 = W*in
   wire signed [14:0] m51_7;
   assign m51_7 =15'b0;

   // m51_8 = W*in
   wire signed [14:0] m51_8;
   assign m51_8 ={ {3{in51[14]}} , in51[14:3] };

   // m51_9 = W*in
   wire signed [14:0] m51_9;
   assign m51_9 =15'b0;

   // m51_10 = W*in
   wire signed [14:0] m51_10;
   assign m51_10 =15'b0;

   // m51_11 = W*in
   wire signed [14:0] m51_11;
   assign m51_11 =15'b0;

   // m51_12 = W*in
   wire signed [14:0] m51_12;
   assign m51_12 =15'b0;

   // m51_13 = W*in
   wire signed [14:0] m51_13;
   assign m51_13 =15'b0;

   // m51_14 = W*in
   wire signed [14:0] m51_14;
   assign m51_14 =15'b0;

   // m51_15 = W*in
   wire signed [14:0] m51_15;
   assign m51_15 =15'b0;

   // m51_16 = W*in
   wire signed [14:0] m51_16;
   assign m51_16 =15'b0;

   // m51_17 = W*in
   wire signed [14:0] m51_17;
   assign m51_17 =15'b0;

   // m51_18 = W*in
   wire signed [14:0] m51_18;
   assign m51_18 =15'b0;

   // m51_19 = W*in
   wire signed [14:0] m51_19;
   assign m51_19 =15'b0;

   // m51_20 = W*in
   wire signed [14:0] m51_20;
   assign m51_20 ={ {4{neg51[14]}} , neg51[14:4] };

   // m51_21 = W*in
   wire signed [14:0] m51_21;
   assign m51_21 =15'b0;

   // m51_22 = W*in
   wire signed [14:0] m51_22;
   assign m51_22 =15'b0;

   // m51_23 = W*in
   wire signed [14:0] m51_23;
   assign m51_23 =15'b0;

   // m51_24 = W*in
   wire signed [14:0] m51_24;
   assign m51_24 =15'b0;

   // m51_25 = W*in
   wire signed [14:0] m51_25;
   assign m51_25 =15'b0;

   // m51_26 = W*in
   wire signed [14:0] m51_26;
   assign m51_26 =15'b0;

   // m51_27 = W*in
   wire signed [14:0] m51_27;
   assign m51_27 =15'b0;

   // m51_28 = W*in
   wire signed [14:0] m51_28;
   assign m51_28 =15'b0;

   // m51_29 = W*in
   wire signed [14:0] m51_29;
   assign m51_29 =15'b0;

   // m51_30 = W*in
   wire signed [14:0] m51_30;
   assign m51_30 =15'b0;

   // m51_31 = W*in
   wire signed [14:0] m51_31;
   assign m51_31 =15'b0;

   // m51_32 = W*in
   wire signed [14:0] m51_32;
   assign m51_32 =15'b0;

   // m51_33 = W*in
   wire signed [14:0] m51_33;
   assign m51_33 =15'b0;

   // m51_34 = W*in
   wire signed [14:0] m51_34;
   assign m51_34 ={ {4{neg51[14]}} , neg51[14:4] };

   // m51_35 = W*in
   wire signed [14:0] m51_35;
   assign m51_35 =15'b0;

   // m51_36 = W*in
   wire signed [14:0] m51_36;
   assign m51_36 =15'b0;

   // m51_37 = W*in
   wire signed [14:0] m51_37;
   assign m51_37 =15'b0;

   // m51_38 = W*in
   wire signed [14:0] m51_38;
   assign m51_38 =15'b0;

   // m51_39 = W*in
   wire signed [14:0] m51_39;
   assign m51_39 =15'b0;

   // m51_40 = W*in
   wire signed [14:0] m51_40;
   assign m51_40 =15'b0;

   // m51_41 = W*in
   wire signed [14:0] m51_41;
   assign m51_41 =15'b0;

   // m51_42 = W*in
   wire signed [14:0] m51_42;
   assign m51_42 =15'b0;

   // m51_43 = W*in
   wire signed [14:0] m51_43;
   assign m51_43 =15'b0;

   // m51_44 = W*in
   wire signed [14:0] m51_44;
   assign m51_44 =15'b0;

   // m51_45 = W*in
   wire signed [14:0] m51_45;
   assign m51_45 ={ {3{neg51[14]}} , neg51[14:3] };

   // m51_46 = W*in
   wire signed [14:0] m51_46;
   assign m51_46 =15'b0;

   // m51_47 = W*in
   wire signed [14:0] m51_47;
   assign m51_47 =15'b0;

   // m51_48 = W*in
   wire signed [14:0] m51_48;
   assign m51_48 =15'b0;

   // m51_49 = W*in
   wire signed [14:0] m51_49;
   assign m51_49 =15'b0;

   // m51_50 = W*in
   wire signed [14:0] m51_50;
   assign m51_50 =15'b0;

   // m51_51 = W*in
   wire signed [14:0] m51_51;
   assign m51_51 ={ {3{in51[14]}} , in51[14:3] };

   // m51_52 = W*in
   wire signed [14:0] m51_52;
   assign m51_52 =15'b0;

   // m51_53 = W*in
   wire signed [14:0] m51_53;
   assign m51_53 =15'b0;

   // m51_54 = W*in
   wire signed [14:0] m51_54;
   assign m51_54 =15'b0;

   // m51_55 = W*in
   wire signed [14:0] m51_55;
   assign m51_55 =15'b0;

   // m51_56 = W*in
   wire signed [14:0] m51_56;
   assign m51_56 =15'b0;

   // m51_57 = W*in
   wire signed [14:0] m51_57;
   assign m51_57 =15'b0;

   // m51_58 = W*in
   wire signed [14:0] m51_58;
   assign m51_58 ={ {3{in51[14]}} , in51[14:3] };

   // m51_59 = W*in
   wire signed [14:0] m51_59;
   assign m51_59 ={ {4{neg51[14]}} , neg51[14:4] };

   // m51_60 = W*in
   wire signed [14:0] m51_60;
   assign m51_60 =15'b0;

   // m51_61 = W*in
   wire signed [14:0] m51_61;
   assign m51_61 =15'b0;

   // m51_62 = W*in
   wire signed [14:0] m51_62;
   assign m51_62 ={ {3{neg51[14]}} , neg51[14:3] };

   // m51_63 = W*in
   wire signed [14:0] m51_63;
   assign m51_63 ={ {3{in51[14]}} , in51[14:3] };

   // m51_64 = W*in
   wire signed [14:0] m51_64;
   assign m51_64 =15'b0;

   // m51_65 = W*in
   wire signed [14:0] m51_65;
   assign m51_65 =15'b0;

   // m51_66 = W*in
   wire signed [14:0] m51_66;
   assign m51_66 =15'b0;

   // m51_67 = W*in
   wire signed [14:0] m51_67;
   assign m51_67 ={ {4{neg51[14]}} , neg51[14:4] };

   // m51_68 = W*in
   wire signed [14:0] m51_68;
   assign m51_68 =15'b0;

   // m51_69 = W*in
   wire signed [14:0] m51_69;
   assign m51_69 =15'b0;

   // m51_70 = W*in
   wire signed [14:0] m51_70;
   assign m51_70 =15'b0;

   // m51_71 = W*in
   wire signed [14:0] m51_71;
   assign m51_71 =15'b0;

   // m51_72 = W*in
   wire signed [14:0] m51_72;
   assign m51_72 =15'b0;

   // m51_73 = W*in
   wire signed [14:0] m51_73;
   assign m51_73 =15'b0;

   // m51_74 = W*in
   wire signed [14:0] m51_74;
   assign m51_74 =15'b0;

   // m51_75 = W*in
   wire signed [14:0] m51_75;
   assign m51_75 ={ {3{neg51[14]}} , neg51[14:3] };

   // m51_76 = W*in
   wire signed [14:0] m51_76;
   assign m51_76 =15'b0;

   // m51_77 = W*in
   wire signed [14:0] m51_77;
   assign m51_77 =15'b0;

   // m51_78 = W*in
   wire signed [14:0] m51_78;
   assign m51_78 =15'b0;

   // m51_79 = W*in
   wire signed [14:0] m51_79;
   assign m51_79 =15'b0;

   // m51_80 = W*in
   wire signed [14:0] m51_80;
   assign m51_80 =15'b0;

   // m51_81 = W*in
   wire signed [14:0] m51_81;
   assign m51_81 =15'b0;

   // m51_82 = W*in
   wire signed [14:0] m51_82;
   assign m51_82 =15'b0;

   // m51_83 = W*in
   wire signed [14:0] m51_83;
   assign m51_83 =15'b0;

   // m51_84 = W*in
   wire signed [14:0] m51_84;
   assign m51_84 =15'b0;

   // m51_85 = W*in
   wire signed [14:0] m51_85;
   assign m51_85 =15'b0;

   // m51_86 = W*in
   wire signed [14:0] m51_86;
   assign m51_86 ={ {3{neg51[14]}} , neg51[14:3] };

   // m51_87 = W*in
   wire signed [14:0] m51_87;
   assign m51_87 =15'b0;

   // m51_88 = W*in
   wire signed [14:0] m51_88;
   assign m51_88 =15'b0;

   // m51_89 = W*in
   wire signed [14:0] m51_89;
   assign m51_89 =15'b0;

   // m51_90 = W*in
   wire signed [14:0] m51_90;
   assign m51_90 ={ {3{neg51[14]}} , neg51[14:3] };

   // m51_91 = W*in
   wire signed [14:0] m51_91;
   assign m51_91 =15'b0;

   // m51_92 = W*in
   wire signed [14:0] m51_92;
   assign m51_92 =15'b0;

   // m51_93 = W*in
   wire signed [14:0] m51_93;
   assign m51_93 =15'b0;

   // m51_94 = W*in
   wire signed [14:0] m51_94;
   assign m51_94 =15'b0;

   // m51_95 = W*in
   wire signed [14:0] m51_95;
   assign m51_95 ={ {4{neg51[14]}} , neg51[14:4] };

   // m51_96 = W*in
   wire signed [14:0] m51_96;
   assign m51_96 =15'b0;

   // m51_97 = W*in
   wire signed [14:0] m51_97;
   assign m51_97 =15'b0;

   // m51_98 = W*in
   wire signed [14:0] m51_98;
   assign m51_98 =15'b0;

   // m51_99 = W*in
   wire signed [14:0] m51_99;
   assign m51_99 =15'b0;

   // m51_100 = W*in
   wire signed [14:0] m51_100;
   assign m51_100 =15'b0;

   // m52_1 = W*in
   wire signed [14:0] m52_1;
   assign m52_1 =15'b0;

   // m52_2 = W*in
   wire signed [14:0] m52_2;
   assign m52_2 =15'b0;

   // m52_3 = W*in
   wire signed [14:0] m52_3;
   assign m52_3 =15'b0;

   // m52_4 = W*in
   wire signed [14:0] m52_4;
   assign m52_4 ={ {3{neg52[14]}} , neg52[14:3] };

   // m52_5 = W*in
   wire signed [14:0] m52_5;
   assign m52_5 =15'b0;

   // m52_6 = W*in
   wire signed [14:0] m52_6;
   assign m52_6 =15'b0;

   // m52_7 = W*in
   wire signed [14:0] m52_7;
   assign m52_7 =15'b0;

   // m52_8 = W*in
   wire signed [14:0] m52_8;
   assign m52_8 =15'b0;

   // m52_9 = W*in
   wire signed [14:0] m52_9;
   assign m52_9 =15'b0;

   // m52_10 = W*in
   wire signed [14:0] m52_10;
   assign m52_10 =15'b0;

   // m52_11 = W*in
   wire signed [14:0] m52_11;
   assign m52_11 =15'b0;

   // m52_12 = W*in
   wire signed [14:0] m52_12;
   assign m52_12 =15'b0;

   // m52_13 = W*in
   wire signed [14:0] m52_13;
   assign m52_13 =15'b0;

   // m52_14 = W*in
   wire signed [14:0] m52_14;
   assign m52_14 =15'b0;

   // m52_15 = W*in
   wire signed [14:0] m52_15;
   assign m52_15 ={ {3{in52[14]}} , in52[14:3] };

   // m52_16 = W*in
   wire signed [14:0] m52_16;
   assign m52_16 =15'b0;

   // m52_17 = W*in
   wire signed [14:0] m52_17;
   assign m52_17 =15'b0;

   // m52_18 = W*in
   wire signed [14:0] m52_18;
   assign m52_18 =15'b0;

   // m52_19 = W*in
   wire signed [14:0] m52_19;
   assign m52_19 ={ {4{neg52[14]}} , neg52[14:4] };

   // m52_20 = W*in
   wire signed [14:0] m52_20;
   assign m52_20 =15'b0;

   // m52_21 = W*in
   wire signed [14:0] m52_21;
   assign m52_21 =15'b0;

   // m52_22 = W*in
   wire signed [14:0] m52_22;
   assign m52_22 ={ {4{in52[14]}} , in52[14:4] };

   // m52_23 = W*in
   wire signed [14:0] m52_23;
   assign m52_23 =15'b0;

   // m52_24 = W*in
   wire signed [14:0] m52_24;
   assign m52_24 =15'b0;

   // m52_25 = W*in
   wire signed [14:0] m52_25;
   assign m52_25 =15'b0;

   // m52_26 = W*in
   wire signed [14:0] m52_26;
   assign m52_26 =15'b0;

   // m52_27 = W*in
   wire signed [14:0] m52_27;
   assign m52_27 =15'b0;

   // m52_28 = W*in
   wire signed [14:0] m52_28;
   assign m52_28 ={ {3{neg52[14]}} , neg52[14:3] };

   // m52_29 = W*in
   wire signed [14:0] m52_29;
   assign m52_29 =15'b0;

   // m52_30 = W*in
   wire signed [14:0] m52_30;
   assign m52_30 =15'b0;

   // m52_31 = W*in
   wire signed [14:0] m52_31;
   assign m52_31 =15'b0;

   // m52_32 = W*in
   wire signed [14:0] m52_32;
   assign m52_32 ={ {4{neg52[14]}} , neg52[14:4] };

   // m52_33 = W*in
   wire signed [14:0] m52_33;
   assign m52_33 ={ {3{neg52[14]}} , neg52[14:3] };

   // m52_34 = W*in
   wire signed [14:0] m52_34;
   assign m52_34 =15'b0;

   // m52_35 = W*in
   wire signed [14:0] m52_35;
   assign m52_35 =15'b0;

   // m52_36 = W*in
   wire signed [14:0] m52_36;
   assign m52_36 =15'b0;

   // m52_37 = W*in
   wire signed [14:0] m52_37;
   assign m52_37 =15'b0;

   // m52_38 = W*in
   wire signed [14:0] m52_38;
   assign m52_38 ={ {3{neg52[14]}} , neg52[14:3] };

   // m52_39 = W*in
   wire signed [14:0] m52_39;
   assign m52_39 =15'b0;

   // m52_40 = W*in
   wire signed [14:0] m52_40;
   assign m52_40 =15'b0;

   // m52_41 = W*in
   wire signed [14:0] m52_41;
   assign m52_41 =15'b0;

   // m52_42 = W*in
   wire signed [14:0] m52_42;
   assign m52_42 =15'b0;

   // m52_43 = W*in
   wire signed [14:0] m52_43;
   assign m52_43 =15'b0;

   // m52_44 = W*in
   wire signed [14:0] m52_44;
   assign m52_44 ={ {3{neg52[14]}} , neg52[14:3] };

   // m52_45 = W*in
   wire signed [14:0] m52_45;
   assign m52_45 =15'b0;

   // m52_46 = W*in
   wire signed [14:0] m52_46;
   assign m52_46 =15'b0;

   // m52_47 = W*in
   wire signed [14:0] m52_47;
   assign m52_47 =15'b0;

   // m52_48 = W*in
   wire signed [14:0] m52_48;
   assign m52_48 =15'b0;

   // m52_49 = W*in
   wire signed [14:0] m52_49;
   assign m52_49 ={ {3{in52[14]}} , in52[14:3] };

   // m52_50 = W*in
   wire signed [14:0] m52_50;
   assign m52_50 =15'b0;

   // m52_51 = W*in
   wire signed [14:0] m52_51;
   assign m52_51 =15'b0;

   // m52_52 = W*in
   wire signed [14:0] m52_52;
   assign m52_52 =15'b0;

   // m52_53 = W*in
   wire signed [14:0] m52_53;
   assign m52_53 =15'b0;

   // m52_54 = W*in
   wire signed [14:0] m52_54;
   assign m52_54 =15'b0;

   // m52_55 = W*in
   wire signed [14:0] m52_55;
   assign m52_55 =15'b0;

   // m52_56 = W*in
   wire signed [14:0] m52_56;
   assign m52_56 =15'b0;

   // m52_57 = W*in
   wire signed [14:0] m52_57;
   assign m52_57 =15'b0;

   // m52_58 = W*in
   wire signed [14:0] m52_58;
   assign m52_58 =15'b0;

   // m52_59 = W*in
   wire signed [14:0] m52_59;
   assign m52_59 =15'b0;

   // m52_60 = W*in
   wire signed [14:0] m52_60;
   assign m52_60 =15'b0;

   // m52_61 = W*in
   wire signed [14:0] m52_61;
   assign m52_61 =15'b0;

   // m52_62 = W*in
   wire signed [14:0] m52_62;
   assign m52_62 =15'b0;

   // m52_63 = W*in
   wire signed [14:0] m52_63;
   assign m52_63 =15'b0;

   // m52_64 = W*in
   wire signed [14:0] m52_64;
   assign m52_64 ={ {4{in52[14]}} , in52[14:4] };

   // m52_65 = W*in
   wire signed [14:0] m52_65;
   assign m52_65 =15'b0;

   // m52_66 = W*in
   wire signed [14:0] m52_66;
   assign m52_66 =15'b0;

   // m52_67 = W*in
   wire signed [14:0] m52_67;
   assign m52_67 ={ {3{in52[14]}} , in52[14:3] };

   // m52_68 = W*in
   wire signed [14:0] m52_68;
   assign m52_68 ={ {4{neg52[14]}} , neg52[14:4] };

   // m52_69 = W*in
   wire signed [14:0] m52_69;
   assign m52_69 ={ {4{in52[14]}} , in52[14:4] };

   // m52_70 = W*in
   wire signed [14:0] m52_70;
   assign m52_70 =15'b0;

   // m52_71 = W*in
   wire signed [14:0] m52_71;
   assign m52_71 =15'b0;

   // m52_72 = W*in
   wire signed [14:0] m52_72;
   assign m52_72 =15'b0;

   // m52_73 = W*in
   wire signed [14:0] m52_73;
   assign m52_73 =15'b0;

   // m52_74 = W*in
   wire signed [14:0] m52_74;
   assign m52_74 =15'b0;

   // m52_75 = W*in
   wire signed [14:0] m52_75;
   assign m52_75 =15'b0;

   // m52_76 = W*in
   wire signed [14:0] m52_76;
   assign m52_76 =15'b0;

   // m52_77 = W*in
   wire signed [14:0] m52_77;
   assign m52_77 =15'b0;

   // m52_78 = W*in
   wire signed [14:0] m52_78;
   assign m52_78 =15'b0;

   // m52_79 = W*in
   wire signed [14:0] m52_79;
   assign m52_79 =15'b0;

   // m52_80 = W*in
   wire signed [14:0] m52_80;
   assign m52_80 =15'b0;

   // m52_81 = W*in
   wire signed [14:0] m52_81;
   assign m52_81 =15'b0;

   // m52_82 = W*in
   wire signed [14:0] m52_82;
   assign m52_82 =15'b0;

   // m52_83 = W*in
   wire signed [14:0] m52_83;
   assign m52_83 =15'b0;

   // m52_84 = W*in
   wire signed [14:0] m52_84;
   assign m52_84 =15'b0;

   // m52_85 = W*in
   wire signed [14:0] m52_85;
   assign m52_85 =15'b0;

   // m52_86 = W*in
   wire signed [14:0] m52_86;
   assign m52_86 =15'b0;

   // m52_87 = W*in
   wire signed [14:0] m52_87;
   assign m52_87 =15'b0;

   // m52_88 = W*in
   wire signed [14:0] m52_88;
   assign m52_88 =15'b0;

   // m52_89 = W*in
   wire signed [14:0] m52_89;
   assign m52_89 =15'b0;

   // m52_90 = W*in
   wire signed [14:0] m52_90;
   assign m52_90 =15'b0;

   // m52_91 = W*in
   wire signed [14:0] m52_91;
   assign m52_91 =15'b0;

   // m52_92 = W*in
   wire signed [14:0] m52_92;
   assign m52_92 ={ {3{in52[14]}} , in52[14:3] };

   // m52_93 = W*in
   wire signed [14:0] m52_93;
   assign m52_93 =15'b0;

   // m52_94 = W*in
   wire signed [14:0] m52_94;
   assign m52_94 ={ {3{neg52[14]}} , neg52[14:3] };

   // m52_95 = W*in
   wire signed [14:0] m52_95;
   assign m52_95 =15'b0;

   // m52_96 = W*in
   wire signed [14:0] m52_96;
   assign m52_96 =15'b0;

   // m52_97 = W*in
   wire signed [14:0] m52_97;
   assign m52_97 =15'b0;

   // m52_98 = W*in
   wire signed [14:0] m52_98;
   assign m52_98 =15'b0;

   // m52_99 = W*in
   wire signed [14:0] m52_99;
   assign m52_99 =15'b0;

   // m52_100 = W*in
   wire signed [14:0] m52_100;
   assign m52_100 =15'b0;

   // m53_1 = W*in
   wire signed [14:0] m53_1;
   assign m53_1 =15'b0;

   // m53_2 = W*in
   wire signed [14:0] m53_2;
   assign m53_2 =15'b0;

   // m53_3 = W*in
   wire signed [14:0] m53_3;
   assign m53_3 =15'b0;

   // m53_4 = W*in
   wire signed [14:0] m53_4;
   assign m53_4 =15'b0;

   // m53_5 = W*in
   wire signed [14:0] m53_5;
   assign m53_5 =15'b0;

   // m53_6 = W*in
   wire signed [14:0] m53_6;
   assign m53_6 =15'b0;

   // m53_7 = W*in
   wire signed [14:0] m53_7;
   assign m53_7 =15'b0;

   // m53_8 = W*in
   wire signed [14:0] m53_8;
   assign m53_8 =15'b0;

   // m53_9 = W*in
   wire signed [14:0] m53_9;
   assign m53_9 =15'b0;

   // m53_10 = W*in
   wire signed [14:0] m53_10;
   assign m53_10 ={ {3{in53[14]}} , in53[14:3] };

   // m53_11 = W*in
   wire signed [14:0] m53_11;
   assign m53_11 =15'b0;

   // m53_12 = W*in
   wire signed [14:0] m53_12;
   assign m53_12 ={ {3{in53[14]}} , in53[14:3] };

   // m53_13 = W*in
   wire signed [14:0] m53_13;
   assign m53_13 =15'b0;

   // m53_14 = W*in
   wire signed [14:0] m53_14;
   assign m53_14 =15'b0;

   // m53_15 = W*in
   wire signed [14:0] m53_15;
   assign m53_15 =15'b0;

   // m53_16 = W*in
   wire signed [14:0] m53_16;
   assign m53_16 ={ {3{in53[14]}} , in53[14:3] };

   // m53_17 = W*in
   wire signed [14:0] m53_17;
   assign m53_17 =15'b0;

   // m53_18 = W*in
   wire signed [14:0] m53_18;
   assign m53_18 =15'b0;

   // m53_19 = W*in
   wire signed [14:0] m53_19;
   assign m53_19 =15'b0;

   // m53_20 = W*in
   wire signed [14:0] m53_20;
   assign m53_20 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_21 = W*in
   wire signed [14:0] m53_21;
   assign m53_21 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_22 = W*in
   wire signed [14:0] m53_22;
   assign m53_22 =15'b0;

   // m53_23 = W*in
   wire signed [14:0] m53_23;
   assign m53_23 =15'b0;

   // m53_24 = W*in
   wire signed [14:0] m53_24;
   assign m53_24 =15'b0;

   // m53_25 = W*in
   wire signed [14:0] m53_25;
   assign m53_25 =15'b0;

   // m53_26 = W*in
   wire signed [14:0] m53_26;
   assign m53_26 ={ {3{in53[14]}} , in53[14:3] };

   // m53_27 = W*in
   wire signed [14:0] m53_27;
   assign m53_27 =15'b0;

   // m53_28 = W*in
   wire signed [14:0] m53_28;
   assign m53_28 ={ {4{neg53[14]}} , neg53[14:4] };

   // m53_29 = W*in
   wire signed [14:0] m53_29;
   assign m53_29 ={ {4{in53[14]}} , in53[14:4] };

   // m53_30 = W*in
   wire signed [14:0] m53_30;
   assign m53_30 ={ {4{in53[14]}} , in53[14:4] };

   // m53_31 = W*in
   wire signed [14:0] m53_31;
   assign m53_31 =15'b0;

   // m53_32 = W*in
   wire signed [14:0] m53_32;
   assign m53_32 =15'b0;

   // m53_33 = W*in
   wire signed [14:0] m53_33;
   assign m53_33 =15'b0;

   // m53_34 = W*in
   wire signed [14:0] m53_34;
   assign m53_34 =15'b0;

   // m53_35 = W*in
   wire signed [14:0] m53_35;
   assign m53_35 =15'b0;

   // m53_36 = W*in
   wire signed [14:0] m53_36;
   assign m53_36 =15'b0;

   // m53_37 = W*in
   wire signed [14:0] m53_37;
   assign m53_37 =15'b0;

   // m53_38 = W*in
   wire signed [14:0] m53_38;
   assign m53_38 =15'b0;

   // m53_39 = W*in
   wire signed [14:0] m53_39;
   assign m53_39 =15'b0;

   // m53_40 = W*in
   wire signed [14:0] m53_40;
   assign m53_40 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_41 = W*in
   wire signed [14:0] m53_41;
   assign m53_41 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_42 = W*in
   wire signed [14:0] m53_42;
   assign m53_42 =15'b0;

   // m53_43 = W*in
   wire signed [14:0] m53_43;
   assign m53_43 =15'b0;

   // m53_44 = W*in
   wire signed [14:0] m53_44;
   assign m53_44 =15'b0;

   // m53_45 = W*in
   wire signed [14:0] m53_45;
   assign m53_45 =15'b0;

   // m53_46 = W*in
   wire signed [14:0] m53_46;
   assign m53_46 ={ {3{in53[14]}} , in53[14:3] };

   // m53_47 = W*in
   wire signed [14:0] m53_47;
   assign m53_47 ={ {4{in53[14]}} , in53[14:4] };

   // m53_48 = W*in
   wire signed [14:0] m53_48;
   assign m53_48 =15'b0;

   // m53_49 = W*in
   wire signed [14:0] m53_49;
   assign m53_49 ={ {3{in53[14]}} , in53[14:3] };

   // m53_50 = W*in
   wire signed [14:0] m53_50;
   assign m53_50 =15'b0;

   // m53_51 = W*in
   wire signed [14:0] m53_51;
   assign m53_51 =15'b0;

   // m53_52 = W*in
   wire signed [14:0] m53_52;
   assign m53_52 =15'b0;

   // m53_53 = W*in
   wire signed [14:0] m53_53;
   assign m53_53 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_54 = W*in
   wire signed [14:0] m53_54;
   assign m53_54 =15'b0;

   // m53_55 = W*in
   wire signed [14:0] m53_55;
   assign m53_55 =15'b0;

   // m53_56 = W*in
   wire signed [14:0] m53_56;
   assign m53_56 =15'b0;

   // m53_57 = W*in
   wire signed [14:0] m53_57;
   assign m53_57 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_58 = W*in
   wire signed [14:0] m53_58;
   assign m53_58 =15'b0;

   // m53_59 = W*in
   wire signed [14:0] m53_59;
   assign m53_59 ={ {4{neg53[14]}} , neg53[14:4] };

   // m53_60 = W*in
   wire signed [14:0] m53_60;
   assign m53_60 =15'b0;

   // m53_61 = W*in
   wire signed [14:0] m53_61;
   assign m53_61 ={ {4{in53[14]}} , in53[14:4] };

   // m53_62 = W*in
   wire signed [14:0] m53_62;
   assign m53_62 =15'b0;

   // m53_63 = W*in
   wire signed [14:0] m53_63;
   assign m53_63 =15'b0;

   // m53_64 = W*in
   wire signed [14:0] m53_64;
   assign m53_64 ={ {4{neg53[14]}} , neg53[14:4] };

   // m53_65 = W*in
   wire signed [14:0] m53_65;
   assign m53_65 ={ {3{in53[14]}} , in53[14:3] };

   // m53_66 = W*in
   wire signed [14:0] m53_66;
   assign m53_66 ={ {3{in53[14]}} , in53[14:3] };

   // m53_67 = W*in
   wire signed [14:0] m53_67;
   assign m53_67 =15'b0;

   // m53_68 = W*in
   wire signed [14:0] m53_68;
   assign m53_68 ={ {4{neg53[14]}} , neg53[14:4] };

   // m53_69 = W*in
   wire signed [14:0] m53_69;
   assign m53_69 =15'b0;

   // m53_70 = W*in
   wire signed [14:0] m53_70;
   assign m53_70 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_71 = W*in
   wire signed [14:0] m53_71;
   assign m53_71 =15'b0;

   // m53_72 = W*in
   wire signed [14:0] m53_72;
   assign m53_72 =15'b0;

   // m53_73 = W*in
   wire signed [14:0] m53_73;
   assign m53_73 =15'b0;

   // m53_74 = W*in
   wire signed [14:0] m53_74;
   assign m53_74 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_75 = W*in
   wire signed [14:0] m53_75;
   assign m53_75 =15'b0;

   // m53_76 = W*in
   wire signed [14:0] m53_76;
   assign m53_76 =15'b0;

   // m53_77 = W*in
   wire signed [14:0] m53_77;
   assign m53_77 ={ {4{in53[14]}} , in53[14:4] };

   // m53_78 = W*in
   wire signed [14:0] m53_78;
   assign m53_78 =15'b0;

   // m53_79 = W*in
   wire signed [14:0] m53_79;
   assign m53_79 =15'b0;

   // m53_80 = W*in
   wire signed [14:0] m53_80;
   assign m53_80 =15'b0;

   // m53_81 = W*in
   wire signed [14:0] m53_81;
   assign m53_81 ={ {3{in53[14]}} , in53[14:3] };

   // m53_82 = W*in
   wire signed [14:0] m53_82;
   assign m53_82 =15'b0;

   // m53_83 = W*in
   wire signed [14:0] m53_83;
   assign m53_83 =15'b0;

   // m53_84 = W*in
   wire signed [14:0] m53_84;
   assign m53_84 ={ {3{in53[14]}} , in53[14:3] };

   // m53_85 = W*in
   wire signed [14:0] m53_85;
   assign m53_85 =15'b0;

   // m53_86 = W*in
   wire signed [14:0] m53_86;
   assign m53_86 =15'b0;

   // m53_87 = W*in
   wire signed [14:0] m53_87;
   assign m53_87 =15'b0;

   // m53_88 = W*in
   wire signed [14:0] m53_88;
   assign m53_88 =15'b0;

   // m53_89 = W*in
   wire signed [14:0] m53_89;
   assign m53_89 =15'b0;

   // m53_90 = W*in
   wire signed [14:0] m53_90;
   assign m53_90 =15'b0;

   // m53_91 = W*in
   wire signed [14:0] m53_91;
   assign m53_91 =15'b0;

   // m53_92 = W*in
   wire signed [14:0] m53_92;
   assign m53_92 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_93 = W*in
   wire signed [14:0] m53_93;
   assign m53_93 ={ {3{in53[14]}} , in53[14:3] };

   // m53_94 = W*in
   wire signed [14:0] m53_94;
   assign m53_94 =15'b0;

   // m53_95 = W*in
   wire signed [14:0] m53_95;
   assign m53_95 =15'b0;

   // m53_96 = W*in
   wire signed [14:0] m53_96;
   assign m53_96 =15'b0;

   // m53_97 = W*in
   wire signed [14:0] m53_97;
   assign m53_97 =15'b0;

   // m53_98 = W*in
   wire signed [14:0] m53_98;
   assign m53_98 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_99 = W*in
   wire signed [14:0] m53_99;
   assign m53_99 ={ {3{neg53[14]}} , neg53[14:3] };

   // m53_100 = W*in
   wire signed [14:0] m53_100;
   assign m53_100 =15'b0;

   // m54_1 = W*in
   wire signed [14:0] m54_1;
   assign m54_1 =15'b0;

   // m54_2 = W*in
   wire signed [14:0] m54_2;
   assign m54_2 =15'b0;

   // m54_3 = W*in
   wire signed [14:0] m54_3;
   assign m54_3 =15'b0;

   // m54_4 = W*in
   wire signed [14:0] m54_4;
   assign m54_4 =15'b0;

   // m54_5 = W*in
   wire signed [14:0] m54_5;
   assign m54_5 =15'b0;

   // m54_6 = W*in
   wire signed [14:0] m54_6;
   assign m54_6 =15'b0;

   // m54_7 = W*in
   wire signed [14:0] m54_7;
   assign m54_7 =15'b0;

   // m54_8 = W*in
   wire signed [14:0] m54_8;
   assign m54_8 =15'b0;

   // m54_9 = W*in
   wire signed [14:0] m54_9;
   assign m54_9 =15'b0;

   // m54_10 = W*in
   wire signed [14:0] m54_10;
   assign m54_10 =15'b0;

   // m54_11 = W*in
   wire signed [14:0] m54_11;
   assign m54_11 =15'b0;

   // m54_12 = W*in
   wire signed [14:0] m54_12;
   assign m54_12 =15'b0;

   // m54_13 = W*in
   wire signed [14:0] m54_13;
   assign m54_13 =15'b0;

   // m54_14 = W*in
   wire signed [14:0] m54_14;
   assign m54_14 =15'b0;

   // m54_15 = W*in
   wire signed [14:0] m54_15;
   assign m54_15 =15'b0;

   // m54_16 = W*in
   wire signed [14:0] m54_16;
   assign m54_16 =15'b0;

   // m54_17 = W*in
   wire signed [14:0] m54_17;
   assign m54_17 =15'b0;

   // m54_18 = W*in
   wire signed [14:0] m54_18;
   assign m54_18 =15'b0;

   // m54_19 = W*in
   wire signed [14:0] m54_19;
   assign m54_19 =15'b0;

   // m54_20 = W*in
   wire signed [14:0] m54_20;
   assign m54_20 =15'b0;

   // m54_21 = W*in
   wire signed [14:0] m54_21;
   assign m54_21 =15'b0;

   // m54_22 = W*in
   wire signed [14:0] m54_22;
   assign m54_22 =15'b0;

   // m54_23 = W*in
   wire signed [14:0] m54_23;
   assign m54_23 =15'b0;

   // m54_24 = W*in
   wire signed [14:0] m54_24;
   assign m54_24 =15'b0;

   // m54_25 = W*in
   wire signed [14:0] m54_25;
   assign m54_25 =15'b0;

   // m54_26 = W*in
   wire signed [14:0] m54_26;
   assign m54_26 =15'b0;

   // m54_27 = W*in
   wire signed [14:0] m54_27;
   assign m54_27 =15'b0;

   // m54_28 = W*in
   wire signed [14:0] m54_28;
   assign m54_28 =15'b0;

   // m54_29 = W*in
   wire signed [14:0] m54_29;
   assign m54_29 =15'b0;

   // m54_30 = W*in
   wire signed [14:0] m54_30;
   assign m54_30 =15'b0;

   // m54_31 = W*in
   wire signed [14:0] m54_31;
   assign m54_31 =15'b0;

   // m54_32 = W*in
   wire signed [14:0] m54_32;
   assign m54_32 =15'b0;

   // m54_33 = W*in
   wire signed [14:0] m54_33;
   assign m54_33 =15'b0;

   // m54_34 = W*in
   wire signed [14:0] m54_34;
   assign m54_34 =15'b0;

   // m54_35 = W*in
   wire signed [14:0] m54_35;
   assign m54_35 =15'b0;

   // m54_36 = W*in
   wire signed [14:0] m54_36;
   assign m54_36 =15'b0;

   // m54_37 = W*in
   wire signed [14:0] m54_37;
   assign m54_37 =15'b0;

   // m54_38 = W*in
   wire signed [14:0] m54_38;
   assign m54_38 =15'b0;

   // m54_39 = W*in
   wire signed [14:0] m54_39;
   assign m54_39 =15'b0;

   // m54_40 = W*in
   wire signed [14:0] m54_40;
   assign m54_40 =15'b0;

   // m54_41 = W*in
   wire signed [14:0] m54_41;
   assign m54_41 =15'b0;

   // m54_42 = W*in
   wire signed [14:0] m54_42;
   assign m54_42 =15'b0;

   // m54_43 = W*in
   wire signed [14:0] m54_43;
   assign m54_43 =15'b0;

   // m54_44 = W*in
   wire signed [14:0] m54_44;
   assign m54_44 =15'b0;

   // m54_45 = W*in
   wire signed [14:0] m54_45;
   assign m54_45 =15'b0;

   // m54_46 = W*in
   wire signed [14:0] m54_46;
   assign m54_46 =15'b0;

   // m54_47 = W*in
   wire signed [14:0] m54_47;
   assign m54_47 ={ {4{in54[14]}} , in54[14:4] };

   // m54_48 = W*in
   wire signed [14:0] m54_48;
   assign m54_48 =15'b0;

   // m54_49 = W*in
   wire signed [14:0] m54_49;
   assign m54_49 =15'b0;

   // m54_50 = W*in
   wire signed [14:0] m54_50;
   assign m54_50 =15'b0;

   // m54_51 = W*in
   wire signed [14:0] m54_51;
   assign m54_51 =15'b0;

   // m54_52 = W*in
   wire signed [14:0] m54_52;
   assign m54_52 =15'b0;

   // m54_53 = W*in
   wire signed [14:0] m54_53;
   assign m54_53 =15'b0;

   // m54_54 = W*in
   wire signed [14:0] m54_54;
   assign m54_54 =15'b0;

   // m54_55 = W*in
   wire signed [14:0] m54_55;
   assign m54_55 =15'b0;

   // m54_56 = W*in
   wire signed [14:0] m54_56;
   assign m54_56 =15'b0;

   // m54_57 = W*in
   wire signed [14:0] m54_57;
   assign m54_57 =15'b0;

   // m54_58 = W*in
   wire signed [14:0] m54_58;
   assign m54_58 =15'b0;

   // m54_59 = W*in
   wire signed [14:0] m54_59;
   assign m54_59 =15'b0;

   // m54_60 = W*in
   wire signed [14:0] m54_60;
   assign m54_60 =15'b0;

   // m54_61 = W*in
   wire signed [14:0] m54_61;
   assign m54_61 =15'b0;

   // m54_62 = W*in
   wire signed [14:0] m54_62;
   assign m54_62 =15'b0;

   // m54_63 = W*in
   wire signed [14:0] m54_63;
   assign m54_63 =15'b0;

   // m54_64 = W*in
   wire signed [14:0] m54_64;
   assign m54_64 =15'b0;

   // m54_65 = W*in
   wire signed [14:0] m54_65;
   assign m54_65 =15'b0;

   // m54_66 = W*in
   wire signed [14:0] m54_66;
   assign m54_66 =15'b0;

   // m54_67 = W*in
   wire signed [14:0] m54_67;
   assign m54_67 =15'b0;

   // m54_68 = W*in
   wire signed [14:0] m54_68;
   assign m54_68 ={ {4{neg54[14]}} , neg54[14:4] };

   // m54_69 = W*in
   wire signed [14:0] m54_69;
   assign m54_69 =15'b0;

   // m54_70 = W*in
   wire signed [14:0] m54_70;
   assign m54_70 =15'b0;

   // m54_71 = W*in
   wire signed [14:0] m54_71;
   assign m54_71 =15'b0;

   // m54_72 = W*in
   wire signed [14:0] m54_72;
   assign m54_72 =15'b0;

   // m54_73 = W*in
   wire signed [14:0] m54_73;
   assign m54_73 =15'b0;

   // m54_74 = W*in
   wire signed [14:0] m54_74;
   assign m54_74 =15'b0;

   // m54_75 = W*in
   wire signed [14:0] m54_75;
   assign m54_75 =15'b0;

   // m54_76 = W*in
   wire signed [14:0] m54_76;
   assign m54_76 =15'b0;

   // m54_77 = W*in
   wire signed [14:0] m54_77;
   assign m54_77 =15'b0;

   // m54_78 = W*in
   wire signed [14:0] m54_78;
   assign m54_78 =15'b0;

   // m54_79 = W*in
   wire signed [14:0] m54_79;
   assign m54_79 =15'b0;

   // m54_80 = W*in
   wire signed [14:0] m54_80;
   assign m54_80 =15'b0;

   // m54_81 = W*in
   wire signed [14:0] m54_81;
   assign m54_81 =15'b0;

   // m54_82 = W*in
   wire signed [14:0] m54_82;
   assign m54_82 =15'b0;

   // m54_83 = W*in
   wire signed [14:0] m54_83;
   assign m54_83 =15'b0;

   // m54_84 = W*in
   wire signed [14:0] m54_84;
   assign m54_84 =15'b0;

   // m54_85 = W*in
   wire signed [14:0] m54_85;
   assign m54_85 =15'b0;

   // m54_86 = W*in
   wire signed [14:0] m54_86;
   assign m54_86 =15'b0;

   // m54_87 = W*in
   wire signed [14:0] m54_87;
   assign m54_87 =15'b0;

   // m54_88 = W*in
   wire signed [14:0] m54_88;
   assign m54_88 =15'b0;

   // m54_89 = W*in
   wire signed [14:0] m54_89;
   assign m54_89 =15'b0;

   // m54_90 = W*in
   wire signed [14:0] m54_90;
   assign m54_90 =15'b0;

   // m54_91 = W*in
   wire signed [14:0] m54_91;
   assign m54_91 =15'b0;

   // m54_92 = W*in
   wire signed [14:0] m54_92;
   assign m54_92 =15'b0;

   // m54_93 = W*in
   wire signed [14:0] m54_93;
   assign m54_93 =15'b0;

   // m54_94 = W*in
   wire signed [14:0] m54_94;
   assign m54_94 =15'b0;

   // m54_95 = W*in
   wire signed [14:0] m54_95;
   assign m54_95 =15'b0;

   // m54_96 = W*in
   wire signed [14:0] m54_96;
   assign m54_96 =15'b0;

   // m54_97 = W*in
   wire signed [14:0] m54_97;
   assign m54_97 =15'b0;

   // m54_98 = W*in
   wire signed [14:0] m54_98;
   assign m54_98 =15'b0;

   // m54_99 = W*in
   wire signed [14:0] m54_99;
   assign m54_99 =15'b0;

   // m54_100 = W*in
   wire signed [14:0] m54_100;
   assign m54_100 =15'b0;

   // m55_1 = W*in
   wire signed [14:0] m55_1;
   assign m55_1 ={ {3{in55[14]}} , in55[14:3] };

   // m55_2 = W*in
   wire signed [14:0] m55_2;
   assign m55_2 =15'b0;

   // m55_3 = W*in
   wire signed [14:0] m55_3;
   assign m55_3 =15'b0;

   // m55_4 = W*in
   wire signed [14:0] m55_4;
   assign m55_4 =15'b0;

   // m55_5 = W*in
   wire signed [14:0] m55_5;
   assign m55_5 =15'b0;

   // m55_6 = W*in
   wire signed [14:0] m55_6;
   assign m55_6 =15'b0;

   // m55_7 = W*in
   wire signed [14:0] m55_7;
   assign m55_7 =15'b0;

   // m55_8 = W*in
   wire signed [14:0] m55_8;
   assign m55_8 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_9 = W*in
   wire signed [14:0] m55_9;
   assign m55_9 =15'b0;

   // m55_10 = W*in
   wire signed [14:0] m55_10;
   assign m55_10 =15'b0;

   // m55_11 = W*in
   wire signed [14:0] m55_11;
   assign m55_11 =15'b0;

   // m55_12 = W*in
   wire signed [14:0] m55_12;
   assign m55_12 ={ {3{in55[14]}} , in55[14:3] };

   // m55_13 = W*in
   wire signed [14:0] m55_13;
   assign m55_13 =15'b0;

   // m55_14 = W*in
   wire signed [14:0] m55_14;
   assign m55_14 =15'b0;

   // m55_15 = W*in
   wire signed [14:0] m55_15;
   assign m55_15 =15'b0;

   // m55_16 = W*in
   wire signed [14:0] m55_16;
   assign m55_16 =15'b0;

   // m55_17 = W*in
   wire signed [14:0] m55_17;
   assign m55_17 =15'b0;

   // m55_18 = W*in
   wire signed [14:0] m55_18;
   assign m55_18 =15'b0;

   // m55_19 = W*in
   wire signed [14:0] m55_19;
   assign m55_19 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_20 = W*in
   wire signed [14:0] m55_20;
   assign m55_20 ={ {4{neg55[14]}} , neg55[14:4] };

   // m55_21 = W*in
   wire signed [14:0] m55_21;
   assign m55_21 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_22 = W*in
   wire signed [14:0] m55_22;
   assign m55_22 ={ {3{in55[14]}} , in55[14:3] };

   // m55_23 = W*in
   wire signed [14:0] m55_23;
   assign m55_23 =15'b0;

   // m55_24 = W*in
   wire signed [14:0] m55_24;
   assign m55_24 ={ {3{in55[14]}} , in55[14:3] };

   // m55_25 = W*in
   wire signed [14:0] m55_25;
   assign m55_25 =15'b0;

   // m55_26 = W*in
   wire signed [14:0] m55_26;
   assign m55_26 ={ {3{in55[14]}} , in55[14:3] };

   // m55_27 = W*in
   wire signed [14:0] m55_27;
   assign m55_27 ={ {3{in55[14]}} , in55[14:3] };

   // m55_28 = W*in
   wire signed [14:0] m55_28;
   assign m55_28 =15'b0;

   // m55_29 = W*in
   wire signed [14:0] m55_29;
   assign m55_29 =15'b0;

   // m55_30 = W*in
   wire signed [14:0] m55_30;
   assign m55_30 ={ {3{in55[14]}} , in55[14:3] };

   // m55_31 = W*in
   wire signed [14:0] m55_31;
   assign m55_31 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_32 = W*in
   wire signed [14:0] m55_32;
   assign m55_32 =15'b0;

   // m55_33 = W*in
   wire signed [14:0] m55_33;
   assign m55_33 =15'b0;

   // m55_34 = W*in
   wire signed [14:0] m55_34;
   assign m55_34 =15'b0;

   // m55_35 = W*in
   wire signed [14:0] m55_35;
   assign m55_35 =15'b0;

   // m55_36 = W*in
   wire signed [14:0] m55_36;
   assign m55_36 =15'b0;

   // m55_37 = W*in
   wire signed [14:0] m55_37;
   assign m55_37 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_38 = W*in
   wire signed [14:0] m55_38;
   assign m55_38 ={ {4{in55[14]}} , in55[14:4] };

   // m55_39 = W*in
   wire signed [14:0] m55_39;
   assign m55_39 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_40 = W*in
   wire signed [14:0] m55_40;
   assign m55_40 =15'b0;

   // m55_41 = W*in
   wire signed [14:0] m55_41;
   assign m55_41 ={ {3{in55[14]}} , in55[14:3] };

   // m55_42 = W*in
   wire signed [14:0] m55_42;
   assign m55_42 ={ {3{in55[14]}} , in55[14:3] };

   // m55_43 = W*in
   wire signed [14:0] m55_43;
   assign m55_43 =15'b0;

   // m55_44 = W*in
   wire signed [14:0] m55_44;
   assign m55_44 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_45 = W*in
   wire signed [14:0] m55_45;
   assign m55_45 =15'b0;

   // m55_46 = W*in
   wire signed [14:0] m55_46;
   assign m55_46 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_47 = W*in
   wire signed [14:0] m55_47;
   assign m55_47 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_48 = W*in
   wire signed [14:0] m55_48;
   assign m55_48 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_49 = W*in
   wire signed [14:0] m55_49;
   assign m55_49 =15'b0;

   // m55_50 = W*in
   wire signed [14:0] m55_50;
   assign m55_50 =15'b0;

   // m55_51 = W*in
   wire signed [14:0] m55_51;
   assign m55_51 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_52 = W*in
   wire signed [14:0] m55_52;
   assign m55_52 =15'b0;

   // m55_53 = W*in
   wire signed [14:0] m55_53;
   assign m55_53 =15'b0;

   // m55_54 = W*in
   wire signed [14:0] m55_54;
   assign m55_54 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_55 = W*in
   wire signed [14:0] m55_55;
   assign m55_55 =15'b0;

   // m55_56 = W*in
   wire signed [14:0] m55_56;
   assign m55_56 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_57 = W*in
   wire signed [14:0] m55_57;
   assign m55_57 =15'b0;

   // m55_58 = W*in
   wire signed [14:0] m55_58;
   assign m55_58 =15'b0;

   // m55_59 = W*in
   wire signed [14:0] m55_59;
   assign m55_59 =15'b0;

   // m55_60 = W*in
   wire signed [14:0] m55_60;
   assign m55_60 =15'b0;

   // m55_61 = W*in
   wire signed [14:0] m55_61;
   assign m55_61 =15'b0;

   // m55_62 = W*in
   wire signed [14:0] m55_62;
   assign m55_62 ={ {3{in55[14]}} , in55[14:3] };

   // m55_63 = W*in
   wire signed [14:0] m55_63;
   assign m55_63 =15'b0;

   // m55_64 = W*in
   wire signed [14:0] m55_64;
   assign m55_64 =15'b0;

   // m55_65 = W*in
   wire signed [14:0] m55_65;
   assign m55_65 =15'b0;

   // m55_66 = W*in
   wire signed [14:0] m55_66;
   assign m55_66 =15'b0;

   // m55_67 = W*in
   wire signed [14:0] m55_67;
   assign m55_67 =15'b0;

   // m55_68 = W*in
   wire signed [14:0] m55_68;
   assign m55_68 =15'b0;

   // m55_69 = W*in
   wire signed [14:0] m55_69;
   assign m55_69 =15'b0;

   // m55_70 = W*in
   wire signed [14:0] m55_70;
   assign m55_70 =15'b0;

   // m55_71 = W*in
   wire signed [14:0] m55_71;
   assign m55_71 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_72 = W*in
   wire signed [14:0] m55_72;
   assign m55_72 =15'b0;

   // m55_73 = W*in
   wire signed [14:0] m55_73;
   assign m55_73 =15'b0;

   // m55_74 = W*in
   wire signed [14:0] m55_74;
   assign m55_74 ={ {4{neg55[14]}} , neg55[14:4] };

   // m55_75 = W*in
   wire signed [14:0] m55_75;
   assign m55_75 =15'b0;

   // m55_76 = W*in
   wire signed [14:0] m55_76;
   assign m55_76 =15'b0;

   // m55_77 = W*in
   wire signed [14:0] m55_77;
   assign m55_77 =15'b0;

   // m55_78 = W*in
   wire signed [14:0] m55_78;
   assign m55_78 =15'b0;

   // m55_79 = W*in
   wire signed [14:0] m55_79;
   assign m55_79 =15'b0;

   // m55_80 = W*in
   wire signed [14:0] m55_80;
   assign m55_80 =15'b0;

   // m55_81 = W*in
   wire signed [14:0] m55_81;
   assign m55_81 ={ {2{in55[14]}} , in55[14:2] };

   // m55_82 = W*in
   wire signed [14:0] m55_82;
   assign m55_82 ={ {3{in55[14]}} , in55[14:3] };

   // m55_83 = W*in
   wire signed [14:0] m55_83;
   assign m55_83 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_84 = W*in
   wire signed [14:0] m55_84;
   assign m55_84 ={ {3{in55[14]}} , in55[14:3] };

   // m55_85 = W*in
   wire signed [14:0] m55_85;
   assign m55_85 =15'b0;

   // m55_86 = W*in
   wire signed [14:0] m55_86;
   assign m55_86 =15'b0;

   // m55_87 = W*in
   wire signed [14:0] m55_87;
   assign m55_87 =15'b0;

   // m55_88 = W*in
   wire signed [14:0] m55_88;
   assign m55_88 ={ {3{in55[14]}} , in55[14:3] };

   // m55_89 = W*in
   wire signed [14:0] m55_89;
   assign m55_89 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_90 = W*in
   wire signed [14:0] m55_90;
   assign m55_90 =15'b0;

   // m55_91 = W*in
   wire signed [14:0] m55_91;
   assign m55_91 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_92 = W*in
   wire signed [14:0] m55_92;
   assign m55_92 =15'b0;

   // m55_93 = W*in
   wire signed [14:0] m55_93;
   assign m55_93 =15'b0;

   // m55_94 = W*in
   wire signed [14:0] m55_94;
   assign m55_94 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_95 = W*in
   wire signed [14:0] m55_95;
   assign m55_95 =15'b0;

   // m55_96 = W*in
   wire signed [14:0] m55_96;
   assign m55_96 =15'b0;

   // m55_97 = W*in
   wire signed [14:0] m55_97;
   assign m55_97 =15'b0;

   // m55_98 = W*in
   wire signed [14:0] m55_98;
   assign m55_98 ={ {3{neg55[14]}} , neg55[14:3] };

   // m55_99 = W*in
   wire signed [14:0] m55_99;
   assign m55_99 =15'b0;

   // m55_100 = W*in
   wire signed [14:0] m55_100;
   assign m55_100 =15'b0;

   // m56_1 = W*in
   wire signed [14:0] m56_1;
   assign m56_1 =15'b0;

   // m56_2 = W*in
   wire signed [14:0] m56_2;
   assign m56_2 =15'b0;

   // m56_3 = W*in
   wire signed [14:0] m56_3;
   assign m56_3 =15'b0;

   // m56_4 = W*in
   wire signed [14:0] m56_4;
   assign m56_4 =15'b0;

   // m56_5 = W*in
   wire signed [14:0] m56_5;
   assign m56_5 =15'b0;

   // m56_6 = W*in
   wire signed [14:0] m56_6;
   assign m56_6 =15'b0;

   // m56_7 = W*in
   wire signed [14:0] m56_7;
   assign m56_7 =15'b0;

   // m56_8 = W*in
   wire signed [14:0] m56_8;
   assign m56_8 =15'b0;

   // m56_9 = W*in
   wire signed [14:0] m56_9;
   assign m56_9 =15'b0;

   // m56_10 = W*in
   wire signed [14:0] m56_10;
   assign m56_10 =15'b0;

   // m56_11 = W*in
   wire signed [14:0] m56_11;
   assign m56_11 =15'b0;

   // m56_12 = W*in
   wire signed [14:0] m56_12;
   assign m56_12 =15'b0;

   // m56_13 = W*in
   wire signed [14:0] m56_13;
   assign m56_13 =15'b0;

   // m56_14 = W*in
   wire signed [14:0] m56_14;
   assign m56_14 =15'b0;

   // m56_15 = W*in
   wire signed [14:0] m56_15;
   assign m56_15 =15'b0;

   // m56_16 = W*in
   wire signed [14:0] m56_16;
   assign m56_16 ={ {3{in56[14]}} , in56[14:3] };

   // m56_17 = W*in
   wire signed [14:0] m56_17;
   assign m56_17 =15'b0;

   // m56_18 = W*in
   wire signed [14:0] m56_18;
   assign m56_18 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_19 = W*in
   wire signed [14:0] m56_19;
   assign m56_19 =15'b0;

   // m56_20 = W*in
   wire signed [14:0] m56_20;
   assign m56_20 ={ {4{neg56[14]}} , neg56[14:4] };

   // m56_21 = W*in
   wire signed [14:0] m56_21;
   assign m56_21 =15'b0;

   // m56_22 = W*in
   wire signed [14:0] m56_22;
   assign m56_22 ={ {4{neg56[14]}} , neg56[14:4] };

   // m56_23 = W*in
   wire signed [14:0] m56_23;
   assign m56_23 =15'b0;

   // m56_24 = W*in
   wire signed [14:0] m56_24;
   assign m56_24 =15'b0;

   // m56_25 = W*in
   wire signed [14:0] m56_25;
   assign m56_25 ={ {3{in56[14]}} , in56[14:3] };

   // m56_26 = W*in
   wire signed [14:0] m56_26;
   assign m56_26 =15'b0;

   // m56_27 = W*in
   wire signed [14:0] m56_27;
   assign m56_27 =15'b0;

   // m56_28 = W*in
   wire signed [14:0] m56_28;
   assign m56_28 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_29 = W*in
   wire signed [14:0] m56_29;
   assign m56_29 =15'b0;

   // m56_30 = W*in
   wire signed [14:0] m56_30;
   assign m56_30 ={ {4{in56[14]}} , in56[14:4] };

   // m56_31 = W*in
   wire signed [14:0] m56_31;
   assign m56_31 =15'b0;

   // m56_32 = W*in
   wire signed [14:0] m56_32;
   assign m56_32 =15'b0;

   // m56_33 = W*in
   wire signed [14:0] m56_33;
   assign m56_33 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_34 = W*in
   wire signed [14:0] m56_34;
   assign m56_34 =15'b0;

   // m56_35 = W*in
   wire signed [14:0] m56_35;
   assign m56_35 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_36 = W*in
   wire signed [14:0] m56_36;
   assign m56_36 =15'b0;

   // m56_37 = W*in
   wire signed [14:0] m56_37;
   assign m56_37 =15'b0;

   // m56_38 = W*in
   wire signed [14:0] m56_38;
   assign m56_38 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_39 = W*in
   wire signed [14:0] m56_39;
   assign m56_39 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_40 = W*in
   wire signed [14:0] m56_40;
   assign m56_40 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_41 = W*in
   wire signed [14:0] m56_41;
   assign m56_41 =15'b0;

   // m56_42 = W*in
   wire signed [14:0] m56_42;
   assign m56_42 =15'b0;

   // m56_43 = W*in
   wire signed [14:0] m56_43;
   assign m56_43 ={ {3{in56[14]}} , in56[14:3] };

   // m56_44 = W*in
   wire signed [14:0] m56_44;
   assign m56_44 =15'b0;

   // m56_45 = W*in
   wire signed [14:0] m56_45;
   assign m56_45 =15'b0;

   // m56_46 = W*in
   wire signed [14:0] m56_46;
   assign m56_46 =15'b0;

   // m56_47 = W*in
   wire signed [14:0] m56_47;
   assign m56_47 ={ {4{in56[14]}} , in56[14:4] };

   // m56_48 = W*in
   wire signed [14:0] m56_48;
   assign m56_48 =15'b0;

   // m56_49 = W*in
   wire signed [14:0] m56_49;
   assign m56_49 ={ {3{in56[14]}} , in56[14:3] };

   // m56_50 = W*in
   wire signed [14:0] m56_50;
   assign m56_50 =15'b0;

   // m56_51 = W*in
   wire signed [14:0] m56_51;
   assign m56_51 =15'b0;

   // m56_52 = W*in
   wire signed [14:0] m56_52;
   assign m56_52 =15'b0;

   // m56_53 = W*in
   wire signed [14:0] m56_53;
   assign m56_53 =15'b0;

   // m56_54 = W*in
   wire signed [14:0] m56_54;
   assign m56_54 =15'b0;

   // m56_55 = W*in
   wire signed [14:0] m56_55;
   assign m56_55 =15'b0;

   // m56_56 = W*in
   wire signed [14:0] m56_56;
   assign m56_56 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_57 = W*in
   wire signed [14:0] m56_57;
   assign m56_57 =15'b0;

   // m56_58 = W*in
   wire signed [14:0] m56_58;
   assign m56_58 ={ {4{in56[14]}} , in56[14:4] };

   // m56_59 = W*in
   wire signed [14:0] m56_59;
   assign m56_59 =15'b0;

   // m56_60 = W*in
   wire signed [14:0] m56_60;
   assign m56_60 =15'b0;

   // m56_61 = W*in
   wire signed [14:0] m56_61;
   assign m56_61 =15'b0;

   // m56_62 = W*in
   wire signed [14:0] m56_62;
   assign m56_62 =15'b0;

   // m56_63 = W*in
   wire signed [14:0] m56_63;
   assign m56_63 =15'b0;

   // m56_64 = W*in
   wire signed [14:0] m56_64;
   assign m56_64 =15'b0;

   // m56_65 = W*in
   wire signed [14:0] m56_65;
   assign m56_65 ={ {2{in56[14]}} , in56[14:2] };

   // m56_66 = W*in
   wire signed [14:0] m56_66;
   assign m56_66 ={ {4{neg56[14]}} , neg56[14:4] };

   // m56_67 = W*in
   wire signed [14:0] m56_67;
   assign m56_67 ={ {4{in56[14]}} , in56[14:4] };

   // m56_68 = W*in
   wire signed [14:0] m56_68;
   assign m56_68 =15'b0;

   // m56_69 = W*in
   wire signed [14:0] m56_69;
   assign m56_69 ={ {2{in56[14]}} , in56[14:2] };

   // m56_70 = W*in
   wire signed [14:0] m56_70;
   assign m56_70 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_71 = W*in
   wire signed [14:0] m56_71;
   assign m56_71 =15'b0;

   // m56_72 = W*in
   wire signed [14:0] m56_72;
   assign m56_72 =15'b0;

   // m56_73 = W*in
   wire signed [14:0] m56_73;
   assign m56_73 =15'b0;

   // m56_74 = W*in
   wire signed [14:0] m56_74;
   assign m56_74 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_75 = W*in
   wire signed [14:0] m56_75;
   assign m56_75 =15'b0;

   // m56_76 = W*in
   wire signed [14:0] m56_76;
   assign m56_76 =15'b0;

   // m56_77 = W*in
   wire signed [14:0] m56_77;
   assign m56_77 ={ {3{in56[14]}} , in56[14:3] };

   // m56_78 = W*in
   wire signed [14:0] m56_78;
   assign m56_78 =15'b0;

   // m56_79 = W*in
   wire signed [14:0] m56_79;
   assign m56_79 =15'b0;

   // m56_80 = W*in
   wire signed [14:0] m56_80;
   assign m56_80 =15'b0;

   // m56_81 = W*in
   wire signed [14:0] m56_81;
   assign m56_81 =15'b0;

   // m56_82 = W*in
   wire signed [14:0] m56_82;
   assign m56_82 =15'b0;

   // m56_83 = W*in
   wire signed [14:0] m56_83;
   assign m56_83 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_84 = W*in
   wire signed [14:0] m56_84;
   assign m56_84 =15'b0;

   // m56_85 = W*in
   wire signed [14:0] m56_85;
   assign m56_85 =15'b0;

   // m56_86 = W*in
   wire signed [14:0] m56_86;
   assign m56_86 =15'b0;

   // m56_87 = W*in
   wire signed [14:0] m56_87;
   assign m56_87 =15'b0;

   // m56_88 = W*in
   wire signed [14:0] m56_88;
   assign m56_88 =15'b0;

   // m56_89 = W*in
   wire signed [14:0] m56_89;
   assign m56_89 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_90 = W*in
   wire signed [14:0] m56_90;
   assign m56_90 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_91 = W*in
   wire signed [14:0] m56_91;
   assign m56_91 =15'b0;

   // m56_92 = W*in
   wire signed [14:0] m56_92;
   assign m56_92 =15'b0;

   // m56_93 = W*in
   wire signed [14:0] m56_93;
   assign m56_93 =15'b0;

   // m56_94 = W*in
   wire signed [14:0] m56_94;
   assign m56_94 ={ {3{neg56[14]}} , neg56[14:3] };

   // m56_95 = W*in
   wire signed [14:0] m56_95;
   assign m56_95 =15'b0;

   // m56_96 = W*in
   wire signed [14:0] m56_96;
   assign m56_96 =15'b0;

   // m56_97 = W*in
   wire signed [14:0] m56_97;
   assign m56_97 =15'b0;

   // m56_98 = W*in
   wire signed [14:0] m56_98;
   assign m56_98 =15'b0;

   // m56_99 = W*in
   wire signed [14:0] m56_99;
   assign m56_99 =15'b0;

   // m56_100 = W*in
   wire signed [14:0] m56_100;
   assign m56_100 =15'b0;

   // m57_1 = W*in
   wire signed [14:0] m57_1;
   assign m57_1 ={ {3{in57[14]}} , in57[14:3] };

   // m57_2 = W*in
   wire signed [14:0] m57_2;
   assign m57_2 =15'b0;

   // m57_3 = W*in
   wire signed [14:0] m57_3;
   assign m57_3 =15'b0;

   // m57_4 = W*in
   wire signed [14:0] m57_4;
   assign m57_4 =15'b0;

   // m57_5 = W*in
   wire signed [14:0] m57_5;
   assign m57_5 =15'b0;

   // m57_6 = W*in
   wire signed [14:0] m57_6;
   assign m57_6 ={ {3{neg57[14]}} , neg57[14:3] };

   // m57_7 = W*in
   wire signed [14:0] m57_7;
   assign m57_7 =15'b0;

   // m57_8 = W*in
   wire signed [14:0] m57_8;
   assign m57_8 =15'b0;

   // m57_9 = W*in
   wire signed [14:0] m57_9;
   assign m57_9 =15'b0;

   // m57_10 = W*in
   wire signed [14:0] m57_10;
   assign m57_10 =15'b0;

   // m57_11 = W*in
   wire signed [14:0] m57_11;
   assign m57_11 =15'b0;

   // m57_12 = W*in
   wire signed [14:0] m57_12;
   assign m57_12 ={ {3{in57[14]}} , in57[14:3] };

   // m57_13 = W*in
   wire signed [14:0] m57_13;
   assign m57_13 =15'b0;

   // m57_14 = W*in
   wire signed [14:0] m57_14;
   assign m57_14 =15'b0;

   // m57_15 = W*in
   wire signed [14:0] m57_15;
   assign m57_15 =15'b0;

   // m57_16 = W*in
   wire signed [14:0] m57_16;
   assign m57_16 =15'b0;

   // m57_17 = W*in
   wire signed [14:0] m57_17;
   assign m57_17 =15'b0;

   // m57_18 = W*in
   wire signed [14:0] m57_18;
   assign m57_18 =15'b0;

   // m57_19 = W*in
   wire signed [14:0] m57_19;
   assign m57_19 =15'b0;

   // m57_20 = W*in
   wire signed [14:0] m57_20;
   assign m57_20 =15'b0;

   // m57_21 = W*in
   wire signed [14:0] m57_21;
   assign m57_21 =15'b0;

   // m57_22 = W*in
   wire signed [14:0] m57_22;
   assign m57_22 =15'b0;

   // m57_23 = W*in
   wire signed [14:0] m57_23;
   assign m57_23 =15'b0;

   // m57_24 = W*in
   wire signed [14:0] m57_24;
   assign m57_24 =15'b0;

   // m57_25 = W*in
   wire signed [14:0] m57_25;
   assign m57_25 =15'b0;

   // m57_26 = W*in
   wire signed [14:0] m57_26;
   assign m57_26 =15'b0;

   // m57_27 = W*in
   wire signed [14:0] m57_27;
   assign m57_27 ={ {3{neg57[14]}} , neg57[14:3] };

   // m57_28 = W*in
   wire signed [14:0] m57_28;
   assign m57_28 =15'b0;

   // m57_29 = W*in
   wire signed [14:0] m57_29;
   assign m57_29 =15'b0;

   // m57_30 = W*in
   wire signed [14:0] m57_30;
   assign m57_30 =15'b0;

   // m57_31 = W*in
   wire signed [14:0] m57_31;
   assign m57_31 =15'b0;

   // m57_32 = W*in
   wire signed [14:0] m57_32;
   assign m57_32 =15'b0;

   // m57_33 = W*in
   wire signed [14:0] m57_33;
   assign m57_33 =15'b0;

   // m57_34 = W*in
   wire signed [14:0] m57_34;
   assign m57_34 =15'b0;

   // m57_35 = W*in
   wire signed [14:0] m57_35;
   assign m57_35 =15'b0;

   // m57_36 = W*in
   wire signed [14:0] m57_36;
   assign m57_36 =15'b0;

   // m57_37 = W*in
   wire signed [14:0] m57_37;
   assign m57_37 =15'b0;

   // m57_38 = W*in
   wire signed [14:0] m57_38;
   assign m57_38 =15'b0;

   // m57_39 = W*in
   wire signed [14:0] m57_39;
   assign m57_39 =15'b0;

   // m57_40 = W*in
   wire signed [14:0] m57_40;
   assign m57_40 ={ {3{in57[14]}} , in57[14:3] };

   // m57_41 = W*in
   wire signed [14:0] m57_41;
   assign m57_41 =15'b0;

   // m57_42 = W*in
   wire signed [14:0] m57_42;
   assign m57_42 =15'b0;

   // m57_43 = W*in
   wire signed [14:0] m57_43;
   assign m57_43 =15'b0;

   // m57_44 = W*in
   wire signed [14:0] m57_44;
   assign m57_44 =15'b0;

   // m57_45 = W*in
   wire signed [14:0] m57_45;
   assign m57_45 =15'b0;

   // m57_46 = W*in
   wire signed [14:0] m57_46;
   assign m57_46 ={ {3{neg57[14]}} , neg57[14:3] };

   // m57_47 = W*in
   wire signed [14:0] m57_47;
   assign m57_47 =15'b0;

   // m57_48 = W*in
   wire signed [14:0] m57_48;
   assign m57_48 ={ {3{neg57[14]}} , neg57[14:3] };

   // m57_49 = W*in
   wire signed [14:0] m57_49;
   assign m57_49 =15'b0;

   // m57_50 = W*in
   wire signed [14:0] m57_50;
   assign m57_50 =15'b0;

   // m57_51 = W*in
   wire signed [14:0] m57_51;
   assign m57_51 =15'b0;

   // m57_52 = W*in
   wire signed [14:0] m57_52;
   assign m57_52 =15'b0;

   // m57_53 = W*in
   wire signed [14:0] m57_53;
   assign m57_53 =15'b0;

   // m57_54 = W*in
   wire signed [14:0] m57_54;
   assign m57_54 =15'b0;

   // m57_55 = W*in
   wire signed [14:0] m57_55;
   assign m57_55 =15'b0;

   // m57_56 = W*in
   wire signed [14:0] m57_56;
   assign m57_56 =15'b0;

   // m57_57 = W*in
   wire signed [14:0] m57_57;
   assign m57_57 =15'b0;

   // m57_58 = W*in
   wire signed [14:0] m57_58;
   assign m57_58 ={ {4{neg57[14]}} , neg57[14:4] };

   // m57_59 = W*in
   wire signed [14:0] m57_59;
   assign m57_59 =15'b0;

   // m57_60 = W*in
   wire signed [14:0] m57_60;
   assign m57_60 =15'b0;

   // m57_61 = W*in
   wire signed [14:0] m57_61;
   assign m57_61 =15'b0;

   // m57_62 = W*in
   wire signed [14:0] m57_62;
   assign m57_62 =15'b0;

   // m57_63 = W*in
   wire signed [14:0] m57_63;
   assign m57_63 =15'b0;

   // m57_64 = W*in
   wire signed [14:0] m57_64;
   assign m57_64 ={ {3{in57[14]}} , in57[14:3] };

   // m57_65 = W*in
   wire signed [14:0] m57_65;
   assign m57_65 =15'b0;

   // m57_66 = W*in
   wire signed [14:0] m57_66;
   assign m57_66 =15'b0;

   // m57_67 = W*in
   wire signed [14:0] m57_67;
   assign m57_67 =15'b0;

   // m57_68 = W*in
   wire signed [14:0] m57_68;
   assign m57_68 ={ {4{in57[14]}} , in57[14:4] };

   // m57_69 = W*in
   wire signed [14:0] m57_69;
   assign m57_69 =15'b0;

   // m57_70 = W*in
   wire signed [14:0] m57_70;
   assign m57_70 =15'b0;

   // m57_71 = W*in
   wire signed [14:0] m57_71;
   assign m57_71 =15'b0;

   // m57_72 = W*in
   wire signed [14:0] m57_72;
   assign m57_72 =15'b0;

   // m57_73 = W*in
   wire signed [14:0] m57_73;
   assign m57_73 =15'b0;

   // m57_74 = W*in
   wire signed [14:0] m57_74;
   assign m57_74 ={ {4{in57[14]}} , in57[14:4] };

   // m57_75 = W*in
   wire signed [14:0] m57_75;
   assign m57_75 =15'b0;

   // m57_76 = W*in
   wire signed [14:0] m57_76;
   assign m57_76 =15'b0;

   // m57_77 = W*in
   wire signed [14:0] m57_77;
   assign m57_77 =15'b0;

   // m57_78 = W*in
   wire signed [14:0] m57_78;
   assign m57_78 =15'b0;

   // m57_79 = W*in
   wire signed [14:0] m57_79;
   assign m57_79 =15'b0;

   // m57_80 = W*in
   wire signed [14:0] m57_80;
   assign m57_80 =15'b0;

   // m57_81 = W*in
   wire signed [14:0] m57_81;
   assign m57_81 =15'b0;

   // m57_82 = W*in
   wire signed [14:0] m57_82;
   assign m57_82 =15'b0;

   // m57_83 = W*in
   wire signed [14:0] m57_83;
   assign m57_83 ={ {3{neg57[14]}} , neg57[14:3] };

   // m57_84 = W*in
   wire signed [14:0] m57_84;
   assign m57_84 =15'b0;

   // m57_85 = W*in
   wire signed [14:0] m57_85;
   assign m57_85 =15'b0;

   // m57_86 = W*in
   wire signed [14:0] m57_86;
   assign m57_86 =15'b0;

   // m57_87 = W*in
   wire signed [14:0] m57_87;
   assign m57_87 ={ {3{in57[14]}} , in57[14:3] };

   // m57_88 = W*in
   wire signed [14:0] m57_88;
   assign m57_88 =15'b0;

   // m57_89 = W*in
   wire signed [14:0] m57_89;
   assign m57_89 =15'b0;

   // m57_90 = W*in
   wire signed [14:0] m57_90;
   assign m57_90 =15'b0;

   // m57_91 = W*in
   wire signed [14:0] m57_91;
   assign m57_91 =15'b0;

   // m57_92 = W*in
   wire signed [14:0] m57_92;
   assign m57_92 =15'b0;

   // m57_93 = W*in
   wire signed [14:0] m57_93;
   assign m57_93 =15'b0;

   // m57_94 = W*in
   wire signed [14:0] m57_94;
   assign m57_94 =15'b0;

   // m57_95 = W*in
   wire signed [14:0] m57_95;
   assign m57_95 =15'b0;

   // m57_96 = W*in
   wire signed [14:0] m57_96;
   assign m57_96 =15'b0;

   // m57_97 = W*in
   wire signed [14:0] m57_97;
   assign m57_97 =15'b0;

   // m57_98 = W*in
   wire signed [14:0] m57_98;
   assign m57_98 =15'b0;

   // m57_99 = W*in
   wire signed [14:0] m57_99;
   assign m57_99 =15'b0;

   // m57_100 = W*in
   wire signed [14:0] m57_100;
   assign m57_100 =15'b0;

   // m58_1 = W*in
   wire signed [14:0] m58_1;
   assign m58_1 =15'b0;

   // m58_2 = W*in
   wire signed [14:0] m58_2;
   assign m58_2 =15'b0;

   // m58_3 = W*in
   wire signed [14:0] m58_3;
   assign m58_3 =15'b0;

   // m58_4 = W*in
   wire signed [14:0] m58_4;
   assign m58_4 =15'b0;

   // m58_5 = W*in
   wire signed [14:0] m58_5;
   assign m58_5 =15'b0;

   // m58_6 = W*in
   wire signed [14:0] m58_6;
   assign m58_6 =15'b0;

   // m58_7 = W*in
   wire signed [14:0] m58_7;
   assign m58_7 =15'b0;

   // m58_8 = W*in
   wire signed [14:0] m58_8;
   assign m58_8 =15'b0;

   // m58_9 = W*in
   wire signed [14:0] m58_9;
   assign m58_9 =15'b0;

   // m58_10 = W*in
   wire signed [14:0] m58_10;
   assign m58_10 =15'b0;

   // m58_11 = W*in
   wire signed [14:0] m58_11;
   assign m58_11 =15'b0;

   // m58_12 = W*in
   wire signed [14:0] m58_12;
   assign m58_12 =15'b0;

   // m58_13 = W*in
   wire signed [14:0] m58_13;
   assign m58_13 =15'b0;

   // m58_14 = W*in
   wire signed [14:0] m58_14;
   assign m58_14 =15'b0;

   // m58_15 = W*in
   wire signed [14:0] m58_15;
   assign m58_15 =15'b0;

   // m58_16 = W*in
   wire signed [14:0] m58_16;
   assign m58_16 =15'b0;

   // m58_17 = W*in
   wire signed [14:0] m58_17;
   assign m58_17 =15'b0;

   // m58_18 = W*in
   wire signed [14:0] m58_18;
   assign m58_18 =15'b0;

   // m58_19 = W*in
   wire signed [14:0] m58_19;
   assign m58_19 =15'b0;

   // m58_20 = W*in
   wire signed [14:0] m58_20;
   assign m58_20 =15'b0;

   // m58_21 = W*in
   wire signed [14:0] m58_21;
   assign m58_21 =15'b0;

   // m58_22 = W*in
   wire signed [14:0] m58_22;
   assign m58_22 =15'b0;

   // m58_23 = W*in
   wire signed [14:0] m58_23;
   assign m58_23 =15'b0;

   // m58_24 = W*in
   wire signed [14:0] m58_24;
   assign m58_24 =15'b0;

   // m58_25 = W*in
   wire signed [14:0] m58_25;
   assign m58_25 =15'b0;

   // m58_26 = W*in
   wire signed [14:0] m58_26;
   assign m58_26 =15'b0;

   // m58_27 = W*in
   wire signed [14:0] m58_27;
   assign m58_27 =15'b0;

   // m58_28 = W*in
   wire signed [14:0] m58_28;
   assign m58_28 =15'b0;

   // m58_29 = W*in
   wire signed [14:0] m58_29;
   assign m58_29 =15'b0;

   // m58_30 = W*in
   wire signed [14:0] m58_30;
   assign m58_30 =15'b0;

   // m58_31 = W*in
   wire signed [14:0] m58_31;
   assign m58_31 =15'b0;

   // m58_32 = W*in
   wire signed [14:0] m58_32;
   assign m58_32 =15'b0;

   // m58_33 = W*in
   wire signed [14:0] m58_33;
   assign m58_33 =15'b0;

   // m58_34 = W*in
   wire signed [14:0] m58_34;
   assign m58_34 =15'b0;

   // m58_35 = W*in
   wire signed [14:0] m58_35;
   assign m58_35 =15'b0;

   // m58_36 = W*in
   wire signed [14:0] m58_36;
   assign m58_36 =15'b0;

   // m58_37 = W*in
   wire signed [14:0] m58_37;
   assign m58_37 =15'b0;

   // m58_38 = W*in
   wire signed [14:0] m58_38;
   assign m58_38 =15'b0;

   // m58_39 = W*in
   wire signed [14:0] m58_39;
   assign m58_39 =15'b0;

   // m58_40 = W*in
   wire signed [14:0] m58_40;
   assign m58_40 ={ {3{in58[14]}} , in58[14:3] };

   // m58_41 = W*in
   wire signed [14:0] m58_41;
   assign m58_41 =15'b0;

   // m58_42 = W*in
   wire signed [14:0] m58_42;
   assign m58_42 =15'b0;

   // m58_43 = W*in
   wire signed [14:0] m58_43;
   assign m58_43 =15'b0;

   // m58_44 = W*in
   wire signed [14:0] m58_44;
   assign m58_44 =15'b0;

   // m58_45 = W*in
   wire signed [14:0] m58_45;
   assign m58_45 =15'b0;

   // m58_46 = W*in
   wire signed [14:0] m58_46;
   assign m58_46 =15'b0;

   // m58_47 = W*in
   wire signed [14:0] m58_47;
   assign m58_47 =15'b0;

   // m58_48 = W*in
   wire signed [14:0] m58_48;
   assign m58_48 =15'b0;

   // m58_49 = W*in
   wire signed [14:0] m58_49;
   assign m58_49 =15'b0;

   // m58_50 = W*in
   wire signed [14:0] m58_50;
   assign m58_50 =15'b0;

   // m58_51 = W*in
   wire signed [14:0] m58_51;
   assign m58_51 =15'b0;

   // m58_52 = W*in
   wire signed [14:0] m58_52;
   assign m58_52 =15'b0;

   // m58_53 = W*in
   wire signed [14:0] m58_53;
   assign m58_53 =15'b0;

   // m58_54 = W*in
   wire signed [14:0] m58_54;
   assign m58_54 =15'b0;

   // m58_55 = W*in
   wire signed [14:0] m58_55;
   assign m58_55 =15'b0;

   // m58_56 = W*in
   wire signed [14:0] m58_56;
   assign m58_56 =15'b0;

   // m58_57 = W*in
   wire signed [14:0] m58_57;
   assign m58_57 =15'b0;

   // m58_58 = W*in
   wire signed [14:0] m58_58;
   assign m58_58 =15'b0;

   // m58_59 = W*in
   wire signed [14:0] m58_59;
   assign m58_59 =15'b0;

   // m58_60 = W*in
   wire signed [14:0] m58_60;
   assign m58_60 =15'b0;

   // m58_61 = W*in
   wire signed [14:0] m58_61;
   assign m58_61 =15'b0;

   // m58_62 = W*in
   wire signed [14:0] m58_62;
   assign m58_62 =15'b0;

   // m58_63 = W*in
   wire signed [14:0] m58_63;
   assign m58_63 =15'b0;

   // m58_64 = W*in
   wire signed [14:0] m58_64;
   assign m58_64 ={ {3{in58[14]}} , in58[14:3] };

   // m58_65 = W*in
   wire signed [14:0] m58_65;
   assign m58_65 =15'b0;

   // m58_66 = W*in
   wire signed [14:0] m58_66;
   assign m58_66 =15'b0;

   // m58_67 = W*in
   wire signed [14:0] m58_67;
   assign m58_67 =15'b0;

   // m58_68 = W*in
   wire signed [14:0] m58_68;
   assign m58_68 =15'b0;

   // m58_69 = W*in
   wire signed [14:0] m58_69;
   assign m58_69 ={ {4{neg58[14]}} , neg58[14:4] };

   // m58_70 = W*in
   wire signed [14:0] m58_70;
   assign m58_70 =15'b0;

   // m58_71 = W*in
   wire signed [14:0] m58_71;
   assign m58_71 =15'b0;

   // m58_72 = W*in
   wire signed [14:0] m58_72;
   assign m58_72 =15'b0;

   // m58_73 = W*in
   wire signed [14:0] m58_73;
   assign m58_73 =15'b0;

   // m58_74 = W*in
   wire signed [14:0] m58_74;
   assign m58_74 =15'b0;

   // m58_75 = W*in
   wire signed [14:0] m58_75;
   assign m58_75 =15'b0;

   // m58_76 = W*in
   wire signed [14:0] m58_76;
   assign m58_76 =15'b0;

   // m58_77 = W*in
   wire signed [14:0] m58_77;
   assign m58_77 =15'b0;

   // m58_78 = W*in
   wire signed [14:0] m58_78;
   assign m58_78 =15'b0;

   // m58_79 = W*in
   wire signed [14:0] m58_79;
   assign m58_79 =15'b0;

   // m58_80 = W*in
   wire signed [14:0] m58_80;
   assign m58_80 =15'b0;

   // m58_81 = W*in
   wire signed [14:0] m58_81;
   assign m58_81 ={ {3{in58[14]}} , in58[14:3] };

   // m58_82 = W*in
   wire signed [14:0] m58_82;
   assign m58_82 =15'b0;

   // m58_83 = W*in
   wire signed [14:0] m58_83;
   assign m58_83 =15'b0;

   // m58_84 = W*in
   wire signed [14:0] m58_84;
   assign m58_84 =15'b0;

   // m58_85 = W*in
   wire signed [14:0] m58_85;
   assign m58_85 ={ {3{neg58[14]}} , neg58[14:3] };

   // m58_86 = W*in
   wire signed [14:0] m58_86;
   assign m58_86 =15'b0;

   // m58_87 = W*in
   wire signed [14:0] m58_87;
   assign m58_87 =15'b0;

   // m58_88 = W*in
   wire signed [14:0] m58_88;
   assign m58_88 =15'b0;

   // m58_89 = W*in
   wire signed [14:0] m58_89;
   assign m58_89 =15'b0;

   // m58_90 = W*in
   wire signed [14:0] m58_90;
   assign m58_90 =15'b0;

   // m58_91 = W*in
   wire signed [14:0] m58_91;
   assign m58_91 =15'b0;

   // m58_92 = W*in
   wire signed [14:0] m58_92;
   assign m58_92 =15'b0;

   // m58_93 = W*in
   wire signed [14:0] m58_93;
   assign m58_93 =15'b0;

   // m58_94 = W*in
   wire signed [14:0] m58_94;
   assign m58_94 =15'b0;

   // m58_95 = W*in
   wire signed [14:0] m58_95;
   assign m58_95 =15'b0;

   // m58_96 = W*in
   wire signed [14:0] m58_96;
   assign m58_96 =15'b0;

   // m58_97 = W*in
   wire signed [14:0] m58_97;
   assign m58_97 =15'b0;

   // m58_98 = W*in
   wire signed [14:0] m58_98;
   assign m58_98 =15'b0;

   // m58_99 = W*in
   wire signed [14:0] m58_99;
   assign m58_99 =15'b0;

   // m58_100 = W*in
   wire signed [14:0] m58_100;
   assign m58_100 =15'b0;

   // m59_1 = W*in
   wire signed [14:0] m59_1;
   assign m59_1 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_2 = W*in
   wire signed [14:0] m59_2;
   assign m59_2 =15'b0;

   // m59_3 = W*in
   wire signed [14:0] m59_3;
   assign m59_3 =15'b0;

   // m59_4 = W*in
   wire signed [14:0] m59_4;
   assign m59_4 =15'b0;

   // m59_5 = W*in
   wire signed [14:0] m59_5;
   assign m59_5 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_6 = W*in
   wire signed [14:0] m59_6;
   assign m59_6 ={ {2{in59[14]}} , in59[14:2] };

   // m59_7 = W*in
   wire signed [14:0] m59_7;
   assign m59_7 =15'b0;

   // m59_8 = W*in
   wire signed [14:0] m59_8;
   assign m59_8 =15'b0;

   // m59_9 = W*in
   wire signed [14:0] m59_9;
   assign m59_9 =15'b0;

   // m59_10 = W*in
   wire signed [14:0] m59_10;
   assign m59_10 =15'b0;

   // m59_11 = W*in
   wire signed [14:0] m59_11;
   assign m59_11 =15'b0;

   // m59_12 = W*in
   wire signed [14:0] m59_12;
   assign m59_12 ={ {3{in59[14]}} , in59[14:3] };

   // m59_13 = W*in
   wire signed [14:0] m59_13;
   assign m59_13 =15'b0;

   // m59_14 = W*in
   wire signed [14:0] m59_14;
   assign m59_14 =15'b0;

   // m59_15 = W*in
   wire signed [14:0] m59_15;
   assign m59_15 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_16 = W*in
   wire signed [14:0] m59_16;
   assign m59_16 =15'b0;

   // m59_17 = W*in
   wire signed [14:0] m59_17;
   assign m59_17 =15'b0;

   // m59_18 = W*in
   wire signed [14:0] m59_18;
   assign m59_18 =15'b0;

   // m59_19 = W*in
   wire signed [14:0] m59_19;
   assign m59_19 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_20 = W*in
   wire signed [14:0] m59_20;
   assign m59_20 =15'b0;

   // m59_21 = W*in
   wire signed [14:0] m59_21;
   assign m59_21 =15'b0;

   // m59_22 = W*in
   wire signed [14:0] m59_22;
   assign m59_22 =15'b0;

   // m59_23 = W*in
   wire signed [14:0] m59_23;
   assign m59_23 =15'b0;

   // m59_24 = W*in
   wire signed [14:0] m59_24;
   assign m59_24 =15'b0;

   // m59_25 = W*in
   wire signed [14:0] m59_25;
   assign m59_25 ={ {3{in59[14]}} , in59[14:3] };

   // m59_26 = W*in
   wire signed [14:0] m59_26;
   assign m59_26 =15'b0;

   // m59_27 = W*in
   wire signed [14:0] m59_27;
   assign m59_27 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_28 = W*in
   wire signed [14:0] m59_28;
   assign m59_28 ={ {4{neg59[14]}} , neg59[14:4] };

   // m59_29 = W*in
   wire signed [14:0] m59_29;
   assign m59_29 ={ {3{in59[14]}} , in59[14:3] };

   // m59_30 = W*in
   wire signed [14:0] m59_30;
   assign m59_30 =15'b0;

   // m59_31 = W*in
   wire signed [14:0] m59_31;
   assign m59_31 ={ {3{in59[14]}} , in59[14:3] };

   // m59_32 = W*in
   wire signed [14:0] m59_32;
   assign m59_32 =15'b0;

   // m59_33 = W*in
   wire signed [14:0] m59_33;
   assign m59_33 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_34 = W*in
   wire signed [14:0] m59_34;
   assign m59_34 ={ {3{in59[14]}} , in59[14:3] };

   // m59_35 = W*in
   wire signed [14:0] m59_35;
   assign m59_35 =15'b0;

   // m59_36 = W*in
   wire signed [14:0] m59_36;
   assign m59_36 =15'b0;

   // m59_37 = W*in
   wire signed [14:0] m59_37;
   assign m59_37 =15'b0;

   // m59_38 = W*in
   wire signed [14:0] m59_38;
   assign m59_38 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_39 = W*in
   wire signed [14:0] m59_39;
   assign m59_39 =15'b0;

   // m59_40 = W*in
   wire signed [14:0] m59_40;
   assign m59_40 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_41 = W*in
   wire signed [14:0] m59_41;
   assign m59_41 =15'b0;

   // m59_42 = W*in
   wire signed [14:0] m59_42;
   assign m59_42 =15'b0;

   // m59_43 = W*in
   wire signed [14:0] m59_43;
   assign m59_43 =15'b0;

   // m59_44 = W*in
   wire signed [14:0] m59_44;
   assign m59_44 =15'b0;

   // m59_45 = W*in
   wire signed [14:0] m59_45;
   assign m59_45 =15'b0;

   // m59_46 = W*in
   wire signed [14:0] m59_46;
   assign m59_46 =15'b0;

   // m59_47 = W*in
   wire signed [14:0] m59_47;
   assign m59_47 =15'b0;

   // m59_48 = W*in
   wire signed [14:0] m59_48;
   assign m59_48 =15'b0;

   // m59_49 = W*in
   wire signed [14:0] m59_49;
   assign m59_49 ={ {3{in59[14]}} , in59[14:3] };

   // m59_50 = W*in
   wire signed [14:0] m59_50;
   assign m59_50 ={ {3{in59[14]}} , in59[14:3] };

   // m59_51 = W*in
   wire signed [14:0] m59_51;
   assign m59_51 =15'b0;

   // m59_52 = W*in
   wire signed [14:0] m59_52;
   assign m59_52 ={ {3{in59[14]}} , in59[14:3] };

   // m59_53 = W*in
   wire signed [14:0] m59_53;
   assign m59_53 =15'b0;

   // m59_54 = W*in
   wire signed [14:0] m59_54;
   assign m59_54 =15'b0;

   // m59_55 = W*in
   wire signed [14:0] m59_55;
   assign m59_55 =15'b0;

   // m59_56 = W*in
   wire signed [14:0] m59_56;
   assign m59_56 =15'b0;

   // m59_57 = W*in
   wire signed [14:0] m59_57;
   assign m59_57 =15'b0;

   // m59_58 = W*in
   wire signed [14:0] m59_58;
   assign m59_58 =15'b0;

   // m59_59 = W*in
   wire signed [14:0] m59_59;
   assign m59_59 =15'b0;

   // m59_60 = W*in
   wire signed [14:0] m59_60;
   assign m59_60 ={ {2{in59[14]}} , in59[14:2] };

   // m59_61 = W*in
   wire signed [14:0] m59_61;
   assign m59_61 ={ {4{neg59[14]}} , neg59[14:4] };

   // m59_62 = W*in
   wire signed [14:0] m59_62;
   assign m59_62 =15'b0;

   // m59_63 = W*in
   wire signed [14:0] m59_63;
   assign m59_63 =15'b0;

   // m59_64 = W*in
   wire signed [14:0] m59_64;
   assign m59_64 =15'b0;

   // m59_65 = W*in
   wire signed [14:0] m59_65;
   assign m59_65 =15'b0;

   // m59_66 = W*in
   wire signed [14:0] m59_66;
   assign m59_66 =15'b0;

   // m59_67 = W*in
   wire signed [14:0] m59_67;
   assign m59_67 =15'b0;

   // m59_68 = W*in
   wire signed [14:0] m59_68;
   assign m59_68 =15'b0;

   // m59_69 = W*in
   wire signed [14:0] m59_69;
   assign m59_69 =15'b0;

   // m59_70 = W*in
   wire signed [14:0] m59_70;
   assign m59_70 =15'b0;

   // m59_71 = W*in
   wire signed [14:0] m59_71;
   assign m59_71 =15'b0;

   // m59_72 = W*in
   wire signed [14:0] m59_72;
   assign m59_72 =15'b0;

   // m59_73 = W*in
   wire signed [14:0] m59_73;
   assign m59_73 =15'b0;

   // m59_74 = W*in
   wire signed [14:0] m59_74;
   assign m59_74 =15'b0;

   // m59_75 = W*in
   wire signed [14:0] m59_75;
   assign m59_75 =15'b0;

   // m59_76 = W*in
   wire signed [14:0] m59_76;
   assign m59_76 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_77 = W*in
   wire signed [14:0] m59_77;
   assign m59_77 ={ {3{in59[14]}} , in59[14:3] };

   // m59_78 = W*in
   wire signed [14:0] m59_78;
   assign m59_78 =15'b0;

   // m59_79 = W*in
   wire signed [14:0] m59_79;
   assign m59_79 =15'b0;

   // m59_80 = W*in
   wire signed [14:0] m59_80;
   assign m59_80 =15'b0;

   // m59_81 = W*in
   wire signed [14:0] m59_81;
   assign m59_81 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_82 = W*in
   wire signed [14:0] m59_82;
   assign m59_82 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_83 = W*in
   wire signed [14:0] m59_83;
   assign m59_83 =15'b0;

   // m59_84 = W*in
   wire signed [14:0] m59_84;
   assign m59_84 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_85 = W*in
   wire signed [14:0] m59_85;
   assign m59_85 =15'b0;

   // m59_86 = W*in
   wire signed [14:0] m59_86;
   assign m59_86 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_87 = W*in
   wire signed [14:0] m59_87;
   assign m59_87 =15'b0;

   // m59_88 = W*in
   wire signed [14:0] m59_88;
   assign m59_88 ={ {3{in59[14]}} , in59[14:3] };

   // m59_89 = W*in
   wire signed [14:0] m59_89;
   assign m59_89 =15'b0;

   // m59_90 = W*in
   wire signed [14:0] m59_90;
   assign m59_90 =15'b0;

   // m59_91 = W*in
   wire signed [14:0] m59_91;
   assign m59_91 =15'b0;

   // m59_92 = W*in
   wire signed [14:0] m59_92;
   assign m59_92 =15'b0;

   // m59_93 = W*in
   wire signed [14:0] m59_93;
   assign m59_93 =15'b0;

   // m59_94 = W*in
   wire signed [14:0] m59_94;
   assign m59_94 ={ {4{neg59[14]}} , neg59[14:4] };

   // m59_95 = W*in
   wire signed [14:0] m59_95;
   assign m59_95 =15'b0;

   // m59_96 = W*in
   wire signed [14:0] m59_96;
   assign m59_96 ={ {2{in59[14]}} , in59[14:2] };

   // m59_97 = W*in
   wire signed [14:0] m59_97;
   assign m59_97 ={ {3{neg59[14]}} , neg59[14:3] };

   // m59_98 = W*in
   wire signed [14:0] m59_98;
   assign m59_98 =15'b0;

   // m59_99 = W*in
   wire signed [14:0] m59_99;
   assign m59_99 =15'b0;

   // m59_100 = W*in
   wire signed [14:0] m59_100;
   assign m59_100 =15'b0;

   // m60_1 = W*in
   wire signed [14:0] m60_1;
   assign m60_1 =15'b0;

   // m60_2 = W*in
   wire signed [14:0] m60_2;
   assign m60_2 =15'b0;

   // m60_3 = W*in
   wire signed [14:0] m60_3;
   assign m60_3 =15'b0;

   // m60_4 = W*in
   wire signed [14:0] m60_4;
   assign m60_4 =15'b0;

   // m60_5 = W*in
   wire signed [14:0] m60_5;
   assign m60_5 =15'b0;

   // m60_6 = W*in
   wire signed [14:0] m60_6;
   assign m60_6 =15'b0;

   // m60_7 = W*in
   wire signed [14:0] m60_7;
   assign m60_7 =15'b0;

   // m60_8 = W*in
   wire signed [14:0] m60_8;
   assign m60_8 ={ {4{neg60[14]}} , neg60[14:4] };

   // m60_9 = W*in
   wire signed [14:0] m60_9;
   assign m60_9 =15'b0;

   // m60_10 = W*in
   wire signed [14:0] m60_10;
   assign m60_10 =15'b0;

   // m60_11 = W*in
   wire signed [14:0] m60_11;
   assign m60_11 =15'b0;

   // m60_12 = W*in
   wire signed [14:0] m60_12;
   assign m60_12 =15'b0;

   // m60_13 = W*in
   wire signed [14:0] m60_13;
   assign m60_13 =15'b0;

   // m60_14 = W*in
   wire signed [14:0] m60_14;
   assign m60_14 =15'b0;

   // m60_15 = W*in
   wire signed [14:0] m60_15;
   assign m60_15 =15'b0;

   // m60_16 = W*in
   wire signed [14:0] m60_16;
   assign m60_16 =15'b0;

   // m60_17 = W*in
   wire signed [14:0] m60_17;
   assign m60_17 =15'b0;

   // m60_18 = W*in
   wire signed [14:0] m60_18;
   assign m60_18 =15'b0;

   // m60_19 = W*in
   wire signed [14:0] m60_19;
   assign m60_19 ={ {4{in60[14]}} , in60[14:4] };

   // m60_20 = W*in
   wire signed [14:0] m60_20;
   assign m60_20 =15'b0;

   // m60_21 = W*in
   wire signed [14:0] m60_21;
   assign m60_21 =15'b0;

   // m60_22 = W*in
   wire signed [14:0] m60_22;
   assign m60_22 ={ {4{in60[14]}} , in60[14:4] };

   // m60_23 = W*in
   wire signed [14:0] m60_23;
   assign m60_23 =15'b0;

   // m60_24 = W*in
   wire signed [14:0] m60_24;
   assign m60_24 =15'b0;

   // m60_25 = W*in
   wire signed [14:0] m60_25;
   assign m60_25 =15'b0;

   // m60_26 = W*in
   wire signed [14:0] m60_26;
   assign m60_26 =15'b0;

   // m60_27 = W*in
   wire signed [14:0] m60_27;
   assign m60_27 =15'b0;

   // m60_28 = W*in
   wire signed [14:0] m60_28;
   assign m60_28 =15'b0;

   // m60_29 = W*in
   wire signed [14:0] m60_29;
   assign m60_29 =15'b0;

   // m60_30 = W*in
   wire signed [14:0] m60_30;
   assign m60_30 =15'b0;

   // m60_31 = W*in
   wire signed [14:0] m60_31;
   assign m60_31 ={ {4{neg60[14]}} , neg60[14:4] };

   // m60_32 = W*in
   wire signed [14:0] m60_32;
   assign m60_32 =15'b0;

   // m60_33 = W*in
   wire signed [14:0] m60_33;
   assign m60_33 =15'b0;

   // m60_34 = W*in
   wire signed [14:0] m60_34;
   assign m60_34 =15'b0;

   // m60_35 = W*in
   wire signed [14:0] m60_35;
   assign m60_35 =15'b0;

   // m60_36 = W*in
   wire signed [14:0] m60_36;
   assign m60_36 =15'b0;

   // m60_37 = W*in
   wire signed [14:0] m60_37;
   assign m60_37 =15'b0;

   // m60_38 = W*in
   wire signed [14:0] m60_38;
   assign m60_38 =15'b0;

   // m60_39 = W*in
   wire signed [14:0] m60_39;
   assign m60_39 =15'b0;

   // m60_40 = W*in
   wire signed [14:0] m60_40;
   assign m60_40 =15'b0;

   // m60_41 = W*in
   wire signed [14:0] m60_41;
   assign m60_41 =15'b0;

   // m60_42 = W*in
   wire signed [14:0] m60_42;
   assign m60_42 =15'b0;

   // m60_43 = W*in
   wire signed [14:0] m60_43;
   assign m60_43 =15'b0;

   // m60_44 = W*in
   wire signed [14:0] m60_44;
   assign m60_44 ={ {4{neg60[14]}} , neg60[14:4] };

   // m60_45 = W*in
   wire signed [14:0] m60_45;
   assign m60_45 =15'b0;

   // m60_46 = W*in
   wire signed [14:0] m60_46;
   assign m60_46 =15'b0;

   // m60_47 = W*in
   wire signed [14:0] m60_47;
   assign m60_47 =15'b0;

   // m60_48 = W*in
   wire signed [14:0] m60_48;
   assign m60_48 =15'b0;

   // m60_49 = W*in
   wire signed [14:0] m60_49;
   assign m60_49 =15'b0;

   // m60_50 = W*in
   wire signed [14:0] m60_50;
   assign m60_50 =15'b0;

   // m60_51 = W*in
   wire signed [14:0] m60_51;
   assign m60_51 =15'b0;

   // m60_52 = W*in
   wire signed [14:0] m60_52;
   assign m60_52 =15'b0;

   // m60_53 = W*in
   wire signed [14:0] m60_53;
   assign m60_53 =15'b0;

   // m60_54 = W*in
   wire signed [14:0] m60_54;
   assign m60_54 =15'b0;

   // m60_55 = W*in
   wire signed [14:0] m60_55;
   assign m60_55 =15'b0;

   // m60_56 = W*in
   wire signed [14:0] m60_56;
   assign m60_56 =15'b0;

   // m60_57 = W*in
   wire signed [14:0] m60_57;
   assign m60_57 =15'b0;

   // m60_58 = W*in
   wire signed [14:0] m60_58;
   assign m60_58 ={ {3{in60[14]}} , in60[14:3] };

   // m60_59 = W*in
   wire signed [14:0] m60_59;
   assign m60_59 =15'b0;

   // m60_60 = W*in
   wire signed [14:0] m60_60;
   assign m60_60 =15'b0;

   // m60_61 = W*in
   wire signed [14:0] m60_61;
   assign m60_61 ={ {4{in60[14]}} , in60[14:4] };

   // m60_62 = W*in
   wire signed [14:0] m60_62;
   assign m60_62 =15'b0;

   // m60_63 = W*in
   wire signed [14:0] m60_63;
   assign m60_63 =15'b0;

   // m60_64 = W*in
   wire signed [14:0] m60_64;
   assign m60_64 =15'b0;

   // m60_65 = W*in
   wire signed [14:0] m60_65;
   assign m60_65 =15'b0;

   // m60_66 = W*in
   wire signed [14:0] m60_66;
   assign m60_66 =15'b0;

   // m60_67 = W*in
   wire signed [14:0] m60_67;
   assign m60_67 =15'b0;

   // m60_68 = W*in
   wire signed [14:0] m60_68;
   assign m60_68 =15'b0;

   // m60_69 = W*in
   wire signed [14:0] m60_69;
   assign m60_69 =15'b0;

   // m60_70 = W*in
   wire signed [14:0] m60_70;
   assign m60_70 =15'b0;

   // m60_71 = W*in
   wire signed [14:0] m60_71;
   assign m60_71 =15'b0;

   // m60_72 = W*in
   wire signed [14:0] m60_72;
   assign m60_72 =15'b0;

   // m60_73 = W*in
   wire signed [14:0] m60_73;
   assign m60_73 =15'b0;

   // m60_74 = W*in
   wire signed [14:0] m60_74;
   assign m60_74 =15'b0;

   // m60_75 = W*in
   wire signed [14:0] m60_75;
   assign m60_75 =15'b0;

   // m60_76 = W*in
   wire signed [14:0] m60_76;
   assign m60_76 ={ {3{neg60[14]}} , neg60[14:3] };

   // m60_77 = W*in
   wire signed [14:0] m60_77;
   assign m60_77 =15'b0;

   // m60_78 = W*in
   wire signed [14:0] m60_78;
   assign m60_78 =15'b0;

   // m60_79 = W*in
   wire signed [14:0] m60_79;
   assign m60_79 ={ {4{neg60[14]}} , neg60[14:4] };

   // m60_80 = W*in
   wire signed [14:0] m60_80;
   assign m60_80 =15'b0;

   // m60_81 = W*in
   wire signed [14:0] m60_81;
   assign m60_81 =15'b0;

   // m60_82 = W*in
   wire signed [14:0] m60_82;
   assign m60_82 =15'b0;

   // m60_83 = W*in
   wire signed [14:0] m60_83;
   assign m60_83 =15'b0;

   // m60_84 = W*in
   wire signed [14:0] m60_84;
   assign m60_84 =15'b0;

   // m60_85 = W*in
   wire signed [14:0] m60_85;
   assign m60_85 =15'b0;

   // m60_86 = W*in
   wire signed [14:0] m60_86;
   assign m60_86 =15'b0;

   // m60_87 = W*in
   wire signed [14:0] m60_87;
   assign m60_87 =15'b0;

   // m60_88 = W*in
   wire signed [14:0] m60_88;
   assign m60_88 =15'b0;

   // m60_89 = W*in
   wire signed [14:0] m60_89;
   assign m60_89 ={ {4{neg60[14]}} , neg60[14:4] };

   // m60_90 = W*in
   wire signed [14:0] m60_90;
   assign m60_90 =15'b0;

   // m60_91 = W*in
   wire signed [14:0] m60_91;
   assign m60_91 ={ {3{in60[14]}} , in60[14:3] };

   // m60_92 = W*in
   wire signed [14:0] m60_92;
   assign m60_92 =15'b0;

   // m60_93 = W*in
   wire signed [14:0] m60_93;
   assign m60_93 =15'b0;

   // m60_94 = W*in
   wire signed [14:0] m60_94;
   assign m60_94 =15'b0;

   // m60_95 = W*in
   wire signed [14:0] m60_95;
   assign m60_95 ={ {4{neg60[14]}} , neg60[14:4] };

   // m60_96 = W*in
   wire signed [14:0] m60_96;
   assign m60_96 =15'b0;

   // m60_97 = W*in
   wire signed [14:0] m60_97;
   assign m60_97 =15'b0;

   // m60_98 = W*in
   wire signed [14:0] m60_98;
   assign m60_98 =15'b0;

   // m60_99 = W*in
   wire signed [14:0] m60_99;
   assign m60_99 =15'b0;

   // m60_100 = W*in
   wire signed [14:0] m60_100;
   assign m60_100 =15'b0;

   // m61_1 = W*in
   wire signed [14:0] m61_1;
   assign m61_1 =15'b0;

   // m61_2 = W*in
   wire signed [14:0] m61_2;
   assign m61_2 ={ {3{in61[14]}} , in61[14:3] };

   // m61_3 = W*in
   wire signed [14:0] m61_3;
   assign m61_3 =15'b0;

   // m61_4 = W*in
   wire signed [14:0] m61_4;
   assign m61_4 =15'b0;

   // m61_5 = W*in
   wire signed [14:0] m61_5;
   assign m61_5 =15'b0;

   // m61_6 = W*in
   wire signed [14:0] m61_6;
   assign m61_6 =15'b0;

   // m61_7 = W*in
   wire signed [14:0] m61_7;
   assign m61_7 =15'b0;

   // m61_8 = W*in
   wire signed [14:0] m61_8;
   assign m61_8 =15'b0;

   // m61_9 = W*in
   wire signed [14:0] m61_9;
   assign m61_9 ={ {3{in61[14]}} , in61[14:3] };

   // m61_10 = W*in
   wire signed [14:0] m61_10;
   assign m61_10 =15'b0;

   // m61_11 = W*in
   wire signed [14:0] m61_11;
   assign m61_11 =15'b0;

   // m61_12 = W*in
   wire signed [14:0] m61_12;
   assign m61_12 =15'b0;

   // m61_13 = W*in
   wire signed [14:0] m61_13;
   assign m61_13 =15'b0;

   // m61_14 = W*in
   wire signed [14:0] m61_14;
   assign m61_14 =15'b0;

   // m61_15 = W*in
   wire signed [14:0] m61_15;
   assign m61_15 =15'b0;

   // m61_16 = W*in
   wire signed [14:0] m61_16;
   assign m61_16 ={ {4{neg61[14]}} , neg61[14:4] };

   // m61_17 = W*in
   wire signed [14:0] m61_17;
   assign m61_17 =15'b0;

   // m61_18 = W*in
   wire signed [14:0] m61_18;
   assign m61_18 =15'b0;

   // m61_19 = W*in
   wire signed [14:0] m61_19;
   assign m61_19 =15'b0;

   // m61_20 = W*in
   wire signed [14:0] m61_20;
   assign m61_20 =15'b0;

   // m61_21 = W*in
   wire signed [14:0] m61_21;
   assign m61_21 =15'b0;

   // m61_22 = W*in
   wire signed [14:0] m61_22;
   assign m61_22 =15'b0;

   // m61_23 = W*in
   wire signed [14:0] m61_23;
   assign m61_23 =15'b0;

   // m61_24 = W*in
   wire signed [14:0] m61_24;
   assign m61_24 =15'b0;

   // m61_25 = W*in
   wire signed [14:0] m61_25;
   assign m61_25 =15'b0;

   // m61_26 = W*in
   wire signed [14:0] m61_26;
   assign m61_26 =15'b0;

   // m61_27 = W*in
   wire signed [14:0] m61_27;
   assign m61_27 =15'b0;

   // m61_28 = W*in
   wire signed [14:0] m61_28;
   assign m61_28 ={ {3{in61[14]}} , in61[14:3] };

   // m61_29 = W*in
   wire signed [14:0] m61_29;
   assign m61_29 =15'b0;

   // m61_30 = W*in
   wire signed [14:0] m61_30;
   assign m61_30 =15'b0;

   // m61_31 = W*in
   wire signed [14:0] m61_31;
   assign m61_31 =15'b0;

   // m61_32 = W*in
   wire signed [14:0] m61_32;
   assign m61_32 =15'b0;

   // m61_33 = W*in
   wire signed [14:0] m61_33;
   assign m61_33 ={ {3{in61[14]}} , in61[14:3] };

   // m61_34 = W*in
   wire signed [14:0] m61_34;
   assign m61_34 =15'b0;

   // m61_35 = W*in
   wire signed [14:0] m61_35;
   assign m61_35 =15'b0;

   // m61_36 = W*in
   wire signed [14:0] m61_36;
   assign m61_36 =15'b0;

   // m61_37 = W*in
   wire signed [14:0] m61_37;
   assign m61_37 =15'b0;

   // m61_38 = W*in
   wire signed [14:0] m61_38;
   assign m61_38 =15'b0;

   // m61_39 = W*in
   wire signed [14:0] m61_39;
   assign m61_39 =15'b0;

   // m61_40 = W*in
   wire signed [14:0] m61_40;
   assign m61_40 =15'b0;

   // m61_41 = W*in
   wire signed [14:0] m61_41;
   assign m61_41 =15'b0;

   // m61_42 = W*in
   wire signed [14:0] m61_42;
   assign m61_42 ={ {3{neg61[14]}} , neg61[14:3] };

   // m61_43 = W*in
   wire signed [14:0] m61_43;
   assign m61_43 =15'b0;

   // m61_44 = W*in
   wire signed [14:0] m61_44;
   assign m61_44 =15'b0;

   // m61_45 = W*in
   wire signed [14:0] m61_45;
   assign m61_45 =15'b0;

   // m61_46 = W*in
   wire signed [14:0] m61_46;
   assign m61_46 =15'b0;

   // m61_47 = W*in
   wire signed [14:0] m61_47;
   assign m61_47 =15'b0;

   // m61_48 = W*in
   wire signed [14:0] m61_48;
   assign m61_48 =15'b0;

   // m61_49 = W*in
   wire signed [14:0] m61_49;
   assign m61_49 =15'b0;

   // m61_50 = W*in
   wire signed [14:0] m61_50;
   assign m61_50 =15'b0;

   // m61_51 = W*in
   wire signed [14:0] m61_51;
   assign m61_51 =15'b0;

   // m61_52 = W*in
   wire signed [14:0] m61_52;
   assign m61_52 =15'b0;

   // m61_53 = W*in
   wire signed [14:0] m61_53;
   assign m61_53 =15'b0;

   // m61_54 = W*in
   wire signed [14:0] m61_54;
   assign m61_54 =15'b0;

   // m61_55 = W*in
   wire signed [14:0] m61_55;
   assign m61_55 =15'b0;

   // m61_56 = W*in
   wire signed [14:0] m61_56;
   assign m61_56 =15'b0;

   // m61_57 = W*in
   wire signed [14:0] m61_57;
   assign m61_57 ={ {3{in61[14]}} , in61[14:3] };

   // m61_58 = W*in
   wire signed [14:0] m61_58;
   assign m61_58 =15'b0;

   // m61_59 = W*in
   wire signed [14:0] m61_59;
   assign m61_59 ={ {3{in61[14]}} , in61[14:3] };

   // m61_60 = W*in
   wire signed [14:0] m61_60;
   assign m61_60 =15'b0;

   // m61_61 = W*in
   wire signed [14:0] m61_61;
   assign m61_61 =15'b0;

   // m61_62 = W*in
   wire signed [14:0] m61_62;
   assign m61_62 =15'b0;

   // m61_63 = W*in
   wire signed [14:0] m61_63;
   assign m61_63 =15'b0;

   // m61_64 = W*in
   wire signed [14:0] m61_64;
   assign m61_64 =15'b0;

   // m61_65 = W*in
   wire signed [14:0] m61_65;
   assign m61_65 =15'b0;

   // m61_66 = W*in
   wire signed [14:0] m61_66;
   assign m61_66 =15'b0;

   // m61_67 = W*in
   wire signed [14:0] m61_67;
   assign m61_67 =15'b0;

   // m61_68 = W*in
   wire signed [14:0] m61_68;
   assign m61_68 =15'b0;

   // m61_69 = W*in
   wire signed [14:0] m61_69;
   assign m61_69 =15'b0;

   // m61_70 = W*in
   wire signed [14:0] m61_70;
   assign m61_70 =15'b0;

   // m61_71 = W*in
   wire signed [14:0] m61_71;
   assign m61_71 =15'b0;

   // m61_72 = W*in
   wire signed [14:0] m61_72;
   assign m61_72 =15'b0;

   // m61_73 = W*in
   wire signed [14:0] m61_73;
   assign m61_73 =15'b0;

   // m61_74 = W*in
   wire signed [14:0] m61_74;
   assign m61_74 ={ {3{in61[14]}} , in61[14:3] };

   // m61_75 = W*in
   wire signed [14:0] m61_75;
   assign m61_75 =15'b0;

   // m61_76 = W*in
   wire signed [14:0] m61_76;
   assign m61_76 =15'b0;

   // m61_77 = W*in
   wire signed [14:0] m61_77;
   assign m61_77 ={ {3{neg61[14]}} , neg61[14:3] };

   // m61_78 = W*in
   wire signed [14:0] m61_78;
   assign m61_78 =15'b0;

   // m61_79 = W*in
   wire signed [14:0] m61_79;
   assign m61_79 =15'b0;

   // m61_80 = W*in
   wire signed [14:0] m61_80;
   assign m61_80 =15'b0;

   // m61_81 = W*in
   wire signed [14:0] m61_81;
   assign m61_81 =15'b0;

   // m61_82 = W*in
   wire signed [14:0] m61_82;
   assign m61_82 ={ {4{in61[14]}} , in61[14:4] };

   // m61_83 = W*in
   wire signed [14:0] m61_83;
   assign m61_83 =15'b0;

   // m61_84 = W*in
   wire signed [14:0] m61_84;
   assign m61_84 =15'b0;

   // m61_85 = W*in
   wire signed [14:0] m61_85;
   assign m61_85 ={ {3{neg61[14]}} , neg61[14:3] };

   // m61_86 = W*in
   wire signed [14:0] m61_86;
   assign m61_86 =15'b0;

   // m61_87 = W*in
   wire signed [14:0] m61_87;
   assign m61_87 ={ {3{neg61[14]}} , neg61[14:3] };

   // m61_88 = W*in
   wire signed [14:0] m61_88;
   assign m61_88 =15'b0;

   // m61_89 = W*in
   wire signed [14:0] m61_89;
   assign m61_89 =15'b0;

   // m61_90 = W*in
   wire signed [14:0] m61_90;
   assign m61_90 ={ {3{in61[14]}} , in61[14:3] };

   // m61_91 = W*in
   wire signed [14:0] m61_91;
   assign m61_91 =15'b0;

   // m61_92 = W*in
   wire signed [14:0] m61_92;
   assign m61_92 ={ {3{in61[14]}} , in61[14:3] };

   // m61_93 = W*in
   wire signed [14:0] m61_93;
   assign m61_93 =15'b0;

   // m61_94 = W*in
   wire signed [14:0] m61_94;
   assign m61_94 ={ {4{in61[14]}} , in61[14:4] };

   // m61_95 = W*in
   wire signed [14:0] m61_95;
   assign m61_95 =15'b0;

   // m61_96 = W*in
   wire signed [14:0] m61_96;
   assign m61_96 ={ {4{neg61[14]}} , neg61[14:4] };

   // m61_97 = W*in
   wire signed [14:0] m61_97;
   assign m61_97 =15'b0;

   // m61_98 = W*in
   wire signed [14:0] m61_98;
   assign m61_98 =15'b0;

   // m61_99 = W*in
   wire signed [14:0] m61_99;
   assign m61_99 ={ {3{in61[14]}} , in61[14:3] };

   // m61_100 = W*in
   wire signed [14:0] m61_100;
   assign m61_100 =15'b0;

   // m62_1 = W*in
   wire signed [14:0] m62_1;
   assign m62_1 =15'b0;

   // m62_2 = W*in
   wire signed [14:0] m62_2;
   assign m62_2 =15'b0;

   // m62_3 = W*in
   wire signed [14:0] m62_3;
   assign m62_3 =15'b0;

   // m62_4 = W*in
   wire signed [14:0] m62_4;
   assign m62_4 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_5 = W*in
   wire signed [14:0] m62_5;
   assign m62_5 =15'b0;

   // m62_6 = W*in
   wire signed [14:0] m62_6;
   assign m62_6 =15'b0;

   // m62_7 = W*in
   wire signed [14:0] m62_7;
   assign m62_7 ={ {3{in62[14]}} , in62[14:3] };

   // m62_8 = W*in
   wire signed [14:0] m62_8;
   assign m62_8 =15'b0;

   // m62_9 = W*in
   wire signed [14:0] m62_9;
   assign m62_9 ={ {2{in62[14]}} , in62[14:2] };

   // m62_10 = W*in
   wire signed [14:0] m62_10;
   assign m62_10 =15'b0;

   // m62_11 = W*in
   wire signed [14:0] m62_11;
   assign m62_11 =15'b0;

   // m62_12 = W*in
   wire signed [14:0] m62_12;
   assign m62_12 =15'b0;

   // m62_13 = W*in
   wire signed [14:0] m62_13;
   assign m62_13 ={ {3{in62[14]}} , in62[14:3] };

   // m62_14 = W*in
   wire signed [14:0] m62_14;
   assign m62_14 =15'b0;

   // m62_15 = W*in
   wire signed [14:0] m62_15;
   assign m62_15 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_16 = W*in
   wire signed [14:0] m62_16;
   assign m62_16 =15'b0;

   // m62_17 = W*in
   wire signed [14:0] m62_17;
   assign m62_17 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_18 = W*in
   wire signed [14:0] m62_18;
   assign m62_18 ={ {3{in62[14]}} , in62[14:3] };

   // m62_19 = W*in
   wire signed [14:0] m62_19;
   assign m62_19 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_20 = W*in
   wire signed [14:0] m62_20;
   assign m62_20 =15'b0;

   // m62_21 = W*in
   wire signed [14:0] m62_21;
   assign m62_21 =15'b0;

   // m62_22 = W*in
   wire signed [14:0] m62_22;
   assign m62_22 =15'b0;

   // m62_23 = W*in
   wire signed [14:0] m62_23;
   assign m62_23 =15'b0;

   // m62_24 = W*in
   wire signed [14:0] m62_24;
   assign m62_24 =15'b0;

   // m62_25 = W*in
   wire signed [14:0] m62_25;
   assign m62_25 =15'b0;

   // m62_26 = W*in
   wire signed [14:0] m62_26;
   assign m62_26 ={ {3{in62[14]}} , in62[14:3] };

   // m62_27 = W*in
   wire signed [14:0] m62_27;
   assign m62_27 =15'b0;

   // m62_28 = W*in
   wire signed [14:0] m62_28;
   assign m62_28 =15'b0;

   // m62_29 = W*in
   wire signed [14:0] m62_29;
   assign m62_29 ={ {3{in62[14]}} , in62[14:3] };

   // m62_30 = W*in
   wire signed [14:0] m62_30;
   assign m62_30 =15'b0;

   // m62_31 = W*in
   wire signed [14:0] m62_31;
   assign m62_31 ={ {2{in62[14]}} , in62[14:2] };

   // m62_32 = W*in
   wire signed [14:0] m62_32;
   assign m62_32 =15'b0;

   // m62_33 = W*in
   wire signed [14:0] m62_33;
   assign m62_33 =15'b0;

   // m62_34 = W*in
   wire signed [14:0] m62_34;
   assign m62_34 ={ {2{in62[14]}} , in62[14:2] };

   // m62_35 = W*in
   wire signed [14:0] m62_35;
   assign m62_35 =15'b0;

   // m62_36 = W*in
   wire signed [14:0] m62_36;
   assign m62_36 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_37 = W*in
   wire signed [14:0] m62_37;
   assign m62_37 =15'b0;

   // m62_38 = W*in
   wire signed [14:0] m62_38;
   assign m62_38 =15'b0;

   // m62_39 = W*in
   wire signed [14:0] m62_39;
   assign m62_39 =15'b0;

   // m62_40 = W*in
   wire signed [14:0] m62_40;
   assign m62_40 =15'b0;

   // m62_41 = W*in
   wire signed [14:0] m62_41;
   assign m62_41 =15'b0;

   // m62_42 = W*in
   wire signed [14:0] m62_42;
   assign m62_42 =15'b0;

   // m62_43 = W*in
   wire signed [14:0] m62_43;
   assign m62_43 =15'b0;

   // m62_44 = W*in
   wire signed [14:0] m62_44;
   assign m62_44 =15'b0;

   // m62_45 = W*in
   wire signed [14:0] m62_45;
   assign m62_45 =15'b0;

   // m62_46 = W*in
   wire signed [14:0] m62_46;
   assign m62_46 =15'b0;

   // m62_47 = W*in
   wire signed [14:0] m62_47;
   assign m62_47 =15'b0;

   // m62_48 = W*in
   wire signed [14:0] m62_48;
   assign m62_48 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_49 = W*in
   wire signed [14:0] m62_49;
   assign m62_49 =15'b0;

   // m62_50 = W*in
   wire signed [14:0] m62_50;
   assign m62_50 =15'b0;

   // m62_51 = W*in
   wire signed [14:0] m62_51;
   assign m62_51 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_52 = W*in
   wire signed [14:0] m62_52;
   assign m62_52 =15'b0;

   // m62_53 = W*in
   wire signed [14:0] m62_53;
   assign m62_53 =15'b0;

   // m62_54 = W*in
   wire signed [14:0] m62_54;
   assign m62_54 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_55 = W*in
   wire signed [14:0] m62_55;
   assign m62_55 =15'b0;

   // m62_56 = W*in
   wire signed [14:0] m62_56;
   assign m62_56 =15'b0;

   // m62_57 = W*in
   wire signed [14:0] m62_57;
   assign m62_57 =15'b0;

   // m62_58 = W*in
   wire signed [14:0] m62_58;
   assign m62_58 =15'b0;

   // m62_59 = W*in
   wire signed [14:0] m62_59;
   assign m62_59 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_60 = W*in
   wire signed [14:0] m62_60;
   assign m62_60 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_61 = W*in
   wire signed [14:0] m62_61;
   assign m62_61 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_62 = W*in
   wire signed [14:0] m62_62;
   assign m62_62 =15'b0;

   // m62_63 = W*in
   wire signed [14:0] m62_63;
   assign m62_63 =15'b0;

   // m62_64 = W*in
   wire signed [14:0] m62_64;
   assign m62_64 =15'b0;

   // m62_65 = W*in
   wire signed [14:0] m62_65;
   assign m62_65 =15'b0;

   // m62_66 = W*in
   wire signed [14:0] m62_66;
   assign m62_66 =15'b0;

   // m62_67 = W*in
   wire signed [14:0] m62_67;
   assign m62_67 =15'b0;

   // m62_68 = W*in
   wire signed [14:0] m62_68;
   assign m62_68 =15'b0;

   // m62_69 = W*in
   wire signed [14:0] m62_69;
   assign m62_69 =15'b0;

   // m62_70 = W*in
   wire signed [14:0] m62_70;
   assign m62_70 =15'b0;

   // m62_71 = W*in
   wire signed [14:0] m62_71;
   assign m62_71 =15'b0;

   // m62_72 = W*in
   wire signed [14:0] m62_72;
   assign m62_72 =15'b0;

   // m62_73 = W*in
   wire signed [14:0] m62_73;
   assign m62_73 =15'b0;

   // m62_74 = W*in
   wire signed [14:0] m62_74;
   assign m62_74 =15'b0;

   // m62_75 = W*in
   wire signed [14:0] m62_75;
   assign m62_75 =15'b0;

   // m62_76 = W*in
   wire signed [14:0] m62_76;
   assign m62_76 =15'b0;

   // m62_77 = W*in
   wire signed [14:0] m62_77;
   assign m62_77 =15'b0;

   // m62_78 = W*in
   wire signed [14:0] m62_78;
   assign m62_78 =15'b0;

   // m62_79 = W*in
   wire signed [14:0] m62_79;
   assign m62_79 =15'b0;

   // m62_80 = W*in
   wire signed [14:0] m62_80;
   assign m62_80 =15'b0;

   // m62_81 = W*in
   wire signed [14:0] m62_81;
   assign m62_81 ={ {2{neg62[14]}} , neg62[14:2] };

   // m62_82 = W*in
   wire signed [14:0] m62_82;
   assign m62_82 =15'b0;

   // m62_83 = W*in
   wire signed [14:0] m62_83;
   assign m62_83 =15'b0;

   // m62_84 = W*in
   wire signed [14:0] m62_84;
   assign m62_84 =15'b0;

   // m62_85 = W*in
   wire signed [14:0] m62_85;
   assign m62_85 =15'b0;

   // m62_86 = W*in
   wire signed [14:0] m62_86;
   assign m62_86 =15'b0;

   // m62_87 = W*in
   wire signed [14:0] m62_87;
   assign m62_87 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_88 = W*in
   wire signed [14:0] m62_88;
   assign m62_88 ={ {3{in62[14]}} , in62[14:3] };

   // m62_89 = W*in
   wire signed [14:0] m62_89;
   assign m62_89 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_90 = W*in
   wire signed [14:0] m62_90;
   assign m62_90 ={ {3{in62[14]}} , in62[14:3] };

   // m62_91 = W*in
   wire signed [14:0] m62_91;
   assign m62_91 ={ {3{neg62[14]}} , neg62[14:3] };

   // m62_92 = W*in
   wire signed [14:0] m62_92;
   assign m62_92 =15'b0;

   // m62_93 = W*in
   wire signed [14:0] m62_93;
   assign m62_93 =15'b0;

   // m62_94 = W*in
   wire signed [14:0] m62_94;
   assign m62_94 =15'b0;

   // m62_95 = W*in
   wire signed [14:0] m62_95;
   assign m62_95 =15'b0;

   // m62_96 = W*in
   wire signed [14:0] m62_96;
   assign m62_96 =15'b0;

   // m62_97 = W*in
   wire signed [14:0] m62_97;
   assign m62_97 =15'b0;

   // m62_98 = W*in
   wire signed [14:0] m62_98;
   assign m62_98 =15'b0;

   // m62_99 = W*in
   wire signed [14:0] m62_99;
   assign m62_99 ={ {3{in62[14]}} , in62[14:3] };

   // m62_100 = W*in
   wire signed [14:0] m62_100;
   assign m62_100 =15'b0;

   // m63_1 = W*in
   wire signed [14:0] m63_1;
   assign m63_1 =15'b0;

   // m63_2 = W*in
   wire signed [14:0] m63_2;
   assign m63_2 =15'b0;

   // m63_3 = W*in
   wire signed [14:0] m63_3;
   assign m63_3 =15'b0;

   // m63_4 = W*in
   wire signed [14:0] m63_4;
   assign m63_4 =15'b0;

   // m63_5 = W*in
   wire signed [14:0] m63_5;
   assign m63_5 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_6 = W*in
   wire signed [14:0] m63_6;
   assign m63_6 ={ {2{in63[14]}} , in63[14:2] };

   // m63_7 = W*in
   wire signed [14:0] m63_7;
   assign m63_7 =15'b0;

   // m63_8 = W*in
   wire signed [14:0] m63_8;
   assign m63_8 =15'b0;

   // m63_9 = W*in
   wire signed [14:0] m63_9;
   assign m63_9 =15'b0;

   // m63_10 = W*in
   wire signed [14:0] m63_10;
   assign m63_10 =15'b0;

   // m63_11 = W*in
   wire signed [14:0] m63_11;
   assign m63_11 =15'b0;

   // m63_12 = W*in
   wire signed [14:0] m63_12;
   assign m63_12 ={ {3{in63[14]}} , in63[14:3] };

   // m63_13 = W*in
   wire signed [14:0] m63_13;
   assign m63_13 =15'b0;

   // m63_14 = W*in
   wire signed [14:0] m63_14;
   assign m63_14 =15'b0;

   // m63_15 = W*in
   wire signed [14:0] m63_15;
   assign m63_15 =15'b0;

   // m63_16 = W*in
   wire signed [14:0] m63_16;
   assign m63_16 =15'b0;

   // m63_17 = W*in
   wire signed [14:0] m63_17;
   assign m63_17 =15'b0;

   // m63_18 = W*in
   wire signed [14:0] m63_18;
   assign m63_18 =15'b0;

   // m63_19 = W*in
   wire signed [14:0] m63_19;
   assign m63_19 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_20 = W*in
   wire signed [14:0] m63_20;
   assign m63_20 =15'b0;

   // m63_21 = W*in
   wire signed [14:0] m63_21;
   assign m63_21 =15'b0;

   // m63_22 = W*in
   wire signed [14:0] m63_22;
   assign m63_22 =15'b0;

   // m63_23 = W*in
   wire signed [14:0] m63_23;
   assign m63_23 =15'b0;

   // m63_24 = W*in
   wire signed [14:0] m63_24;
   assign m63_24 =15'b0;

   // m63_25 = W*in
   wire signed [14:0] m63_25;
   assign m63_25 ={ {4{neg63[14]}} , neg63[14:4] };

   // m63_26 = W*in
   wire signed [14:0] m63_26;
   assign m63_26 ={ {3{in63[14]}} , in63[14:3] };

   // m63_27 = W*in
   wire signed [14:0] m63_27;
   assign m63_27 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_28 = W*in
   wire signed [14:0] m63_28;
   assign m63_28 =15'b0;

   // m63_29 = W*in
   wire signed [14:0] m63_29;
   assign m63_29 ={ {3{in63[14]}} , in63[14:3] };

   // m63_30 = W*in
   wire signed [14:0] m63_30;
   assign m63_30 =15'b0;

   // m63_31 = W*in
   wire signed [14:0] m63_31;
   assign m63_31 ={ {3{in63[14]}} , in63[14:3] };

   // m63_32 = W*in
   wire signed [14:0] m63_32;
   assign m63_32 =15'b0;

   // m63_33 = W*in
   wire signed [14:0] m63_33;
   assign m63_33 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_34 = W*in
   wire signed [14:0] m63_34;
   assign m63_34 ={ {3{in63[14]}} , in63[14:3] };

   // m63_35 = W*in
   wire signed [14:0] m63_35;
   assign m63_35 =15'b0;

   // m63_36 = W*in
   wire signed [14:0] m63_36;
   assign m63_36 =15'b0;

   // m63_37 = W*in
   wire signed [14:0] m63_37;
   assign m63_37 =15'b0;

   // m63_38 = W*in
   wire signed [14:0] m63_38;
   assign m63_38 =15'b0;

   // m63_39 = W*in
   wire signed [14:0] m63_39;
   assign m63_39 =15'b0;

   // m63_40 = W*in
   wire signed [14:0] m63_40;
   assign m63_40 =15'b0;

   // m63_41 = W*in
   wire signed [14:0] m63_41;
   assign m63_41 =15'b0;

   // m63_42 = W*in
   wire signed [14:0] m63_42;
   assign m63_42 =15'b0;

   // m63_43 = W*in
   wire signed [14:0] m63_43;
   assign m63_43 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_44 = W*in
   wire signed [14:0] m63_44;
   assign m63_44 =15'b0;

   // m63_45 = W*in
   wire signed [14:0] m63_45;
   assign m63_45 =15'b0;

   // m63_46 = W*in
   wire signed [14:0] m63_46;
   assign m63_46 =15'b0;

   // m63_47 = W*in
   wire signed [14:0] m63_47;
   assign m63_47 =15'b0;

   // m63_48 = W*in
   wire signed [14:0] m63_48;
   assign m63_48 =15'b0;

   // m63_49 = W*in
   wire signed [14:0] m63_49;
   assign m63_49 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_50 = W*in
   wire signed [14:0] m63_50;
   assign m63_50 =15'b0;

   // m63_51 = W*in
   wire signed [14:0] m63_51;
   assign m63_51 =15'b0;

   // m63_52 = W*in
   wire signed [14:0] m63_52;
   assign m63_52 ={ {3{in63[14]}} , in63[14:3] };

   // m63_53 = W*in
   wire signed [14:0] m63_53;
   assign m63_53 =15'b0;

   // m63_54 = W*in
   wire signed [14:0] m63_54;
   assign m63_54 =15'b0;

   // m63_55 = W*in
   wire signed [14:0] m63_55;
   assign m63_55 =15'b0;

   // m63_56 = W*in
   wire signed [14:0] m63_56;
   assign m63_56 =15'b0;

   // m63_57 = W*in
   wire signed [14:0] m63_57;
   assign m63_57 =15'b0;

   // m63_58 = W*in
   wire signed [14:0] m63_58;
   assign m63_58 =15'b0;

   // m63_59 = W*in
   wire signed [14:0] m63_59;
   assign m63_59 =15'b0;

   // m63_60 = W*in
   wire signed [14:0] m63_60;
   assign m63_60 ={ {2{in63[14]}} , in63[14:2] };

   // m63_61 = W*in
   wire signed [14:0] m63_61;
   assign m63_61 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_62 = W*in
   wire signed [14:0] m63_62;
   assign m63_62 =15'b0;

   // m63_63 = W*in
   wire signed [14:0] m63_63;
   assign m63_63 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_64 = W*in
   wire signed [14:0] m63_64;
   assign m63_64 =15'b0;

   // m63_65 = W*in
   wire signed [14:0] m63_65;
   assign m63_65 =15'b0;

   // m63_66 = W*in
   wire signed [14:0] m63_66;
   assign m63_66 =15'b0;

   // m63_67 = W*in
   wire signed [14:0] m63_67;
   assign m63_67 =15'b0;

   // m63_68 = W*in
   wire signed [14:0] m63_68;
   assign m63_68 =15'b0;

   // m63_69 = W*in
   wire signed [14:0] m63_69;
   assign m63_69 =15'b0;

   // m63_70 = W*in
   wire signed [14:0] m63_70;
   assign m63_70 =15'b0;

   // m63_71 = W*in
   wire signed [14:0] m63_71;
   assign m63_71 =15'b0;

   // m63_72 = W*in
   wire signed [14:0] m63_72;
   assign m63_72 =15'b0;

   // m63_73 = W*in
   wire signed [14:0] m63_73;
   assign m63_73 =15'b0;

   // m63_74 = W*in
   wire signed [14:0] m63_74;
   assign m63_74 ={ {4{neg63[14]}} , neg63[14:4] };

   // m63_75 = W*in
   wire signed [14:0] m63_75;
   assign m63_75 =15'b0;

   // m63_76 = W*in
   wire signed [14:0] m63_76;
   assign m63_76 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_77 = W*in
   wire signed [14:0] m63_77;
   assign m63_77 ={ {3{in63[14]}} , in63[14:3] };

   // m63_78 = W*in
   wire signed [14:0] m63_78;
   assign m63_78 =15'b0;

   // m63_79 = W*in
   wire signed [14:0] m63_79;
   assign m63_79 =15'b0;

   // m63_80 = W*in
   wire signed [14:0] m63_80;
   assign m63_80 ={ {3{in63[14]}} , in63[14:3] };

   // m63_81 = W*in
   wire signed [14:0] m63_81;
   assign m63_81 =15'b0;

   // m63_82 = W*in
   wire signed [14:0] m63_82;
   assign m63_82 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_83 = W*in
   wire signed [14:0] m63_83;
   assign m63_83 =15'b0;

   // m63_84 = W*in
   wire signed [14:0] m63_84;
   assign m63_84 =15'b0;

   // m63_85 = W*in
   wire signed [14:0] m63_85;
   assign m63_85 =15'b0;

   // m63_86 = W*in
   wire signed [14:0] m63_86;
   assign m63_86 =15'b0;

   // m63_87 = W*in
   wire signed [14:0] m63_87;
   assign m63_87 =15'b0;

   // m63_88 = W*in
   wire signed [14:0] m63_88;
   assign m63_88 =15'b0;

   // m63_89 = W*in
   wire signed [14:0] m63_89;
   assign m63_89 =15'b0;

   // m63_90 = W*in
   wire signed [14:0] m63_90;
   assign m63_90 =15'b0;

   // m63_91 = W*in
   wire signed [14:0] m63_91;
   assign m63_91 =15'b0;

   // m63_92 = W*in
   wire signed [14:0] m63_92;
   assign m63_92 =15'b0;

   // m63_93 = W*in
   wire signed [14:0] m63_93;
   assign m63_93 =15'b0;

   // m63_94 = W*in
   wire signed [14:0] m63_94;
   assign m63_94 ={ {3{neg63[14]}} , neg63[14:3] };

   // m63_95 = W*in
   wire signed [14:0] m63_95;
   assign m63_95 =15'b0;

   // m63_96 = W*in
   wire signed [14:0] m63_96;
   assign m63_96 ={ {2{in63[14]}} , in63[14:2] };

   // m63_97 = W*in
   wire signed [14:0] m63_97;
   assign m63_97 =15'b0;

   // m63_98 = W*in
   wire signed [14:0] m63_98;
   assign m63_98 =15'b0;

   // m63_99 = W*in
   wire signed [14:0] m63_99;
   assign m63_99 =15'b0;

   // m63_100 = W*in
   wire signed [14:0] m63_100;
   assign m63_100 =15'b0;

   // m64_1 = W*in
   wire signed [14:0] m64_1;
   assign m64_1 ={ {3{in64[14]}} , in64[14:3] };

   // m64_2 = W*in
   wire signed [14:0] m64_2;
   assign m64_2 =15'b0;

   // m64_3 = W*in
   wire signed [14:0] m64_3;
   assign m64_3 ={ {3{in64[14]}} , in64[14:3] };

   // m64_4 = W*in
   wire signed [14:0] m64_4;
   assign m64_4 ={ {2{in64[14]}} , in64[14:2] };

   // m64_5 = W*in
   wire signed [14:0] m64_5;
   assign m64_5 =15'b0;

   // m64_6 = W*in
   wire signed [14:0] m64_6;
   assign m64_6 ={ {3{in64[14]}} , in64[14:3] };

   // m64_7 = W*in
   wire signed [14:0] m64_7;
   assign m64_7 =15'b0;

   // m64_8 = W*in
   wire signed [14:0] m64_8;
   assign m64_8 ={ {3{in64[14]}} , in64[14:3] };

   // m64_9 = W*in
   wire signed [14:0] m64_9;
   assign m64_9 =15'b0;

   // m64_10 = W*in
   wire signed [14:0] m64_10;
   assign m64_10 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_11 = W*in
   wire signed [14:0] m64_11;
   assign m64_11 =15'b0;

   // m64_12 = W*in
   wire signed [14:0] m64_12;
   assign m64_12 =15'b0;

   // m64_13 = W*in
   wire signed [14:0] m64_13;
   assign m64_13 ={ {3{in64[14]}} , in64[14:3] };

   // m64_14 = W*in
   wire signed [14:0] m64_14;
   assign m64_14 =15'b0;

   // m64_15 = W*in
   wire signed [14:0] m64_15;
   assign m64_15 =15'b0;

   // m64_16 = W*in
   wire signed [14:0] m64_16;
   assign m64_16 =15'b0;

   // m64_17 = W*in
   wire signed [14:0] m64_17;
   assign m64_17 =15'b0;

   // m64_18 = W*in
   wire signed [14:0] m64_18;
   assign m64_18 ={ {3{in64[14]}} , in64[14:3] };

   // m64_19 = W*in
   wire signed [14:0] m64_19;
   assign m64_19 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_20 = W*in
   wire signed [14:0] m64_20;
   assign m64_20 =15'b0;

   // m64_21 = W*in
   wire signed [14:0] m64_21;
   assign m64_21 =15'b0;

   // m64_22 = W*in
   wire signed [14:0] m64_22;
   assign m64_22 =15'b0;

   // m64_23 = W*in
   wire signed [14:0] m64_23;
   assign m64_23 =15'b0;

   // m64_24 = W*in
   wire signed [14:0] m64_24;
   assign m64_24 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_25 = W*in
   wire signed [14:0] m64_25;
   assign m64_25 =15'b0;

   // m64_26 = W*in
   wire signed [14:0] m64_26;
   assign m64_26 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_27 = W*in
   wire signed [14:0] m64_27;
   assign m64_27 =15'b0;

   // m64_28 = W*in
   wire signed [14:0] m64_28;
   assign m64_28 ={ {4{in64[14]}} , in64[14:4] };

   // m64_29 = W*in
   wire signed [14:0] m64_29;
   assign m64_29 ={ {3{in64[14]}} , in64[14:3] };

   // m64_30 = W*in
   wire signed [14:0] m64_30;
   assign m64_30 =15'b0;

   // m64_31 = W*in
   wire signed [14:0] m64_31;
   assign m64_31 =15'b0;

   // m64_32 = W*in
   wire signed [14:0] m64_32;
   assign m64_32 =15'b0;

   // m64_33 = W*in
   wire signed [14:0] m64_33;
   assign m64_33 ={ {4{neg64[14]}} , neg64[14:4] };

   // m64_34 = W*in
   wire signed [14:0] m64_34;
   assign m64_34 ={ {3{in64[14]}} , in64[14:3] };

   // m64_35 = W*in
   wire signed [14:0] m64_35;
   assign m64_35 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_36 = W*in
   wire signed [14:0] m64_36;
   assign m64_36 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_37 = W*in
   wire signed [14:0] m64_37;
   assign m64_37 =15'b0;

   // m64_38 = W*in
   wire signed [14:0] m64_38;
   assign m64_38 =15'b0;

   // m64_39 = W*in
   wire signed [14:0] m64_39;
   assign m64_39 =15'b0;

   // m64_40 = W*in
   wire signed [14:0] m64_40;
   assign m64_40 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_41 = W*in
   wire signed [14:0] m64_41;
   assign m64_41 =15'b0;

   // m64_42 = W*in
   wire signed [14:0] m64_42;
   assign m64_42 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_43 = W*in
   wire signed [14:0] m64_43;
   assign m64_43 =15'b0;

   // m64_44 = W*in
   wire signed [14:0] m64_44;
   assign m64_44 =15'b0;

   // m64_45 = W*in
   wire signed [14:0] m64_45;
   assign m64_45 =15'b0;

   // m64_46 = W*in
   wire signed [14:0] m64_46;
   assign m64_46 =15'b0;

   // m64_47 = W*in
   wire signed [14:0] m64_47;
   assign m64_47 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_48 = W*in
   wire signed [14:0] m64_48;
   assign m64_48 =15'b0;

   // m64_49 = W*in
   wire signed [14:0] m64_49;
   assign m64_49 =15'b0;

   // m64_50 = W*in
   wire signed [14:0] m64_50;
   assign m64_50 =15'b0;

   // m64_51 = W*in
   wire signed [14:0] m64_51;
   assign m64_51 =15'b0;

   // m64_52 = W*in
   wire signed [14:0] m64_52;
   assign m64_52 =15'b0;

   // m64_53 = W*in
   wire signed [14:0] m64_53;
   assign m64_53 =15'b0;

   // m64_54 = W*in
   wire signed [14:0] m64_54;
   assign m64_54 =15'b0;

   // m64_55 = W*in
   wire signed [14:0] m64_55;
   assign m64_55 =15'b0;

   // m64_56 = W*in
   wire signed [14:0] m64_56;
   assign m64_56 =15'b0;

   // m64_57 = W*in
   wire signed [14:0] m64_57;
   assign m64_57 =15'b0;

   // m64_58 = W*in
   wire signed [14:0] m64_58;
   assign m64_58 ={ {3{in64[14]}} , in64[14:3] };

   // m64_59 = W*in
   wire signed [14:0] m64_59;
   assign m64_59 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_60 = W*in
   wire signed [14:0] m64_60;
   assign m64_60 ={ {3{in64[14]}} , in64[14:3] };

   // m64_61 = W*in
   wire signed [14:0] m64_61;
   assign m64_61 =15'b0;

   // m64_62 = W*in
   wire signed [14:0] m64_62;
   assign m64_62 =15'b0;

   // m64_63 = W*in
   wire signed [14:0] m64_63;
   assign m64_63 =15'b0;

   // m64_64 = W*in
   wire signed [14:0] m64_64;
   assign m64_64 =15'b0;

   // m64_65 = W*in
   wire signed [14:0] m64_65;
   assign m64_65 =15'b0;

   // m64_66 = W*in
   wire signed [14:0] m64_66;
   assign m64_66 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_67 = W*in
   wire signed [14:0] m64_67;
   assign m64_67 =15'b0;

   // m64_68 = W*in
   wire signed [14:0] m64_68;
   assign m64_68 ={ {2{in64[14]}} , in64[14:2] };

   // m64_69 = W*in
   wire signed [14:0] m64_69;
   assign m64_69 ={ {3{in64[14]}} , in64[14:3] };

   // m64_70 = W*in
   wire signed [14:0] m64_70;
   assign m64_70 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_71 = W*in
   wire signed [14:0] m64_71;
   assign m64_71 =15'b0;

   // m64_72 = W*in
   wire signed [14:0] m64_72;
   assign m64_72 ={ {3{in64[14]}} , in64[14:3] };

   // m64_73 = W*in
   wire signed [14:0] m64_73;
   assign m64_73 =15'b0;

   // m64_74 = W*in
   wire signed [14:0] m64_74;
   assign m64_74 =15'b0;

   // m64_75 = W*in
   wire signed [14:0] m64_75;
   assign m64_75 =15'b0;

   // m64_76 = W*in
   wire signed [14:0] m64_76;
   assign m64_76 =15'b0;

   // m64_77 = W*in
   wire signed [14:0] m64_77;
   assign m64_77 =15'b0;

   // m64_78 = W*in
   wire signed [14:0] m64_78;
   assign m64_78 ={ {3{in64[14]}} , in64[14:3] };

   // m64_79 = W*in
   wire signed [14:0] m64_79;
   assign m64_79 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_80 = W*in
   wire signed [14:0] m64_80;
   assign m64_80 ={ {3{in64[14]}} , in64[14:3] };

   // m64_81 = W*in
   wire signed [14:0] m64_81;
   assign m64_81 =15'b0;

   // m64_82 = W*in
   wire signed [14:0] m64_82;
   assign m64_82 =15'b0;

   // m64_83 = W*in
   wire signed [14:0] m64_83;
   assign m64_83 =15'b0;

   // m64_84 = W*in
   wire signed [14:0] m64_84;
   assign m64_84 =15'b0;

   // m64_85 = W*in
   wire signed [14:0] m64_85;
   assign m64_85 =15'b0;

   // m64_86 = W*in
   wire signed [14:0] m64_86;
   assign m64_86 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_87 = W*in
   wire signed [14:0] m64_87;
   assign m64_87 =15'b0;

   // m64_88 = W*in
   wire signed [14:0] m64_88;
   assign m64_88 =15'b0;

   // m64_89 = W*in
   wire signed [14:0] m64_89;
   assign m64_89 =15'b0;

   // m64_90 = W*in
   wire signed [14:0] m64_90;
   assign m64_90 =15'b0;

   // m64_91 = W*in
   wire signed [14:0] m64_91;
   assign m64_91 =15'b0;

   // m64_92 = W*in
   wire signed [14:0] m64_92;
   assign m64_92 =15'b0;

   // m64_93 = W*in
   wire signed [14:0] m64_93;
   assign m64_93 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_94 = W*in
   wire signed [14:0] m64_94;
   assign m64_94 ={ {3{neg64[14]}} , neg64[14:3] };

   // m64_95 = W*in
   wire signed [14:0] m64_95;
   assign m64_95 =15'b0;

   // m64_96 = W*in
   wire signed [14:0] m64_96;
   assign m64_96 ={ {3{in64[14]}} , in64[14:3] };

   // m64_97 = W*in
   wire signed [14:0] m64_97;
   assign m64_97 =15'b0;

   // m64_98 = W*in
   wire signed [14:0] m64_98;
   assign m64_98 =15'b0;

   // m64_99 = W*in
   wire signed [14:0] m64_99;
   assign m64_99 =15'b0;

   // m64_100 = W*in
   wire signed [14:0] m64_100;
   assign m64_100 =15'b0;

   // m65_1 = W*in
   wire signed [14:0] m65_1;
   assign m65_1 =15'b0;

   // m65_2 = W*in
   wire signed [14:0] m65_2;
   assign m65_2 =15'b0;

   // m65_3 = W*in
   wire signed [14:0] m65_3;
   assign m65_3 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_4 = W*in
   wire signed [14:0] m65_4;
   assign m65_4 ={ {3{in65[14]}} , in65[14:3] };

   // m65_5 = W*in
   wire signed [14:0] m65_5;
   assign m65_5 =15'b0;

   // m65_6 = W*in
   wire signed [14:0] m65_6;
   assign m65_6 =15'b0;

   // m65_7 = W*in
   wire signed [14:0] m65_7;
   assign m65_7 =15'b0;

   // m65_8 = W*in
   wire signed [14:0] m65_8;
   assign m65_8 =15'b0;

   // m65_9 = W*in
   wire signed [14:0] m65_9;
   assign m65_9 =15'b0;

   // m65_10 = W*in
   wire signed [14:0] m65_10;
   assign m65_10 =15'b0;

   // m65_11 = W*in
   wire signed [14:0] m65_11;
   assign m65_11 =15'b0;

   // m65_12 = W*in
   wire signed [14:0] m65_12;
   assign m65_12 =15'b0;

   // m65_13 = W*in
   wire signed [14:0] m65_13;
   assign m65_13 =15'b0;

   // m65_14 = W*in
   wire signed [14:0] m65_14;
   assign m65_14 =15'b0;

   // m65_15 = W*in
   wire signed [14:0] m65_15;
   assign m65_15 =15'b0;

   // m65_16 = W*in
   wire signed [14:0] m65_16;
   assign m65_16 =15'b0;

   // m65_17 = W*in
   wire signed [14:0] m65_17;
   assign m65_17 =15'b0;

   // m65_18 = W*in
   wire signed [14:0] m65_18;
   assign m65_18 ={ {3{in65[14]}} , in65[14:3] };

   // m65_19 = W*in
   wire signed [14:0] m65_19;
   assign m65_19 =15'b0;

   // m65_20 = W*in
   wire signed [14:0] m65_20;
   assign m65_20 =15'b0;

   // m65_21 = W*in
   wire signed [14:0] m65_21;
   assign m65_21 =15'b0;

   // m65_22 = W*in
   wire signed [14:0] m65_22;
   assign m65_22 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_23 = W*in
   wire signed [14:0] m65_23;
   assign m65_23 =15'b0;

   // m65_24 = W*in
   wire signed [14:0] m65_24;
   assign m65_24 =15'b0;

   // m65_25 = W*in
   wire signed [14:0] m65_25;
   assign m65_25 =15'b0;

   // m65_26 = W*in
   wire signed [14:0] m65_26;
   assign m65_26 =15'b0;

   // m65_27 = W*in
   wire signed [14:0] m65_27;
   assign m65_27 =15'b0;

   // m65_28 = W*in
   wire signed [14:0] m65_28;
   assign m65_28 =15'b0;

   // m65_29 = W*in
   wire signed [14:0] m65_29;
   assign m65_29 =15'b0;

   // m65_30 = W*in
   wire signed [14:0] m65_30;
   assign m65_30 =15'b0;

   // m65_31 = W*in
   wire signed [14:0] m65_31;
   assign m65_31 ={ {3{in65[14]}} , in65[14:3] };

   // m65_32 = W*in
   wire signed [14:0] m65_32;
   assign m65_32 =15'b0;

   // m65_33 = W*in
   wire signed [14:0] m65_33;
   assign m65_33 =15'b0;

   // m65_34 = W*in
   wire signed [14:0] m65_34;
   assign m65_34 =15'b0;

   // m65_35 = W*in
   wire signed [14:0] m65_35;
   assign m65_35 =15'b0;

   // m65_36 = W*in
   wire signed [14:0] m65_36;
   assign m65_36 =15'b0;

   // m65_37 = W*in
   wire signed [14:0] m65_37;
   assign m65_37 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_38 = W*in
   wire signed [14:0] m65_38;
   assign m65_38 =15'b0;

   // m65_39 = W*in
   wire signed [14:0] m65_39;
   assign m65_39 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_40 = W*in
   wire signed [14:0] m65_40;
   assign m65_40 =15'b0;

   // m65_41 = W*in
   wire signed [14:0] m65_41;
   assign m65_41 ={ {3{in65[14]}} , in65[14:3] };

   // m65_42 = W*in
   wire signed [14:0] m65_42;
   assign m65_42 =15'b0;

   // m65_43 = W*in
   wire signed [14:0] m65_43;
   assign m65_43 =15'b0;

   // m65_44 = W*in
   wire signed [14:0] m65_44;
   assign m65_44 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_45 = W*in
   wire signed [14:0] m65_45;
   assign m65_45 =15'b0;

   // m65_46 = W*in
   wire signed [14:0] m65_46;
   assign m65_46 =15'b0;

   // m65_47 = W*in
   wire signed [14:0] m65_47;
   assign m65_47 =15'b0;

   // m65_48 = W*in
   wire signed [14:0] m65_48;
   assign m65_48 =15'b0;

   // m65_49 = W*in
   wire signed [14:0] m65_49;
   assign m65_49 =15'b0;

   // m65_50 = W*in
   wire signed [14:0] m65_50;
   assign m65_50 =15'b0;

   // m65_51 = W*in
   wire signed [14:0] m65_51;
   assign m65_51 =15'b0;

   // m65_52 = W*in
   wire signed [14:0] m65_52;
   assign m65_52 ={ {3{in65[14]}} , in65[14:3] };

   // m65_53 = W*in
   wire signed [14:0] m65_53;
   assign m65_53 =15'b0;

   // m65_54 = W*in
   wire signed [14:0] m65_54;
   assign m65_54 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_55 = W*in
   wire signed [14:0] m65_55;
   assign m65_55 =15'b0;

   // m65_56 = W*in
   wire signed [14:0] m65_56;
   assign m65_56 =15'b0;

   // m65_57 = W*in
   wire signed [14:0] m65_57;
   assign m65_57 =15'b0;

   // m65_58 = W*in
   wire signed [14:0] m65_58;
   assign m65_58 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_59 = W*in
   wire signed [14:0] m65_59;
   assign m65_59 ={ {4{neg65[14]}} , neg65[14:4] };

   // m65_60 = W*in
   wire signed [14:0] m65_60;
   assign m65_60 =15'b0;

   // m65_61 = W*in
   wire signed [14:0] m65_61;
   assign m65_61 ={ {4{in65[14]}} , in65[14:4] };

   // m65_62 = W*in
   wire signed [14:0] m65_62;
   assign m65_62 =15'b0;

   // m65_63 = W*in
   wire signed [14:0] m65_63;
   assign m65_63 =15'b0;

   // m65_64 = W*in
   wire signed [14:0] m65_64;
   assign m65_64 =15'b0;

   // m65_65 = W*in
   wire signed [14:0] m65_65;
   assign m65_65 =15'b0;

   // m65_66 = W*in
   wire signed [14:0] m65_66;
   assign m65_66 =15'b0;

   // m65_67 = W*in
   wire signed [14:0] m65_67;
   assign m65_67 =15'b0;

   // m65_68 = W*in
   wire signed [14:0] m65_68;
   assign m65_68 =15'b0;

   // m65_69 = W*in
   wire signed [14:0] m65_69;
   assign m65_69 ={ {4{neg65[14]}} , neg65[14:4] };

   // m65_70 = W*in
   wire signed [14:0] m65_70;
   assign m65_70 =15'b0;

   // m65_71 = W*in
   wire signed [14:0] m65_71;
   assign m65_71 =15'b0;

   // m65_72 = W*in
   wire signed [14:0] m65_72;
   assign m65_72 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_73 = W*in
   wire signed [14:0] m65_73;
   assign m65_73 =15'b0;

   // m65_74 = W*in
   wire signed [14:0] m65_74;
   assign m65_74 ={ {4{neg65[14]}} , neg65[14:4] };

   // m65_75 = W*in
   wire signed [14:0] m65_75;
   assign m65_75 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_76 = W*in
   wire signed [14:0] m65_76;
   assign m65_76 =15'b0;

   // m65_77 = W*in
   wire signed [14:0] m65_77;
   assign m65_77 =15'b0;

   // m65_78 = W*in
   wire signed [14:0] m65_78;
   assign m65_78 ={ {3{in65[14]}} , in65[14:3] };

   // m65_79 = W*in
   wire signed [14:0] m65_79;
   assign m65_79 =15'b0;

   // m65_80 = W*in
   wire signed [14:0] m65_80;
   assign m65_80 =15'b0;

   // m65_81 = W*in
   wire signed [14:0] m65_81;
   assign m65_81 =15'b0;

   // m65_82 = W*in
   wire signed [14:0] m65_82;
   assign m65_82 =15'b0;

   // m65_83 = W*in
   wire signed [14:0] m65_83;
   assign m65_83 =15'b0;

   // m65_84 = W*in
   wire signed [14:0] m65_84;
   assign m65_84 =15'b0;

   // m65_85 = W*in
   wire signed [14:0] m65_85;
   assign m65_85 =15'b0;

   // m65_86 = W*in
   wire signed [14:0] m65_86;
   assign m65_86 =15'b0;

   // m65_87 = W*in
   wire signed [14:0] m65_87;
   assign m65_87 =15'b0;

   // m65_88 = W*in
   wire signed [14:0] m65_88;
   assign m65_88 =15'b0;

   // m65_89 = W*in
   wire signed [14:0] m65_89;
   assign m65_89 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_90 = W*in
   wire signed [14:0] m65_90;
   assign m65_90 =15'b0;

   // m65_91 = W*in
   wire signed [14:0] m65_91;
   assign m65_91 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_92 = W*in
   wire signed [14:0] m65_92;
   assign m65_92 =15'b0;

   // m65_93 = W*in
   wire signed [14:0] m65_93;
   assign m65_93 ={ {3{neg65[14]}} , neg65[14:3] };

   // m65_94 = W*in
   wire signed [14:0] m65_94;
   assign m65_94 =15'b0;

   // m65_95 = W*in
   wire signed [14:0] m65_95;
   assign m65_95 ={ {4{neg65[14]}} , neg65[14:4] };

   // m65_96 = W*in
   wire signed [14:0] m65_96;
   assign m65_96 =15'b0;

   // m65_97 = W*in
   wire signed [14:0] m65_97;
   assign m65_97 =15'b0;

   // m65_98 = W*in
   wire signed [14:0] m65_98;
   assign m65_98 =15'b0;

   // m65_99 = W*in
   wire signed [14:0] m65_99;
   assign m65_99 =15'b0;

   // m65_100 = W*in
   wire signed [14:0] m65_100;
   assign m65_100 =15'b0;

   // m66_1 = W*in
   wire signed [14:0] m66_1;
   assign m66_1 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_2 = W*in
   wire signed [14:0] m66_2;
   assign m66_2 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_3 = W*in
   wire signed [14:0] m66_3;
   assign m66_3 =15'b0;

   // m66_4 = W*in
   wire signed [14:0] m66_4;
   assign m66_4 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_5 = W*in
   wire signed [14:0] m66_5;
   assign m66_5 =15'b0;

   // m66_6 = W*in
   wire signed [14:0] m66_6;
   assign m66_6 =15'b0;

   // m66_7 = W*in
   wire signed [14:0] m66_7;
   assign m66_7 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_8 = W*in
   wire signed [14:0] m66_8;
   assign m66_8 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_9 = W*in
   wire signed [14:0] m66_9;
   assign m66_9 =15'b0;

   // m66_10 = W*in
   wire signed [14:0] m66_10;
   assign m66_10 =15'b0;

   // m66_11 = W*in
   wire signed [14:0] m66_11;
   assign m66_11 =15'b0;

   // m66_12 = W*in
   wire signed [14:0] m66_12;
   assign m66_12 =15'b0;

   // m66_13 = W*in
   wire signed [14:0] m66_13;
   assign m66_13 =15'b0;

   // m66_14 = W*in
   wire signed [14:0] m66_14;
   assign m66_14 =15'b0;

   // m66_15 = W*in
   wire signed [14:0] m66_15;
   assign m66_15 ={ {3{in66[14]}} , in66[14:3] };

   // m66_16 = W*in
   wire signed [14:0] m66_16;
   assign m66_16 =15'b0;

   // m66_17 = W*in
   wire signed [14:0] m66_17;
   assign m66_17 ={ {3{in66[14]}} , in66[14:3] };

   // m66_18 = W*in
   wire signed [14:0] m66_18;
   assign m66_18 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_19 = W*in
   wire signed [14:0] m66_19;
   assign m66_19 =15'b0;

   // m66_20 = W*in
   wire signed [14:0] m66_20;
   assign m66_20 =15'b0;

   // m66_21 = W*in
   wire signed [14:0] m66_21;
   assign m66_21 ={ {4{neg66[14]}} , neg66[14:4] };

   // m66_22 = W*in
   wire signed [14:0] m66_22;
   assign m66_22 =15'b0;

   // m66_23 = W*in
   wire signed [14:0] m66_23;
   assign m66_23 =15'b0;

   // m66_24 = W*in
   wire signed [14:0] m66_24;
   assign m66_24 =15'b0;

   // m66_25 = W*in
   wire signed [14:0] m66_25;
   assign m66_25 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_26 = W*in
   wire signed [14:0] m66_26;
   assign m66_26 =15'b0;

   // m66_27 = W*in
   wire signed [14:0] m66_27;
   assign m66_27 =15'b0;

   // m66_28 = W*in
   wire signed [14:0] m66_28;
   assign m66_28 =15'b0;

   // m66_29 = W*in
   wire signed [14:0] m66_29;
   assign m66_29 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_30 = W*in
   wire signed [14:0] m66_30;
   assign m66_30 =15'b0;

   // m66_31 = W*in
   wire signed [14:0] m66_31;
   assign m66_31 ={ {4{neg66[14]}} , neg66[14:4] };

   // m66_32 = W*in
   wire signed [14:0] m66_32;
   assign m66_32 ={ {4{neg66[14]}} , neg66[14:4] };

   // m66_33 = W*in
   wire signed [14:0] m66_33;
   assign m66_33 =15'b0;

   // m66_34 = W*in
   wire signed [14:0] m66_34;
   assign m66_34 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_35 = W*in
   wire signed [14:0] m66_35;
   assign m66_35 =15'b0;

   // m66_36 = W*in
   wire signed [14:0] m66_36;
   assign m66_36 =15'b0;

   // m66_37 = W*in
   wire signed [14:0] m66_37;
   assign m66_37 =15'b0;

   // m66_38 = W*in
   wire signed [14:0] m66_38;
   assign m66_38 =15'b0;

   // m66_39 = W*in
   wire signed [14:0] m66_39;
   assign m66_39 =15'b0;

   // m66_40 = W*in
   wire signed [14:0] m66_40;
   assign m66_40 =15'b0;

   // m66_41 = W*in
   wire signed [14:0] m66_41;
   assign m66_41 =15'b0;

   // m66_42 = W*in
   wire signed [14:0] m66_42;
   assign m66_42 =15'b0;

   // m66_43 = W*in
   wire signed [14:0] m66_43;
   assign m66_43 =15'b0;

   // m66_44 = W*in
   wire signed [14:0] m66_44;
   assign m66_44 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_45 = W*in
   wire signed [14:0] m66_45;
   assign m66_45 =15'b0;

   // m66_46 = W*in
   wire signed [14:0] m66_46;
   assign m66_46 =15'b0;

   // m66_47 = W*in
   wire signed [14:0] m66_47;
   assign m66_47 =15'b0;

   // m66_48 = W*in
   wire signed [14:0] m66_48;
   assign m66_48 =15'b0;

   // m66_49 = W*in
   wire signed [14:0] m66_49;
   assign m66_49 =15'b0;

   // m66_50 = W*in
   wire signed [14:0] m66_50;
   assign m66_50 =15'b0;

   // m66_51 = W*in
   wire signed [14:0] m66_51;
   assign m66_51 =15'b0;

   // m66_52 = W*in
   wire signed [14:0] m66_52;
   assign m66_52 =15'b0;

   // m66_53 = W*in
   wire signed [14:0] m66_53;
   assign m66_53 =15'b0;

   // m66_54 = W*in
   wire signed [14:0] m66_54;
   assign m66_54 =15'b0;

   // m66_55 = W*in
   wire signed [14:0] m66_55;
   assign m66_55 =15'b0;

   // m66_56 = W*in
   wire signed [14:0] m66_56;
   assign m66_56 ={ {2{in66[14]}} , in66[14:2] };

   // m66_57 = W*in
   wire signed [14:0] m66_57;
   assign m66_57 ={ {4{in66[14]}} , in66[14:4] };

   // m66_58 = W*in
   wire signed [14:0] m66_58;
   assign m66_58 ={ {4{in66[14]}} , in66[14:4] };

   // m66_59 = W*in
   wire signed [14:0] m66_59;
   assign m66_59 ={ {3{in66[14]}} , in66[14:3] };

   // m66_60 = W*in
   wire signed [14:0] m66_60;
   assign m66_60 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_61 = W*in
   wire signed [14:0] m66_61;
   assign m66_61 ={ {3{in66[14]}} , in66[14:3] };

   // m66_62 = W*in
   wire signed [14:0] m66_62;
   assign m66_62 ={ {3{in66[14]}} , in66[14:3] };

   // m66_63 = W*in
   wire signed [14:0] m66_63;
   assign m66_63 =15'b0;

   // m66_64 = W*in
   wire signed [14:0] m66_64;
   assign m66_64 ={ {3{in66[14]}} , in66[14:3] };

   // m66_65 = W*in
   wire signed [14:0] m66_65;
   assign m66_65 =15'b0;

   // m66_66 = W*in
   wire signed [14:0] m66_66;
   assign m66_66 ={ {4{neg66[14]}} , neg66[14:4] };

   // m66_67 = W*in
   wire signed [14:0] m66_67;
   assign m66_67 =15'b0;

   // m66_68 = W*in
   wire signed [14:0] m66_68;
   assign m66_68 =15'b0;

   // m66_69 = W*in
   wire signed [14:0] m66_69;
   assign m66_69 ={ {4{neg66[14]}} , neg66[14:4] };

   // m66_70 = W*in
   wire signed [14:0] m66_70;
   assign m66_70 ={ {3{in66[14]}} , in66[14:3] };

   // m66_71 = W*in
   wire signed [14:0] m66_71;
   assign m66_71 =15'b0;

   // m66_72 = W*in
   wire signed [14:0] m66_72;
   assign m66_72 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_73 = W*in
   wire signed [14:0] m66_73;
   assign m66_73 =15'b0;

   // m66_74 = W*in
   wire signed [14:0] m66_74;
   assign m66_74 ={ {4{in66[14]}} , in66[14:4] };

   // m66_75 = W*in
   wire signed [14:0] m66_75;
   assign m66_75 ={ {4{in66[14]}} , in66[14:4] };

   // m66_76 = W*in
   wire signed [14:0] m66_76;
   assign m66_76 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_77 = W*in
   wire signed [14:0] m66_77;
   assign m66_77 =15'b0;

   // m66_78 = W*in
   wire signed [14:0] m66_78;
   assign m66_78 =15'b0;

   // m66_79 = W*in
   wire signed [14:0] m66_79;
   assign m66_79 =15'b0;

   // m66_80 = W*in
   wire signed [14:0] m66_80;
   assign m66_80 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_81 = W*in
   wire signed [14:0] m66_81;
   assign m66_81 ={ {3{in66[14]}} , in66[14:3] };

   // m66_82 = W*in
   wire signed [14:0] m66_82;
   assign m66_82 =15'b0;

   // m66_83 = W*in
   wire signed [14:0] m66_83;
   assign m66_83 =15'b0;

   // m66_84 = W*in
   wire signed [14:0] m66_84;
   assign m66_84 =15'b0;

   // m66_85 = W*in
   wire signed [14:0] m66_85;
   assign m66_85 =15'b0;

   // m66_86 = W*in
   wire signed [14:0] m66_86;
   assign m66_86 =15'b0;

   // m66_87 = W*in
   wire signed [14:0] m66_87;
   assign m66_87 =15'b0;

   // m66_88 = W*in
   wire signed [14:0] m66_88;
   assign m66_88 =15'b0;

   // m66_89 = W*in
   wire signed [14:0] m66_89;
   assign m66_89 =15'b0;

   // m66_90 = W*in
   wire signed [14:0] m66_90;
   assign m66_90 =15'b0;

   // m66_91 = W*in
   wire signed [14:0] m66_91;
   assign m66_91 =15'b0;

   // m66_92 = W*in
   wire signed [14:0] m66_92;
   assign m66_92 ={ {3{in66[14]}} , in66[14:3] };

   // m66_93 = W*in
   wire signed [14:0] m66_93;
   assign m66_93 =15'b0;

   // m66_94 = W*in
   wire signed [14:0] m66_94;
   assign m66_94 =15'b0;

   // m66_95 = W*in
   wire signed [14:0] m66_95;
   assign m66_95 =15'b0;

   // m66_96 = W*in
   wire signed [14:0] m66_96;
   assign m66_96 ={ {3{neg66[14]}} , neg66[14:3] };

   // m66_97 = W*in
   wire signed [14:0] m66_97;
   assign m66_97 =15'b0;

   // m66_98 = W*in
   wire signed [14:0] m66_98;
   assign m66_98 =15'b0;

   // m66_99 = W*in
   wire signed [14:0] m66_99;
   assign m66_99 =15'b0;

   // m66_100 = W*in
   wire signed [14:0] m66_100;
   assign m66_100 =15'b0;

   // m67_1 = W*in
   wire signed [14:0] m67_1;
   assign m67_1 ={ {3{in67[14]}} , in67[14:3] };

   // m67_2 = W*in
   wire signed [14:0] m67_2;
   assign m67_2 ={ {3{in67[14]}} , in67[14:3] };

   // m67_3 = W*in
   wire signed [14:0] m67_3;
   assign m67_3 =15'b0;

   // m67_4 = W*in
   wire signed [14:0] m67_4;
   assign m67_4 =15'b0;

   // m67_5 = W*in
   wire signed [14:0] m67_5;
   assign m67_5 =15'b0;

   // m67_6 = W*in
   wire signed [14:0] m67_6;
   assign m67_6 =15'b0;

   // m67_7 = W*in
   wire signed [14:0] m67_7;
   assign m67_7 =15'b0;

   // m67_8 = W*in
   wire signed [14:0] m67_8;
   assign m67_8 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_9 = W*in
   wire signed [14:0] m67_9;
   assign m67_9 ={ {3{in67[14]}} , in67[14:3] };

   // m67_10 = W*in
   wire signed [14:0] m67_10;
   assign m67_10 =15'b0;

   // m67_11 = W*in
   wire signed [14:0] m67_11;
   assign m67_11 =15'b0;

   // m67_12 = W*in
   wire signed [14:0] m67_12;
   assign m67_12 =15'b0;

   // m67_13 = W*in
   wire signed [14:0] m67_13;
   assign m67_13 ={ {3{in67[14]}} , in67[14:3] };

   // m67_14 = W*in
   wire signed [14:0] m67_14;
   assign m67_14 =15'b0;

   // m67_15 = W*in
   wire signed [14:0] m67_15;
   assign m67_15 =15'b0;

   // m67_16 = W*in
   wire signed [14:0] m67_16;
   assign m67_16 =15'b0;

   // m67_17 = W*in
   wire signed [14:0] m67_17;
   assign m67_17 =15'b0;

   // m67_18 = W*in
   wire signed [14:0] m67_18;
   assign m67_18 =15'b0;

   // m67_19 = W*in
   wire signed [14:0] m67_19;
   assign m67_19 =15'b0;

   // m67_20 = W*in
   wire signed [14:0] m67_20;
   assign m67_20 =15'b0;

   // m67_21 = W*in
   wire signed [14:0] m67_21;
   assign m67_21 =15'b0;

   // m67_22 = W*in
   wire signed [14:0] m67_22;
   assign m67_22 =15'b0;

   // m67_23 = W*in
   wire signed [14:0] m67_23;
   assign m67_23 =15'b0;

   // m67_24 = W*in
   wire signed [14:0] m67_24;
   assign m67_24 =15'b0;

   // m67_25 = W*in
   wire signed [14:0] m67_25;
   assign m67_25 =15'b0;

   // m67_26 = W*in
   wire signed [14:0] m67_26;
   assign m67_26 ={ {3{in67[14]}} , in67[14:3] };

   // m67_27 = W*in
   wire signed [14:0] m67_27;
   assign m67_27 ={ {3{in67[14]}} , in67[14:3] };

   // m67_28 = W*in
   wire signed [14:0] m67_28;
   assign m67_28 =15'b0;

   // m67_29 = W*in
   wire signed [14:0] m67_29;
   assign m67_29 =15'b0;

   // m67_30 = W*in
   wire signed [14:0] m67_30;
   assign m67_30 =15'b0;

   // m67_31 = W*in
   wire signed [14:0] m67_31;
   assign m67_31 =15'b0;

   // m67_32 = W*in
   wire signed [14:0] m67_32;
   assign m67_32 =15'b0;

   // m67_33 = W*in
   wire signed [14:0] m67_33;
   assign m67_33 ={ {3{in67[14]}} , in67[14:3] };

   // m67_34 = W*in
   wire signed [14:0] m67_34;
   assign m67_34 =15'b0;

   // m67_35 = W*in
   wire signed [14:0] m67_35;
   assign m67_35 =15'b0;

   // m67_36 = W*in
   wire signed [14:0] m67_36;
   assign m67_36 =15'b0;

   // m67_37 = W*in
   wire signed [14:0] m67_37;
   assign m67_37 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_38 = W*in
   wire signed [14:0] m67_38;
   assign m67_38 ={ {3{in67[14]}} , in67[14:3] };

   // m67_39 = W*in
   wire signed [14:0] m67_39;
   assign m67_39 =15'b0;

   // m67_40 = W*in
   wire signed [14:0] m67_40;
   assign m67_40 ={ {3{in67[14]}} , in67[14:3] };

   // m67_41 = W*in
   wire signed [14:0] m67_41;
   assign m67_41 =15'b0;

   // m67_42 = W*in
   wire signed [14:0] m67_42;
   assign m67_42 ={ {3{in67[14]}} , in67[14:3] };

   // m67_43 = W*in
   wire signed [14:0] m67_43;
   assign m67_43 =15'b0;

   // m67_44 = W*in
   wire signed [14:0] m67_44;
   assign m67_44 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_45 = W*in
   wire signed [14:0] m67_45;
   assign m67_45 =15'b0;

   // m67_46 = W*in
   wire signed [14:0] m67_46;
   assign m67_46 =15'b0;

   // m67_47 = W*in
   wire signed [14:0] m67_47;
   assign m67_47 =15'b0;

   // m67_48 = W*in
   wire signed [14:0] m67_48;
   assign m67_48 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_49 = W*in
   wire signed [14:0] m67_49;
   assign m67_49 =15'b0;

   // m67_50 = W*in
   wire signed [14:0] m67_50;
   assign m67_50 =15'b0;

   // m67_51 = W*in
   wire signed [14:0] m67_51;
   assign m67_51 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_52 = W*in
   wire signed [14:0] m67_52;
   assign m67_52 =15'b0;

   // m67_53 = W*in
   wire signed [14:0] m67_53;
   assign m67_53 =15'b0;

   // m67_54 = W*in
   wire signed [14:0] m67_54;
   assign m67_54 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_55 = W*in
   wire signed [14:0] m67_55;
   assign m67_55 =15'b0;

   // m67_56 = W*in
   wire signed [14:0] m67_56;
   assign m67_56 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_57 = W*in
   wire signed [14:0] m67_57;
   assign m67_57 =15'b0;

   // m67_58 = W*in
   wire signed [14:0] m67_58;
   assign m67_58 =15'b0;

   // m67_59 = W*in
   wire signed [14:0] m67_59;
   assign m67_59 ={ {4{neg67[14]}} , neg67[14:4] };

   // m67_60 = W*in
   wire signed [14:0] m67_60;
   assign m67_60 =15'b0;

   // m67_61 = W*in
   wire signed [14:0] m67_61;
   assign m67_61 =15'b0;

   // m67_62 = W*in
   wire signed [14:0] m67_62;
   assign m67_62 =15'b0;

   // m67_63 = W*in
   wire signed [14:0] m67_63;
   assign m67_63 =15'b0;

   // m67_64 = W*in
   wire signed [14:0] m67_64;
   assign m67_64 =15'b0;

   // m67_65 = W*in
   wire signed [14:0] m67_65;
   assign m67_65 =15'b0;

   // m67_66 = W*in
   wire signed [14:0] m67_66;
   assign m67_66 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_67 = W*in
   wire signed [14:0] m67_67;
   assign m67_67 =15'b0;

   // m67_68 = W*in
   wire signed [14:0] m67_68;
   assign m67_68 =15'b0;

   // m67_69 = W*in
   wire signed [14:0] m67_69;
   assign m67_69 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_70 = W*in
   wire signed [14:0] m67_70;
   assign m67_70 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_71 = W*in
   wire signed [14:0] m67_71;
   assign m67_71 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_72 = W*in
   wire signed [14:0] m67_72;
   assign m67_72 =15'b0;

   // m67_73 = W*in
   wire signed [14:0] m67_73;
   assign m67_73 =15'b0;

   // m67_74 = W*in
   wire signed [14:0] m67_74;
   assign m67_74 =15'b0;

   // m67_75 = W*in
   wire signed [14:0] m67_75;
   assign m67_75 =15'b0;

   // m67_76 = W*in
   wire signed [14:0] m67_76;
   assign m67_76 =15'b0;

   // m67_77 = W*in
   wire signed [14:0] m67_77;
   assign m67_77 =15'b0;

   // m67_78 = W*in
   wire signed [14:0] m67_78;
   assign m67_78 =15'b0;

   // m67_79 = W*in
   wire signed [14:0] m67_79;
   assign m67_79 =15'b0;

   // m67_80 = W*in
   wire signed [14:0] m67_80;
   assign m67_80 =15'b0;

   // m67_81 = W*in
   wire signed [14:0] m67_81;
   assign m67_81 =15'b0;

   // m67_82 = W*in
   wire signed [14:0] m67_82;
   assign m67_82 =15'b0;

   // m67_83 = W*in
   wire signed [14:0] m67_83;
   assign m67_83 =15'b0;

   // m67_84 = W*in
   wire signed [14:0] m67_84;
   assign m67_84 =15'b0;

   // m67_85 = W*in
   wire signed [14:0] m67_85;
   assign m67_85 =15'b0;

   // m67_86 = W*in
   wire signed [14:0] m67_86;
   assign m67_86 =15'b0;

   // m67_87 = W*in
   wire signed [14:0] m67_87;
   assign m67_87 =15'b0;

   // m67_88 = W*in
   wire signed [14:0] m67_88;
   assign m67_88 =15'b0;

   // m67_89 = W*in
   wire signed [14:0] m67_89;
   assign m67_89 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_90 = W*in
   wire signed [14:0] m67_90;
   assign m67_90 =15'b0;

   // m67_91 = W*in
   wire signed [14:0] m67_91;
   assign m67_91 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_92 = W*in
   wire signed [14:0] m67_92;
   assign m67_92 =15'b0;

   // m67_93 = W*in
   wire signed [14:0] m67_93;
   assign m67_93 ={ {3{neg67[14]}} , neg67[14:3] };

   // m67_94 = W*in
   wire signed [14:0] m67_94;
   assign m67_94 =15'b0;

   // m67_95 = W*in
   wire signed [14:0] m67_95;
   assign m67_95 =15'b0;

   // m67_96 = W*in
   wire signed [14:0] m67_96;
   assign m67_96 =15'b0;

   // m67_97 = W*in
   wire signed [14:0] m67_97;
   assign m67_97 =15'b0;

   // m67_98 = W*in
   wire signed [14:0] m67_98;
   assign m67_98 =15'b0;

   // m67_99 = W*in
   wire signed [14:0] m67_99;
   assign m67_99 =15'b0;

   // m67_100 = W*in
   wire signed [14:0] m67_100;
   assign m67_100 ={ {3{neg67[14]}} , neg67[14:3] };

   // m68_1 = W*in
   wire signed [14:0] m68_1;
   assign m68_1 =15'b0;

   // m68_2 = W*in
   wire signed [14:0] m68_2;
   assign m68_2 ={ {3{in68[14]}} , in68[14:3] };

   // m68_3 = W*in
   wire signed [14:0] m68_3;
   assign m68_3 =15'b0;

   // m68_4 = W*in
   wire signed [14:0] m68_4;
   assign m68_4 =15'b0;

   // m68_5 = W*in
   wire signed [14:0] m68_5;
   assign m68_5 =15'b0;

   // m68_6 = W*in
   wire signed [14:0] m68_6;
   assign m68_6 ={ {4{neg68[14]}} , neg68[14:4] };

   // m68_7 = W*in
   wire signed [14:0] m68_7;
   assign m68_7 =15'b0;

   // m68_8 = W*in
   wire signed [14:0] m68_8;
   assign m68_8 =15'b0;

   // m68_9 = W*in
   wire signed [14:0] m68_9;
   assign m68_9 =15'b0;

   // m68_10 = W*in
   wire signed [14:0] m68_10;
   assign m68_10 =15'b0;

   // m68_11 = W*in
   wire signed [14:0] m68_11;
   assign m68_11 =15'b0;

   // m68_12 = W*in
   wire signed [14:0] m68_12;
   assign m68_12 =15'b0;

   // m68_13 = W*in
   wire signed [14:0] m68_13;
   assign m68_13 ={ {3{in68[14]}} , in68[14:3] };

   // m68_14 = W*in
   wire signed [14:0] m68_14;
   assign m68_14 =15'b0;

   // m68_15 = W*in
   wire signed [14:0] m68_15;
   assign m68_15 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_16 = W*in
   wire signed [14:0] m68_16;
   assign m68_16 =15'b0;

   // m68_17 = W*in
   wire signed [14:0] m68_17;
   assign m68_17 =15'b0;

   // m68_18 = W*in
   wire signed [14:0] m68_18;
   assign m68_18 ={ {3{in68[14]}} , in68[14:3] };

   // m68_19 = W*in
   wire signed [14:0] m68_19;
   assign m68_19 =15'b0;

   // m68_20 = W*in
   wire signed [14:0] m68_20;
   assign m68_20 =15'b0;

   // m68_21 = W*in
   wire signed [14:0] m68_21;
   assign m68_21 =15'b0;

   // m68_22 = W*in
   wire signed [14:0] m68_22;
   assign m68_22 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_23 = W*in
   wire signed [14:0] m68_23;
   assign m68_23 =15'b0;

   // m68_24 = W*in
   wire signed [14:0] m68_24;
   assign m68_24 =15'b0;

   // m68_25 = W*in
   wire signed [14:0] m68_25;
   assign m68_25 ={ {3{in68[14]}} , in68[14:3] };

   // m68_26 = W*in
   wire signed [14:0] m68_26;
   assign m68_26 =15'b0;

   // m68_27 = W*in
   wire signed [14:0] m68_27;
   assign m68_27 =15'b0;

   // m68_28 = W*in
   wire signed [14:0] m68_28;
   assign m68_28 =15'b0;

   // m68_29 = W*in
   wire signed [14:0] m68_29;
   assign m68_29 ={ {4{in68[14]}} , in68[14:4] };

   // m68_30 = W*in
   wire signed [14:0] m68_30;
   assign m68_30 =15'b0;

   // m68_31 = W*in
   wire signed [14:0] m68_31;
   assign m68_31 ={ {3{in68[14]}} , in68[14:3] };

   // m68_32 = W*in
   wire signed [14:0] m68_32;
   assign m68_32 ={ {3{in68[14]}} , in68[14:3] };

   // m68_33 = W*in
   wire signed [14:0] m68_33;
   assign m68_33 ={ {3{in68[14]}} , in68[14:3] };

   // m68_34 = W*in
   wire signed [14:0] m68_34;
   assign m68_34 =15'b0;

   // m68_35 = W*in
   wire signed [14:0] m68_35;
   assign m68_35 =15'b0;

   // m68_36 = W*in
   wire signed [14:0] m68_36;
   assign m68_36 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_37 = W*in
   wire signed [14:0] m68_37;
   assign m68_37 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_38 = W*in
   wire signed [14:0] m68_38;
   assign m68_38 ={ {3{in68[14]}} , in68[14:3] };

   // m68_39 = W*in
   wire signed [14:0] m68_39;
   assign m68_39 =15'b0;

   // m68_40 = W*in
   wire signed [14:0] m68_40;
   assign m68_40 =15'b0;

   // m68_41 = W*in
   wire signed [14:0] m68_41;
   assign m68_41 =15'b0;

   // m68_42 = W*in
   wire signed [14:0] m68_42;
   assign m68_42 =15'b0;

   // m68_43 = W*in
   wire signed [14:0] m68_43;
   assign m68_43 ={ {3{in68[14]}} , in68[14:3] };

   // m68_44 = W*in
   wire signed [14:0] m68_44;
   assign m68_44 =15'b0;

   // m68_45 = W*in
   wire signed [14:0] m68_45;
   assign m68_45 =15'b0;

   // m68_46 = W*in
   wire signed [14:0] m68_46;
   assign m68_46 =15'b0;

   // m68_47 = W*in
   wire signed [14:0] m68_47;
   assign m68_47 =15'b0;

   // m68_48 = W*in
   wire signed [14:0] m68_48;
   assign m68_48 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_49 = W*in
   wire signed [14:0] m68_49;
   assign m68_49 =15'b0;

   // m68_50 = W*in
   wire signed [14:0] m68_50;
   assign m68_50 =15'b0;

   // m68_51 = W*in
   wire signed [14:0] m68_51;
   assign m68_51 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_52 = W*in
   wire signed [14:0] m68_52;
   assign m68_52 =15'b0;

   // m68_53 = W*in
   wire signed [14:0] m68_53;
   assign m68_53 =15'b0;

   // m68_54 = W*in
   wire signed [14:0] m68_54;
   assign m68_54 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_55 = W*in
   wire signed [14:0] m68_55;
   assign m68_55 =15'b0;

   // m68_56 = W*in
   wire signed [14:0] m68_56;
   assign m68_56 =15'b0;

   // m68_57 = W*in
   wire signed [14:0] m68_57;
   assign m68_57 =15'b0;

   // m68_58 = W*in
   wire signed [14:0] m68_58;
   assign m68_58 ={ {2{neg68[14]}} , neg68[14:2] };

   // m68_59 = W*in
   wire signed [14:0] m68_59;
   assign m68_59 =15'b0;

   // m68_60 = W*in
   wire signed [14:0] m68_60;
   assign m68_60 ={ {4{neg68[14]}} , neg68[14:4] };

   // m68_61 = W*in
   wire signed [14:0] m68_61;
   assign m68_61 ={ {4{neg68[14]}} , neg68[14:4] };

   // m68_62 = W*in
   wire signed [14:0] m68_62;
   assign m68_62 ={ {2{neg68[14]}} , neg68[14:2] };

   // m68_63 = W*in
   wire signed [14:0] m68_63;
   assign m68_63 =15'b0;

   // m68_64 = W*in
   wire signed [14:0] m68_64;
   assign m68_64 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_65 = W*in
   wire signed [14:0] m68_65;
   assign m68_65 =15'b0;

   // m68_66 = W*in
   wire signed [14:0] m68_66;
   assign m68_66 ={ {4{neg68[14]}} , neg68[14:4] };

   // m68_67 = W*in
   wire signed [14:0] m68_67;
   assign m68_67 =15'b0;

   // m68_68 = W*in
   wire signed [14:0] m68_68;
   assign m68_68 ={ {3{in68[14]}} , in68[14:3] };

   // m68_69 = W*in
   wire signed [14:0] m68_69;
   assign m68_69 =15'b0;

   // m68_70 = W*in
   wire signed [14:0] m68_70;
   assign m68_70 =15'b0;

   // m68_71 = W*in
   wire signed [14:0] m68_71;
   assign m68_71 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_72 = W*in
   wire signed [14:0] m68_72;
   assign m68_72 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_73 = W*in
   wire signed [14:0] m68_73;
   assign m68_73 ={ {3{in68[14]}} , in68[14:3] };

   // m68_74 = W*in
   wire signed [14:0] m68_74;
   assign m68_74 =15'b0;

   // m68_75 = W*in
   wire signed [14:0] m68_75;
   assign m68_75 ={ {4{in68[14]}} , in68[14:4] };

   // m68_76 = W*in
   wire signed [14:0] m68_76;
   assign m68_76 =15'b0;

   // m68_77 = W*in
   wire signed [14:0] m68_77;
   assign m68_77 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_78 = W*in
   wire signed [14:0] m68_78;
   assign m68_78 =15'b0;

   // m68_79 = W*in
   wire signed [14:0] m68_79;
   assign m68_79 =15'b0;

   // m68_80 = W*in
   wire signed [14:0] m68_80;
   assign m68_80 =15'b0;

   // m68_81 = W*in
   wire signed [14:0] m68_81;
   assign m68_81 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_82 = W*in
   wire signed [14:0] m68_82;
   assign m68_82 ={ {3{in68[14]}} , in68[14:3] };

   // m68_83 = W*in
   wire signed [14:0] m68_83;
   assign m68_83 =15'b0;

   // m68_84 = W*in
   wire signed [14:0] m68_84;
   assign m68_84 =15'b0;

   // m68_85 = W*in
   wire signed [14:0] m68_85;
   assign m68_85 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_86 = W*in
   wire signed [14:0] m68_86;
   assign m68_86 =15'b0;

   // m68_87 = W*in
   wire signed [14:0] m68_87;
   assign m68_87 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_88 = W*in
   wire signed [14:0] m68_88;
   assign m68_88 =15'b0;

   // m68_89 = W*in
   wire signed [14:0] m68_89;
   assign m68_89 ={ {2{neg68[14]}} , neg68[14:2] };

   // m68_90 = W*in
   wire signed [14:0] m68_90;
   assign m68_90 ={ {3{in68[14]}} , in68[14:3] };

   // m68_91 = W*in
   wire signed [14:0] m68_91;
   assign m68_91 ={ {2{neg68[14]}} , neg68[14:2] };

   // m68_92 = W*in
   wire signed [14:0] m68_92;
   assign m68_92 =15'b0;

   // m68_93 = W*in
   wire signed [14:0] m68_93;
   assign m68_93 ={ {3{neg68[14]}} , neg68[14:3] };

   // m68_94 = W*in
   wire signed [14:0] m68_94;
   assign m68_94 ={ {3{in68[14]}} , in68[14:3] };

   // m68_95 = W*in
   wire signed [14:0] m68_95;
   assign m68_95 =15'b0;

   // m68_96 = W*in
   wire signed [14:0] m68_96;
   assign m68_96 =15'b0;

   // m68_97 = W*in
   wire signed [14:0] m68_97;
   assign m68_97 ={ {3{in68[14]}} , in68[14:3] };

   // m68_98 = W*in
   wire signed [14:0] m68_98;
   assign m68_98 =15'b0;

   // m68_99 = W*in
   wire signed [14:0] m68_99;
   assign m68_99 =15'b0;

   // m68_100 = W*in
   wire signed [14:0] m68_100;
   assign m68_100 ={ {3{neg68[14]}} , neg68[14:3] };

   // m69_1 = W*in
   wire signed [14:0] m69_1;
   assign m69_1 =15'b0;

   // m69_2 = W*in
   wire signed [14:0] m69_2;
   assign m69_2 =15'b0;

   // m69_3 = W*in
   wire signed [14:0] m69_3;
   assign m69_3 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_4 = W*in
   wire signed [14:0] m69_4;
   assign m69_4 =15'b0;

   // m69_5 = W*in
   wire signed [14:0] m69_5;
   assign m69_5 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_6 = W*in
   wire signed [14:0] m69_6;
   assign m69_6 =15'b0;

   // m69_7 = W*in
   wire signed [14:0] m69_7;
   assign m69_7 ={ {4{in69[14]}} , in69[14:4] };

   // m69_8 = W*in
   wire signed [14:0] m69_8;
   assign m69_8 =15'b0;

   // m69_9 = W*in
   wire signed [14:0] m69_9;
   assign m69_9 =15'b0;

   // m69_10 = W*in
   wire signed [14:0] m69_10;
   assign m69_10 =15'b0;

   // m69_11 = W*in
   wire signed [14:0] m69_11;
   assign m69_11 =15'b0;

   // m69_12 = W*in
   wire signed [14:0] m69_12;
   assign m69_12 =15'b0;

   // m69_13 = W*in
   wire signed [14:0] m69_13;
   assign m69_13 =15'b0;

   // m69_14 = W*in
   wire signed [14:0] m69_14;
   assign m69_14 =15'b0;

   // m69_15 = W*in
   wire signed [14:0] m69_15;
   assign m69_15 =15'b0;

   // m69_16 = W*in
   wire signed [14:0] m69_16;
   assign m69_16 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_17 = W*in
   wire signed [14:0] m69_17;
   assign m69_17 =15'b0;

   // m69_18 = W*in
   wire signed [14:0] m69_18;
   assign m69_18 ={ {4{in69[14]}} , in69[14:4] };

   // m69_19 = W*in
   wire signed [14:0] m69_19;
   assign m69_19 =15'b0;

   // m69_20 = W*in
   wire signed [14:0] m69_20;
   assign m69_20 =15'b0;

   // m69_21 = W*in
   wire signed [14:0] m69_21;
   assign m69_21 =15'b0;

   // m69_22 = W*in
   wire signed [14:0] m69_22;
   assign m69_22 =15'b0;

   // m69_23 = W*in
   wire signed [14:0] m69_23;
   assign m69_23 ={ {3{in69[14]}} , in69[14:3] };

   // m69_24 = W*in
   wire signed [14:0] m69_24;
   assign m69_24 =15'b0;

   // m69_25 = W*in
   wire signed [14:0] m69_25;
   assign m69_25 ={ {3{in69[14]}} , in69[14:3] };

   // m69_26 = W*in
   wire signed [14:0] m69_26;
   assign m69_26 =15'b0;

   // m69_27 = W*in
   wire signed [14:0] m69_27;
   assign m69_27 ={ {4{neg69[14]}} , neg69[14:4] };

   // m69_28 = W*in
   wire signed [14:0] m69_28;
   assign m69_28 =15'b0;

   // m69_29 = W*in
   wire signed [14:0] m69_29;
   assign m69_29 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_30 = W*in
   wire signed [14:0] m69_30;
   assign m69_30 =15'b0;

   // m69_31 = W*in
   wire signed [14:0] m69_31;
   assign m69_31 =15'b0;

   // m69_32 = W*in
   wire signed [14:0] m69_32;
   assign m69_32 ={ {3{in69[14]}} , in69[14:3] };

   // m69_33 = W*in
   wire signed [14:0] m69_33;
   assign m69_33 =15'b0;

   // m69_34 = W*in
   wire signed [14:0] m69_34;
   assign m69_34 =15'b0;

   // m69_35 = W*in
   wire signed [14:0] m69_35;
   assign m69_35 =15'b0;

   // m69_36 = W*in
   wire signed [14:0] m69_36;
   assign m69_36 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_37 = W*in
   wire signed [14:0] m69_37;
   assign m69_37 =15'b0;

   // m69_38 = W*in
   wire signed [14:0] m69_38;
   assign m69_38 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_39 = W*in
   wire signed [14:0] m69_39;
   assign m69_39 =15'b0;

   // m69_40 = W*in
   wire signed [14:0] m69_40;
   assign m69_40 =15'b0;

   // m69_41 = W*in
   wire signed [14:0] m69_41;
   assign m69_41 =15'b0;

   // m69_42 = W*in
   wire signed [14:0] m69_42;
   assign m69_42 =15'b0;

   // m69_43 = W*in
   wire signed [14:0] m69_43;
   assign m69_43 =15'b0;

   // m69_44 = W*in
   wire signed [14:0] m69_44;
   assign m69_44 =15'b0;

   // m69_45 = W*in
   wire signed [14:0] m69_45;
   assign m69_45 =15'b0;

   // m69_46 = W*in
   wire signed [14:0] m69_46;
   assign m69_46 ={ {4{neg69[14]}} , neg69[14:4] };

   // m69_47 = W*in
   wire signed [14:0] m69_47;
   assign m69_47 ={ {3{in69[14]}} , in69[14:3] };

   // m69_48 = W*in
   wire signed [14:0] m69_48;
   assign m69_48 =15'b0;

   // m69_49 = W*in
   wire signed [14:0] m69_49;
   assign m69_49 =15'b0;

   // m69_50 = W*in
   wire signed [14:0] m69_50;
   assign m69_50 =15'b0;

   // m69_51 = W*in
   wire signed [14:0] m69_51;
   assign m69_51 =15'b0;

   // m69_52 = W*in
   wire signed [14:0] m69_52;
   assign m69_52 =15'b0;

   // m69_53 = W*in
   wire signed [14:0] m69_53;
   assign m69_53 =15'b0;

   // m69_54 = W*in
   wire signed [14:0] m69_54;
   assign m69_54 =15'b0;

   // m69_55 = W*in
   wire signed [14:0] m69_55;
   assign m69_55 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_56 = W*in
   wire signed [14:0] m69_56;
   assign m69_56 =15'b0;

   // m69_57 = W*in
   wire signed [14:0] m69_57;
   assign m69_57 =15'b0;

   // m69_58 = W*in
   wire signed [14:0] m69_58;
   assign m69_58 =15'b0;

   // m69_59 = W*in
   wire signed [14:0] m69_59;
   assign m69_59 ={ {3{in69[14]}} , in69[14:3] };

   // m69_60 = W*in
   wire signed [14:0] m69_60;
   assign m69_60 =15'b0;

   // m69_61 = W*in
   wire signed [14:0] m69_61;
   assign m69_61 =15'b0;

   // m69_62 = W*in
   wire signed [14:0] m69_62;
   assign m69_62 =15'b0;

   // m69_63 = W*in
   wire signed [14:0] m69_63;
   assign m69_63 =15'b0;

   // m69_64 = W*in
   wire signed [14:0] m69_64;
   assign m69_64 =15'b0;

   // m69_65 = W*in
   wire signed [14:0] m69_65;
   assign m69_65 =15'b0;

   // m69_66 = W*in
   wire signed [14:0] m69_66;
   assign m69_66 =15'b0;

   // m69_67 = W*in
   wire signed [14:0] m69_67;
   assign m69_67 =15'b0;

   // m69_68 = W*in
   wire signed [14:0] m69_68;
   assign m69_68 =15'b0;

   // m69_69 = W*in
   wire signed [14:0] m69_69;
   assign m69_69 =15'b0;

   // m69_70 = W*in
   wire signed [14:0] m69_70;
   assign m69_70 =15'b0;

   // m69_71 = W*in
   wire signed [14:0] m69_71;
   assign m69_71 =15'b0;

   // m69_72 = W*in
   wire signed [14:0] m69_72;
   assign m69_72 =15'b0;

   // m69_73 = W*in
   wire signed [14:0] m69_73;
   assign m69_73 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_74 = W*in
   wire signed [14:0] m69_74;
   assign m69_74 =15'b0;

   // m69_75 = W*in
   wire signed [14:0] m69_75;
   assign m69_75 =15'b0;

   // m69_76 = W*in
   wire signed [14:0] m69_76;
   assign m69_76 =15'b0;

   // m69_77 = W*in
   wire signed [14:0] m69_77;
   assign m69_77 =15'b0;

   // m69_78 = W*in
   wire signed [14:0] m69_78;
   assign m69_78 =15'b0;

   // m69_79 = W*in
   wire signed [14:0] m69_79;
   assign m69_79 =15'b0;

   // m69_80 = W*in
   wire signed [14:0] m69_80;
   assign m69_80 =15'b0;

   // m69_81 = W*in
   wire signed [14:0] m69_81;
   assign m69_81 =15'b0;

   // m69_82 = W*in
   wire signed [14:0] m69_82;
   assign m69_82 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_83 = W*in
   wire signed [14:0] m69_83;
   assign m69_83 =15'b0;

   // m69_84 = W*in
   wire signed [14:0] m69_84;
   assign m69_84 =15'b0;

   // m69_85 = W*in
   wire signed [14:0] m69_85;
   assign m69_85 =15'b0;

   // m69_86 = W*in
   wire signed [14:0] m69_86;
   assign m69_86 =15'b0;

   // m69_87 = W*in
   wire signed [14:0] m69_87;
   assign m69_87 =15'b0;

   // m69_88 = W*in
   wire signed [14:0] m69_88;
   assign m69_88 =15'b0;

   // m69_89 = W*in
   wire signed [14:0] m69_89;
   assign m69_89 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_90 = W*in
   wire signed [14:0] m69_90;
   assign m69_90 =15'b0;

   // m69_91 = W*in
   wire signed [14:0] m69_91;
   assign m69_91 =15'b0;

   // m69_92 = W*in
   wire signed [14:0] m69_92;
   assign m69_92 =15'b0;

   // m69_93 = W*in
   wire signed [14:0] m69_93;
   assign m69_93 =15'b0;

   // m69_94 = W*in
   wire signed [14:0] m69_94;
   assign m69_94 =15'b0;

   // m69_95 = W*in
   wire signed [14:0] m69_95;
   assign m69_95 =15'b0;

   // m69_96 = W*in
   wire signed [14:0] m69_96;
   assign m69_96 =15'b0;

   // m69_97 = W*in
   wire signed [14:0] m69_97;
   assign m69_97 ={ {3{neg69[14]}} , neg69[14:3] };

   // m69_98 = W*in
   wire signed [14:0] m69_98;
   assign m69_98 =15'b0;

   // m69_99 = W*in
   wire signed [14:0] m69_99;
   assign m69_99 =15'b0;

   // m69_100 = W*in
   wire signed [14:0] m69_100;
   assign m69_100 ={ {3{neg69[14]}} , neg69[14:3] };

   // m70_1 = W*in
   wire signed [14:0] m70_1;
   assign m70_1 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_2 = W*in
   wire signed [14:0] m70_2;
   assign m70_2 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_3 = W*in
   wire signed [14:0] m70_3;
   assign m70_3 =15'b0;

   // m70_4 = W*in
   wire signed [14:0] m70_4;
   assign m70_4 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_5 = W*in
   wire signed [14:0] m70_5;
   assign m70_5 =15'b0;

   // m70_6 = W*in
   wire signed [14:0] m70_6;
   assign m70_6 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_7 = W*in
   wire signed [14:0] m70_7;
   assign m70_7 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_8 = W*in
   wire signed [14:0] m70_8;
   assign m70_8 =15'b0;

   // m70_9 = W*in
   wire signed [14:0] m70_9;
   assign m70_9 =15'b0;

   // m70_10 = W*in
   wire signed [14:0] m70_10;
   assign m70_10 =15'b0;

   // m70_11 = W*in
   wire signed [14:0] m70_11;
   assign m70_11 =15'b0;

   // m70_12 = W*in
   wire signed [14:0] m70_12;
   assign m70_12 =15'b0;

   // m70_13 = W*in
   wire signed [14:0] m70_13;
   assign m70_13 =15'b0;

   // m70_14 = W*in
   wire signed [14:0] m70_14;
   assign m70_14 =15'b0;

   // m70_15 = W*in
   wire signed [14:0] m70_15;
   assign m70_15 ={ {3{in70[14]}} , in70[14:3] };

   // m70_16 = W*in
   wire signed [14:0] m70_16;
   assign m70_16 =15'b0;

   // m70_17 = W*in
   wire signed [14:0] m70_17;
   assign m70_17 =15'b0;

   // m70_18 = W*in
   wire signed [14:0] m70_18;
   assign m70_18 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_19 = W*in
   wire signed [14:0] m70_19;
   assign m70_19 ={ {4{in70[14]}} , in70[14:4] };

   // m70_20 = W*in
   wire signed [14:0] m70_20;
   assign m70_20 =15'b0;

   // m70_21 = W*in
   wire signed [14:0] m70_21;
   assign m70_21 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_22 = W*in
   wire signed [14:0] m70_22;
   assign m70_22 =15'b0;

   // m70_23 = W*in
   wire signed [14:0] m70_23;
   assign m70_23 =15'b0;

   // m70_24 = W*in
   wire signed [14:0] m70_24;
   assign m70_24 =15'b0;

   // m70_25 = W*in
   wire signed [14:0] m70_25;
   assign m70_25 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_26 = W*in
   wire signed [14:0] m70_26;
   assign m70_26 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_27 = W*in
   wire signed [14:0] m70_27;
   assign m70_27 =15'b0;

   // m70_28 = W*in
   wire signed [14:0] m70_28;
   assign m70_28 =15'b0;

   // m70_29 = W*in
   wire signed [14:0] m70_29;
   assign m70_29 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_30 = W*in
   wire signed [14:0] m70_30;
   assign m70_30 =15'b0;

   // m70_31 = W*in
   wire signed [14:0] m70_31;
   assign m70_31 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_32 = W*in
   wire signed [14:0] m70_32;
   assign m70_32 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_33 = W*in
   wire signed [14:0] m70_33;
   assign m70_33 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_34 = W*in
   wire signed [14:0] m70_34;
   assign m70_34 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_35 = W*in
   wire signed [14:0] m70_35;
   assign m70_35 =15'b0;

   // m70_36 = W*in
   wire signed [14:0] m70_36;
   assign m70_36 =15'b0;

   // m70_37 = W*in
   wire signed [14:0] m70_37;
   assign m70_37 =15'b0;

   // m70_38 = W*in
   wire signed [14:0] m70_38;
   assign m70_38 =15'b0;

   // m70_39 = W*in
   wire signed [14:0] m70_39;
   assign m70_39 =15'b0;

   // m70_40 = W*in
   wire signed [14:0] m70_40;
   assign m70_40 =15'b0;

   // m70_41 = W*in
   wire signed [14:0] m70_41;
   assign m70_41 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_42 = W*in
   wire signed [14:0] m70_42;
   assign m70_42 =15'b0;

   // m70_43 = W*in
   wire signed [14:0] m70_43;
   assign m70_43 =15'b0;

   // m70_44 = W*in
   wire signed [14:0] m70_44;
   assign m70_44 =15'b0;

   // m70_45 = W*in
   wire signed [14:0] m70_45;
   assign m70_45 =15'b0;

   // m70_46 = W*in
   wire signed [14:0] m70_46;
   assign m70_46 =15'b0;

   // m70_47 = W*in
   wire signed [14:0] m70_47;
   assign m70_47 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_48 = W*in
   wire signed [14:0] m70_48;
   assign m70_48 =15'b0;

   // m70_49 = W*in
   wire signed [14:0] m70_49;
   assign m70_49 =15'b0;

   // m70_50 = W*in
   wire signed [14:0] m70_50;
   assign m70_50 =15'b0;

   // m70_51 = W*in
   wire signed [14:0] m70_51;
   assign m70_51 =15'b0;

   // m70_52 = W*in
   wire signed [14:0] m70_52;
   assign m70_52 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_53 = W*in
   wire signed [14:0] m70_53;
   assign m70_53 =15'b0;

   // m70_54 = W*in
   wire signed [14:0] m70_54;
   assign m70_54 =15'b0;

   // m70_55 = W*in
   wire signed [14:0] m70_55;
   assign m70_55 =15'b0;

   // m70_56 = W*in
   wire signed [14:0] m70_56;
   assign m70_56 =15'b0;

   // m70_57 = W*in
   wire signed [14:0] m70_57;
   assign m70_57 ={ {3{in70[14]}} , in70[14:3] };

   // m70_58 = W*in
   wire signed [14:0] m70_58;
   assign m70_58 ={ {3{in70[14]}} , in70[14:3] };

   // m70_59 = W*in
   wire signed [14:0] m70_59;
   assign m70_59 ={ {4{in70[14]}} , in70[14:4] };

   // m70_60 = W*in
   wire signed [14:0] m70_60;
   assign m70_60 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_61 = W*in
   wire signed [14:0] m70_61;
   assign m70_61 ={ {3{in70[14]}} , in70[14:3] };

   // m70_62 = W*in
   wire signed [14:0] m70_62;
   assign m70_62 =15'b0;

   // m70_63 = W*in
   wire signed [14:0] m70_63;
   assign m70_63 =15'b0;

   // m70_64 = W*in
   wire signed [14:0] m70_64;
   assign m70_64 ={ {3{in70[14]}} , in70[14:3] };

   // m70_65 = W*in
   wire signed [14:0] m70_65;
   assign m70_65 =15'b0;

   // m70_66 = W*in
   wire signed [14:0] m70_66;
   assign m70_66 =15'b0;

   // m70_67 = W*in
   wire signed [14:0] m70_67;
   assign m70_67 =15'b0;

   // m70_68 = W*in
   wire signed [14:0] m70_68;
   assign m70_68 =15'b0;

   // m70_69 = W*in
   wire signed [14:0] m70_69;
   assign m70_69 =15'b0;

   // m70_70 = W*in
   wire signed [14:0] m70_70;
   assign m70_70 ={ {4{in70[14]}} , in70[14:4] };

   // m70_71 = W*in
   wire signed [14:0] m70_71;
   assign m70_71 =15'b0;

   // m70_72 = W*in
   wire signed [14:0] m70_72;
   assign m70_72 =15'b0;

   // m70_73 = W*in
   wire signed [14:0] m70_73;
   assign m70_73 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_74 = W*in
   wire signed [14:0] m70_74;
   assign m70_74 ={ {4{in70[14]}} , in70[14:4] };

   // m70_75 = W*in
   wire signed [14:0] m70_75;
   assign m70_75 ={ {4{neg70[14]}} , neg70[14:4] };

   // m70_76 = W*in
   wire signed [14:0] m70_76;
   assign m70_76 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_77 = W*in
   wire signed [14:0] m70_77;
   assign m70_77 =15'b0;

   // m70_78 = W*in
   wire signed [14:0] m70_78;
   assign m70_78 =15'b0;

   // m70_79 = W*in
   wire signed [14:0] m70_79;
   assign m70_79 ={ {3{in70[14]}} , in70[14:3] };

   // m70_80 = W*in
   wire signed [14:0] m70_80;
   assign m70_80 =15'b0;

   // m70_81 = W*in
   wire signed [14:0] m70_81;
   assign m70_81 =15'b0;

   // m70_82 = W*in
   wire signed [14:0] m70_82;
   assign m70_82 =15'b0;

   // m70_83 = W*in
   wire signed [14:0] m70_83;
   assign m70_83 =15'b0;

   // m70_84 = W*in
   wire signed [14:0] m70_84;
   assign m70_84 =15'b0;

   // m70_85 = W*in
   wire signed [14:0] m70_85;
   assign m70_85 =15'b0;

   // m70_86 = W*in
   wire signed [14:0] m70_86;
   assign m70_86 =15'b0;

   // m70_87 = W*in
   wire signed [14:0] m70_87;
   assign m70_87 =15'b0;

   // m70_88 = W*in
   wire signed [14:0] m70_88;
   assign m70_88 =15'b0;

   // m70_89 = W*in
   wire signed [14:0] m70_89;
   assign m70_89 =15'b0;

   // m70_90 = W*in
   wire signed [14:0] m70_90;
   assign m70_90 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_91 = W*in
   wire signed [14:0] m70_91;
   assign m70_91 =15'b0;

   // m70_92 = W*in
   wire signed [14:0] m70_92;
   assign m70_92 ={ {3{in70[14]}} , in70[14:3] };

   // m70_93 = W*in
   wire signed [14:0] m70_93;
   assign m70_93 =15'b0;

   // m70_94 = W*in
   wire signed [14:0] m70_94;
   assign m70_94 =15'b0;

   // m70_95 = W*in
   wire signed [14:0] m70_95;
   assign m70_95 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_96 = W*in
   wire signed [14:0] m70_96;
   assign m70_96 ={ {3{neg70[14]}} , neg70[14:3] };

   // m70_97 = W*in
   wire signed [14:0] m70_97;
   assign m70_97 ={ {3{in70[14]}} , in70[14:3] };

   // m70_98 = W*in
   wire signed [14:0] m70_98;
   assign m70_98 =15'b0;

   // m70_99 = W*in
   wire signed [14:0] m70_99;
   assign m70_99 =15'b0;

   // m70_100 = W*in
   wire signed [14:0] m70_100;
   assign m70_100 =15'b0;

   // m71_1 = W*in
   wire signed [14:0] m71_1;
   assign m71_1 =15'b0;

   // m71_2 = W*in
   wire signed [14:0] m71_2;
   assign m71_2 =15'b0;

   // m71_3 = W*in
   wire signed [14:0] m71_3;
   assign m71_3 =15'b0;

   // m71_4 = W*in
   wire signed [14:0] m71_4;
   assign m71_4 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_5 = W*in
   wire signed [14:0] m71_5;
   assign m71_5 =15'b0;

   // m71_6 = W*in
   wire signed [14:0] m71_6;
   assign m71_6 =15'b0;

   // m71_7 = W*in
   wire signed [14:0] m71_7;
   assign m71_7 =15'b0;

   // m71_8 = W*in
   wire signed [14:0] m71_8;
   assign m71_8 =15'b0;

   // m71_9 = W*in
   wire signed [14:0] m71_9;
   assign m71_9 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_10 = W*in
   wire signed [14:0] m71_10;
   assign m71_10 ={ {2{in71[14]}} , in71[14:2] };

   // m71_11 = W*in
   wire signed [14:0] m71_11;
   assign m71_11 =15'b0;

   // m71_12 = W*in
   wire signed [14:0] m71_12;
   assign m71_12 =15'b0;

   // m71_13 = W*in
   wire signed [14:0] m71_13;
   assign m71_13 =15'b0;

   // m71_14 = W*in
   wire signed [14:0] m71_14;
   assign m71_14 =15'b0;

   // m71_15 = W*in
   wire signed [14:0] m71_15;
   assign m71_15 =15'b0;

   // m71_16 = W*in
   wire signed [14:0] m71_16;
   assign m71_16 =15'b0;

   // m71_17 = W*in
   wire signed [14:0] m71_17;
   assign m71_17 =15'b0;

   // m71_18 = W*in
   wire signed [14:0] m71_18;
   assign m71_18 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_19 = W*in
   wire signed [14:0] m71_19;
   assign m71_19 ={ {3{in71[14]}} , in71[14:3] };

   // m71_20 = W*in
   wire signed [14:0] m71_20;
   assign m71_20 =15'b0;

   // m71_21 = W*in
   wire signed [14:0] m71_21;
   assign m71_21 =15'b0;

   // m71_22 = W*in
   wire signed [14:0] m71_22;
   assign m71_22 =15'b0;

   // m71_23 = W*in
   wire signed [14:0] m71_23;
   assign m71_23 =15'b0;

   // m71_24 = W*in
   wire signed [14:0] m71_24;
   assign m71_24 =15'b0;

   // m71_25 = W*in
   wire signed [14:0] m71_25;
   assign m71_25 =15'b0;

   // m71_26 = W*in
   wire signed [14:0] m71_26;
   assign m71_26 =15'b0;

   // m71_27 = W*in
   wire signed [14:0] m71_27;
   assign m71_27 =15'b0;

   // m71_28 = W*in
   wire signed [14:0] m71_28;
   assign m71_28 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_29 = W*in
   wire signed [14:0] m71_29;
   assign m71_29 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_30 = W*in
   wire signed [14:0] m71_30;
   assign m71_30 =15'b0;

   // m71_31 = W*in
   wire signed [14:0] m71_31;
   assign m71_31 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_32 = W*in
   wire signed [14:0] m71_32;
   assign m71_32 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_33 = W*in
   wire signed [14:0] m71_33;
   assign m71_33 =15'b0;

   // m71_34 = W*in
   wire signed [14:0] m71_34;
   assign m71_34 =15'b0;

   // m71_35 = W*in
   wire signed [14:0] m71_35;
   assign m71_35 =15'b0;

   // m71_36 = W*in
   wire signed [14:0] m71_36;
   assign m71_36 =15'b0;

   // m71_37 = W*in
   wire signed [14:0] m71_37;
   assign m71_37 =15'b0;

   // m71_38 = W*in
   wire signed [14:0] m71_38;
   assign m71_38 =15'b0;

   // m71_39 = W*in
   wire signed [14:0] m71_39;
   assign m71_39 ={ {3{in71[14]}} , in71[14:3] };

   // m71_40 = W*in
   wire signed [14:0] m71_40;
   assign m71_40 =15'b0;

   // m71_41 = W*in
   wire signed [14:0] m71_41;
   assign m71_41 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_42 = W*in
   wire signed [14:0] m71_42;
   assign m71_42 =15'b0;

   // m71_43 = W*in
   wire signed [14:0] m71_43;
   assign m71_43 =15'b0;

   // m71_44 = W*in
   wire signed [14:0] m71_44;
   assign m71_44 =15'b0;

   // m71_45 = W*in
   wire signed [14:0] m71_45;
   assign m71_45 =15'b0;

   // m71_46 = W*in
   wire signed [14:0] m71_46;
   assign m71_46 ={ {2{in71[14]}} , in71[14:2] };

   // m71_47 = W*in
   wire signed [14:0] m71_47;
   assign m71_47 =15'b0;

   // m71_48 = W*in
   wire signed [14:0] m71_48;
   assign m71_48 =15'b0;

   // m71_49 = W*in
   wire signed [14:0] m71_49;
   assign m71_49 =15'b0;

   // m71_50 = W*in
   wire signed [14:0] m71_50;
   assign m71_50 =15'b0;

   // m71_51 = W*in
   wire signed [14:0] m71_51;
   assign m71_51 =15'b0;

   // m71_52 = W*in
   wire signed [14:0] m71_52;
   assign m71_52 =15'b0;

   // m71_53 = W*in
   wire signed [14:0] m71_53;
   assign m71_53 =15'b0;

   // m71_54 = W*in
   wire signed [14:0] m71_54;
   assign m71_54 ={ {3{in71[14]}} , in71[14:3] };

   // m71_55 = W*in
   wire signed [14:0] m71_55;
   assign m71_55 =15'b0;

   // m71_56 = W*in
   wire signed [14:0] m71_56;
   assign m71_56 =15'b0;

   // m71_57 = W*in
   wire signed [14:0] m71_57;
   assign m71_57 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_58 = W*in
   wire signed [14:0] m71_58;
   assign m71_58 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_59 = W*in
   wire signed [14:0] m71_59;
   assign m71_59 =15'b0;

   // m71_60 = W*in
   wire signed [14:0] m71_60;
   assign m71_60 =15'b0;

   // m71_61 = W*in
   wire signed [14:0] m71_61;
   assign m71_61 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_62 = W*in
   wire signed [14:0] m71_62;
   assign m71_62 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_63 = W*in
   wire signed [14:0] m71_63;
   assign m71_63 =15'b0;

   // m71_64 = W*in
   wire signed [14:0] m71_64;
   assign m71_64 =15'b0;

   // m71_65 = W*in
   wire signed [14:0] m71_65;
   assign m71_65 ={ {3{in71[14]}} , in71[14:3] };

   // m71_66 = W*in
   wire signed [14:0] m71_66;
   assign m71_66 ={ {3{in71[14]}} , in71[14:3] };

   // m71_67 = W*in
   wire signed [14:0] m71_67;
   assign m71_67 =15'b0;

   // m71_68 = W*in
   wire signed [14:0] m71_68;
   assign m71_68 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_69 = W*in
   wire signed [14:0] m71_69;
   assign m71_69 ={ {4{in71[14]}} , in71[14:4] };

   // m71_70 = W*in
   wire signed [14:0] m71_70;
   assign m71_70 =15'b0;

   // m71_71 = W*in
   wire signed [14:0] m71_71;
   assign m71_71 =15'b0;

   // m71_72 = W*in
   wire signed [14:0] m71_72;
   assign m71_72 =15'b0;

   // m71_73 = W*in
   wire signed [14:0] m71_73;
   assign m71_73 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_74 = W*in
   wire signed [14:0] m71_74;
   assign m71_74 ={ {4{neg71[14]}} , neg71[14:4] };

   // m71_75 = W*in
   wire signed [14:0] m71_75;
   assign m71_75 =15'b0;

   // m71_76 = W*in
   wire signed [14:0] m71_76;
   assign m71_76 =15'b0;

   // m71_77 = W*in
   wire signed [14:0] m71_77;
   assign m71_77 =15'b0;

   // m71_78 = W*in
   wire signed [14:0] m71_78;
   assign m71_78 =15'b0;

   // m71_79 = W*in
   wire signed [14:0] m71_79;
   assign m71_79 ={ {3{in71[14]}} , in71[14:3] };

   // m71_80 = W*in
   wire signed [14:0] m71_80;
   assign m71_80 =15'b0;

   // m71_81 = W*in
   wire signed [14:0] m71_81;
   assign m71_81 =15'b0;

   // m71_82 = W*in
   wire signed [14:0] m71_82;
   assign m71_82 =15'b0;

   // m71_83 = W*in
   wire signed [14:0] m71_83;
   assign m71_83 =15'b0;

   // m71_84 = W*in
   wire signed [14:0] m71_84;
   assign m71_84 =15'b0;

   // m71_85 = W*in
   wire signed [14:0] m71_85;
   assign m71_85 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_86 = W*in
   wire signed [14:0] m71_86;
   assign m71_86 ={ {3{in71[14]}} , in71[14:3] };

   // m71_87 = W*in
   wire signed [14:0] m71_87;
   assign m71_87 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_88 = W*in
   wire signed [14:0] m71_88;
   assign m71_88 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_89 = W*in
   wire signed [14:0] m71_89;
   assign m71_89 =15'b0;

   // m71_90 = W*in
   wire signed [14:0] m71_90;
   assign m71_90 =15'b0;

   // m71_91 = W*in
   wire signed [14:0] m71_91;
   assign m71_91 =15'b0;

   // m71_92 = W*in
   wire signed [14:0] m71_92;
   assign m71_92 =15'b0;

   // m71_93 = W*in
   wire signed [14:0] m71_93;
   assign m71_93 =15'b0;

   // m71_94 = W*in
   wire signed [14:0] m71_94;
   assign m71_94 =15'b0;

   // m71_95 = W*in
   wire signed [14:0] m71_95;
   assign m71_95 =15'b0;

   // m71_96 = W*in
   wire signed [14:0] m71_96;
   assign m71_96 =15'b0;

   // m71_97 = W*in
   wire signed [14:0] m71_97;
   assign m71_97 =15'b0;

   // m71_98 = W*in
   wire signed [14:0] m71_98;
   assign m71_98 =15'b0;

   // m71_99 = W*in
   wire signed [14:0] m71_99;
   assign m71_99 ={ {3{neg71[14]}} , neg71[14:3] };

   // m71_100 = W*in
   wire signed [14:0] m71_100;
   assign m71_100 =15'b0;

   // m72_1 = W*in
   wire signed [14:0] m72_1;
   assign m72_1 ={ {3{in72[14]}} , in72[14:3] };

   // m72_2 = W*in
   wire signed [14:0] m72_2;
   assign m72_2 =15'b0;

   // m72_3 = W*in
   wire signed [14:0] m72_3;
   assign m72_3 =15'b0;

   // m72_4 = W*in
   wire signed [14:0] m72_4;
   assign m72_4 =15'b0;

   // m72_5 = W*in
   wire signed [14:0] m72_5;
   assign m72_5 =15'b0;

   // m72_6 = W*in
   wire signed [14:0] m72_6;
   assign m72_6 =15'b0;

   // m72_7 = W*in
   wire signed [14:0] m72_7;
   assign m72_7 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_8 = W*in
   wire signed [14:0] m72_8;
   assign m72_8 =15'b0;

   // m72_9 = W*in
   wire signed [14:0] m72_9;
   assign m72_9 =15'b0;

   // m72_10 = W*in
   wire signed [14:0] m72_10;
   assign m72_10 =15'b0;

   // m72_11 = W*in
   wire signed [14:0] m72_11;
   assign m72_11 =15'b0;

   // m72_12 = W*in
   wire signed [14:0] m72_12;
   assign m72_12 =15'b0;

   // m72_13 = W*in
   wire signed [14:0] m72_13;
   assign m72_13 ={ {3{in72[14]}} , in72[14:3] };

   // m72_14 = W*in
   wire signed [14:0] m72_14;
   assign m72_14 =15'b0;

   // m72_15 = W*in
   wire signed [14:0] m72_15;
   assign m72_15 =15'b0;

   // m72_16 = W*in
   wire signed [14:0] m72_16;
   assign m72_16 =15'b0;

   // m72_17 = W*in
   wire signed [14:0] m72_17;
   assign m72_17 =15'b0;

   // m72_18 = W*in
   wire signed [14:0] m72_18;
   assign m72_18 =15'b0;

   // m72_19 = W*in
   wire signed [14:0] m72_19;
   assign m72_19 =15'b0;

   // m72_20 = W*in
   wire signed [14:0] m72_20;
   assign m72_20 =15'b0;

   // m72_21 = W*in
   wire signed [14:0] m72_21;
   assign m72_21 ={ {3{in72[14]}} , in72[14:3] };

   // m72_22 = W*in
   wire signed [14:0] m72_22;
   assign m72_22 ={ {4{in72[14]}} , in72[14:4] };

   // m72_23 = W*in
   wire signed [14:0] m72_23;
   assign m72_23 =15'b0;

   // m72_24 = W*in
   wire signed [14:0] m72_24;
   assign m72_24 ={ {3{in72[14]}} , in72[14:3] };

   // m72_25 = W*in
   wire signed [14:0] m72_25;
   assign m72_25 =15'b0;

   // m72_26 = W*in
   wire signed [14:0] m72_26;
   assign m72_26 =15'b0;

   // m72_27 = W*in
   wire signed [14:0] m72_27;
   assign m72_27 ={ {4{in72[14]}} , in72[14:4] };

   // m72_28 = W*in
   wire signed [14:0] m72_28;
   assign m72_28 =15'b0;

   // m72_29 = W*in
   wire signed [14:0] m72_29;
   assign m72_29 ={ {4{neg72[14]}} , neg72[14:4] };

   // m72_30 = W*in
   wire signed [14:0] m72_30;
   assign m72_30 =15'b0;

   // m72_31 = W*in
   wire signed [14:0] m72_31;
   assign m72_31 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_32 = W*in
   wire signed [14:0] m72_32;
   assign m72_32 ={ {4{neg72[14]}} , neg72[14:4] };

   // m72_33 = W*in
   wire signed [14:0] m72_33;
   assign m72_33 ={ {4{neg72[14]}} , neg72[14:4] };

   // m72_34 = W*in
   wire signed [14:0] m72_34;
   assign m72_34 =15'b0;

   // m72_35 = W*in
   wire signed [14:0] m72_35;
   assign m72_35 =15'b0;

   // m72_36 = W*in
   wire signed [14:0] m72_36;
   assign m72_36 =15'b0;

   // m72_37 = W*in
   wire signed [14:0] m72_37;
   assign m72_37 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_38 = W*in
   wire signed [14:0] m72_38;
   assign m72_38 =15'b0;

   // m72_39 = W*in
   wire signed [14:0] m72_39;
   assign m72_39 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_40 = W*in
   wire signed [14:0] m72_40;
   assign m72_40 =15'b0;

   // m72_41 = W*in
   wire signed [14:0] m72_41;
   assign m72_41 =15'b0;

   // m72_42 = W*in
   wire signed [14:0] m72_42;
   assign m72_42 =15'b0;

   // m72_43 = W*in
   wire signed [14:0] m72_43;
   assign m72_43 =15'b0;

   // m72_44 = W*in
   wire signed [14:0] m72_44;
   assign m72_44 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_45 = W*in
   wire signed [14:0] m72_45;
   assign m72_45 =15'b0;

   // m72_46 = W*in
   wire signed [14:0] m72_46;
   assign m72_46 =15'b0;

   // m72_47 = W*in
   wire signed [14:0] m72_47;
   assign m72_47 =15'b0;

   // m72_48 = W*in
   wire signed [14:0] m72_48;
   assign m72_48 =15'b0;

   // m72_49 = W*in
   wire signed [14:0] m72_49;
   assign m72_49 =15'b0;

   // m72_50 = W*in
   wire signed [14:0] m72_50;
   assign m72_50 =15'b0;

   // m72_51 = W*in
   wire signed [14:0] m72_51;
   assign m72_51 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_52 = W*in
   wire signed [14:0] m72_52;
   assign m72_52 =15'b0;

   // m72_53 = W*in
   wire signed [14:0] m72_53;
   assign m72_53 =15'b0;

   // m72_54 = W*in
   wire signed [14:0] m72_54;
   assign m72_54 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_55 = W*in
   wire signed [14:0] m72_55;
   assign m72_55 =15'b0;

   // m72_56 = W*in
   wire signed [14:0] m72_56;
   assign m72_56 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_57 = W*in
   wire signed [14:0] m72_57;
   assign m72_57 ={ {3{in72[14]}} , in72[14:3] };

   // m72_58 = W*in
   wire signed [14:0] m72_58;
   assign m72_58 ={ {4{in72[14]}} , in72[14:4] };

   // m72_59 = W*in
   wire signed [14:0] m72_59;
   assign m72_59 =15'b0;

   // m72_60 = W*in
   wire signed [14:0] m72_60;
   assign m72_60 =15'b0;

   // m72_61 = W*in
   wire signed [14:0] m72_61;
   assign m72_61 ={ {3{in72[14]}} , in72[14:3] };

   // m72_62 = W*in
   wire signed [14:0] m72_62;
   assign m72_62 =15'b0;

   // m72_63 = W*in
   wire signed [14:0] m72_63;
   assign m72_63 =15'b0;

   // m72_64 = W*in
   wire signed [14:0] m72_64;
   assign m72_64 ={ {3{in72[14]}} , in72[14:3] };

   // m72_65 = W*in
   wire signed [14:0] m72_65;
   assign m72_65 ={ {3{in72[14]}} , in72[14:3] };

   // m72_66 = W*in
   wire signed [14:0] m72_66;
   assign m72_66 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_67 = W*in
   wire signed [14:0] m72_67;
   assign m72_67 ={ {4{in72[14]}} , in72[14:4] };

   // m72_68 = W*in
   wire signed [14:0] m72_68;
   assign m72_68 ={ {3{in72[14]}} , in72[14:3] };

   // m72_69 = W*in
   wire signed [14:0] m72_69;
   assign m72_69 ={ {4{in72[14]}} , in72[14:4] };

   // m72_70 = W*in
   wire signed [14:0] m72_70;
   assign m72_70 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_71 = W*in
   wire signed [14:0] m72_71;
   assign m72_71 =15'b0;

   // m72_72 = W*in
   wire signed [14:0] m72_72;
   assign m72_72 =15'b0;

   // m72_73 = W*in
   wire signed [14:0] m72_73;
   assign m72_73 ={ {3{in72[14]}} , in72[14:3] };

   // m72_74 = W*in
   wire signed [14:0] m72_74;
   assign m72_74 =15'b0;

   // m72_75 = W*in
   wire signed [14:0] m72_75;
   assign m72_75 =15'b0;

   // m72_76 = W*in
   wire signed [14:0] m72_76;
   assign m72_76 =15'b0;

   // m72_77 = W*in
   wire signed [14:0] m72_77;
   assign m72_77 =15'b0;

   // m72_78 = W*in
   wire signed [14:0] m72_78;
   assign m72_78 =15'b0;

   // m72_79 = W*in
   wire signed [14:0] m72_79;
   assign m72_79 =15'b0;

   // m72_80 = W*in
   wire signed [14:0] m72_80;
   assign m72_80 =15'b0;

   // m72_81 = W*in
   wire signed [14:0] m72_81;
   assign m72_81 =15'b0;

   // m72_82 = W*in
   wire signed [14:0] m72_82;
   assign m72_82 ={ {3{in72[14]}} , in72[14:3] };

   // m72_83 = W*in
   wire signed [14:0] m72_83;
   assign m72_83 =15'b0;

   // m72_84 = W*in
   wire signed [14:0] m72_84;
   assign m72_84 ={ {3{neg72[14]}} , neg72[14:3] };

   // m72_85 = W*in
   wire signed [14:0] m72_85;
   assign m72_85 =15'b0;

   // m72_86 = W*in
   wire signed [14:0] m72_86;
   assign m72_86 =15'b0;

   // m72_87 = W*in
   wire signed [14:0] m72_87;
   assign m72_87 =15'b0;

   // m72_88 = W*in
   wire signed [14:0] m72_88;
   assign m72_88 =15'b0;

   // m72_89 = W*in
   wire signed [14:0] m72_89;
   assign m72_89 =15'b0;

   // m72_90 = W*in
   wire signed [14:0] m72_90;
   assign m72_90 =15'b0;

   // m72_91 = W*in
   wire signed [14:0] m72_91;
   assign m72_91 =15'b0;

   // m72_92 = W*in
   wire signed [14:0] m72_92;
   assign m72_92 ={ {3{in72[14]}} , in72[14:3] };

   // m72_93 = W*in
   wire signed [14:0] m72_93;
   assign m72_93 =15'b0;

   // m72_94 = W*in
   wire signed [14:0] m72_94;
   assign m72_94 =15'b0;

   // m72_95 = W*in
   wire signed [14:0] m72_95;
   assign m72_95 =15'b0;

   // m72_96 = W*in
   wire signed [14:0] m72_96;
   assign m72_96 =15'b0;

   // m72_97 = W*in
   wire signed [14:0] m72_97;
   assign m72_97 ={ {3{in72[14]}} , in72[14:3] };

   // m72_98 = W*in
   wire signed [14:0] m72_98;
   assign m72_98 =15'b0;

   // m72_99 = W*in
   wire signed [14:0] m72_99;
   assign m72_99 =15'b0;

   // m72_100 = W*in
   wire signed [14:0] m72_100;
   assign m72_100 =15'b0;

   // m73_1 = W*in
   wire signed [14:0] m73_1;
   assign m73_1 =15'b0;

   // m73_2 = W*in
   wire signed [14:0] m73_2;
   assign m73_2 =15'b0;

   // m73_3 = W*in
   wire signed [14:0] m73_3;
   assign m73_3 =15'b0;

   // m73_4 = W*in
   wire signed [14:0] m73_4;
   assign m73_4 =15'b0;

   // m73_5 = W*in
   wire signed [14:0] m73_5;
   assign m73_5 ={ {3{in73[14]}} , in73[14:3] };

   // m73_6 = W*in
   wire signed [14:0] m73_6;
   assign m73_6 =15'b0;

   // m73_7 = W*in
   wire signed [14:0] m73_7;
   assign m73_7 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_8 = W*in
   wire signed [14:0] m73_8;
   assign m73_8 =15'b0;

   // m73_9 = W*in
   wire signed [14:0] m73_9;
   assign m73_9 =15'b0;

   // m73_10 = W*in
   wire signed [14:0] m73_10;
   assign m73_10 =15'b0;

   // m73_11 = W*in
   wire signed [14:0] m73_11;
   assign m73_11 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_12 = W*in
   wire signed [14:0] m73_12;
   assign m73_12 =15'b0;

   // m73_13 = W*in
   wire signed [14:0] m73_13;
   assign m73_13 =15'b0;

   // m73_14 = W*in
   wire signed [14:0] m73_14;
   assign m73_14 =15'b0;

   // m73_15 = W*in
   wire signed [14:0] m73_15;
   assign m73_15 =15'b0;

   // m73_16 = W*in
   wire signed [14:0] m73_16;
   assign m73_16 =15'b0;

   // m73_17 = W*in
   wire signed [14:0] m73_17;
   assign m73_17 =15'b0;

   // m73_18 = W*in
   wire signed [14:0] m73_18;
   assign m73_18 =15'b0;

   // m73_19 = W*in
   wire signed [14:0] m73_19;
   assign m73_19 ={ {4{in73[14]}} , in73[14:4] };

   // m73_20 = W*in
   wire signed [14:0] m73_20;
   assign m73_20 =15'b0;

   // m73_21 = W*in
   wire signed [14:0] m73_21;
   assign m73_21 =15'b0;

   // m73_22 = W*in
   wire signed [14:0] m73_22;
   assign m73_22 ={ {3{in73[14]}} , in73[14:3] };

   // m73_23 = W*in
   wire signed [14:0] m73_23;
   assign m73_23 =15'b0;

   // m73_24 = W*in
   wire signed [14:0] m73_24;
   assign m73_24 =15'b0;

   // m73_25 = W*in
   wire signed [14:0] m73_25;
   assign m73_25 =15'b0;

   // m73_26 = W*in
   wire signed [14:0] m73_26;
   assign m73_26 =15'b0;

   // m73_27 = W*in
   wire signed [14:0] m73_27;
   assign m73_27 =15'b0;

   // m73_28 = W*in
   wire signed [14:0] m73_28;
   assign m73_28 =15'b0;

   // m73_29 = W*in
   wire signed [14:0] m73_29;
   assign m73_29 =15'b0;

   // m73_30 = W*in
   wire signed [14:0] m73_30;
   assign m73_30 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_31 = W*in
   wire signed [14:0] m73_31;
   assign m73_31 =15'b0;

   // m73_32 = W*in
   wire signed [14:0] m73_32;
   assign m73_32 ={ {4{neg73[14]}} , neg73[14:4] };

   // m73_33 = W*in
   wire signed [14:0] m73_33;
   assign m73_33 =15'b0;

   // m73_34 = W*in
   wire signed [14:0] m73_34;
   assign m73_34 =15'b0;

   // m73_35 = W*in
   wire signed [14:0] m73_35;
   assign m73_35 =15'b0;

   // m73_36 = W*in
   wire signed [14:0] m73_36;
   assign m73_36 =15'b0;

   // m73_37 = W*in
   wire signed [14:0] m73_37;
   assign m73_37 =15'b0;

   // m73_38 = W*in
   wire signed [14:0] m73_38;
   assign m73_38 =15'b0;

   // m73_39 = W*in
   wire signed [14:0] m73_39;
   assign m73_39 =15'b0;

   // m73_40 = W*in
   wire signed [14:0] m73_40;
   assign m73_40 ={ {3{in73[14]}} , in73[14:3] };

   // m73_41 = W*in
   wire signed [14:0] m73_41;
   assign m73_41 =15'b0;

   // m73_42 = W*in
   wire signed [14:0] m73_42;
   assign m73_42 =15'b0;

   // m73_43 = W*in
   wire signed [14:0] m73_43;
   assign m73_43 =15'b0;

   // m73_44 = W*in
   wire signed [14:0] m73_44;
   assign m73_44 =15'b0;

   // m73_45 = W*in
   wire signed [14:0] m73_45;
   assign m73_45 =15'b0;

   // m73_46 = W*in
   wire signed [14:0] m73_46;
   assign m73_46 =15'b0;

   // m73_47 = W*in
   wire signed [14:0] m73_47;
   assign m73_47 =15'b0;

   // m73_48 = W*in
   wire signed [14:0] m73_48;
   assign m73_48 =15'b0;

   // m73_49 = W*in
   wire signed [14:0] m73_49;
   assign m73_49 =15'b0;

   // m73_50 = W*in
   wire signed [14:0] m73_50;
   assign m73_50 =15'b0;

   // m73_51 = W*in
   wire signed [14:0] m73_51;
   assign m73_51 =15'b0;

   // m73_52 = W*in
   wire signed [14:0] m73_52;
   assign m73_52 =15'b0;

   // m73_53 = W*in
   wire signed [14:0] m73_53;
   assign m73_53 =15'b0;

   // m73_54 = W*in
   wire signed [14:0] m73_54;
   assign m73_54 =15'b0;

   // m73_55 = W*in
   wire signed [14:0] m73_55;
   assign m73_55 =15'b0;

   // m73_56 = W*in
   wire signed [14:0] m73_56;
   assign m73_56 =15'b0;

   // m73_57 = W*in
   wire signed [14:0] m73_57;
   assign m73_57 ={ {3{in73[14]}} , in73[14:3] };

   // m73_58 = W*in
   wire signed [14:0] m73_58;
   assign m73_58 =15'b0;

   // m73_59 = W*in
   wire signed [14:0] m73_59;
   assign m73_59 =15'b0;

   // m73_60 = W*in
   wire signed [14:0] m73_60;
   assign m73_60 =15'b0;

   // m73_61 = W*in
   wire signed [14:0] m73_61;
   assign m73_61 =15'b0;

   // m73_62 = W*in
   wire signed [14:0] m73_62;
   assign m73_62 =15'b0;

   // m73_63 = W*in
   wire signed [14:0] m73_63;
   assign m73_63 =15'b0;

   // m73_64 = W*in
   wire signed [14:0] m73_64;
   assign m73_64 =15'b0;

   // m73_65 = W*in
   wire signed [14:0] m73_65;
   assign m73_65 =15'b0;

   // m73_66 = W*in
   wire signed [14:0] m73_66;
   assign m73_66 =15'b0;

   // m73_67 = W*in
   wire signed [14:0] m73_67;
   assign m73_67 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_68 = W*in
   wire signed [14:0] m73_68;
   assign m73_68 =15'b0;

   // m73_69 = W*in
   wire signed [14:0] m73_69;
   assign m73_69 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_70 = W*in
   wire signed [14:0] m73_70;
   assign m73_70 =15'b0;

   // m73_71 = W*in
   wire signed [14:0] m73_71;
   assign m73_71 =15'b0;

   // m73_72 = W*in
   wire signed [14:0] m73_72;
   assign m73_72 =15'b0;

   // m73_73 = W*in
   wire signed [14:0] m73_73;
   assign m73_73 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_74 = W*in
   wire signed [14:0] m73_74;
   assign m73_74 ={ {4{in73[14]}} , in73[14:4] };

   // m73_75 = W*in
   wire signed [14:0] m73_75;
   assign m73_75 =15'b0;

   // m73_76 = W*in
   wire signed [14:0] m73_76;
   assign m73_76 =15'b0;

   // m73_77 = W*in
   wire signed [14:0] m73_77;
   assign m73_77 =15'b0;

   // m73_78 = W*in
   wire signed [14:0] m73_78;
   assign m73_78 =15'b0;

   // m73_79 = W*in
   wire signed [14:0] m73_79;
   assign m73_79 =15'b0;

   // m73_80 = W*in
   wire signed [14:0] m73_80;
   assign m73_80 =15'b0;

   // m73_81 = W*in
   wire signed [14:0] m73_81;
   assign m73_81 =15'b0;

   // m73_82 = W*in
   wire signed [14:0] m73_82;
   assign m73_82 =15'b0;

   // m73_83 = W*in
   wire signed [14:0] m73_83;
   assign m73_83 =15'b0;

   // m73_84 = W*in
   wire signed [14:0] m73_84;
   assign m73_84 =15'b0;

   // m73_85 = W*in
   wire signed [14:0] m73_85;
   assign m73_85 =15'b0;

   // m73_86 = W*in
   wire signed [14:0] m73_86;
   assign m73_86 =15'b0;

   // m73_87 = W*in
   wire signed [14:0] m73_87;
   assign m73_87 =15'b0;

   // m73_88 = W*in
   wire signed [14:0] m73_88;
   assign m73_88 =15'b0;

   // m73_89 = W*in
   wire signed [14:0] m73_89;
   assign m73_89 =15'b0;

   // m73_90 = W*in
   wire signed [14:0] m73_90;
   assign m73_90 =15'b0;

   // m73_91 = W*in
   wire signed [14:0] m73_91;
   assign m73_91 ={ {3{in73[14]}} , in73[14:3] };

   // m73_92 = W*in
   wire signed [14:0] m73_92;
   assign m73_92 ={ {3{in73[14]}} , in73[14:3] };

   // m73_93 = W*in
   wire signed [14:0] m73_93;
   assign m73_93 =15'b0;

   // m73_94 = W*in
   wire signed [14:0] m73_94;
   assign m73_94 =15'b0;

   // m73_95 = W*in
   wire signed [14:0] m73_95;
   assign m73_95 ={ {3{neg73[14]}} , neg73[14:3] };

   // m73_96 = W*in
   wire signed [14:0] m73_96;
   assign m73_96 =15'b0;

   // m73_97 = W*in
   wire signed [14:0] m73_97;
   assign m73_97 =15'b0;

   // m73_98 = W*in
   wire signed [14:0] m73_98;
   assign m73_98 =15'b0;

   // m73_99 = W*in
   wire signed [14:0] m73_99;
   assign m73_99 =15'b0;

   // m73_100 = W*in
   wire signed [14:0] m73_100;
   assign m73_100 =15'b0;

   // m74_1 = W*in
   wire signed [14:0] m74_1;
   assign m74_1 =15'b0;

   // m74_2 = W*in
   wire signed [14:0] m74_2;
   assign m74_2 =15'b0;

   // m74_3 = W*in
   wire signed [14:0] m74_3;
   assign m74_3 =15'b0;

   // m74_4 = W*in
   wire signed [14:0] m74_4;
   assign m74_4 =15'b0;

   // m74_5 = W*in
   wire signed [14:0] m74_5;
   assign m74_5 =15'b0;

   // m74_6 = W*in
   wire signed [14:0] m74_6;
   assign m74_6 =15'b0;

   // m74_7 = W*in
   wire signed [14:0] m74_7;
   assign m74_7 =15'b0;

   // m74_8 = W*in
   wire signed [14:0] m74_8;
   assign m74_8 =15'b0;

   // m74_9 = W*in
   wire signed [14:0] m74_9;
   assign m74_9 =15'b0;

   // m74_10 = W*in
   wire signed [14:0] m74_10;
   assign m74_10 =15'b0;

   // m74_11 = W*in
   wire signed [14:0] m74_11;
   assign m74_11 =15'b0;

   // m74_12 = W*in
   wire signed [14:0] m74_12;
   assign m74_12 =15'b0;

   // m74_13 = W*in
   wire signed [14:0] m74_13;
   assign m74_13 =15'b0;

   // m74_14 = W*in
   wire signed [14:0] m74_14;
   assign m74_14 =15'b0;

   // m74_15 = W*in
   wire signed [14:0] m74_15;
   assign m74_15 =15'b0;

   // m74_16 = W*in
   wire signed [14:0] m74_16;
   assign m74_16 =15'b0;

   // m74_17 = W*in
   wire signed [14:0] m74_17;
   assign m74_17 =15'b0;

   // m74_18 = W*in
   wire signed [14:0] m74_18;
   assign m74_18 =15'b0;

   // m74_19 = W*in
   wire signed [14:0] m74_19;
   assign m74_19 =15'b0;

   // m74_20 = W*in
   wire signed [14:0] m74_20;
   assign m74_20 =15'b0;

   // m74_21 = W*in
   wire signed [14:0] m74_21;
   assign m74_21 =15'b0;

   // m74_22 = W*in
   wire signed [14:0] m74_22;
   assign m74_22 =15'b0;

   // m74_23 = W*in
   wire signed [14:0] m74_23;
   assign m74_23 =15'b0;

   // m74_24 = W*in
   wire signed [14:0] m74_24;
   assign m74_24 =15'b0;

   // m74_25 = W*in
   wire signed [14:0] m74_25;
   assign m74_25 =15'b0;

   // m74_26 = W*in
   wire signed [14:0] m74_26;
   assign m74_26 =15'b0;

   // m74_27 = W*in
   wire signed [14:0] m74_27;
   assign m74_27 =15'b0;

   // m74_28 = W*in
   wire signed [14:0] m74_28;
   assign m74_28 =15'b0;

   // m74_29 = W*in
   wire signed [14:0] m74_29;
   assign m74_29 =15'b0;

   // m74_30 = W*in
   wire signed [14:0] m74_30;
   assign m74_30 =15'b0;

   // m74_31 = W*in
   wire signed [14:0] m74_31;
   assign m74_31 ={ {4{neg74[14]}} , neg74[14:4] };

   // m74_32 = W*in
   wire signed [14:0] m74_32;
   assign m74_32 =15'b0;

   // m74_33 = W*in
   wire signed [14:0] m74_33;
   assign m74_33 =15'b0;

   // m74_34 = W*in
   wire signed [14:0] m74_34;
   assign m74_34 =15'b0;

   // m74_35 = W*in
   wire signed [14:0] m74_35;
   assign m74_35 =15'b0;

   // m74_36 = W*in
   wire signed [14:0] m74_36;
   assign m74_36 =15'b0;

   // m74_37 = W*in
   wire signed [14:0] m74_37;
   assign m74_37 =15'b0;

   // m74_38 = W*in
   wire signed [14:0] m74_38;
   assign m74_38 =15'b0;

   // m74_39 = W*in
   wire signed [14:0] m74_39;
   assign m74_39 =15'b0;

   // m74_40 = W*in
   wire signed [14:0] m74_40;
   assign m74_40 =15'b0;

   // m74_41 = W*in
   wire signed [14:0] m74_41;
   assign m74_41 =15'b0;

   // m74_42 = W*in
   wire signed [14:0] m74_42;
   assign m74_42 ={ {4{neg74[14]}} , neg74[14:4] };

   // m74_43 = W*in
   wire signed [14:0] m74_43;
   assign m74_43 =15'b0;

   // m74_44 = W*in
   wire signed [14:0] m74_44;
   assign m74_44 =15'b0;

   // m74_45 = W*in
   wire signed [14:0] m74_45;
   assign m74_45 =15'b0;

   // m74_46 = W*in
   wire signed [14:0] m74_46;
   assign m74_46 =15'b0;

   // m74_47 = W*in
   wire signed [14:0] m74_47;
   assign m74_47 =15'b0;

   // m74_48 = W*in
   wire signed [14:0] m74_48;
   assign m74_48 =15'b0;

   // m74_49 = W*in
   wire signed [14:0] m74_49;
   assign m74_49 =15'b0;

   // m74_50 = W*in
   wire signed [14:0] m74_50;
   assign m74_50 =15'b0;

   // m74_51 = W*in
   wire signed [14:0] m74_51;
   assign m74_51 =15'b0;

   // m74_52 = W*in
   wire signed [14:0] m74_52;
   assign m74_52 =15'b0;

   // m74_53 = W*in
   wire signed [14:0] m74_53;
   assign m74_53 =15'b0;

   // m74_54 = W*in
   wire signed [14:0] m74_54;
   assign m74_54 =15'b0;

   // m74_55 = W*in
   wire signed [14:0] m74_55;
   assign m74_55 =15'b0;

   // m74_56 = W*in
   wire signed [14:0] m74_56;
   assign m74_56 =15'b0;

   // m74_57 = W*in
   wire signed [14:0] m74_57;
   assign m74_57 =15'b0;

   // m74_58 = W*in
   wire signed [14:0] m74_58;
   assign m74_58 =15'b0;

   // m74_59 = W*in
   wire signed [14:0] m74_59;
   assign m74_59 =15'b0;

   // m74_60 = W*in
   wire signed [14:0] m74_60;
   assign m74_60 =15'b0;

   // m74_61 = W*in
   wire signed [14:0] m74_61;
   assign m74_61 =15'b0;

   // m74_62 = W*in
   wire signed [14:0] m74_62;
   assign m74_62 =15'b0;

   // m74_63 = W*in
   wire signed [14:0] m74_63;
   assign m74_63 =15'b0;

   // m74_64 = W*in
   wire signed [14:0] m74_64;
   assign m74_64 ={ {4{neg74[14]}} , neg74[14:4] };

   // m74_65 = W*in
   wire signed [14:0] m74_65;
   assign m74_65 =15'b0;

   // m74_66 = W*in
   wire signed [14:0] m74_66;
   assign m74_66 =15'b0;

   // m74_67 = W*in
   wire signed [14:0] m74_67;
   assign m74_67 ={ {3{neg74[14]}} , neg74[14:3] };

   // m74_68 = W*in
   wire signed [14:0] m74_68;
   assign m74_68 =15'b0;

   // m74_69 = W*in
   wire signed [14:0] m74_69;
   assign m74_69 =15'b0;

   // m74_70 = W*in
   wire signed [14:0] m74_70;
   assign m74_70 =15'b0;

   // m74_71 = W*in
   wire signed [14:0] m74_71;
   assign m74_71 =15'b0;

   // m74_72 = W*in
   wire signed [14:0] m74_72;
   assign m74_72 =15'b0;

   // m74_73 = W*in
   wire signed [14:0] m74_73;
   assign m74_73 =15'b0;

   // m74_74 = W*in
   wire signed [14:0] m74_74;
   assign m74_74 ={ {4{neg74[14]}} , neg74[14:4] };

   // m74_75 = W*in
   wire signed [14:0] m74_75;
   assign m74_75 ={ {4{in74[14]}} , in74[14:4] };

   // m74_76 = W*in
   wire signed [14:0] m74_76;
   assign m74_76 ={ {3{neg74[14]}} , neg74[14:3] };

   // m74_77 = W*in
   wire signed [14:0] m74_77;
   assign m74_77 =15'b0;

   // m74_78 = W*in
   wire signed [14:0] m74_78;
   assign m74_78 =15'b0;

   // m74_79 = W*in
   wire signed [14:0] m74_79;
   assign m74_79 =15'b0;

   // m74_80 = W*in
   wire signed [14:0] m74_80;
   assign m74_80 =15'b0;

   // m74_81 = W*in
   wire signed [14:0] m74_81;
   assign m74_81 =15'b0;

   // m74_82 = W*in
   wire signed [14:0] m74_82;
   assign m74_82 =15'b0;

   // m74_83 = W*in
   wire signed [14:0] m74_83;
   assign m74_83 =15'b0;

   // m74_84 = W*in
   wire signed [14:0] m74_84;
   assign m74_84 =15'b0;

   // m74_85 = W*in
   wire signed [14:0] m74_85;
   assign m74_85 =15'b0;

   // m74_86 = W*in
   wire signed [14:0] m74_86;
   assign m74_86 =15'b0;

   // m74_87 = W*in
   wire signed [14:0] m74_87;
   assign m74_87 =15'b0;

   // m74_88 = W*in
   wire signed [14:0] m74_88;
   assign m74_88 =15'b0;

   // m74_89 = W*in
   wire signed [14:0] m74_89;
   assign m74_89 =15'b0;

   // m74_90 = W*in
   wire signed [14:0] m74_90;
   assign m74_90 =15'b0;

   // m74_91 = W*in
   wire signed [14:0] m74_91;
   assign m74_91 ={ {3{in74[14]}} , in74[14:3] };

   // m74_92 = W*in
   wire signed [14:0] m74_92;
   assign m74_92 ={ {3{in74[14]}} , in74[14:3] };

   // m74_93 = W*in
   wire signed [14:0] m74_93;
   assign m74_93 =15'b0;

   // m74_94 = W*in
   wire signed [14:0] m74_94;
   assign m74_94 =15'b0;

   // m74_95 = W*in
   wire signed [14:0] m74_95;
   assign m74_95 =15'b0;

   // m74_96 = W*in
   wire signed [14:0] m74_96;
   assign m74_96 =15'b0;

   // m74_97 = W*in
   wire signed [14:0] m74_97;
   assign m74_97 =15'b0;

   // m74_98 = W*in
   wire signed [14:0] m74_98;
   assign m74_98 ={ {4{neg74[14]}} , neg74[14:4] };

   // m74_99 = W*in
   wire signed [14:0] m74_99;
   assign m74_99 =15'b0;

   // m74_100 = W*in
   wire signed [14:0] m74_100;
   assign m74_100 =15'b0;

   // m75_1 = W*in
   wire signed [14:0] m75_1;
   assign m75_1 =15'b0;

   // m75_2 = W*in
   wire signed [14:0] m75_2;
   assign m75_2 =15'b0;

   // m75_3 = W*in
   wire signed [14:0] m75_3;
   assign m75_3 =15'b0;

   // m75_4 = W*in
   wire signed [14:0] m75_4;
   assign m75_4 =15'b0;

   // m75_5 = W*in
   wire signed [14:0] m75_5;
   assign m75_5 =15'b0;

   // m75_6 = W*in
   wire signed [14:0] m75_6;
   assign m75_6 =15'b0;

   // m75_7 = W*in
   wire signed [14:0] m75_7;
   assign m75_7 =15'b0;

   // m75_8 = W*in
   wire signed [14:0] m75_8;
   assign m75_8 =15'b0;

   // m75_9 = W*in
   wire signed [14:0] m75_9;
   assign m75_9 =15'b0;

   // m75_10 = W*in
   wire signed [14:0] m75_10;
   assign m75_10 =15'b0;

   // m75_11 = W*in
   wire signed [14:0] m75_11;
   assign m75_11 =15'b0;

   // m75_12 = W*in
   wire signed [14:0] m75_12;
   assign m75_12 =15'b0;

   // m75_13 = W*in
   wire signed [14:0] m75_13;
   assign m75_13 =15'b0;

   // m75_14 = W*in
   wire signed [14:0] m75_14;
   assign m75_14 =15'b0;

   // m75_15 = W*in
   wire signed [14:0] m75_15;
   assign m75_15 =15'b0;

   // m75_16 = W*in
   wire signed [14:0] m75_16;
   assign m75_16 =15'b0;

   // m75_17 = W*in
   wire signed [14:0] m75_17;
   assign m75_17 =15'b0;

   // m75_18 = W*in
   wire signed [14:0] m75_18;
   assign m75_18 =15'b0;

   // m75_19 = W*in
   wire signed [14:0] m75_19;
   assign m75_19 =15'b0;

   // m75_20 = W*in
   wire signed [14:0] m75_20;
   assign m75_20 =15'b0;

   // m75_21 = W*in
   wire signed [14:0] m75_21;
   assign m75_21 ={ {4{neg75[14]}} , neg75[14:4] };

   // m75_22 = W*in
   wire signed [14:0] m75_22;
   assign m75_22 ={ {4{neg75[14]}} , neg75[14:4] };

   // m75_23 = W*in
   wire signed [14:0] m75_23;
   assign m75_23 =15'b0;

   // m75_24 = W*in
   wire signed [14:0] m75_24;
   assign m75_24 =15'b0;

   // m75_25 = W*in
   wire signed [14:0] m75_25;
   assign m75_25 =15'b0;

   // m75_26 = W*in
   wire signed [14:0] m75_26;
   assign m75_26 ={ {3{neg75[14]}} , neg75[14:3] };

   // m75_27 = W*in
   wire signed [14:0] m75_27;
   assign m75_27 =15'b0;

   // m75_28 = W*in
   wire signed [14:0] m75_28;
   assign m75_28 =15'b0;

   // m75_29 = W*in
   wire signed [14:0] m75_29;
   assign m75_29 ={ {3{neg75[14]}} , neg75[14:3] };

   // m75_30 = W*in
   wire signed [14:0] m75_30;
   assign m75_30 =15'b0;

   // m75_31 = W*in
   wire signed [14:0] m75_31;
   assign m75_31 =15'b0;

   // m75_32 = W*in
   wire signed [14:0] m75_32;
   assign m75_32 =15'b0;

   // m75_33 = W*in
   wire signed [14:0] m75_33;
   assign m75_33 =15'b0;

   // m75_34 = W*in
   wire signed [14:0] m75_34;
   assign m75_34 =15'b0;

   // m75_35 = W*in
   wire signed [14:0] m75_35;
   assign m75_35 ={ {2{in75[14]}} , in75[14:2] };

   // m75_36 = W*in
   wire signed [14:0] m75_36;
   assign m75_36 =15'b0;

   // m75_37 = W*in
   wire signed [14:0] m75_37;
   assign m75_37 =15'b0;

   // m75_38 = W*in
   wire signed [14:0] m75_38;
   assign m75_38 =15'b0;

   // m75_39 = W*in
   wire signed [14:0] m75_39;
   assign m75_39 =15'b0;

   // m75_40 = W*in
   wire signed [14:0] m75_40;
   assign m75_40 =15'b0;

   // m75_41 = W*in
   wire signed [14:0] m75_41;
   assign m75_41 =15'b0;

   // m75_42 = W*in
   wire signed [14:0] m75_42;
   assign m75_42 =15'b0;

   // m75_43 = W*in
   wire signed [14:0] m75_43;
   assign m75_43 =15'b0;

   // m75_44 = W*in
   wire signed [14:0] m75_44;
   assign m75_44 =15'b0;

   // m75_45 = W*in
   wire signed [14:0] m75_45;
   assign m75_45 =15'b0;

   // m75_46 = W*in
   wire signed [14:0] m75_46;
   assign m75_46 =15'b0;

   // m75_47 = W*in
   wire signed [14:0] m75_47;
   assign m75_47 =15'b0;

   // m75_48 = W*in
   wire signed [14:0] m75_48;
   assign m75_48 ={ {3{in75[14]}} , in75[14:3] };

   // m75_49 = W*in
   wire signed [14:0] m75_49;
   assign m75_49 =15'b0;

   // m75_50 = W*in
   wire signed [14:0] m75_50;
   assign m75_50 =15'b0;

   // m75_51 = W*in
   wire signed [14:0] m75_51;
   assign m75_51 =15'b0;

   // m75_52 = W*in
   wire signed [14:0] m75_52;
   assign m75_52 =15'b0;

   // m75_53 = W*in
   wire signed [14:0] m75_53;
   assign m75_53 =15'b0;

   // m75_54 = W*in
   wire signed [14:0] m75_54;
   assign m75_54 =15'b0;

   // m75_55 = W*in
   wire signed [14:0] m75_55;
   assign m75_55 =15'b0;

   // m75_56 = W*in
   wire signed [14:0] m75_56;
   assign m75_56 =15'b0;

   // m75_57 = W*in
   wire signed [14:0] m75_57;
   assign m75_57 =15'b0;

   // m75_58 = W*in
   wire signed [14:0] m75_58;
   assign m75_58 =15'b0;

   // m75_59 = W*in
   wire signed [14:0] m75_59;
   assign m75_59 =15'b0;

   // m75_60 = W*in
   wire signed [14:0] m75_60;
   assign m75_60 ={ {3{neg75[14]}} , neg75[14:3] };

   // m75_61 = W*in
   wire signed [14:0] m75_61;
   assign m75_61 =15'b0;

   // m75_62 = W*in
   wire signed [14:0] m75_62;
   assign m75_62 =15'b0;

   // m75_63 = W*in
   wire signed [14:0] m75_63;
   assign m75_63 =15'b0;

   // m75_64 = W*in
   wire signed [14:0] m75_64;
   assign m75_64 =15'b0;

   // m75_65 = W*in
   wire signed [14:0] m75_65;
   assign m75_65 ={ {3{neg75[14]}} , neg75[14:3] };

   // m75_66 = W*in
   wire signed [14:0] m75_66;
   assign m75_66 ={ {3{in75[14]}} , in75[14:3] };

   // m75_67 = W*in
   wire signed [14:0] m75_67;
   assign m75_67 =15'b0;

   // m75_68 = W*in
   wire signed [14:0] m75_68;
   assign m75_68 =15'b0;

   // m75_69 = W*in
   wire signed [14:0] m75_69;
   assign m75_69 =15'b0;

   // m75_70 = W*in
   wire signed [14:0] m75_70;
   assign m75_70 =15'b0;

   // m75_71 = W*in
   wire signed [14:0] m75_71;
   assign m75_71 =15'b0;

   // m75_72 = W*in
   wire signed [14:0] m75_72;
   assign m75_72 =15'b0;

   // m75_73 = W*in
   wire signed [14:0] m75_73;
   assign m75_73 =15'b0;

   // m75_74 = W*in
   wire signed [14:0] m75_74;
   assign m75_74 =15'b0;

   // m75_75 = W*in
   wire signed [14:0] m75_75;
   assign m75_75 =15'b0;

   // m75_76 = W*in
   wire signed [14:0] m75_76;
   assign m75_76 =15'b0;

   // m75_77 = W*in
   wire signed [14:0] m75_77;
   assign m75_77 =15'b0;

   // m75_78 = W*in
   wire signed [14:0] m75_78;
   assign m75_78 =15'b0;

   // m75_79 = W*in
   wire signed [14:0] m75_79;
   assign m75_79 =15'b0;

   // m75_80 = W*in
   wire signed [14:0] m75_80;
   assign m75_80 =15'b0;

   // m75_81 = W*in
   wire signed [14:0] m75_81;
   assign m75_81 =15'b0;

   // m75_82 = W*in
   wire signed [14:0] m75_82;
   assign m75_82 =15'b0;

   // m75_83 = W*in
   wire signed [14:0] m75_83;
   assign m75_83 =15'b0;

   // m75_84 = W*in
   wire signed [14:0] m75_84;
   assign m75_84 =15'b0;

   // m75_85 = W*in
   wire signed [14:0] m75_85;
   assign m75_85 =15'b0;

   // m75_86 = W*in
   wire signed [14:0] m75_86;
   assign m75_86 =15'b0;

   // m75_87 = W*in
   wire signed [14:0] m75_87;
   assign m75_87 =15'b0;

   // m75_88 = W*in
   wire signed [14:0] m75_88;
   assign m75_88 =15'b0;

   // m75_89 = W*in
   wire signed [14:0] m75_89;
   assign m75_89 =15'b0;

   // m75_90 = W*in
   wire signed [14:0] m75_90;
   assign m75_90 =15'b0;

   // m75_91 = W*in
   wire signed [14:0] m75_91;
   assign m75_91 =15'b0;

   // m75_92 = W*in
   wire signed [14:0] m75_92;
   assign m75_92 =15'b0;

   // m75_93 = W*in
   wire signed [14:0] m75_93;
   assign m75_93 ={ {3{neg75[14]}} , neg75[14:3] };

   // m75_94 = W*in
   wire signed [14:0] m75_94;
   assign m75_94 =15'b0;

   // m75_95 = W*in
   wire signed [14:0] m75_95;
   assign m75_95 =15'b0;

   // m75_96 = W*in
   wire signed [14:0] m75_96;
   assign m75_96 =15'b0;

   // m75_97 = W*in
   wire signed [14:0] m75_97;
   assign m75_97 ={ {3{neg75[14]}} , neg75[14:3] };

   // m75_98 = W*in
   wire signed [14:0] m75_98;
   assign m75_98 =15'b0;

   // m75_99 = W*in
   wire signed [14:0] m75_99;
   assign m75_99 =15'b0;

   // m75_100 = W*in
   wire signed [14:0] m75_100;
   assign m75_100 =15'b0;

   // m76_1 = W*in
   wire signed [14:0] m76_1;
   assign m76_1 =15'b0;

   // m76_2 = W*in
   wire signed [14:0] m76_2;
   assign m76_2 =15'b0;

   // m76_3 = W*in
   wire signed [14:0] m76_3;
   assign m76_3 =15'b0;

   // m76_4 = W*in
   wire signed [14:0] m76_4;
   assign m76_4 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_5 = W*in
   wire signed [14:0] m76_5;
   assign m76_5 =15'b0;

   // m76_6 = W*in
   wire signed [14:0] m76_6;
   assign m76_6 ={ {4{neg76[14]}} , neg76[14:4] };

   // m76_7 = W*in
   wire signed [14:0] m76_7;
   assign m76_7 =15'b0;

   // m76_8 = W*in
   wire signed [14:0] m76_8;
   assign m76_8 =15'b0;

   // m76_9 = W*in
   wire signed [14:0] m76_9;
   assign m76_9 =15'b0;

   // m76_10 = W*in
   wire signed [14:0] m76_10;
   assign m76_10 =15'b0;

   // m76_11 = W*in
   wire signed [14:0] m76_11;
   assign m76_11 =15'b0;

   // m76_12 = W*in
   wire signed [14:0] m76_12;
   assign m76_12 =15'b0;

   // m76_13 = W*in
   wire signed [14:0] m76_13;
   assign m76_13 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_14 = W*in
   wire signed [14:0] m76_14;
   assign m76_14 =15'b0;

   // m76_15 = W*in
   wire signed [14:0] m76_15;
   assign m76_15 =15'b0;

   // m76_16 = W*in
   wire signed [14:0] m76_16;
   assign m76_16 =15'b0;

   // m76_17 = W*in
   wire signed [14:0] m76_17;
   assign m76_17 ={ {4{in76[14]}} , in76[14:4] };

   // m76_18 = W*in
   wire signed [14:0] m76_18;
   assign m76_18 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_19 = W*in
   wire signed [14:0] m76_19;
   assign m76_19 ={ {3{in76[14]}} , in76[14:3] };

   // m76_20 = W*in
   wire signed [14:0] m76_20;
   assign m76_20 =15'b0;

   // m76_21 = W*in
   wire signed [14:0] m76_21;
   assign m76_21 =15'b0;

   // m76_22 = W*in
   wire signed [14:0] m76_22;
   assign m76_22 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_23 = W*in
   wire signed [14:0] m76_23;
   assign m76_23 =15'b0;

   // m76_24 = W*in
   wire signed [14:0] m76_24;
   assign m76_24 ={ {3{in76[14]}} , in76[14:3] };

   // m76_25 = W*in
   wire signed [14:0] m76_25;
   assign m76_25 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_26 = W*in
   wire signed [14:0] m76_26;
   assign m76_26 =15'b0;

   // m76_27 = W*in
   wire signed [14:0] m76_27;
   assign m76_27 =15'b0;

   // m76_28 = W*in
   wire signed [14:0] m76_28;
   assign m76_28 =15'b0;

   // m76_29 = W*in
   wire signed [14:0] m76_29;
   assign m76_29 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_30 = W*in
   wire signed [14:0] m76_30;
   assign m76_30 =15'b0;

   // m76_31 = W*in
   wire signed [14:0] m76_31;
   assign m76_31 =15'b0;

   // m76_32 = W*in
   wire signed [14:0] m76_32;
   assign m76_32 ={ {3{in76[14]}} , in76[14:3] };

   // m76_33 = W*in
   wire signed [14:0] m76_33;
   assign m76_33 ={ {4{in76[14]}} , in76[14:4] };

   // m76_34 = W*in
   wire signed [14:0] m76_34;
   assign m76_34 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_35 = W*in
   wire signed [14:0] m76_35;
   assign m76_35 ={ {3{in76[14]}} , in76[14:3] };

   // m76_36 = W*in
   wire signed [14:0] m76_36;
   assign m76_36 =15'b0;

   // m76_37 = W*in
   wire signed [14:0] m76_37;
   assign m76_37 =15'b0;

   // m76_38 = W*in
   wire signed [14:0] m76_38;
   assign m76_38 =15'b0;

   // m76_39 = W*in
   wire signed [14:0] m76_39;
   assign m76_39 =15'b0;

   // m76_40 = W*in
   wire signed [14:0] m76_40;
   assign m76_40 ={ {3{in76[14]}} , in76[14:3] };

   // m76_41 = W*in
   wire signed [14:0] m76_41;
   assign m76_41 =15'b0;

   // m76_42 = W*in
   wire signed [14:0] m76_42;
   assign m76_42 ={ {2{in76[14]}} , in76[14:2] };

   // m76_43 = W*in
   wire signed [14:0] m76_43;
   assign m76_43 =15'b0;

   // m76_44 = W*in
   wire signed [14:0] m76_44;
   assign m76_44 =15'b0;

   // m76_45 = W*in
   wire signed [14:0] m76_45;
   assign m76_45 =15'b0;

   // m76_46 = W*in
   wire signed [14:0] m76_46;
   assign m76_46 =15'b0;

   // m76_47 = W*in
   wire signed [14:0] m76_47;
   assign m76_47 ={ {4{in76[14]}} , in76[14:4] };

   // m76_48 = W*in
   wire signed [14:0] m76_48;
   assign m76_48 =15'b0;

   // m76_49 = W*in
   wire signed [14:0] m76_49;
   assign m76_49 =15'b0;

   // m76_50 = W*in
   wire signed [14:0] m76_50;
   assign m76_50 =15'b0;

   // m76_51 = W*in
   wire signed [14:0] m76_51;
   assign m76_51 =15'b0;

   // m76_52 = W*in
   wire signed [14:0] m76_52;
   assign m76_52 =15'b0;

   // m76_53 = W*in
   wire signed [14:0] m76_53;
   assign m76_53 =15'b0;

   // m76_54 = W*in
   wire signed [14:0] m76_54;
   assign m76_54 =15'b0;

   // m76_55 = W*in
   wire signed [14:0] m76_55;
   assign m76_55 =15'b0;

   // m76_56 = W*in
   wire signed [14:0] m76_56;
   assign m76_56 ={ {3{in76[14]}} , in76[14:3] };

   // m76_57 = W*in
   wire signed [14:0] m76_57;
   assign m76_57 ={ {3{in76[14]}} , in76[14:3] };

   // m76_58 = W*in
   wire signed [14:0] m76_58;
   assign m76_58 ={ {4{neg76[14]}} , neg76[14:4] };

   // m76_59 = W*in
   wire signed [14:0] m76_59;
   assign m76_59 ={ {4{in76[14]}} , in76[14:4] };

   // m76_60 = W*in
   wire signed [14:0] m76_60;
   assign m76_60 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_61 = W*in
   wire signed [14:0] m76_61;
   assign m76_61 ={ {4{neg76[14]}} , neg76[14:4] };

   // m76_62 = W*in
   wire signed [14:0] m76_62;
   assign m76_62 =15'b0;

   // m76_63 = W*in
   wire signed [14:0] m76_63;
   assign m76_63 =15'b0;

   // m76_64 = W*in
   wire signed [14:0] m76_64;
   assign m76_64 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_65 = W*in
   wire signed [14:0] m76_65;
   assign m76_65 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_66 = W*in
   wire signed [14:0] m76_66;
   assign m76_66 ={ {4{in76[14]}} , in76[14:4] };

   // m76_67 = W*in
   wire signed [14:0] m76_67;
   assign m76_67 ={ {4{in76[14]}} , in76[14:4] };

   // m76_68 = W*in
   wire signed [14:0] m76_68;
   assign m76_68 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_69 = W*in
   wire signed [14:0] m76_69;
   assign m76_69 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_70 = W*in
   wire signed [14:0] m76_70;
   assign m76_70 ={ {3{in76[14]}} , in76[14:3] };

   // m76_71 = W*in
   wire signed [14:0] m76_71;
   assign m76_71 =15'b0;

   // m76_72 = W*in
   wire signed [14:0] m76_72;
   assign m76_72 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_73 = W*in
   wire signed [14:0] m76_73;
   assign m76_73 =15'b0;

   // m76_74 = W*in
   wire signed [14:0] m76_74;
   assign m76_74 =15'b0;

   // m76_75 = W*in
   wire signed [14:0] m76_75;
   assign m76_75 =15'b0;

   // m76_76 = W*in
   wire signed [14:0] m76_76;
   assign m76_76 =15'b0;

   // m76_77 = W*in
   wire signed [14:0] m76_77;
   assign m76_77 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_78 = W*in
   wire signed [14:0] m76_78;
   assign m76_78 =15'b0;

   // m76_79 = W*in
   wire signed [14:0] m76_79;
   assign m76_79 =15'b0;

   // m76_80 = W*in
   wire signed [14:0] m76_80;
   assign m76_80 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_81 = W*in
   wire signed [14:0] m76_81;
   assign m76_81 =15'b0;

   // m76_82 = W*in
   wire signed [14:0] m76_82;
   assign m76_82 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_83 = W*in
   wire signed [14:0] m76_83;
   assign m76_83 =15'b0;

   // m76_84 = W*in
   wire signed [14:0] m76_84;
   assign m76_84 =15'b0;

   // m76_85 = W*in
   wire signed [14:0] m76_85;
   assign m76_85 =15'b0;

   // m76_86 = W*in
   wire signed [14:0] m76_86;
   assign m76_86 =15'b0;

   // m76_87 = W*in
   wire signed [14:0] m76_87;
   assign m76_87 =15'b0;

   // m76_88 = W*in
   wire signed [14:0] m76_88;
   assign m76_88 =15'b0;

   // m76_89 = W*in
   wire signed [14:0] m76_89;
   assign m76_89 ={ {3{in76[14]}} , in76[14:3] };

   // m76_90 = W*in
   wire signed [14:0] m76_90;
   assign m76_90 =15'b0;

   // m76_91 = W*in
   wire signed [14:0] m76_91;
   assign m76_91 =15'b0;

   // m76_92 = W*in
   wire signed [14:0] m76_92;
   assign m76_92 ={ {3{neg76[14]}} , neg76[14:3] };

   // m76_93 = W*in
   wire signed [14:0] m76_93;
   assign m76_93 =15'b0;

   // m76_94 = W*in
   wire signed [14:0] m76_94;
   assign m76_94 =15'b0;

   // m76_95 = W*in
   wire signed [14:0] m76_95;
   assign m76_95 =15'b0;

   // m76_96 = W*in
   wire signed [14:0] m76_96;
   assign m76_96 =15'b0;

   // m76_97 = W*in
   wire signed [14:0] m76_97;
   assign m76_97 =15'b0;

   // m76_98 = W*in
   wire signed [14:0] m76_98;
   assign m76_98 ={ {3{in76[14]}} , in76[14:3] };

   // m76_99 = W*in
   wire signed [14:0] m76_99;
   assign m76_99 =15'b0;

   // m76_100 = W*in
   wire signed [14:0] m76_100;
   assign m76_100 =15'b0;

   // m77_1 = W*in
   wire signed [14:0] m77_1;
   assign m77_1 =15'b0;

   // m77_2 = W*in
   wire signed [14:0] m77_2;
   assign m77_2 =15'b0;

   // m77_3 = W*in
   wire signed [14:0] m77_3;
   assign m77_3 =15'b0;

   // m77_4 = W*in
   wire signed [14:0] m77_4;
   assign m77_4 =15'b0;

   // m77_5 = W*in
   wire signed [14:0] m77_5;
   assign m77_5 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_6 = W*in
   wire signed [14:0] m77_6;
   assign m77_6 =15'b0;

   // m77_7 = W*in
   wire signed [14:0] m77_7;
   assign m77_7 =15'b0;

   // m77_8 = W*in
   wire signed [14:0] m77_8;
   assign m77_8 =15'b0;

   // m77_9 = W*in
   wire signed [14:0] m77_9;
   assign m77_9 =15'b0;

   // m77_10 = W*in
   wire signed [14:0] m77_10;
   assign m77_10 =15'b0;

   // m77_11 = W*in
   wire signed [14:0] m77_11;
   assign m77_11 =15'b0;

   // m77_12 = W*in
   wire signed [14:0] m77_12;
   assign m77_12 =15'b0;

   // m77_13 = W*in
   wire signed [14:0] m77_13;
   assign m77_13 =15'b0;

   // m77_14 = W*in
   wire signed [14:0] m77_14;
   assign m77_14 =15'b0;

   // m77_15 = W*in
   wire signed [14:0] m77_15;
   assign m77_15 =15'b0;

   // m77_16 = W*in
   wire signed [14:0] m77_16;
   assign m77_16 =15'b0;

   // m77_17 = W*in
   wire signed [14:0] m77_17;
   assign m77_17 ={ {3{in77[14]}} , in77[14:3] };

   // m77_18 = W*in
   wire signed [14:0] m77_18;
   assign m77_18 =15'b0;

   // m77_19 = W*in
   wire signed [14:0] m77_19;
   assign m77_19 =15'b0;

   // m77_20 = W*in
   wire signed [14:0] m77_20;
   assign m77_20 =15'b0;

   // m77_21 = W*in
   wire signed [14:0] m77_21;
   assign m77_21 =15'b0;

   // m77_22 = W*in
   wire signed [14:0] m77_22;
   assign m77_22 =15'b0;

   // m77_23 = W*in
   wire signed [14:0] m77_23;
   assign m77_23 ={ {4{in77[14]}} , in77[14:4] };

   // m77_24 = W*in
   wire signed [14:0] m77_24;
   assign m77_24 =15'b0;

   // m77_25 = W*in
   wire signed [14:0] m77_25;
   assign m77_25 =15'b0;

   // m77_26 = W*in
   wire signed [14:0] m77_26;
   assign m77_26 =15'b0;

   // m77_27 = W*in
   wire signed [14:0] m77_27;
   assign m77_27 =15'b0;

   // m77_28 = W*in
   wire signed [14:0] m77_28;
   assign m77_28 =15'b0;

   // m77_29 = W*in
   wire signed [14:0] m77_29;
   assign m77_29 =15'b0;

   // m77_30 = W*in
   wire signed [14:0] m77_30;
   assign m77_30 =15'b0;

   // m77_31 = W*in
   wire signed [14:0] m77_31;
   assign m77_31 =15'b0;

   // m77_32 = W*in
   wire signed [14:0] m77_32;
   assign m77_32 =15'b0;

   // m77_33 = W*in
   wire signed [14:0] m77_33;
   assign m77_33 =15'b0;

   // m77_34 = W*in
   wire signed [14:0] m77_34;
   assign m77_34 =15'b0;

   // m77_35 = W*in
   wire signed [14:0] m77_35;
   assign m77_35 =15'b0;

   // m77_36 = W*in
   wire signed [14:0] m77_36;
   assign m77_36 =15'b0;

   // m77_37 = W*in
   wire signed [14:0] m77_37;
   assign m77_37 =15'b0;

   // m77_38 = W*in
   wire signed [14:0] m77_38;
   assign m77_38 =15'b0;

   // m77_39 = W*in
   wire signed [14:0] m77_39;
   assign m77_39 =15'b0;

   // m77_40 = W*in
   wire signed [14:0] m77_40;
   assign m77_40 ={ {4{neg77[14]}} , neg77[14:4] };

   // m77_41 = W*in
   wire signed [14:0] m77_41;
   assign m77_41 =15'b0;

   // m77_42 = W*in
   wire signed [14:0] m77_42;
   assign m77_42 =15'b0;

   // m77_43 = W*in
   wire signed [14:0] m77_43;
   assign m77_43 =15'b0;

   // m77_44 = W*in
   wire signed [14:0] m77_44;
   assign m77_44 =15'b0;

   // m77_45 = W*in
   wire signed [14:0] m77_45;
   assign m77_45 =15'b0;

   // m77_46 = W*in
   wire signed [14:0] m77_46;
   assign m77_46 =15'b0;

   // m77_47 = W*in
   wire signed [14:0] m77_47;
   assign m77_47 =15'b0;

   // m77_48 = W*in
   wire signed [14:0] m77_48;
   assign m77_48 =15'b0;

   // m77_49 = W*in
   wire signed [14:0] m77_49;
   assign m77_49 =15'b0;

   // m77_50 = W*in
   wire signed [14:0] m77_50;
   assign m77_50 =15'b0;

   // m77_51 = W*in
   wire signed [14:0] m77_51;
   assign m77_51 =15'b0;

   // m77_52 = W*in
   wire signed [14:0] m77_52;
   assign m77_52 =15'b0;

   // m77_53 = W*in
   wire signed [14:0] m77_53;
   assign m77_53 =15'b0;

   // m77_54 = W*in
   wire signed [14:0] m77_54;
   assign m77_54 =15'b0;

   // m77_55 = W*in
   wire signed [14:0] m77_55;
   assign m77_55 =15'b0;

   // m77_56 = W*in
   wire signed [14:0] m77_56;
   assign m77_56 ={ {3{in77[14]}} , in77[14:3] };

   // m77_57 = W*in
   wire signed [14:0] m77_57;
   assign m77_57 ={ {4{neg77[14]}} , neg77[14:4] };

   // m77_58 = W*in
   wire signed [14:0] m77_58;
   assign m77_58 =15'b0;

   // m77_59 = W*in
   wire signed [14:0] m77_59;
   assign m77_59 =15'b0;

   // m77_60 = W*in
   wire signed [14:0] m77_60;
   assign m77_60 =15'b0;

   // m77_61 = W*in
   wire signed [14:0] m77_61;
   assign m77_61 =15'b0;

   // m77_62 = W*in
   wire signed [14:0] m77_62;
   assign m77_62 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_63 = W*in
   wire signed [14:0] m77_63;
   assign m77_63 =15'b0;

   // m77_64 = W*in
   wire signed [14:0] m77_64;
   assign m77_64 ={ {4{in77[14]}} , in77[14:4] };

   // m77_65 = W*in
   wire signed [14:0] m77_65;
   assign m77_65 =15'b0;

   // m77_66 = W*in
   wire signed [14:0] m77_66;
   assign m77_66 =15'b0;

   // m77_67 = W*in
   wire signed [14:0] m77_67;
   assign m77_67 =15'b0;

   // m77_68 = W*in
   wire signed [14:0] m77_68;
   assign m77_68 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_69 = W*in
   wire signed [14:0] m77_69;
   assign m77_69 =15'b0;

   // m77_70 = W*in
   wire signed [14:0] m77_70;
   assign m77_70 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_71 = W*in
   wire signed [14:0] m77_71;
   assign m77_71 =15'b0;

   // m77_72 = W*in
   wire signed [14:0] m77_72;
   assign m77_72 =15'b0;

   // m77_73 = W*in
   wire signed [14:0] m77_73;
   assign m77_73 =15'b0;

   // m77_74 = W*in
   wire signed [14:0] m77_74;
   assign m77_74 =15'b0;

   // m77_75 = W*in
   wire signed [14:0] m77_75;
   assign m77_75 =15'b0;

   // m77_76 = W*in
   wire signed [14:0] m77_76;
   assign m77_76 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_77 = W*in
   wire signed [14:0] m77_77;
   assign m77_77 =15'b0;

   // m77_78 = W*in
   wire signed [14:0] m77_78;
   assign m77_78 =15'b0;

   // m77_79 = W*in
   wire signed [14:0] m77_79;
   assign m77_79 ={ {4{neg77[14]}} , neg77[14:4] };

   // m77_80 = W*in
   wire signed [14:0] m77_80;
   assign m77_80 =15'b0;

   // m77_81 = W*in
   wire signed [14:0] m77_81;
   assign m77_81 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_82 = W*in
   wire signed [14:0] m77_82;
   assign m77_82 =15'b0;

   // m77_83 = W*in
   wire signed [14:0] m77_83;
   assign m77_83 =15'b0;

   // m77_84 = W*in
   wire signed [14:0] m77_84;
   assign m77_84 =15'b0;

   // m77_85 = W*in
   wire signed [14:0] m77_85;
   assign m77_85 =15'b0;

   // m77_86 = W*in
   wire signed [14:0] m77_86;
   assign m77_86 ={ {3{neg77[14]}} , neg77[14:3] };

   // m77_87 = W*in
   wire signed [14:0] m77_87;
   assign m77_87 =15'b0;

   // m77_88 = W*in
   wire signed [14:0] m77_88;
   assign m77_88 =15'b0;

   // m77_89 = W*in
   wire signed [14:0] m77_89;
   assign m77_89 =15'b0;

   // m77_90 = W*in
   wire signed [14:0] m77_90;
   assign m77_90 =15'b0;

   // m77_91 = W*in
   wire signed [14:0] m77_91;
   assign m77_91 =15'b0;

   // m77_92 = W*in
   wire signed [14:0] m77_92;
   assign m77_92 =15'b0;

   // m77_93 = W*in
   wire signed [14:0] m77_93;
   assign m77_93 =15'b0;

   // m77_94 = W*in
   wire signed [14:0] m77_94;
   assign m77_94 =15'b0;

   // m77_95 = W*in
   wire signed [14:0] m77_95;
   assign m77_95 =15'b0;

   // m77_96 = W*in
   wire signed [14:0] m77_96;
   assign m77_96 =15'b0;

   // m77_97 = W*in
   wire signed [14:0] m77_97;
   assign m77_97 =15'b0;

   // m77_98 = W*in
   wire signed [14:0] m77_98;
   assign m77_98 =15'b0;

   // m77_99 = W*in
   wire signed [14:0] m77_99;
   assign m77_99 =15'b0;

   // m77_100 = W*in
   wire signed [14:0] m77_100;
   assign m77_100 =15'b0;

   // m78_1 = W*in
   wire signed [14:0] m78_1;
   assign m78_1 =15'b0;

   // m78_2 = W*in
   wire signed [14:0] m78_2;
   assign m78_2 =15'b0;

   // m78_3 = W*in
   wire signed [14:0] m78_3;
   assign m78_3 =15'b0;

   // m78_4 = W*in
   wire signed [14:0] m78_4;
   assign m78_4 =15'b0;

   // m78_5 = W*in
   wire signed [14:0] m78_5;
   assign m78_5 =15'b0;

   // m78_6 = W*in
   wire signed [14:0] m78_6;
   assign m78_6 =15'b0;

   // m78_7 = W*in
   wire signed [14:0] m78_7;
   assign m78_7 =15'b0;

   // m78_8 = W*in
   wire signed [14:0] m78_8;
   assign m78_8 =15'b0;

   // m78_9 = W*in
   wire signed [14:0] m78_9;
   assign m78_9 =15'b0;

   // m78_10 = W*in
   wire signed [14:0] m78_10;
   assign m78_10 =15'b0;

   // m78_11 = W*in
   wire signed [14:0] m78_11;
   assign m78_11 =15'b0;

   // m78_12 = W*in
   wire signed [14:0] m78_12;
   assign m78_12 =15'b0;

   // m78_13 = W*in
   wire signed [14:0] m78_13;
   assign m78_13 =15'b0;

   // m78_14 = W*in
   wire signed [14:0] m78_14;
   assign m78_14 =15'b0;

   // m78_15 = W*in
   wire signed [14:0] m78_15;
   assign m78_15 ={ {3{in78[14]}} , in78[14:3] };

   // m78_16 = W*in
   wire signed [14:0] m78_16;
   assign m78_16 =15'b0;

   // m78_17 = W*in
   wire signed [14:0] m78_17;
   assign m78_17 =15'b0;

   // m78_18 = W*in
   wire signed [14:0] m78_18;
   assign m78_18 =15'b0;

   // m78_19 = W*in
   wire signed [14:0] m78_19;
   assign m78_19 =15'b0;

   // m78_20 = W*in
   wire signed [14:0] m78_20;
   assign m78_20 ={ {3{neg78[14]}} , neg78[14:3] };

   // m78_21 = W*in
   wire signed [14:0] m78_21;
   assign m78_21 =15'b0;

   // m78_22 = W*in
   wire signed [14:0] m78_22;
   assign m78_22 =15'b0;

   // m78_23 = W*in
   wire signed [14:0] m78_23;
   assign m78_23 =15'b0;

   // m78_24 = W*in
   wire signed [14:0] m78_24;
   assign m78_24 =15'b0;

   // m78_25 = W*in
   wire signed [14:0] m78_25;
   assign m78_25 =15'b0;

   // m78_26 = W*in
   wire signed [14:0] m78_26;
   assign m78_26 =15'b0;

   // m78_27 = W*in
   wire signed [14:0] m78_27;
   assign m78_27 =15'b0;

   // m78_28 = W*in
   wire signed [14:0] m78_28;
   assign m78_28 =15'b0;

   // m78_29 = W*in
   wire signed [14:0] m78_29;
   assign m78_29 =15'b0;

   // m78_30 = W*in
   wire signed [14:0] m78_30;
   assign m78_30 =15'b0;

   // m78_31 = W*in
   wire signed [14:0] m78_31;
   assign m78_31 =15'b0;

   // m78_32 = W*in
   wire signed [14:0] m78_32;
   assign m78_32 =15'b0;

   // m78_33 = W*in
   wire signed [14:0] m78_33;
   assign m78_33 =15'b0;

   // m78_34 = W*in
   wire signed [14:0] m78_34;
   assign m78_34 =15'b0;

   // m78_35 = W*in
   wire signed [14:0] m78_35;
   assign m78_35 =15'b0;

   // m78_36 = W*in
   wire signed [14:0] m78_36;
   assign m78_36 =15'b0;

   // m78_37 = W*in
   wire signed [14:0] m78_37;
   assign m78_37 =15'b0;

   // m78_38 = W*in
   wire signed [14:0] m78_38;
   assign m78_38 =15'b0;

   // m78_39 = W*in
   wire signed [14:0] m78_39;
   assign m78_39 =15'b0;

   // m78_40 = W*in
   wire signed [14:0] m78_40;
   assign m78_40 =15'b0;

   // m78_41 = W*in
   wire signed [14:0] m78_41;
   assign m78_41 ={ {3{neg78[14]}} , neg78[14:3] };

   // m78_42 = W*in
   wire signed [14:0] m78_42;
   assign m78_42 =15'b0;

   // m78_43 = W*in
   wire signed [14:0] m78_43;
   assign m78_43 =15'b0;

   // m78_44 = W*in
   wire signed [14:0] m78_44;
   assign m78_44 =15'b0;

   // m78_45 = W*in
   wire signed [14:0] m78_45;
   assign m78_45 =15'b0;

   // m78_46 = W*in
   wire signed [14:0] m78_46;
   assign m78_46 =15'b0;

   // m78_47 = W*in
   wire signed [14:0] m78_47;
   assign m78_47 =15'b0;

   // m78_48 = W*in
   wire signed [14:0] m78_48;
   assign m78_48 ={ {3{in78[14]}} , in78[14:3] };

   // m78_49 = W*in
   wire signed [14:0] m78_49;
   assign m78_49 ={ {4{in78[14]}} , in78[14:4] };

   // m78_50 = W*in
   wire signed [14:0] m78_50;
   assign m78_50 ={ {4{in78[14]}} , in78[14:4] };

   // m78_51 = W*in
   wire signed [14:0] m78_51;
   assign m78_51 =15'b0;

   // m78_52 = W*in
   wire signed [14:0] m78_52;
   assign m78_52 =15'b0;

   // m78_53 = W*in
   wire signed [14:0] m78_53;
   assign m78_53 =15'b0;

   // m78_54 = W*in
   wire signed [14:0] m78_54;
   assign m78_54 =15'b0;

   // m78_55 = W*in
   wire signed [14:0] m78_55;
   assign m78_55 =15'b0;

   // m78_56 = W*in
   wire signed [14:0] m78_56;
   assign m78_56 =15'b0;

   // m78_57 = W*in
   wire signed [14:0] m78_57;
   assign m78_57 =15'b0;

   // m78_58 = W*in
   wire signed [14:0] m78_58;
   assign m78_58 =15'b0;

   // m78_59 = W*in
   wire signed [14:0] m78_59;
   assign m78_59 =15'b0;

   // m78_60 = W*in
   wire signed [14:0] m78_60;
   assign m78_60 =15'b0;

   // m78_61 = W*in
   wire signed [14:0] m78_61;
   assign m78_61 ={ {4{neg78[14]}} , neg78[14:4] };

   // m78_62 = W*in
   wire signed [14:0] m78_62;
   assign m78_62 =15'b0;

   // m78_63 = W*in
   wire signed [14:0] m78_63;
   assign m78_63 =15'b0;

   // m78_64 = W*in
   wire signed [14:0] m78_64;
   assign m78_64 =15'b0;

   // m78_65 = W*in
   wire signed [14:0] m78_65;
   assign m78_65 =15'b0;

   // m78_66 = W*in
   wire signed [14:0] m78_66;
   assign m78_66 =15'b0;

   // m78_67 = W*in
   wire signed [14:0] m78_67;
   assign m78_67 =15'b0;

   // m78_68 = W*in
   wire signed [14:0] m78_68;
   assign m78_68 =15'b0;

   // m78_69 = W*in
   wire signed [14:0] m78_69;
   assign m78_69 =15'b0;

   // m78_70 = W*in
   wire signed [14:0] m78_70;
   assign m78_70 =15'b0;

   // m78_71 = W*in
   wire signed [14:0] m78_71;
   assign m78_71 =15'b0;

   // m78_72 = W*in
   wire signed [14:0] m78_72;
   assign m78_72 =15'b0;

   // m78_73 = W*in
   wire signed [14:0] m78_73;
   assign m78_73 =15'b0;

   // m78_74 = W*in
   wire signed [14:0] m78_74;
   assign m78_74 ={ {3{neg78[14]}} , neg78[14:3] };

   // m78_75 = W*in
   wire signed [14:0] m78_75;
   assign m78_75 =15'b0;

   // m78_76 = W*in
   wire signed [14:0] m78_76;
   assign m78_76 ={ {3{neg78[14]}} , neg78[14:3] };

   // m78_77 = W*in
   wire signed [14:0] m78_77;
   assign m78_77 =15'b0;

   // m78_78 = W*in
   wire signed [14:0] m78_78;
   assign m78_78 =15'b0;

   // m78_79 = W*in
   wire signed [14:0] m78_79;
   assign m78_79 ={ {4{in78[14]}} , in78[14:4] };

   // m78_80 = W*in
   wire signed [14:0] m78_80;
   assign m78_80 =15'b0;

   // m78_81 = W*in
   wire signed [14:0] m78_81;
   assign m78_81 ={ {3{in78[14]}} , in78[14:3] };

   // m78_82 = W*in
   wire signed [14:0] m78_82;
   assign m78_82 =15'b0;

   // m78_83 = W*in
   wire signed [14:0] m78_83;
   assign m78_83 =15'b0;

   // m78_84 = W*in
   wire signed [14:0] m78_84;
   assign m78_84 =15'b0;

   // m78_85 = W*in
   wire signed [14:0] m78_85;
   assign m78_85 ={ {3{in78[14]}} , in78[14:3] };

   // m78_86 = W*in
   wire signed [14:0] m78_86;
   assign m78_86 =15'b0;

   // m78_87 = W*in
   wire signed [14:0] m78_87;
   assign m78_87 ={ {3{in78[14]}} , in78[14:3] };

   // m78_88 = W*in
   wire signed [14:0] m78_88;
   assign m78_88 =15'b0;

   // m78_89 = W*in
   wire signed [14:0] m78_89;
   assign m78_89 =15'b0;

   // m78_90 = W*in
   wire signed [14:0] m78_90;
   assign m78_90 =15'b0;

   // m78_91 = W*in
   wire signed [14:0] m78_91;
   assign m78_91 =15'b0;

   // m78_92 = W*in
   wire signed [14:0] m78_92;
   assign m78_92 =15'b0;

   // m78_93 = W*in
   wire signed [14:0] m78_93;
   assign m78_93 =15'b0;

   // m78_94 = W*in
   wire signed [14:0] m78_94;
   assign m78_94 =15'b0;

   // m78_95 = W*in
   wire signed [14:0] m78_95;
   assign m78_95 =15'b0;

   // m78_96 = W*in
   wire signed [14:0] m78_96;
   assign m78_96 =15'b0;

   // m78_97 = W*in
   wire signed [14:0] m78_97;
   assign m78_97 =15'b0;

   // m78_98 = W*in
   wire signed [14:0] m78_98;
   assign m78_98 =15'b0;

   // m78_99 = W*in
   wire signed [14:0] m78_99;
   assign m78_99 =15'b0;

   // m78_100 = W*in
   wire signed [14:0] m78_100;
   assign m78_100 =15'b0;

   // m79_1 = W*in
   wire signed [14:0] m79_1;
   assign m79_1 =15'b0;

   // m79_2 = W*in
   wire signed [14:0] m79_2;
   assign m79_2 =15'b0;

   // m79_3 = W*in
   wire signed [14:0] m79_3;
   assign m79_3 =15'b0;

   // m79_4 = W*in
   wire signed [14:0] m79_4;
   assign m79_4 =15'b0;

   // m79_5 = W*in
   wire signed [14:0] m79_5;
   assign m79_5 =15'b0;

   // m79_6 = W*in
   wire signed [14:0] m79_6;
   assign m79_6 =15'b0;

   // m79_7 = W*in
   wire signed [14:0] m79_7;
   assign m79_7 =15'b0;

   // m79_8 = W*in
   wire signed [14:0] m79_8;
   assign m79_8 =15'b0;

   // m79_9 = W*in
   wire signed [14:0] m79_9;
   assign m79_9 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_10 = W*in
   wire signed [14:0] m79_10;
   assign m79_10 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_11 = W*in
   wire signed [14:0] m79_11;
   assign m79_11 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_12 = W*in
   wire signed [14:0] m79_12;
   assign m79_12 ={ {4{neg79[14]}} , neg79[14:4] };

   // m79_13 = W*in
   wire signed [14:0] m79_13;
   assign m79_13 =15'b0;

   // m79_14 = W*in
   wire signed [14:0] m79_14;
   assign m79_14 =15'b0;

   // m79_15 = W*in
   wire signed [14:0] m79_15;
   assign m79_15 =15'b0;

   // m79_16 = W*in
   wire signed [14:0] m79_16;
   assign m79_16 =15'b0;

   // m79_17 = W*in
   wire signed [14:0] m79_17;
   assign m79_17 =15'b0;

   // m79_18 = W*in
   wire signed [14:0] m79_18;
   assign m79_18 =15'b0;

   // m79_19 = W*in
   wire signed [14:0] m79_19;
   assign m79_19 =15'b0;

   // m79_20 = W*in
   wire signed [14:0] m79_20;
   assign m79_20 =15'b0;

   // m79_21 = W*in
   wire signed [14:0] m79_21;
   assign m79_21 =15'b0;

   // m79_22 = W*in
   wire signed [14:0] m79_22;
   assign m79_22 =15'b0;

   // m79_23 = W*in
   wire signed [14:0] m79_23;
   assign m79_23 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_24 = W*in
   wire signed [14:0] m79_24;
   assign m79_24 =15'b0;

   // m79_25 = W*in
   wire signed [14:0] m79_25;
   assign m79_25 =15'b0;

   // m79_26 = W*in
   wire signed [14:0] m79_26;
   assign m79_26 =15'b0;

   // m79_27 = W*in
   wire signed [14:0] m79_27;
   assign m79_27 =15'b0;

   // m79_28 = W*in
   wire signed [14:0] m79_28;
   assign m79_28 =15'b0;

   // m79_29 = W*in
   wire signed [14:0] m79_29;
   assign m79_29 =15'b0;

   // m79_30 = W*in
   wire signed [14:0] m79_30;
   assign m79_30 ={ {3{in79[14]}} , in79[14:3] };

   // m79_31 = W*in
   wire signed [14:0] m79_31;
   assign m79_31 =15'b0;

   // m79_32 = W*in
   wire signed [14:0] m79_32;
   assign m79_32 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_33 = W*in
   wire signed [14:0] m79_33;
   assign m79_33 =15'b0;

   // m79_34 = W*in
   wire signed [14:0] m79_34;
   assign m79_34 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_35 = W*in
   wire signed [14:0] m79_35;
   assign m79_35 =15'b0;

   // m79_36 = W*in
   wire signed [14:0] m79_36;
   assign m79_36 =15'b0;

   // m79_37 = W*in
   wire signed [14:0] m79_37;
   assign m79_37 =15'b0;

   // m79_38 = W*in
   wire signed [14:0] m79_38;
   assign m79_38 ={ {4{neg79[14]}} , neg79[14:4] };

   // m79_39 = W*in
   wire signed [14:0] m79_39;
   assign m79_39 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_40 = W*in
   wire signed [14:0] m79_40;
   assign m79_40 =15'b0;

   // m79_41 = W*in
   wire signed [14:0] m79_41;
   assign m79_41 =15'b0;

   // m79_42 = W*in
   wire signed [14:0] m79_42;
   assign m79_42 =15'b0;

   // m79_43 = W*in
   wire signed [14:0] m79_43;
   assign m79_43 =15'b0;

   // m79_44 = W*in
   wire signed [14:0] m79_44;
   assign m79_44 =15'b0;

   // m79_45 = W*in
   wire signed [14:0] m79_45;
   assign m79_45 ={ {4{neg79[14]}} , neg79[14:4] };

   // m79_46 = W*in
   wire signed [14:0] m79_46;
   assign m79_46 =15'b0;

   // m79_47 = W*in
   wire signed [14:0] m79_47;
   assign m79_47 ={ {3{in79[14]}} , in79[14:3] };

   // m79_48 = W*in
   wire signed [14:0] m79_48;
   assign m79_48 =15'b0;

   // m79_49 = W*in
   wire signed [14:0] m79_49;
   assign m79_49 =15'b0;

   // m79_50 = W*in
   wire signed [14:0] m79_50;
   assign m79_50 =15'b0;

   // m79_51 = W*in
   wire signed [14:0] m79_51;
   assign m79_51 =15'b0;

   // m79_52 = W*in
   wire signed [14:0] m79_52;
   assign m79_52 =15'b0;

   // m79_53 = W*in
   wire signed [14:0] m79_53;
   assign m79_53 =15'b0;

   // m79_54 = W*in
   wire signed [14:0] m79_54;
   assign m79_54 =15'b0;

   // m79_55 = W*in
   wire signed [14:0] m79_55;
   assign m79_55 =15'b0;

   // m79_56 = W*in
   wire signed [14:0] m79_56;
   assign m79_56 =15'b0;

   // m79_57 = W*in
   wire signed [14:0] m79_57;
   assign m79_57 =15'b0;

   // m79_58 = W*in
   wire signed [14:0] m79_58;
   assign m79_58 =15'b0;

   // m79_59 = W*in
   wire signed [14:0] m79_59;
   assign m79_59 =15'b0;

   // m79_60 = W*in
   wire signed [14:0] m79_60;
   assign m79_60 =15'b0;

   // m79_61 = W*in
   wire signed [14:0] m79_61;
   assign m79_61 =15'b0;

   // m79_62 = W*in
   wire signed [14:0] m79_62;
   assign m79_62 =15'b0;

   // m79_63 = W*in
   wire signed [14:0] m79_63;
   assign m79_63 ={ {4{neg79[14]}} , neg79[14:4] };

   // m79_64 = W*in
   wire signed [14:0] m79_64;
   assign m79_64 =15'b0;

   // m79_65 = W*in
   wire signed [14:0] m79_65;
   assign m79_65 =15'b0;

   // m79_66 = W*in
   wire signed [14:0] m79_66;
   assign m79_66 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_67 = W*in
   wire signed [14:0] m79_67;
   assign m79_67 =15'b0;

   // m79_68 = W*in
   wire signed [14:0] m79_68;
   assign m79_68 =15'b0;

   // m79_69 = W*in
   wire signed [14:0] m79_69;
   assign m79_69 =15'b0;

   // m79_70 = W*in
   wire signed [14:0] m79_70;
   assign m79_70 =15'b0;

   // m79_71 = W*in
   wire signed [14:0] m79_71;
   assign m79_71 =15'b0;

   // m79_72 = W*in
   wire signed [14:0] m79_72;
   assign m79_72 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_73 = W*in
   wire signed [14:0] m79_73;
   assign m79_73 ={ {3{in79[14]}} , in79[14:3] };

   // m79_74 = W*in
   wire signed [14:0] m79_74;
   assign m79_74 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_75 = W*in
   wire signed [14:0] m79_75;
   assign m79_75 =15'b0;

   // m79_76 = W*in
   wire signed [14:0] m79_76;
   assign m79_76 =15'b0;

   // m79_77 = W*in
   wire signed [14:0] m79_77;
   assign m79_77 =15'b0;

   // m79_78 = W*in
   wire signed [14:0] m79_78;
   assign m79_78 =15'b0;

   // m79_79 = W*in
   wire signed [14:0] m79_79;
   assign m79_79 =15'b0;

   // m79_80 = W*in
   wire signed [14:0] m79_80;
   assign m79_80 ={ {4{neg79[14]}} , neg79[14:4] };

   // m79_81 = W*in
   wire signed [14:0] m79_81;
   assign m79_81 =15'b0;

   // m79_82 = W*in
   wire signed [14:0] m79_82;
   assign m79_82 =15'b0;

   // m79_83 = W*in
   wire signed [14:0] m79_83;
   assign m79_83 =15'b0;

   // m79_84 = W*in
   wire signed [14:0] m79_84;
   assign m79_84 =15'b0;

   // m79_85 = W*in
   wire signed [14:0] m79_85;
   assign m79_85 =15'b0;

   // m79_86 = W*in
   wire signed [14:0] m79_86;
   assign m79_86 =15'b0;

   // m79_87 = W*in
   wire signed [14:0] m79_87;
   assign m79_87 =15'b0;

   // m79_88 = W*in
   wire signed [14:0] m79_88;
   assign m79_88 =15'b0;

   // m79_89 = W*in
   wire signed [14:0] m79_89;
   assign m79_89 =15'b0;

   // m79_90 = W*in
   wire signed [14:0] m79_90;
   assign m79_90 ={ {3{neg79[14]}} , neg79[14:3] };

   // m79_91 = W*in
   wire signed [14:0] m79_91;
   assign m79_91 =15'b0;

   // m79_92 = W*in
   wire signed [14:0] m79_92;
   assign m79_92 =15'b0;

   // m79_93 = W*in
   wire signed [14:0] m79_93;
   assign m79_93 =15'b0;

   // m79_94 = W*in
   wire signed [14:0] m79_94;
   assign m79_94 =15'b0;

   // m79_95 = W*in
   wire signed [14:0] m79_95;
   assign m79_95 =15'b0;

   // m79_96 = W*in
   wire signed [14:0] m79_96;
   assign m79_96 =15'b0;

   // m79_97 = W*in
   wire signed [14:0] m79_97;
   assign m79_97 =15'b0;

   // m79_98 = W*in
   wire signed [14:0] m79_98;
   assign m79_98 ={ {3{in79[14]}} , in79[14:3] };

   // m79_99 = W*in
   wire signed [14:0] m79_99;
   assign m79_99 =15'b0;

   // m79_100 = W*in
   wire signed [14:0] m79_100;
   assign m79_100 =15'b0;

   // m80_1 = W*in
   wire signed [14:0] m80_1;
   assign m80_1 =15'b0;

   // m80_2 = W*in
   wire signed [14:0] m80_2;
   assign m80_2 =15'b0;

   // m80_3 = W*in
   wire signed [14:0] m80_3;
   assign m80_3 =15'b0;

   // m80_4 = W*in
   wire signed [14:0] m80_4;
   assign m80_4 =15'b0;

   // m80_5 = W*in
   wire signed [14:0] m80_5;
   assign m80_5 =15'b0;

   // m80_6 = W*in
   wire signed [14:0] m80_6;
   assign m80_6 =15'b0;

   // m80_7 = W*in
   wire signed [14:0] m80_7;
   assign m80_7 =15'b0;

   // m80_8 = W*in
   wire signed [14:0] m80_8;
   assign m80_8 =15'b0;

   // m80_9 = W*in
   wire signed [14:0] m80_9;
   assign m80_9 =15'b0;

   // m80_10 = W*in
   wire signed [14:0] m80_10;
   assign m80_10 =15'b0;

   // m80_11 = W*in
   wire signed [14:0] m80_11;
   assign m80_11 =15'b0;

   // m80_12 = W*in
   wire signed [14:0] m80_12;
   assign m80_12 =15'b0;

   // m80_13 = W*in
   wire signed [14:0] m80_13;
   assign m80_13 =15'b0;

   // m80_14 = W*in
   wire signed [14:0] m80_14;
   assign m80_14 =15'b0;

   // m80_15 = W*in
   wire signed [14:0] m80_15;
   assign m80_15 =15'b0;

   // m80_16 = W*in
   wire signed [14:0] m80_16;
   assign m80_16 =15'b0;

   // m80_17 = W*in
   wire signed [14:0] m80_17;
   assign m80_17 =15'b0;

   // m80_18 = W*in
   wire signed [14:0] m80_18;
   assign m80_18 =15'b0;

   // m80_19 = W*in
   wire signed [14:0] m80_19;
   assign m80_19 =15'b0;

   // m80_20 = W*in
   wire signed [14:0] m80_20;
   assign m80_20 =15'b0;

   // m80_21 = W*in
   wire signed [14:0] m80_21;
   assign m80_21 =15'b0;

   // m80_22 = W*in
   wire signed [14:0] m80_22;
   assign m80_22 =15'b0;

   // m80_23 = W*in
   wire signed [14:0] m80_23;
   assign m80_23 =15'b0;

   // m80_24 = W*in
   wire signed [14:0] m80_24;
   assign m80_24 =15'b0;

   // m80_25 = W*in
   wire signed [14:0] m80_25;
   assign m80_25 =15'b0;

   // m80_26 = W*in
   wire signed [14:0] m80_26;
   assign m80_26 ={ {4{neg80[14]}} , neg80[14:4] };

   // m80_27 = W*in
   wire signed [14:0] m80_27;
   assign m80_27 =15'b0;

   // m80_28 = W*in
   wire signed [14:0] m80_28;
   assign m80_28 =15'b0;

   // m80_29 = W*in
   wire signed [14:0] m80_29;
   assign m80_29 =15'b0;

   // m80_30 = W*in
   wire signed [14:0] m80_30;
   assign m80_30 =15'b0;

   // m80_31 = W*in
   wire signed [14:0] m80_31;
   assign m80_31 =15'b0;

   // m80_32 = W*in
   wire signed [14:0] m80_32;
   assign m80_32 =15'b0;

   // m80_33 = W*in
   wire signed [14:0] m80_33;
   assign m80_33 =15'b0;

   // m80_34 = W*in
   wire signed [14:0] m80_34;
   assign m80_34 =15'b0;

   // m80_35 = W*in
   wire signed [14:0] m80_35;
   assign m80_35 =15'b0;

   // m80_36 = W*in
   wire signed [14:0] m80_36;
   assign m80_36 =15'b0;

   // m80_37 = W*in
   wire signed [14:0] m80_37;
   assign m80_37 =15'b0;

   // m80_38 = W*in
   wire signed [14:0] m80_38;
   assign m80_38 =15'b0;

   // m80_39 = W*in
   wire signed [14:0] m80_39;
   assign m80_39 =15'b0;

   // m80_40 = W*in
   wire signed [14:0] m80_40;
   assign m80_40 =15'b0;

   // m80_41 = W*in
   wire signed [14:0] m80_41;
   assign m80_41 =15'b0;

   // m80_42 = W*in
   wire signed [14:0] m80_42;
   assign m80_42 =15'b0;

   // m80_43 = W*in
   wire signed [14:0] m80_43;
   assign m80_43 =15'b0;

   // m80_44 = W*in
   wire signed [14:0] m80_44;
   assign m80_44 =15'b0;

   // m80_45 = W*in
   wire signed [14:0] m80_45;
   assign m80_45 =15'b0;

   // m80_46 = W*in
   wire signed [14:0] m80_46;
   assign m80_46 =15'b0;

   // m80_47 = W*in
   wire signed [14:0] m80_47;
   assign m80_47 ={ {4{in80[14]}} , in80[14:4] };

   // m80_48 = W*in
   wire signed [14:0] m80_48;
   assign m80_48 =15'b0;

   // m80_49 = W*in
   wire signed [14:0] m80_49;
   assign m80_49 =15'b0;

   // m80_50 = W*in
   wire signed [14:0] m80_50;
   assign m80_50 =15'b0;

   // m80_51 = W*in
   wire signed [14:0] m80_51;
   assign m80_51 =15'b0;

   // m80_52 = W*in
   wire signed [14:0] m80_52;
   assign m80_52 =15'b0;

   // m80_53 = W*in
   wire signed [14:0] m80_53;
   assign m80_53 =15'b0;

   // m80_54 = W*in
   wire signed [14:0] m80_54;
   assign m80_54 =15'b0;

   // m80_55 = W*in
   wire signed [14:0] m80_55;
   assign m80_55 =15'b0;

   // m80_56 = W*in
   wire signed [14:0] m80_56;
   assign m80_56 =15'b0;

   // m80_57 = W*in
   wire signed [14:0] m80_57;
   assign m80_57 =15'b0;

   // m80_58 = W*in
   wire signed [14:0] m80_58;
   assign m80_58 =15'b0;

   // m80_59 = W*in
   wire signed [14:0] m80_59;
   assign m80_59 =15'b0;

   // m80_60 = W*in
   wire signed [14:0] m80_60;
   assign m80_60 =15'b0;

   // m80_61 = W*in
   wire signed [14:0] m80_61;
   assign m80_61 =15'b0;

   // m80_62 = W*in
   wire signed [14:0] m80_62;
   assign m80_62 =15'b0;

   // m80_63 = W*in
   wire signed [14:0] m80_63;
   assign m80_63 =15'b0;

   // m80_64 = W*in
   wire signed [14:0] m80_64;
   assign m80_64 =15'b0;

   // m80_65 = W*in
   wire signed [14:0] m80_65;
   assign m80_65 =15'b0;

   // m80_66 = W*in
   wire signed [14:0] m80_66;
   assign m80_66 =15'b0;

   // m80_67 = W*in
   wire signed [14:0] m80_67;
   assign m80_67 =15'b0;

   // m80_68 = W*in
   wire signed [14:0] m80_68;
   assign m80_68 =15'b0;

   // m80_69 = W*in
   wire signed [14:0] m80_69;
   assign m80_69 =15'b0;

   // m80_70 = W*in
   wire signed [14:0] m80_70;
   assign m80_70 =15'b0;

   // m80_71 = W*in
   wire signed [14:0] m80_71;
   assign m80_71 =15'b0;

   // m80_72 = W*in
   wire signed [14:0] m80_72;
   assign m80_72 =15'b0;

   // m80_73 = W*in
   wire signed [14:0] m80_73;
   assign m80_73 =15'b0;

   // m80_74 = W*in
   wire signed [14:0] m80_74;
   assign m80_74 =15'b0;

   // m80_75 = W*in
   wire signed [14:0] m80_75;
   assign m80_75 =15'b0;

   // m80_76 = W*in
   wire signed [14:0] m80_76;
   assign m80_76 =15'b0;

   // m80_77 = W*in
   wire signed [14:0] m80_77;
   assign m80_77 =15'b0;

   // m80_78 = W*in
   wire signed [14:0] m80_78;
   assign m80_78 =15'b0;

   // m80_79 = W*in
   wire signed [14:0] m80_79;
   assign m80_79 =15'b0;

   // m80_80 = W*in
   wire signed [14:0] m80_80;
   assign m80_80 =15'b0;

   // m80_81 = W*in
   wire signed [14:0] m80_81;
   assign m80_81 =15'b0;

   // m80_82 = W*in
   wire signed [14:0] m80_82;
   assign m80_82 =15'b0;

   // m80_83 = W*in
   wire signed [14:0] m80_83;
   assign m80_83 =15'b0;

   // m80_84 = W*in
   wire signed [14:0] m80_84;
   assign m80_84 =15'b0;

   // m80_85 = W*in
   wire signed [14:0] m80_85;
   assign m80_85 =15'b0;

   // m80_86 = W*in
   wire signed [14:0] m80_86;
   assign m80_86 =15'b0;

   // m80_87 = W*in
   wire signed [14:0] m80_87;
   assign m80_87 =15'b0;

   // m80_88 = W*in
   wire signed [14:0] m80_88;
   assign m80_88 =15'b0;

   // m80_89 = W*in
   wire signed [14:0] m80_89;
   assign m80_89 =15'b0;

   // m80_90 = W*in
   wire signed [14:0] m80_90;
   assign m80_90 =15'b0;

   // m80_91 = W*in
   wire signed [14:0] m80_91;
   assign m80_91 =15'b0;

   // m80_92 = W*in
   wire signed [14:0] m80_92;
   assign m80_92 =15'b0;

   // m80_93 = W*in
   wire signed [14:0] m80_93;
   assign m80_93 =15'b0;

   // m80_94 = W*in
   wire signed [14:0] m80_94;
   assign m80_94 =15'b0;

   // m80_95 = W*in
   wire signed [14:0] m80_95;
   assign m80_95 =15'b0;

   // m80_96 = W*in
   wire signed [14:0] m80_96;
   assign m80_96 =15'b0;

   // m80_97 = W*in
   wire signed [14:0] m80_97;
   assign m80_97 =15'b0;

   // m80_98 = W*in
   wire signed [14:0] m80_98;
   assign m80_98 =15'b0;

   // m80_99 = W*in
   wire signed [14:0] m80_99;
   assign m80_99 =15'b0;

   // m80_100 = W*in
   wire signed [14:0] m80_100;
   assign m80_100 =15'b0;

   // m81_1 = W*in
   wire signed [14:0] m81_1;
   assign m81_1 =15'b0;

   // m81_2 = W*in
   wire signed [14:0] m81_2;
   assign m81_2 =15'b0;

   // m81_3 = W*in
   wire signed [14:0] m81_3;
   assign m81_3 =15'b0;

   // m81_4 = W*in
   wire signed [14:0] m81_4;
   assign m81_4 =15'b0;

   // m81_5 = W*in
   wire signed [14:0] m81_5;
   assign m81_5 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_6 = W*in
   wire signed [14:0] m81_6;
   assign m81_6 =15'b0;

   // m81_7 = W*in
   wire signed [14:0] m81_7;
   assign m81_7 ={ {3{in81[14]}} , in81[14:3] };

   // m81_8 = W*in
   wire signed [14:0] m81_8;
   assign m81_8 =15'b0;

   // m81_9 = W*in
   wire signed [14:0] m81_9;
   assign m81_9 ={ {3{in81[14]}} , in81[14:3] };

   // m81_10 = W*in
   wire signed [14:0] m81_10;
   assign m81_10 =15'b0;

   // m81_11 = W*in
   wire signed [14:0] m81_11;
   assign m81_11 =15'b0;

   // m81_12 = W*in
   wire signed [14:0] m81_12;
   assign m81_12 =15'b0;

   // m81_13 = W*in
   wire signed [14:0] m81_13;
   assign m81_13 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_14 = W*in
   wire signed [14:0] m81_14;
   assign m81_14 =15'b0;

   // m81_15 = W*in
   wire signed [14:0] m81_15;
   assign m81_15 =15'b0;

   // m81_16 = W*in
   wire signed [14:0] m81_16;
   assign m81_16 =15'b0;

   // m81_17 = W*in
   wire signed [14:0] m81_17;
   assign m81_17 =15'b0;

   // m81_18 = W*in
   wire signed [14:0] m81_18;
   assign m81_18 =15'b0;

   // m81_19 = W*in
   wire signed [14:0] m81_19;
   assign m81_19 =15'b0;

   // m81_20 = W*in
   wire signed [14:0] m81_20;
   assign m81_20 =15'b0;

   // m81_21 = W*in
   wire signed [14:0] m81_21;
   assign m81_21 =15'b0;

   // m81_22 = W*in
   wire signed [14:0] m81_22;
   assign m81_22 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_23 = W*in
   wire signed [14:0] m81_23;
   assign m81_23 =15'b0;

   // m81_24 = W*in
   wire signed [14:0] m81_24;
   assign m81_24 =15'b0;

   // m81_25 = W*in
   wire signed [14:0] m81_25;
   assign m81_25 =15'b0;

   // m81_26 = W*in
   wire signed [14:0] m81_26;
   assign m81_26 ={ {3{in81[14]}} , in81[14:3] };

   // m81_27 = W*in
   wire signed [14:0] m81_27;
   assign m81_27 =15'b0;

   // m81_28 = W*in
   wire signed [14:0] m81_28;
   assign m81_28 =15'b0;

   // m81_29 = W*in
   wire signed [14:0] m81_29;
   assign m81_29 =15'b0;

   // m81_30 = W*in
   wire signed [14:0] m81_30;
   assign m81_30 =15'b0;

   // m81_31 = W*in
   wire signed [14:0] m81_31;
   assign m81_31 =15'b0;

   // m81_32 = W*in
   wire signed [14:0] m81_32;
   assign m81_32 =15'b0;

   // m81_33 = W*in
   wire signed [14:0] m81_33;
   assign m81_33 =15'b0;

   // m81_34 = W*in
   wire signed [14:0] m81_34;
   assign m81_34 =15'b0;

   // m81_35 = W*in
   wire signed [14:0] m81_35;
   assign m81_35 =15'b0;

   // m81_36 = W*in
   wire signed [14:0] m81_36;
   assign m81_36 =15'b0;

   // m81_37 = W*in
   wire signed [14:0] m81_37;
   assign m81_37 =15'b0;

   // m81_38 = W*in
   wire signed [14:0] m81_38;
   assign m81_38 =15'b0;

   // m81_39 = W*in
   wire signed [14:0] m81_39;
   assign m81_39 =15'b0;

   // m81_40 = W*in
   wire signed [14:0] m81_40;
   assign m81_40 =15'b0;

   // m81_41 = W*in
   wire signed [14:0] m81_41;
   assign m81_41 =15'b0;

   // m81_42 = W*in
   wire signed [14:0] m81_42;
   assign m81_42 ={ {3{in81[14]}} , in81[14:3] };

   // m81_43 = W*in
   wire signed [14:0] m81_43;
   assign m81_43 =15'b0;

   // m81_44 = W*in
   wire signed [14:0] m81_44;
   assign m81_44 =15'b0;

   // m81_45 = W*in
   wire signed [14:0] m81_45;
   assign m81_45 =15'b0;

   // m81_46 = W*in
   wire signed [14:0] m81_46;
   assign m81_46 =15'b0;

   // m81_47 = W*in
   wire signed [14:0] m81_47;
   assign m81_47 =15'b0;

   // m81_48 = W*in
   wire signed [14:0] m81_48;
   assign m81_48 =15'b0;

   // m81_49 = W*in
   wire signed [14:0] m81_49;
   assign m81_49 ={ {3{in81[14]}} , in81[14:3] };

   // m81_50 = W*in
   wire signed [14:0] m81_50;
   assign m81_50 =15'b0;

   // m81_51 = W*in
   wire signed [14:0] m81_51;
   assign m81_51 =15'b0;

   // m81_52 = W*in
   wire signed [14:0] m81_52;
   assign m81_52 =15'b0;

   // m81_53 = W*in
   wire signed [14:0] m81_53;
   assign m81_53 =15'b0;

   // m81_54 = W*in
   wire signed [14:0] m81_54;
   assign m81_54 ={ {3{in81[14]}} , in81[14:3] };

   // m81_55 = W*in
   wire signed [14:0] m81_55;
   assign m81_55 =15'b0;

   // m81_56 = W*in
   wire signed [14:0] m81_56;
   assign m81_56 =15'b0;

   // m81_57 = W*in
   wire signed [14:0] m81_57;
   assign m81_57 =15'b0;

   // m81_58 = W*in
   wire signed [14:0] m81_58;
   assign m81_58 =15'b0;

   // m81_59 = W*in
   wire signed [14:0] m81_59;
   assign m81_59 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_60 = W*in
   wire signed [14:0] m81_60;
   assign m81_60 =15'b0;

   // m81_61 = W*in
   wire signed [14:0] m81_61;
   assign m81_61 ={ {4{neg81[14]}} , neg81[14:4] };

   // m81_62 = W*in
   wire signed [14:0] m81_62;
   assign m81_62 =15'b0;

   // m81_63 = W*in
   wire signed [14:0] m81_63;
   assign m81_63 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_64 = W*in
   wire signed [14:0] m81_64;
   assign m81_64 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_65 = W*in
   wire signed [14:0] m81_65;
   assign m81_65 =15'b0;

   // m81_66 = W*in
   wire signed [14:0] m81_66;
   assign m81_66 ={ {3{in81[14]}} , in81[14:3] };

   // m81_67 = W*in
   wire signed [14:0] m81_67;
   assign m81_67 ={ {4{in81[14]}} , in81[14:4] };

   // m81_68 = W*in
   wire signed [14:0] m81_68;
   assign m81_68 =15'b0;

   // m81_69 = W*in
   wire signed [14:0] m81_69;
   assign m81_69 =15'b0;

   // m81_70 = W*in
   wire signed [14:0] m81_70;
   assign m81_70 =15'b0;

   // m81_71 = W*in
   wire signed [14:0] m81_71;
   assign m81_71 =15'b0;

   // m81_72 = W*in
   wire signed [14:0] m81_72;
   assign m81_72 ={ {3{in81[14]}} , in81[14:3] };

   // m81_73 = W*in
   wire signed [14:0] m81_73;
   assign m81_73 =15'b0;

   // m81_74 = W*in
   wire signed [14:0] m81_74;
   assign m81_74 ={ {4{neg81[14]}} , neg81[14:4] };

   // m81_75 = W*in
   wire signed [14:0] m81_75;
   assign m81_75 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_76 = W*in
   wire signed [14:0] m81_76;
   assign m81_76 =15'b0;

   // m81_77 = W*in
   wire signed [14:0] m81_77;
   assign m81_77 =15'b0;

   // m81_78 = W*in
   wire signed [14:0] m81_78;
   assign m81_78 =15'b0;

   // m81_79 = W*in
   wire signed [14:0] m81_79;
   assign m81_79 =15'b0;

   // m81_80 = W*in
   wire signed [14:0] m81_80;
   assign m81_80 ={ {4{neg81[14]}} , neg81[14:4] };

   // m81_81 = W*in
   wire signed [14:0] m81_81;
   assign m81_81 =15'b0;

   // m81_82 = W*in
   wire signed [14:0] m81_82;
   assign m81_82 =15'b0;

   // m81_83 = W*in
   wire signed [14:0] m81_83;
   assign m81_83 =15'b0;

   // m81_84 = W*in
   wire signed [14:0] m81_84;
   assign m81_84 =15'b0;

   // m81_85 = W*in
   wire signed [14:0] m81_85;
   assign m81_85 =15'b0;

   // m81_86 = W*in
   wire signed [14:0] m81_86;
   assign m81_86 =15'b0;

   // m81_87 = W*in
   wire signed [14:0] m81_87;
   assign m81_87 =15'b0;

   // m81_88 = W*in
   wire signed [14:0] m81_88;
   assign m81_88 =15'b0;

   // m81_89 = W*in
   wire signed [14:0] m81_89;
   assign m81_89 =15'b0;

   // m81_90 = W*in
   wire signed [14:0] m81_90;
   assign m81_90 ={ {4{neg81[14]}} , neg81[14:4] };

   // m81_91 = W*in
   wire signed [14:0] m81_91;
   assign m81_91 =15'b0;

   // m81_92 = W*in
   wire signed [14:0] m81_92;
   assign m81_92 =15'b0;

   // m81_93 = W*in
   wire signed [14:0] m81_93;
   assign m81_93 =15'b0;

   // m81_94 = W*in
   wire signed [14:0] m81_94;
   assign m81_94 ={ {3{in81[14]}} , in81[14:3] };

   // m81_95 = W*in
   wire signed [14:0] m81_95;
   assign m81_95 =15'b0;

   // m81_96 = W*in
   wire signed [14:0] m81_96;
   assign m81_96 =15'b0;

   // m81_97 = W*in
   wire signed [14:0] m81_97;
   assign m81_97 =15'b0;

   // m81_98 = W*in
   wire signed [14:0] m81_98;
   assign m81_98 ={ {4{in81[14]}} , in81[14:4] };

   // m81_99 = W*in
   wire signed [14:0] m81_99;
   assign m81_99 ={ {3{neg81[14]}} , neg81[14:3] };

   // m81_100 = W*in
   wire signed [14:0] m81_100;
   assign m81_100 =15'b0;

   // m82_1 = W*in
   wire signed [14:0] m82_1;
   assign m82_1 =15'b0;

   // m82_2 = W*in
   wire signed [14:0] m82_2;
   assign m82_2 =15'b0;

   // m82_3 = W*in
   wire signed [14:0] m82_3;
   assign m82_3 =15'b0;

   // m82_4 = W*in
   wire signed [14:0] m82_4;
   assign m82_4 =15'b0;

   // m82_5 = W*in
   wire signed [14:0] m82_5;
   assign m82_5 =15'b0;

   // m82_6 = W*in
   wire signed [14:0] m82_6;
   assign m82_6 =15'b0;

   // m82_7 = W*in
   wire signed [14:0] m82_7;
   assign m82_7 =15'b0;

   // m82_8 = W*in
   wire signed [14:0] m82_8;
   assign m82_8 =15'b0;

   // m82_9 = W*in
   wire signed [14:0] m82_9;
   assign m82_9 =15'b0;

   // m82_10 = W*in
   wire signed [14:0] m82_10;
   assign m82_10 ={ {3{in82[14]}} , in82[14:3] };

   // m82_11 = W*in
   wire signed [14:0] m82_11;
   assign m82_11 =15'b0;

   // m82_12 = W*in
   wire signed [14:0] m82_12;
   assign m82_12 =15'b0;

   // m82_13 = W*in
   wire signed [14:0] m82_13;
   assign m82_13 =15'b0;

   // m82_14 = W*in
   wire signed [14:0] m82_14;
   assign m82_14 =15'b0;

   // m82_15 = W*in
   wire signed [14:0] m82_15;
   assign m82_15 =15'b0;

   // m82_16 = W*in
   wire signed [14:0] m82_16;
   assign m82_16 =15'b0;

   // m82_17 = W*in
   wire signed [14:0] m82_17;
   assign m82_17 =15'b0;

   // m82_18 = W*in
   wire signed [14:0] m82_18;
   assign m82_18 ={ {3{neg82[14]}} , neg82[14:3] };

   // m82_19 = W*in
   wire signed [14:0] m82_19;
   assign m82_19 =15'b0;

   // m82_20 = W*in
   wire signed [14:0] m82_20;
   assign m82_20 ={ {4{neg82[14]}} , neg82[14:4] };

   // m82_21 = W*in
   wire signed [14:0] m82_21;
   assign m82_21 =15'b0;

   // m82_22 = W*in
   wire signed [14:0] m82_22;
   assign m82_22 =15'b0;

   // m82_23 = W*in
   wire signed [14:0] m82_23;
   assign m82_23 =15'b0;

   // m82_24 = W*in
   wire signed [14:0] m82_24;
   assign m82_24 ={ {4{neg82[14]}} , neg82[14:4] };

   // m82_25 = W*in
   wire signed [14:0] m82_25;
   assign m82_25 =15'b0;

   // m82_26 = W*in
   wire signed [14:0] m82_26;
   assign m82_26 =15'b0;

   // m82_27 = W*in
   wire signed [14:0] m82_27;
   assign m82_27 =15'b0;

   // m82_28 = W*in
   wire signed [14:0] m82_28;
   assign m82_28 =15'b0;

   // m82_29 = W*in
   wire signed [14:0] m82_29;
   assign m82_29 =15'b0;

   // m82_30 = W*in
   wire signed [14:0] m82_30;
   assign m82_30 =15'b0;

   // m82_31 = W*in
   wire signed [14:0] m82_31;
   assign m82_31 =15'b0;

   // m82_32 = W*in
   wire signed [14:0] m82_32;
   assign m82_32 =15'b0;

   // m82_33 = W*in
   wire signed [14:0] m82_33;
   assign m82_33 ={ {3{in82[14]}} , in82[14:3] };

   // m82_34 = W*in
   wire signed [14:0] m82_34;
   assign m82_34 =15'b0;

   // m82_35 = W*in
   wire signed [14:0] m82_35;
   assign m82_35 =15'b0;

   // m82_36 = W*in
   wire signed [14:0] m82_36;
   assign m82_36 =15'b0;

   // m82_37 = W*in
   wire signed [14:0] m82_37;
   assign m82_37 =15'b0;

   // m82_38 = W*in
   wire signed [14:0] m82_38;
   assign m82_38 =15'b0;

   // m82_39 = W*in
   wire signed [14:0] m82_39;
   assign m82_39 =15'b0;

   // m82_40 = W*in
   wire signed [14:0] m82_40;
   assign m82_40 =15'b0;

   // m82_41 = W*in
   wire signed [14:0] m82_41;
   assign m82_41 ={ {3{neg82[14]}} , neg82[14:3] };

   // m82_42 = W*in
   wire signed [14:0] m82_42;
   assign m82_42 =15'b0;

   // m82_43 = W*in
   wire signed [14:0] m82_43;
   assign m82_43 =15'b0;

   // m82_44 = W*in
   wire signed [14:0] m82_44;
   assign m82_44 =15'b0;

   // m82_45 = W*in
   wire signed [14:0] m82_45;
   assign m82_45 =15'b0;

   // m82_46 = W*in
   wire signed [14:0] m82_46;
   assign m82_46 =15'b0;

   // m82_47 = W*in
   wire signed [14:0] m82_47;
   assign m82_47 =15'b0;

   // m82_48 = W*in
   wire signed [14:0] m82_48;
   assign m82_48 =15'b0;

   // m82_49 = W*in
   wire signed [14:0] m82_49;
   assign m82_49 =15'b0;

   // m82_50 = W*in
   wire signed [14:0] m82_50;
   assign m82_50 =15'b0;

   // m82_51 = W*in
   wire signed [14:0] m82_51;
   assign m82_51 ={ {4{in82[14]}} , in82[14:4] };

   // m82_52 = W*in
   wire signed [14:0] m82_52;
   assign m82_52 =15'b0;

   // m82_53 = W*in
   wire signed [14:0] m82_53;
   assign m82_53 =15'b0;

   // m82_54 = W*in
   wire signed [14:0] m82_54;
   assign m82_54 =15'b0;

   // m82_55 = W*in
   wire signed [14:0] m82_55;
   assign m82_55 =15'b0;

   // m82_56 = W*in
   wire signed [14:0] m82_56;
   assign m82_56 =15'b0;

   // m82_57 = W*in
   wire signed [14:0] m82_57;
   assign m82_57 ={ {4{neg82[14]}} , neg82[14:4] };

   // m82_58 = W*in
   wire signed [14:0] m82_58;
   assign m82_58 =15'b0;

   // m82_59 = W*in
   wire signed [14:0] m82_59;
   assign m82_59 =15'b0;

   // m82_60 = W*in
   wire signed [14:0] m82_60;
   assign m82_60 =15'b0;

   // m82_61 = W*in
   wire signed [14:0] m82_61;
   assign m82_61 =15'b0;

   // m82_62 = W*in
   wire signed [14:0] m82_62;
   assign m82_62 =15'b0;

   // m82_63 = W*in
   wire signed [14:0] m82_63;
   assign m82_63 ={ {3{in82[14]}} , in82[14:3] };

   // m82_64 = W*in
   wire signed [14:0] m82_64;
   assign m82_64 =15'b0;

   // m82_65 = W*in
   wire signed [14:0] m82_65;
   assign m82_65 =15'b0;

   // m82_66 = W*in
   wire signed [14:0] m82_66;
   assign m82_66 ={ {3{in82[14]}} , in82[14:3] };

   // m82_67 = W*in
   wire signed [14:0] m82_67;
   assign m82_67 =15'b0;

   // m82_68 = W*in
   wire signed [14:0] m82_68;
   assign m82_68 =15'b0;

   // m82_69 = W*in
   wire signed [14:0] m82_69;
   assign m82_69 =15'b0;

   // m82_70 = W*in
   wire signed [14:0] m82_70;
   assign m82_70 =15'b0;

   // m82_71 = W*in
   wire signed [14:0] m82_71;
   assign m82_71 =15'b0;

   // m82_72 = W*in
   wire signed [14:0] m82_72;
   assign m82_72 =15'b0;

   // m82_73 = W*in
   wire signed [14:0] m82_73;
   assign m82_73 =15'b0;

   // m82_74 = W*in
   wire signed [14:0] m82_74;
   assign m82_74 ={ {4{neg82[14]}} , neg82[14:4] };

   // m82_75 = W*in
   wire signed [14:0] m82_75;
   assign m82_75 =15'b0;

   // m82_76 = W*in
   wire signed [14:0] m82_76;
   assign m82_76 =15'b0;

   // m82_77 = W*in
   wire signed [14:0] m82_77;
   assign m82_77 =15'b0;

   // m82_78 = W*in
   wire signed [14:0] m82_78;
   assign m82_78 =15'b0;

   // m82_79 = W*in
   wire signed [14:0] m82_79;
   assign m82_79 ={ {3{in82[14]}} , in82[14:3] };

   // m82_80 = W*in
   wire signed [14:0] m82_80;
   assign m82_80 =15'b0;

   // m82_81 = W*in
   wire signed [14:0] m82_81;
   assign m82_81 =15'b0;

   // m82_82 = W*in
   wire signed [14:0] m82_82;
   assign m82_82 =15'b0;

   // m82_83 = W*in
   wire signed [14:0] m82_83;
   assign m82_83 ={ {3{in82[14]}} , in82[14:3] };

   // m82_84 = W*in
   wire signed [14:0] m82_84;
   assign m82_84 =15'b0;

   // m82_85 = W*in
   wire signed [14:0] m82_85;
   assign m82_85 =15'b0;

   // m82_86 = W*in
   wire signed [14:0] m82_86;
   assign m82_86 =15'b0;

   // m82_87 = W*in
   wire signed [14:0] m82_87;
   assign m82_87 =15'b0;

   // m82_88 = W*in
   wire signed [14:0] m82_88;
   assign m82_88 =15'b0;

   // m82_89 = W*in
   wire signed [14:0] m82_89;
   assign m82_89 =15'b0;

   // m82_90 = W*in
   wire signed [14:0] m82_90;
   assign m82_90 =15'b0;

   // m82_91 = W*in
   wire signed [14:0] m82_91;
   assign m82_91 =15'b0;

   // m82_92 = W*in
   wire signed [14:0] m82_92;
   assign m82_92 =15'b0;

   // m82_93 = W*in
   wire signed [14:0] m82_93;
   assign m82_93 =15'b0;

   // m82_94 = W*in
   wire signed [14:0] m82_94;
   assign m82_94 =15'b0;

   // m82_95 = W*in
   wire signed [14:0] m82_95;
   assign m82_95 =15'b0;

   // m82_96 = W*in
   wire signed [14:0] m82_96;
   assign m82_96 =15'b0;

   // m82_97 = W*in
   wire signed [14:0] m82_97;
   assign m82_97 =15'b0;

   // m82_98 = W*in
   wire signed [14:0] m82_98;
   assign m82_98 =15'b0;

   // m82_99 = W*in
   wire signed [14:0] m82_99;
   assign m82_99 =15'b0;

   // m82_100 = W*in
   wire signed [14:0] m82_100;
   assign m82_100 ={ {3{in82[14]}} , in82[14:3] };

   // m83_1 = W*in
   wire signed [14:0] m83_1;
   assign m83_1 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_2 = W*in
   wire signed [14:0] m83_2;
   assign m83_2 =15'b0;

   // m83_3 = W*in
   wire signed [14:0] m83_3;
   assign m83_3 =15'b0;

   // m83_4 = W*in
   wire signed [14:0] m83_4;
   assign m83_4 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_5 = W*in
   wire signed [14:0] m83_5;
   assign m83_5 =15'b0;

   // m83_6 = W*in
   wire signed [14:0] m83_6;
   assign m83_6 =15'b0;

   // m83_7 = W*in
   wire signed [14:0] m83_7;
   assign m83_7 =15'b0;

   // m83_8 = W*in
   wire signed [14:0] m83_8;
   assign m83_8 =15'b0;

   // m83_9 = W*in
   wire signed [14:0] m83_9;
   assign m83_9 =15'b0;

   // m83_10 = W*in
   wire signed [14:0] m83_10;
   assign m83_10 =15'b0;

   // m83_11 = W*in
   wire signed [14:0] m83_11;
   assign m83_11 =15'b0;

   // m83_12 = W*in
   wire signed [14:0] m83_12;
   assign m83_12 =15'b0;

   // m83_13 = W*in
   wire signed [14:0] m83_13;
   assign m83_13 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_14 = W*in
   wire signed [14:0] m83_14;
   assign m83_14 =15'b0;

   // m83_15 = W*in
   wire signed [14:0] m83_15;
   assign m83_15 =15'b0;

   // m83_16 = W*in
   wire signed [14:0] m83_16;
   assign m83_16 ={ {3{in83[14]}} , in83[14:3] };

   // m83_17 = W*in
   wire signed [14:0] m83_17;
   assign m83_17 =15'b0;

   // m83_18 = W*in
   wire signed [14:0] m83_18;
   assign m83_18 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_19 = W*in
   wire signed [14:0] m83_19;
   assign m83_19 =15'b0;

   // m83_20 = W*in
   wire signed [14:0] m83_20;
   assign m83_20 =15'b0;

   // m83_21 = W*in
   wire signed [14:0] m83_21;
   assign m83_21 =15'b0;

   // m83_22 = W*in
   wire signed [14:0] m83_22;
   assign m83_22 =15'b0;

   // m83_23 = W*in
   wire signed [14:0] m83_23;
   assign m83_23 =15'b0;

   // m83_24 = W*in
   wire signed [14:0] m83_24;
   assign m83_24 =15'b0;

   // m83_25 = W*in
   wire signed [14:0] m83_25;
   assign m83_25 ={ {3{in83[14]}} , in83[14:3] };

   // m83_26 = W*in
   wire signed [14:0] m83_26;
   assign m83_26 =15'b0;

   // m83_27 = W*in
   wire signed [14:0] m83_27;
   assign m83_27 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_28 = W*in
   wire signed [14:0] m83_28;
   assign m83_28 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_29 = W*in
   wire signed [14:0] m83_29;
   assign m83_29 =15'b0;

   // m83_30 = W*in
   wire signed [14:0] m83_30;
   assign m83_30 =15'b0;

   // m83_31 = W*in
   wire signed [14:0] m83_31;
   assign m83_31 =15'b0;

   // m83_32 = W*in
   wire signed [14:0] m83_32;
   assign m83_32 =15'b0;

   // m83_33 = W*in
   wire signed [14:0] m83_33;
   assign m83_33 =15'b0;

   // m83_34 = W*in
   wire signed [14:0] m83_34;
   assign m83_34 =15'b0;

   // m83_35 = W*in
   wire signed [14:0] m83_35;
   assign m83_35 =15'b0;

   // m83_36 = W*in
   wire signed [14:0] m83_36;
   assign m83_36 =15'b0;

   // m83_37 = W*in
   wire signed [14:0] m83_37;
   assign m83_37 =15'b0;

   // m83_38 = W*in
   wire signed [14:0] m83_38;
   assign m83_38 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_39 = W*in
   wire signed [14:0] m83_39;
   assign m83_39 =15'b0;

   // m83_40 = W*in
   wire signed [14:0] m83_40;
   assign m83_40 =15'b0;

   // m83_41 = W*in
   wire signed [14:0] m83_41;
   assign m83_41 =15'b0;

   // m83_42 = W*in
   wire signed [14:0] m83_42;
   assign m83_42 =15'b0;

   // m83_43 = W*in
   wire signed [14:0] m83_43;
   assign m83_43 =15'b0;

   // m83_44 = W*in
   wire signed [14:0] m83_44;
   assign m83_44 =15'b0;

   // m83_45 = W*in
   wire signed [14:0] m83_45;
   assign m83_45 =15'b0;

   // m83_46 = W*in
   wire signed [14:0] m83_46;
   assign m83_46 =15'b0;

   // m83_47 = W*in
   wire signed [14:0] m83_47;
   assign m83_47 ={ {3{in83[14]}} , in83[14:3] };

   // m83_48 = W*in
   wire signed [14:0] m83_48;
   assign m83_48 =15'b0;

   // m83_49 = W*in
   wire signed [14:0] m83_49;
   assign m83_49 =15'b0;

   // m83_50 = W*in
   wire signed [14:0] m83_50;
   assign m83_50 =15'b0;

   // m83_51 = W*in
   wire signed [14:0] m83_51;
   assign m83_51 =15'b0;

   // m83_52 = W*in
   wire signed [14:0] m83_52;
   assign m83_52 =15'b0;

   // m83_53 = W*in
   wire signed [14:0] m83_53;
   assign m83_53 =15'b0;

   // m83_54 = W*in
   wire signed [14:0] m83_54;
   assign m83_54 =15'b0;

   // m83_55 = W*in
   wire signed [14:0] m83_55;
   assign m83_55 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_56 = W*in
   wire signed [14:0] m83_56;
   assign m83_56 =15'b0;

   // m83_57 = W*in
   wire signed [14:0] m83_57;
   assign m83_57 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_58 = W*in
   wire signed [14:0] m83_58;
   assign m83_58 =15'b0;

   // m83_59 = W*in
   wire signed [14:0] m83_59;
   assign m83_59 ={ {3{in83[14]}} , in83[14:3] };

   // m83_60 = W*in
   wire signed [14:0] m83_60;
   assign m83_60 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_61 = W*in
   wire signed [14:0] m83_61;
   assign m83_61 =15'b0;

   // m83_62 = W*in
   wire signed [14:0] m83_62;
   assign m83_62 =15'b0;

   // m83_63 = W*in
   wire signed [14:0] m83_63;
   assign m83_63 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_64 = W*in
   wire signed [14:0] m83_64;
   assign m83_64 =15'b0;

   // m83_65 = W*in
   wire signed [14:0] m83_65;
   assign m83_65 ={ {3{in83[14]}} , in83[14:3] };

   // m83_66 = W*in
   wire signed [14:0] m83_66;
   assign m83_66 =15'b0;

   // m83_67 = W*in
   wire signed [14:0] m83_67;
   assign m83_67 =15'b0;

   // m83_68 = W*in
   wire signed [14:0] m83_68;
   assign m83_68 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_69 = W*in
   wire signed [14:0] m83_69;
   assign m83_69 =15'b0;

   // m83_70 = W*in
   wire signed [14:0] m83_70;
   assign m83_70 =15'b0;

   // m83_71 = W*in
   wire signed [14:0] m83_71;
   assign m83_71 =15'b0;

   // m83_72 = W*in
   wire signed [14:0] m83_72;
   assign m83_72 =15'b0;

   // m83_73 = W*in
   wire signed [14:0] m83_73;
   assign m83_73 =15'b0;

   // m83_74 = W*in
   wire signed [14:0] m83_74;
   assign m83_74 =15'b0;

   // m83_75 = W*in
   wire signed [14:0] m83_75;
   assign m83_75 ={ {4{in83[14]}} , in83[14:4] };

   // m83_76 = W*in
   wire signed [14:0] m83_76;
   assign m83_76 =15'b0;

   // m83_77 = W*in
   wire signed [14:0] m83_77;
   assign m83_77 ={ {4{neg83[14]}} , neg83[14:4] };

   // m83_78 = W*in
   wire signed [14:0] m83_78;
   assign m83_78 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_79 = W*in
   wire signed [14:0] m83_79;
   assign m83_79 =15'b0;

   // m83_80 = W*in
   wire signed [14:0] m83_80;
   assign m83_80 =15'b0;

   // m83_81 = W*in
   wire signed [14:0] m83_81;
   assign m83_81 =15'b0;

   // m83_82 = W*in
   wire signed [14:0] m83_82;
   assign m83_82 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_83 = W*in
   wire signed [14:0] m83_83;
   assign m83_83 =15'b0;

   // m83_84 = W*in
   wire signed [14:0] m83_84;
   assign m83_84 =15'b0;

   // m83_85 = W*in
   wire signed [14:0] m83_85;
   assign m83_85 =15'b0;

   // m83_86 = W*in
   wire signed [14:0] m83_86;
   assign m83_86 =15'b0;

   // m83_87 = W*in
   wire signed [14:0] m83_87;
   assign m83_87 ={ {3{neg83[14]}} , neg83[14:3] };

   // m83_88 = W*in
   wire signed [14:0] m83_88;
   assign m83_88 =15'b0;

   // m83_89 = W*in
   wire signed [14:0] m83_89;
   assign m83_89 =15'b0;

   // m83_90 = W*in
   wire signed [14:0] m83_90;
   assign m83_90 ={ {3{in83[14]}} , in83[14:3] };

   // m83_91 = W*in
   wire signed [14:0] m83_91;
   assign m83_91 =15'b0;

   // m83_92 = W*in
   wire signed [14:0] m83_92;
   assign m83_92 =15'b0;

   // m83_93 = W*in
   wire signed [14:0] m83_93;
   assign m83_93 =15'b0;

   // m83_94 = W*in
   wire signed [14:0] m83_94;
   assign m83_94 =15'b0;

   // m83_95 = W*in
   wire signed [14:0] m83_95;
   assign m83_95 =15'b0;

   // m83_96 = W*in
   wire signed [14:0] m83_96;
   assign m83_96 =15'b0;

   // m83_97 = W*in
   wire signed [14:0] m83_97;
   assign m83_97 =15'b0;

   // m83_98 = W*in
   wire signed [14:0] m83_98;
   assign m83_98 =15'b0;

   // m83_99 = W*in
   wire signed [14:0] m83_99;
   assign m83_99 =15'b0;

   // m83_100 = W*in
   wire signed [14:0] m83_100;
   assign m83_100 =15'b0;

   // m84_1 = W*in
   wire signed [14:0] m84_1;
   assign m84_1 =15'b0;

   // m84_2 = W*in
   wire signed [14:0] m84_2;
   assign m84_2 =15'b0;

   // m84_3 = W*in
   wire signed [14:0] m84_3;
   assign m84_3 =15'b0;

   // m84_4 = W*in
   wire signed [14:0] m84_4;
   assign m84_4 =15'b0;

   // m84_5 = W*in
   wire signed [14:0] m84_5;
   assign m84_5 =15'b0;

   // m84_6 = W*in
   wire signed [14:0] m84_6;
   assign m84_6 =15'b0;

   // m84_7 = W*in
   wire signed [14:0] m84_7;
   assign m84_7 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_8 = W*in
   wire signed [14:0] m84_8;
   assign m84_8 =15'b0;

   // m84_9 = W*in
   wire signed [14:0] m84_9;
   assign m84_9 =15'b0;

   // m84_10 = W*in
   wire signed [14:0] m84_10;
   assign m84_10 =15'b0;

   // m84_11 = W*in
   wire signed [14:0] m84_11;
   assign m84_11 =15'b0;

   // m84_12 = W*in
   wire signed [14:0] m84_12;
   assign m84_12 =15'b0;

   // m84_13 = W*in
   wire signed [14:0] m84_13;
   assign m84_13 =15'b0;

   // m84_14 = W*in
   wire signed [14:0] m84_14;
   assign m84_14 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_15 = W*in
   wire signed [14:0] m84_15;
   assign m84_15 =15'b0;

   // m84_16 = W*in
   wire signed [14:0] m84_16;
   assign m84_16 =15'b0;

   // m84_17 = W*in
   wire signed [14:0] m84_17;
   assign m84_17 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_18 = W*in
   wire signed [14:0] m84_18;
   assign m84_18 =15'b0;

   // m84_19 = W*in
   wire signed [14:0] m84_19;
   assign m84_19 =15'b0;

   // m84_20 = W*in
   wire signed [14:0] m84_20;
   assign m84_20 =15'b0;

   // m84_21 = W*in
   wire signed [14:0] m84_21;
   assign m84_21 ={ {4{in84[14]}} , in84[14:4] };

   // m84_22 = W*in
   wire signed [14:0] m84_22;
   assign m84_22 =15'b0;

   // m84_23 = W*in
   wire signed [14:0] m84_23;
   assign m84_23 =15'b0;

   // m84_24 = W*in
   wire signed [14:0] m84_24;
   assign m84_24 =15'b0;

   // m84_25 = W*in
   wire signed [14:0] m84_25;
   assign m84_25 =15'b0;

   // m84_26 = W*in
   wire signed [14:0] m84_26;
   assign m84_26 =15'b0;

   // m84_27 = W*in
   wire signed [14:0] m84_27;
   assign m84_27 =15'b0;

   // m84_28 = W*in
   wire signed [14:0] m84_28;
   assign m84_28 ={ {4{neg84[14]}} , neg84[14:4] };

   // m84_29 = W*in
   wire signed [14:0] m84_29;
   assign m84_29 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_30 = W*in
   wire signed [14:0] m84_30;
   assign m84_30 =15'b0;

   // m84_31 = W*in
   wire signed [14:0] m84_31;
   assign m84_31 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_32 = W*in
   wire signed [14:0] m84_32;
   assign m84_32 ={ {4{neg84[14]}} , neg84[14:4] };

   // m84_33 = W*in
   wire signed [14:0] m84_33;
   assign m84_33 ={ {4{neg84[14]}} , neg84[14:4] };

   // m84_34 = W*in
   wire signed [14:0] m84_34;
   assign m84_34 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_35 = W*in
   wire signed [14:0] m84_35;
   assign m84_35 =15'b0;

   // m84_36 = W*in
   wire signed [14:0] m84_36;
   assign m84_36 ={ {3{in84[14]}} , in84[14:3] };

   // m84_37 = W*in
   wire signed [14:0] m84_37;
   assign m84_37 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_38 = W*in
   wire signed [14:0] m84_38;
   assign m84_38 =15'b0;

   // m84_39 = W*in
   wire signed [14:0] m84_39;
   assign m84_39 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_40 = W*in
   wire signed [14:0] m84_40;
   assign m84_40 =15'b0;

   // m84_41 = W*in
   wire signed [14:0] m84_41;
   assign m84_41 =15'b0;

   // m84_42 = W*in
   wire signed [14:0] m84_42;
   assign m84_42 =15'b0;

   // m84_43 = W*in
   wire signed [14:0] m84_43;
   assign m84_43 ={ {3{in84[14]}} , in84[14:3] };

   // m84_44 = W*in
   wire signed [14:0] m84_44;
   assign m84_44 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_45 = W*in
   wire signed [14:0] m84_45;
   assign m84_45 =15'b0;

   // m84_46 = W*in
   wire signed [14:0] m84_46;
   assign m84_46 =15'b0;

   // m84_47 = W*in
   wire signed [14:0] m84_47;
   assign m84_47 =15'b0;

   // m84_48 = W*in
   wire signed [14:0] m84_48;
   assign m84_48 =15'b0;

   // m84_49 = W*in
   wire signed [14:0] m84_49;
   assign m84_49 ={ {3{in84[14]}} , in84[14:3] };

   // m84_50 = W*in
   wire signed [14:0] m84_50;
   assign m84_50 =15'b0;

   // m84_51 = W*in
   wire signed [14:0] m84_51;
   assign m84_51 =15'b0;

   // m84_52 = W*in
   wire signed [14:0] m84_52;
   assign m84_52 =15'b0;

   // m84_53 = W*in
   wire signed [14:0] m84_53;
   assign m84_53 =15'b0;

   // m84_54 = W*in
   wire signed [14:0] m84_54;
   assign m84_54 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_55 = W*in
   wire signed [14:0] m84_55;
   assign m84_55 =15'b0;

   // m84_56 = W*in
   wire signed [14:0] m84_56;
   assign m84_56 =15'b0;

   // m84_57 = W*in
   wire signed [14:0] m84_57;
   assign m84_57 ={ {4{in84[14]}} , in84[14:4] };

   // m84_58 = W*in
   wire signed [14:0] m84_58;
   assign m84_58 ={ {4{in84[14]}} , in84[14:4] };

   // m84_59 = W*in
   wire signed [14:0] m84_59;
   assign m84_59 ={ {4{in84[14]}} , in84[14:4] };

   // m84_60 = W*in
   wire signed [14:0] m84_60;
   assign m84_60 =15'b0;

   // m84_61 = W*in
   wire signed [14:0] m84_61;
   assign m84_61 ={ {3{in84[14]}} , in84[14:3] };

   // m84_62 = W*in
   wire signed [14:0] m84_62;
   assign m84_62 =15'b0;

   // m84_63 = W*in
   wire signed [14:0] m84_63;
   assign m84_63 =15'b0;

   // m84_64 = W*in
   wire signed [14:0] m84_64;
   assign m84_64 ={ {3{in84[14]}} , in84[14:3] };

   // m84_65 = W*in
   wire signed [14:0] m84_65;
   assign m84_65 =15'b0;

   // m84_66 = W*in
   wire signed [14:0] m84_66;
   assign m84_66 ={ {4{neg84[14]}} , neg84[14:4] };

   // m84_67 = W*in
   wire signed [14:0] m84_67;
   assign m84_67 ={ {3{in84[14]}} , in84[14:3] };

   // m84_68 = W*in
   wire signed [14:0] m84_68;
   assign m84_68 ={ {4{in84[14]}} , in84[14:4] };

   // m84_69 = W*in
   wire signed [14:0] m84_69;
   assign m84_69 =15'b0;

   // m84_70 = W*in
   wire signed [14:0] m84_70;
   assign m84_70 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_71 = W*in
   wire signed [14:0] m84_71;
   assign m84_71 =15'b0;

   // m84_72 = W*in
   wire signed [14:0] m84_72;
   assign m84_72 =15'b0;

   // m84_73 = W*in
   wire signed [14:0] m84_73;
   assign m84_73 ={ {3{in84[14]}} , in84[14:3] };

   // m84_74 = W*in
   wire signed [14:0] m84_74;
   assign m84_74 =15'b0;

   // m84_75 = W*in
   wire signed [14:0] m84_75;
   assign m84_75 =15'b0;

   // m84_76 = W*in
   wire signed [14:0] m84_76;
   assign m84_76 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_77 = W*in
   wire signed [14:0] m84_77;
   assign m84_77 ={ {3{in84[14]}} , in84[14:3] };

   // m84_78 = W*in
   wire signed [14:0] m84_78;
   assign m84_78 =15'b0;

   // m84_79 = W*in
   wire signed [14:0] m84_79;
   assign m84_79 =15'b0;

   // m84_80 = W*in
   wire signed [14:0] m84_80;
   assign m84_80 ={ {3{neg84[14]}} , neg84[14:3] };

   // m84_81 = W*in
   wire signed [14:0] m84_81;
   assign m84_81 =15'b0;

   // m84_82 = W*in
   wire signed [14:0] m84_82;
   assign m84_82 =15'b0;

   // m84_83 = W*in
   wire signed [14:0] m84_83;
   assign m84_83 =15'b0;

   // m84_84 = W*in
   wire signed [14:0] m84_84;
   assign m84_84 =15'b0;

   // m84_85 = W*in
   wire signed [14:0] m84_85;
   assign m84_85 =15'b0;

   // m84_86 = W*in
   wire signed [14:0] m84_86;
   assign m84_86 =15'b0;

   // m84_87 = W*in
   wire signed [14:0] m84_87;
   assign m84_87 =15'b0;

   // m84_88 = W*in
   wire signed [14:0] m84_88;
   assign m84_88 =15'b0;

   // m84_89 = W*in
   wire signed [14:0] m84_89;
   assign m84_89 =15'b0;

   // m84_90 = W*in
   wire signed [14:0] m84_90;
   assign m84_90 =15'b0;

   // m84_91 = W*in
   wire signed [14:0] m84_91;
   assign m84_91 =15'b0;

   // m84_92 = W*in
   wire signed [14:0] m84_92;
   assign m84_92 ={ {3{in84[14]}} , in84[14:3] };

   // m84_93 = W*in
   wire signed [14:0] m84_93;
   assign m84_93 =15'b0;

   // m84_94 = W*in
   wire signed [14:0] m84_94;
   assign m84_94 =15'b0;

   // m84_95 = W*in
   wire signed [14:0] m84_95;
   assign m84_95 =15'b0;

   // m84_96 = W*in
   wire signed [14:0] m84_96;
   assign m84_96 ={ {4{neg84[14]}} , neg84[14:4] };

   // m84_97 = W*in
   wire signed [14:0] m84_97;
   assign m84_97 =15'b0;

   // m84_98 = W*in
   wire signed [14:0] m84_98;
   assign m84_98 =15'b0;

   // m84_99 = W*in
   wire signed [14:0] m84_99;
   assign m84_99 =15'b0;

   // m84_100 = W*in
   wire signed [14:0] m84_100;
   assign m84_100 ={ {3{neg84[14]}} , neg84[14:3] };

   // m85_1 = W*in
   wire signed [14:0] m85_1;
   assign m85_1 =15'b0;

   // m85_2 = W*in
   wire signed [14:0] m85_2;
   assign m85_2 =15'b0;

   // m85_3 = W*in
   wire signed [14:0] m85_3;
   assign m85_3 =15'b0;

   // m85_4 = W*in
   wire signed [14:0] m85_4;
   assign m85_4 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_5 = W*in
   wire signed [14:0] m85_5;
   assign m85_5 =15'b0;

   // m85_6 = W*in
   wire signed [14:0] m85_6;
   assign m85_6 =15'b0;

   // m85_7 = W*in
   wire signed [14:0] m85_7;
   assign m85_7 =15'b0;

   // m85_8 = W*in
   wire signed [14:0] m85_8;
   assign m85_8 =15'b0;

   // m85_9 = W*in
   wire signed [14:0] m85_9;
   assign m85_9 =15'b0;

   // m85_10 = W*in
   wire signed [14:0] m85_10;
   assign m85_10 =15'b0;

   // m85_11 = W*in
   wire signed [14:0] m85_11;
   assign m85_11 =15'b0;

   // m85_12 = W*in
   wire signed [14:0] m85_12;
   assign m85_12 =15'b0;

   // m85_13 = W*in
   wire signed [14:0] m85_13;
   assign m85_13 =15'b0;

   // m85_14 = W*in
   wire signed [14:0] m85_14;
   assign m85_14 =15'b0;

   // m85_15 = W*in
   wire signed [14:0] m85_15;
   assign m85_15 =15'b0;

   // m85_16 = W*in
   wire signed [14:0] m85_16;
   assign m85_16 =15'b0;

   // m85_17 = W*in
   wire signed [14:0] m85_17;
   assign m85_17 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_18 = W*in
   wire signed [14:0] m85_18;
   assign m85_18 =15'b0;

   // m85_19 = W*in
   wire signed [14:0] m85_19;
   assign m85_19 =15'b0;

   // m85_20 = W*in
   wire signed [14:0] m85_20;
   assign m85_20 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_21 = W*in
   wire signed [14:0] m85_21;
   assign m85_21 =15'b0;

   // m85_22 = W*in
   wire signed [14:0] m85_22;
   assign m85_22 =15'b0;

   // m85_23 = W*in
   wire signed [14:0] m85_23;
   assign m85_23 =15'b0;

   // m85_24 = W*in
   wire signed [14:0] m85_24;
   assign m85_24 =15'b0;

   // m85_25 = W*in
   wire signed [14:0] m85_25;
   assign m85_25 =15'b0;

   // m85_26 = W*in
   wire signed [14:0] m85_26;
   assign m85_26 ={ {3{in85[14]}} , in85[14:3] };

   // m85_27 = W*in
   wire signed [14:0] m85_27;
   assign m85_27 =15'b0;

   // m85_28 = W*in
   wire signed [14:0] m85_28;
   assign m85_28 =15'b0;

   // m85_29 = W*in
   wire signed [14:0] m85_29;
   assign m85_29 ={ {3{in85[14]}} , in85[14:3] };

   // m85_30 = W*in
   wire signed [14:0] m85_30;
   assign m85_30 =15'b0;

   // m85_31 = W*in
   wire signed [14:0] m85_31;
   assign m85_31 =15'b0;

   // m85_32 = W*in
   wire signed [14:0] m85_32;
   assign m85_32 =15'b0;

   // m85_33 = W*in
   wire signed [14:0] m85_33;
   assign m85_33 =15'b0;

   // m85_34 = W*in
   wire signed [14:0] m85_34;
   assign m85_34 ={ {3{in85[14]}} , in85[14:3] };

   // m85_35 = W*in
   wire signed [14:0] m85_35;
   assign m85_35 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_36 = W*in
   wire signed [14:0] m85_36;
   assign m85_36 =15'b0;

   // m85_37 = W*in
   wire signed [14:0] m85_37;
   assign m85_37 =15'b0;

   // m85_38 = W*in
   wire signed [14:0] m85_38;
   assign m85_38 =15'b0;

   // m85_39 = W*in
   wire signed [14:0] m85_39;
   assign m85_39 =15'b0;

   // m85_40 = W*in
   wire signed [14:0] m85_40;
   assign m85_40 =15'b0;

   // m85_41 = W*in
   wire signed [14:0] m85_41;
   assign m85_41 =15'b0;

   // m85_42 = W*in
   wire signed [14:0] m85_42;
   assign m85_42 =15'b0;

   // m85_43 = W*in
   wire signed [14:0] m85_43;
   assign m85_43 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_44 = W*in
   wire signed [14:0] m85_44;
   assign m85_44 ={ {4{neg85[14]}} , neg85[14:4] };

   // m85_45 = W*in
   wire signed [14:0] m85_45;
   assign m85_45 =15'b0;

   // m85_46 = W*in
   wire signed [14:0] m85_46;
   assign m85_46 =15'b0;

   // m85_47 = W*in
   wire signed [14:0] m85_47;
   assign m85_47 =15'b0;

   // m85_48 = W*in
   wire signed [14:0] m85_48;
   assign m85_48 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_49 = W*in
   wire signed [14:0] m85_49;
   assign m85_49 ={ {3{in85[14]}} , in85[14:3] };

   // m85_50 = W*in
   wire signed [14:0] m85_50;
   assign m85_50 ={ {4{in85[14]}} , in85[14:4] };

   // m85_51 = W*in
   wire signed [14:0] m85_51;
   assign m85_51 =15'b0;

   // m85_52 = W*in
   wire signed [14:0] m85_52;
   assign m85_52 ={ {3{in85[14]}} , in85[14:3] };

   // m85_53 = W*in
   wire signed [14:0] m85_53;
   assign m85_53 =15'b0;

   // m85_54 = W*in
   wire signed [14:0] m85_54;
   assign m85_54 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_55 = W*in
   wire signed [14:0] m85_55;
   assign m85_55 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_56 = W*in
   wire signed [14:0] m85_56;
   assign m85_56 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_57 = W*in
   wire signed [14:0] m85_57;
   assign m85_57 =15'b0;

   // m85_58 = W*in
   wire signed [14:0] m85_58;
   assign m85_58 =15'b0;

   // m85_59 = W*in
   wire signed [14:0] m85_59;
   assign m85_59 =15'b0;

   // m85_60 = W*in
   wire signed [14:0] m85_60;
   assign m85_60 =15'b0;

   // m85_61 = W*in
   wire signed [14:0] m85_61;
   assign m85_61 =15'b0;

   // m85_62 = W*in
   wire signed [14:0] m85_62;
   assign m85_62 =15'b0;

   // m85_63 = W*in
   wire signed [14:0] m85_63;
   assign m85_63 =15'b0;

   // m85_64 = W*in
   wire signed [14:0] m85_64;
   assign m85_64 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_65 = W*in
   wire signed [14:0] m85_65;
   assign m85_65 =15'b0;

   // m85_66 = W*in
   wire signed [14:0] m85_66;
   assign m85_66 =15'b0;

   // m85_67 = W*in
   wire signed [14:0] m85_67;
   assign m85_67 =15'b0;

   // m85_68 = W*in
   wire signed [14:0] m85_68;
   assign m85_68 =15'b0;

   // m85_69 = W*in
   wire signed [14:0] m85_69;
   assign m85_69 =15'b0;

   // m85_70 = W*in
   wire signed [14:0] m85_70;
   assign m85_70 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_71 = W*in
   wire signed [14:0] m85_71;
   assign m85_71 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_72 = W*in
   wire signed [14:0] m85_72;
   assign m85_72 =15'b0;

   // m85_73 = W*in
   wire signed [14:0] m85_73;
   assign m85_73 =15'b0;

   // m85_74 = W*in
   wire signed [14:0] m85_74;
   assign m85_74 =15'b0;

   // m85_75 = W*in
   wire signed [14:0] m85_75;
   assign m85_75 =15'b0;

   // m85_76 = W*in
   wire signed [14:0] m85_76;
   assign m85_76 =15'b0;

   // m85_77 = W*in
   wire signed [14:0] m85_77;
   assign m85_77 =15'b0;

   // m85_78 = W*in
   wire signed [14:0] m85_78;
   assign m85_78 =15'b0;

   // m85_79 = W*in
   wire signed [14:0] m85_79;
   assign m85_79 =15'b0;

   // m85_80 = W*in
   wire signed [14:0] m85_80;
   assign m85_80 =15'b0;

   // m85_81 = W*in
   wire signed [14:0] m85_81;
   assign m85_81 =15'b0;

   // m85_82 = W*in
   wire signed [14:0] m85_82;
   assign m85_82 =15'b0;

   // m85_83 = W*in
   wire signed [14:0] m85_83;
   assign m85_83 =15'b0;

   // m85_84 = W*in
   wire signed [14:0] m85_84;
   assign m85_84 =15'b0;

   // m85_85 = W*in
   wire signed [14:0] m85_85;
   assign m85_85 =15'b0;

   // m85_86 = W*in
   wire signed [14:0] m85_86;
   assign m85_86 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_87 = W*in
   wire signed [14:0] m85_87;
   assign m85_87 =15'b0;

   // m85_88 = W*in
   wire signed [14:0] m85_88;
   assign m85_88 =15'b0;

   // m85_89 = W*in
   wire signed [14:0] m85_89;
   assign m85_89 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_90 = W*in
   wire signed [14:0] m85_90;
   assign m85_90 ={ {4{neg85[14]}} , neg85[14:4] };

   // m85_91 = W*in
   wire signed [14:0] m85_91;
   assign m85_91 =15'b0;

   // m85_92 = W*in
   wire signed [14:0] m85_92;
   assign m85_92 =15'b0;

   // m85_93 = W*in
   wire signed [14:0] m85_93;
   assign m85_93 =15'b0;

   // m85_94 = W*in
   wire signed [14:0] m85_94;
   assign m85_94 ={ {3{neg85[14]}} , neg85[14:3] };

   // m85_95 = W*in
   wire signed [14:0] m85_95;
   assign m85_95 ={ {4{neg85[14]}} , neg85[14:4] };

   // m85_96 = W*in
   wire signed [14:0] m85_96;
   assign m85_96 =15'b0;

   // m85_97 = W*in
   wire signed [14:0] m85_97;
   assign m85_97 =15'b0;

   // m85_98 = W*in
   wire signed [14:0] m85_98;
   assign m85_98 =15'b0;

   // m85_99 = W*in
   wire signed [14:0] m85_99;
   assign m85_99 =15'b0;

   // m85_100 = W*in
   wire signed [14:0] m85_100;
   assign m85_100 =15'b0;

   // m86_1 = W*in
   wire signed [14:0] m86_1;
   assign m86_1 =15'b0;

   // m86_2 = W*in
   wire signed [14:0] m86_2;
   assign m86_2 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_3 = W*in
   wire signed [14:0] m86_3;
   assign m86_3 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_4 = W*in
   wire signed [14:0] m86_4;
   assign m86_4 =15'b0;

   // m86_5 = W*in
   wire signed [14:0] m86_5;
   assign m86_5 =15'b0;

   // m86_6 = W*in
   wire signed [14:0] m86_6;
   assign m86_6 =15'b0;

   // m86_7 = W*in
   wire signed [14:0] m86_7;
   assign m86_7 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_8 = W*in
   wire signed [14:0] m86_8;
   assign m86_8 =15'b0;

   // m86_9 = W*in
   wire signed [14:0] m86_9;
   assign m86_9 =15'b0;

   // m86_10 = W*in
   wire signed [14:0] m86_10;
   assign m86_10 =15'b0;

   // m86_11 = W*in
   wire signed [14:0] m86_11;
   assign m86_11 ={ {3{in86[14]}} , in86[14:3] };

   // m86_12 = W*in
   wire signed [14:0] m86_12;
   assign m86_12 =15'b0;

   // m86_13 = W*in
   wire signed [14:0] m86_13;
   assign m86_13 =15'b0;

   // m86_14 = W*in
   wire signed [14:0] m86_14;
   assign m86_14 =15'b0;

   // m86_15 = W*in
   wire signed [14:0] m86_15;
   assign m86_15 =15'b0;

   // m86_16 = W*in
   wire signed [14:0] m86_16;
   assign m86_16 =15'b0;

   // m86_17 = W*in
   wire signed [14:0] m86_17;
   assign m86_17 ={ {3{in86[14]}} , in86[14:3] };

   // m86_18 = W*in
   wire signed [14:0] m86_18;
   assign m86_18 =15'b0;

   // m86_19 = W*in
   wire signed [14:0] m86_19;
   assign m86_19 =15'b0;

   // m86_20 = W*in
   wire signed [14:0] m86_20;
   assign m86_20 =15'b0;

   // m86_21 = W*in
   wire signed [14:0] m86_21;
   assign m86_21 ={ {3{in86[14]}} , in86[14:3] };

   // m86_22 = W*in
   wire signed [14:0] m86_22;
   assign m86_22 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_23 = W*in
   wire signed [14:0] m86_23;
   assign m86_23 =15'b0;

   // m86_24 = W*in
   wire signed [14:0] m86_24;
   assign m86_24 =15'b0;

   // m86_25 = W*in
   wire signed [14:0] m86_25;
   assign m86_25 ={ {3{in86[14]}} , in86[14:3] };

   // m86_26 = W*in
   wire signed [14:0] m86_26;
   assign m86_26 ={ {4{neg86[14]}} , neg86[14:4] };

   // m86_27 = W*in
   wire signed [14:0] m86_27;
   assign m86_27 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_28 = W*in
   wire signed [14:0] m86_28;
   assign m86_28 =15'b0;

   // m86_29 = W*in
   wire signed [14:0] m86_29;
   assign m86_29 ={ {4{neg86[14]}} , neg86[14:4] };

   // m86_30 = W*in
   wire signed [14:0] m86_30;
   assign m86_30 =15'b0;

   // m86_31 = W*in
   wire signed [14:0] m86_31;
   assign m86_31 =15'b0;

   // m86_32 = W*in
   wire signed [14:0] m86_32;
   assign m86_32 =15'b0;

   // m86_33 = W*in
   wire signed [14:0] m86_33;
   assign m86_33 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_34 = W*in
   wire signed [14:0] m86_34;
   assign m86_34 =15'b0;

   // m86_35 = W*in
   wire signed [14:0] m86_35;
   assign m86_35 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_36 = W*in
   wire signed [14:0] m86_36;
   assign m86_36 =15'b0;

   // m86_37 = W*in
   wire signed [14:0] m86_37;
   assign m86_37 =15'b0;

   // m86_38 = W*in
   wire signed [14:0] m86_38;
   assign m86_38 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_39 = W*in
   wire signed [14:0] m86_39;
   assign m86_39 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_40 = W*in
   wire signed [14:0] m86_40;
   assign m86_40 =15'b0;

   // m86_41 = W*in
   wire signed [14:0] m86_41;
   assign m86_41 ={ {4{in86[14]}} , in86[14:4] };

   // m86_42 = W*in
   wire signed [14:0] m86_42;
   assign m86_42 =15'b0;

   // m86_43 = W*in
   wire signed [14:0] m86_43;
   assign m86_43 =15'b0;

   // m86_44 = W*in
   wire signed [14:0] m86_44;
   assign m86_44 =15'b0;

   // m86_45 = W*in
   wire signed [14:0] m86_45;
   assign m86_45 =15'b0;

   // m86_46 = W*in
   wire signed [14:0] m86_46;
   assign m86_46 =15'b0;

   // m86_47 = W*in
   wire signed [14:0] m86_47;
   assign m86_47 ={ {4{in86[14]}} , in86[14:4] };

   // m86_48 = W*in
   wire signed [14:0] m86_48;
   assign m86_48 =15'b0;

   // m86_49 = W*in
   wire signed [14:0] m86_49;
   assign m86_49 ={ {3{in86[14]}} , in86[14:3] };

   // m86_50 = W*in
   wire signed [14:0] m86_50;
   assign m86_50 =15'b0;

   // m86_51 = W*in
   wire signed [14:0] m86_51;
   assign m86_51 =15'b0;

   // m86_52 = W*in
   wire signed [14:0] m86_52;
   assign m86_52 =15'b0;

   // m86_53 = W*in
   wire signed [14:0] m86_53;
   assign m86_53 =15'b0;

   // m86_54 = W*in
   wire signed [14:0] m86_54;
   assign m86_54 =15'b0;

   // m86_55 = W*in
   wire signed [14:0] m86_55;
   assign m86_55 =15'b0;

   // m86_56 = W*in
   wire signed [14:0] m86_56;
   assign m86_56 =15'b0;

   // m86_57 = W*in
   wire signed [14:0] m86_57;
   assign m86_57 ={ {4{neg86[14]}} , neg86[14:4] };

   // m86_58 = W*in
   wire signed [14:0] m86_58;
   assign m86_58 ={ {4{neg86[14]}} , neg86[14:4] };

   // m86_59 = W*in
   wire signed [14:0] m86_59;
   assign m86_59 ={ {4{in86[14]}} , in86[14:4] };

   // m86_60 = W*in
   wire signed [14:0] m86_60;
   assign m86_60 =15'b0;

   // m86_61 = W*in
   wire signed [14:0] m86_61;
   assign m86_61 =15'b0;

   // m86_62 = W*in
   wire signed [14:0] m86_62;
   assign m86_62 =15'b0;

   // m86_63 = W*in
   wire signed [14:0] m86_63;
   assign m86_63 =15'b0;

   // m86_64 = W*in
   wire signed [14:0] m86_64;
   assign m86_64 ={ {4{in86[14]}} , in86[14:4] };

   // m86_65 = W*in
   wire signed [14:0] m86_65;
   assign m86_65 =15'b0;

   // m86_66 = W*in
   wire signed [14:0] m86_66;
   assign m86_66 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_67 = W*in
   wire signed [14:0] m86_67;
   assign m86_67 ={ {4{in86[14]}} , in86[14:4] };

   // m86_68 = W*in
   wire signed [14:0] m86_68;
   assign m86_68 =15'b0;

   // m86_69 = W*in
   wire signed [14:0] m86_69;
   assign m86_69 ={ {3{in86[14]}} , in86[14:3] };

   // m86_70 = W*in
   wire signed [14:0] m86_70;
   assign m86_70 ={ {3{in86[14]}} , in86[14:3] };

   // m86_71 = W*in
   wire signed [14:0] m86_71;
   assign m86_71 =15'b0;

   // m86_72 = W*in
   wire signed [14:0] m86_72;
   assign m86_72 =15'b0;

   // m86_73 = W*in
   wire signed [14:0] m86_73;
   assign m86_73 ={ {3{in86[14]}} , in86[14:3] };

   // m86_74 = W*in
   wire signed [14:0] m86_74;
   assign m86_74 ={ {4{neg86[14]}} , neg86[14:4] };

   // m86_75 = W*in
   wire signed [14:0] m86_75;
   assign m86_75 =15'b0;

   // m86_76 = W*in
   wire signed [14:0] m86_76;
   assign m86_76 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_77 = W*in
   wire signed [14:0] m86_77;
   assign m86_77 ={ {3{in86[14]}} , in86[14:3] };

   // m86_78 = W*in
   wire signed [14:0] m86_78;
   assign m86_78 =15'b0;

   // m86_79 = W*in
   wire signed [14:0] m86_79;
   assign m86_79 =15'b0;

   // m86_80 = W*in
   wire signed [14:0] m86_80;
   assign m86_80 =15'b0;

   // m86_81 = W*in
   wire signed [14:0] m86_81;
   assign m86_81 =15'b0;

   // m86_82 = W*in
   wire signed [14:0] m86_82;
   assign m86_82 =15'b0;

   // m86_83 = W*in
   wire signed [14:0] m86_83;
   assign m86_83 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_84 = W*in
   wire signed [14:0] m86_84;
   assign m86_84 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_85 = W*in
   wire signed [14:0] m86_85;
   assign m86_85 =15'b0;

   // m86_86 = W*in
   wire signed [14:0] m86_86;
   assign m86_86 =15'b0;

   // m86_87 = W*in
   wire signed [14:0] m86_87;
   assign m86_87 =15'b0;

   // m86_88 = W*in
   wire signed [14:0] m86_88;
   assign m86_88 =15'b0;

   // m86_89 = W*in
   wire signed [14:0] m86_89;
   assign m86_89 =15'b0;

   // m86_90 = W*in
   wire signed [14:0] m86_90;
   assign m86_90 =15'b0;

   // m86_91 = W*in
   wire signed [14:0] m86_91;
   assign m86_91 =15'b0;

   // m86_92 = W*in
   wire signed [14:0] m86_92;
   assign m86_92 =15'b0;

   // m86_93 = W*in
   wire signed [14:0] m86_93;
   assign m86_93 =15'b0;

   // m86_94 = W*in
   wire signed [14:0] m86_94;
   assign m86_94 =15'b0;

   // m86_95 = W*in
   wire signed [14:0] m86_95;
   assign m86_95 ={ {3{in86[14]}} , in86[14:3] };

   // m86_96 = W*in
   wire signed [14:0] m86_96;
   assign m86_96 =15'b0;

   // m86_97 = W*in
   wire signed [14:0] m86_97;
   assign m86_97 ={ {3{neg86[14]}} , neg86[14:3] };

   // m86_98 = W*in
   wire signed [14:0] m86_98;
   assign m86_98 ={ {3{in86[14]}} , in86[14:3] };

   // m86_99 = W*in
   wire signed [14:0] m86_99;
   assign m86_99 =15'b0;

   // m86_100 = W*in
   wire signed [14:0] m86_100;
   assign m86_100 ={ {3{neg86[14]}} , neg86[14:3] };

   // m87_1 = W*in
   wire signed [14:0] m87_1;
   assign m87_1 =15'b0;

   // m87_2 = W*in
   wire signed [14:0] m87_2;
   assign m87_2 =15'b0;

   // m87_3 = W*in
   wire signed [14:0] m87_3;
   assign m87_3 =15'b0;

   // m87_4 = W*in
   wire signed [14:0] m87_4;
   assign m87_4 =15'b0;

   // m87_5 = W*in
   wire signed [14:0] m87_5;
   assign m87_5 =15'b0;

   // m87_6 = W*in
   wire signed [14:0] m87_6;
   assign m87_6 =15'b0;

   // m87_7 = W*in
   wire signed [14:0] m87_7;
   assign m87_7 =15'b0;

   // m87_8 = W*in
   wire signed [14:0] m87_8;
   assign m87_8 =15'b0;

   // m87_9 = W*in
   wire signed [14:0] m87_9;
   assign m87_9 =15'b0;

   // m87_10 = W*in
   wire signed [14:0] m87_10;
   assign m87_10 =15'b0;

   // m87_11 = W*in
   wire signed [14:0] m87_11;
   assign m87_11 =15'b0;

   // m87_12 = W*in
   wire signed [14:0] m87_12;
   assign m87_12 =15'b0;

   // m87_13 = W*in
   wire signed [14:0] m87_13;
   assign m87_13 =15'b0;

   // m87_14 = W*in
   wire signed [14:0] m87_14;
   assign m87_14 =15'b0;

   // m87_15 = W*in
   wire signed [14:0] m87_15;
   assign m87_15 =15'b0;

   // m87_16 = W*in
   wire signed [14:0] m87_16;
   assign m87_16 =15'b0;

   // m87_17 = W*in
   wire signed [14:0] m87_17;
   assign m87_17 =15'b0;

   // m87_18 = W*in
   wire signed [14:0] m87_18;
   assign m87_18 =15'b0;

   // m87_19 = W*in
   wire signed [14:0] m87_19;
   assign m87_19 =15'b0;

   // m87_20 = W*in
   wire signed [14:0] m87_20;
   assign m87_20 =15'b0;

   // m87_21 = W*in
   wire signed [14:0] m87_21;
   assign m87_21 =15'b0;

   // m87_22 = W*in
   wire signed [14:0] m87_22;
   assign m87_22 =15'b0;

   // m87_23 = W*in
   wire signed [14:0] m87_23;
   assign m87_23 ={ {3{in87[14]}} , in87[14:3] };

   // m87_24 = W*in
   wire signed [14:0] m87_24;
   assign m87_24 =15'b0;

   // m87_25 = W*in
   wire signed [14:0] m87_25;
   assign m87_25 =15'b0;

   // m87_26 = W*in
   wire signed [14:0] m87_26;
   assign m87_26 =15'b0;

   // m87_27 = W*in
   wire signed [14:0] m87_27;
   assign m87_27 =15'b0;

   // m87_28 = W*in
   wire signed [14:0] m87_28;
   assign m87_28 =15'b0;

   // m87_29 = W*in
   wire signed [14:0] m87_29;
   assign m87_29 =15'b0;

   // m87_30 = W*in
   wire signed [14:0] m87_30;
   assign m87_30 =15'b0;

   // m87_31 = W*in
   wire signed [14:0] m87_31;
   assign m87_31 =15'b0;

   // m87_32 = W*in
   wire signed [14:0] m87_32;
   assign m87_32 =15'b0;

   // m87_33 = W*in
   wire signed [14:0] m87_33;
   assign m87_33 =15'b0;

   // m87_34 = W*in
   wire signed [14:0] m87_34;
   assign m87_34 =15'b0;

   // m87_35 = W*in
   wire signed [14:0] m87_35;
   assign m87_35 =15'b0;

   // m87_36 = W*in
   wire signed [14:0] m87_36;
   assign m87_36 =15'b0;

   // m87_37 = W*in
   wire signed [14:0] m87_37;
   assign m87_37 =15'b0;

   // m87_38 = W*in
   wire signed [14:0] m87_38;
   assign m87_38 =15'b0;

   // m87_39 = W*in
   wire signed [14:0] m87_39;
   assign m87_39 =15'b0;

   // m87_40 = W*in
   wire signed [14:0] m87_40;
   assign m87_40 =15'b0;

   // m87_41 = W*in
   wire signed [14:0] m87_41;
   assign m87_41 =15'b0;

   // m87_42 = W*in
   wire signed [14:0] m87_42;
   assign m87_42 =15'b0;

   // m87_43 = W*in
   wire signed [14:0] m87_43;
   assign m87_43 =15'b0;

   // m87_44 = W*in
   wire signed [14:0] m87_44;
   assign m87_44 =15'b0;

   // m87_45 = W*in
   wire signed [14:0] m87_45;
   assign m87_45 =15'b0;

   // m87_46 = W*in
   wire signed [14:0] m87_46;
   assign m87_46 =15'b0;

   // m87_47 = W*in
   wire signed [14:0] m87_47;
   assign m87_47 =15'b0;

   // m87_48 = W*in
   wire signed [14:0] m87_48;
   assign m87_48 =15'b0;

   // m87_49 = W*in
   wire signed [14:0] m87_49;
   assign m87_49 =15'b0;

   // m87_50 = W*in
   wire signed [14:0] m87_50;
   assign m87_50 =15'b0;

   // m87_51 = W*in
   wire signed [14:0] m87_51;
   assign m87_51 =15'b0;

   // m87_52 = W*in
   wire signed [14:0] m87_52;
   assign m87_52 ={ {3{neg87[14]}} , neg87[14:3] };

   // m87_53 = W*in
   wire signed [14:0] m87_53;
   assign m87_53 =15'b0;

   // m87_54 = W*in
   wire signed [14:0] m87_54;
   assign m87_54 =15'b0;

   // m87_55 = W*in
   wire signed [14:0] m87_55;
   assign m87_55 =15'b0;

   // m87_56 = W*in
   wire signed [14:0] m87_56;
   assign m87_56 =15'b0;

   // m87_57 = W*in
   wire signed [14:0] m87_57;
   assign m87_57 =15'b0;

   // m87_58 = W*in
   wire signed [14:0] m87_58;
   assign m87_58 ={ {4{neg87[14]}} , neg87[14:4] };

   // m87_59 = W*in
   wire signed [14:0] m87_59;
   assign m87_59 =15'b0;

   // m87_60 = W*in
   wire signed [14:0] m87_60;
   assign m87_60 =15'b0;

   // m87_61 = W*in
   wire signed [14:0] m87_61;
   assign m87_61 =15'b0;

   // m87_62 = W*in
   wire signed [14:0] m87_62;
   assign m87_62 =15'b0;

   // m87_63 = W*in
   wire signed [14:0] m87_63;
   assign m87_63 =15'b0;

   // m87_64 = W*in
   wire signed [14:0] m87_64;
   assign m87_64 =15'b0;

   // m87_65 = W*in
   wire signed [14:0] m87_65;
   assign m87_65 =15'b0;

   // m87_66 = W*in
   wire signed [14:0] m87_66;
   assign m87_66 =15'b0;

   // m87_67 = W*in
   wire signed [14:0] m87_67;
   assign m87_67 =15'b0;

   // m87_68 = W*in
   wire signed [14:0] m87_68;
   assign m87_68 =15'b0;

   // m87_69 = W*in
   wire signed [14:0] m87_69;
   assign m87_69 =15'b0;

   // m87_70 = W*in
   wire signed [14:0] m87_70;
   assign m87_70 ={ {4{in87[14]}} , in87[14:4] };

   // m87_71 = W*in
   wire signed [14:0] m87_71;
   assign m87_71 =15'b0;

   // m87_72 = W*in
   wire signed [14:0] m87_72;
   assign m87_72 =15'b0;

   // m87_73 = W*in
   wire signed [14:0] m87_73;
   assign m87_73 =15'b0;

   // m87_74 = W*in
   wire signed [14:0] m87_74;
   assign m87_74 ={ {4{in87[14]}} , in87[14:4] };

   // m87_75 = W*in
   wire signed [14:0] m87_75;
   assign m87_75 ={ {4{neg87[14]}} , neg87[14:4] };

   // m87_76 = W*in
   wire signed [14:0] m87_76;
   assign m87_76 =15'b0;

   // m87_77 = W*in
   wire signed [14:0] m87_77;
   assign m87_77 =15'b0;

   // m87_78 = W*in
   wire signed [14:0] m87_78;
   assign m87_78 =15'b0;

   // m87_79 = W*in
   wire signed [14:0] m87_79;
   assign m87_79 =15'b0;

   // m87_80 = W*in
   wire signed [14:0] m87_80;
   assign m87_80 =15'b0;

   // m87_81 = W*in
   wire signed [14:0] m87_81;
   assign m87_81 =15'b0;

   // m87_82 = W*in
   wire signed [14:0] m87_82;
   assign m87_82 =15'b0;

   // m87_83 = W*in
   wire signed [14:0] m87_83;
   assign m87_83 =15'b0;

   // m87_84 = W*in
   wire signed [14:0] m87_84;
   assign m87_84 =15'b0;

   // m87_85 = W*in
   wire signed [14:0] m87_85;
   assign m87_85 =15'b0;

   // m87_86 = W*in
   wire signed [14:0] m87_86;
   assign m87_86 =15'b0;

   // m87_87 = W*in
   wire signed [14:0] m87_87;
   assign m87_87 =15'b0;

   // m87_88 = W*in
   wire signed [14:0] m87_88;
   assign m87_88 =15'b0;

   // m87_89 = W*in
   wire signed [14:0] m87_89;
   assign m87_89 =15'b0;

   // m87_90 = W*in
   wire signed [14:0] m87_90;
   assign m87_90 =15'b0;

   // m87_91 = W*in
   wire signed [14:0] m87_91;
   assign m87_91 =15'b0;

   // m87_92 = W*in
   wire signed [14:0] m87_92;
   assign m87_92 =15'b0;

   // m87_93 = W*in
   wire signed [14:0] m87_93;
   assign m87_93 =15'b0;

   // m87_94 = W*in
   wire signed [14:0] m87_94;
   assign m87_94 =15'b0;

   // m87_95 = W*in
   wire signed [14:0] m87_95;
   assign m87_95 =15'b0;

   // m87_96 = W*in
   wire signed [14:0] m87_96;
   assign m87_96 =15'b0;

   // m87_97 = W*in
   wire signed [14:0] m87_97;
   assign m87_97 ={ {4{in87[14]}} , in87[14:4] };

   // m87_98 = W*in
   wire signed [14:0] m87_98;
   assign m87_98 =15'b0;

   // m87_99 = W*in
   wire signed [14:0] m87_99;
   assign m87_99 =15'b0;

   // m87_100 = W*in
   wire signed [14:0] m87_100;
   assign m87_100 =15'b0;

   // m88_1 = W*in
   wire signed [14:0] m88_1;
   assign m88_1 =15'b0;

   // m88_2 = W*in
   wire signed [14:0] m88_2;
   assign m88_2 =15'b0;

   // m88_3 = W*in
   wire signed [14:0] m88_3;
   assign m88_3 =15'b0;

   // m88_4 = W*in
   wire signed [14:0] m88_4;
   assign m88_4 =15'b0;

   // m88_5 = W*in
   wire signed [14:0] m88_5;
   assign m88_5 =15'b0;

   // m88_6 = W*in
   wire signed [14:0] m88_6;
   assign m88_6 =15'b0;

   // m88_7 = W*in
   wire signed [14:0] m88_7;
   assign m88_7 =15'b0;

   // m88_8 = W*in
   wire signed [14:0] m88_8;
   assign m88_8 ={ {3{in88[14]}} , in88[14:3] };

   // m88_9 = W*in
   wire signed [14:0] m88_9;
   assign m88_9 =15'b0;

   // m88_10 = W*in
   wire signed [14:0] m88_10;
   assign m88_10 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_11 = W*in
   wire signed [14:0] m88_11;
   assign m88_11 =15'b0;

   // m88_12 = W*in
   wire signed [14:0] m88_12;
   assign m88_12 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_13 = W*in
   wire signed [14:0] m88_13;
   assign m88_13 ={ {3{in88[14]}} , in88[14:3] };

   // m88_14 = W*in
   wire signed [14:0] m88_14;
   assign m88_14 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_15 = W*in
   wire signed [14:0] m88_15;
   assign m88_15 =15'b0;

   // m88_16 = W*in
   wire signed [14:0] m88_16;
   assign m88_16 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_17 = W*in
   wire signed [14:0] m88_17;
   assign m88_17 ={ {3{in88[14]}} , in88[14:3] };

   // m88_18 = W*in
   wire signed [14:0] m88_18;
   assign m88_18 =15'b0;

   // m88_19 = W*in
   wire signed [14:0] m88_19;
   assign m88_19 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_20 = W*in
   wire signed [14:0] m88_20;
   assign m88_20 =15'b0;

   // m88_21 = W*in
   wire signed [14:0] m88_21;
   assign m88_21 =15'b0;

   // m88_22 = W*in
   wire signed [14:0] m88_22;
   assign m88_22 =15'b0;

   // m88_23 = W*in
   wire signed [14:0] m88_23;
   assign m88_23 =15'b0;

   // m88_24 = W*in
   wire signed [14:0] m88_24;
   assign m88_24 =15'b0;

   // m88_25 = W*in
   wire signed [14:0] m88_25;
   assign m88_25 ={ {3{in88[14]}} , in88[14:3] };

   // m88_26 = W*in
   wire signed [14:0] m88_26;
   assign m88_26 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_27 = W*in
   wire signed [14:0] m88_27;
   assign m88_27 =15'b0;

   // m88_28 = W*in
   wire signed [14:0] m88_28;
   assign m88_28 =15'b0;

   // m88_29 = W*in
   wire signed [14:0] m88_29;
   assign m88_29 =15'b0;

   // m88_30 = W*in
   wire signed [14:0] m88_30;
   assign m88_30 =15'b0;

   // m88_31 = W*in
   wire signed [14:0] m88_31;
   assign m88_31 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_32 = W*in
   wire signed [14:0] m88_32;
   assign m88_32 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_33 = W*in
   wire signed [14:0] m88_33;
   assign m88_33 =15'b0;

   // m88_34 = W*in
   wire signed [14:0] m88_34;
   assign m88_34 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_35 = W*in
   wire signed [14:0] m88_35;
   assign m88_35 =15'b0;

   // m88_36 = W*in
   wire signed [14:0] m88_36;
   assign m88_36 =15'b0;

   // m88_37 = W*in
   wire signed [14:0] m88_37;
   assign m88_37 =15'b0;

   // m88_38 = W*in
   wire signed [14:0] m88_38;
   assign m88_38 ={ {4{in88[14]}} , in88[14:4] };

   // m88_39 = W*in
   wire signed [14:0] m88_39;
   assign m88_39 =15'b0;

   // m88_40 = W*in
   wire signed [14:0] m88_40;
   assign m88_40 =15'b0;

   // m88_41 = W*in
   wire signed [14:0] m88_41;
   assign m88_41 =15'b0;

   // m88_42 = W*in
   wire signed [14:0] m88_42;
   assign m88_42 =15'b0;

   // m88_43 = W*in
   wire signed [14:0] m88_43;
   assign m88_43 =15'b0;

   // m88_44 = W*in
   wire signed [14:0] m88_44;
   assign m88_44 =15'b0;

   // m88_45 = W*in
   wire signed [14:0] m88_45;
   assign m88_45 =15'b0;

   // m88_46 = W*in
   wire signed [14:0] m88_46;
   assign m88_46 =15'b0;

   // m88_47 = W*in
   wire signed [14:0] m88_47;
   assign m88_47 =15'b0;

   // m88_48 = W*in
   wire signed [14:0] m88_48;
   assign m88_48 =15'b0;

   // m88_49 = W*in
   wire signed [14:0] m88_49;
   assign m88_49 =15'b0;

   // m88_50 = W*in
   wire signed [14:0] m88_50;
   assign m88_50 =15'b0;

   // m88_51 = W*in
   wire signed [14:0] m88_51;
   assign m88_51 =15'b0;

   // m88_52 = W*in
   wire signed [14:0] m88_52;
   assign m88_52 ={ {3{in88[14]}} , in88[14:3] };

   // m88_53 = W*in
   wire signed [14:0] m88_53;
   assign m88_53 =15'b0;

   // m88_54 = W*in
   wire signed [14:0] m88_54;
   assign m88_54 =15'b0;

   // m88_55 = W*in
   wire signed [14:0] m88_55;
   assign m88_55 =15'b0;

   // m88_56 = W*in
   wire signed [14:0] m88_56;
   assign m88_56 =15'b0;

   // m88_57 = W*in
   wire signed [14:0] m88_57;
   assign m88_57 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_58 = W*in
   wire signed [14:0] m88_58;
   assign m88_58 =15'b0;

   // m88_59 = W*in
   wire signed [14:0] m88_59;
   assign m88_59 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_60 = W*in
   wire signed [14:0] m88_60;
   assign m88_60 =15'b0;

   // m88_61 = W*in
   wire signed [14:0] m88_61;
   assign m88_61 =15'b0;

   // m88_62 = W*in
   wire signed [14:0] m88_62;
   assign m88_62 =15'b0;

   // m88_63 = W*in
   wire signed [14:0] m88_63;
   assign m88_63 =15'b0;

   // m88_64 = W*in
   wire signed [14:0] m88_64;
   assign m88_64 =15'b0;

   // m88_65 = W*in
   wire signed [14:0] m88_65;
   assign m88_65 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_66 = W*in
   wire signed [14:0] m88_66;
   assign m88_66 =15'b0;

   // m88_67 = W*in
   wire signed [14:0] m88_67;
   assign m88_67 =15'b0;

   // m88_68 = W*in
   wire signed [14:0] m88_68;
   assign m88_68 =15'b0;

   // m88_69 = W*in
   wire signed [14:0] m88_69;
   assign m88_69 ={ {3{in88[14]}} , in88[14:3] };

   // m88_70 = W*in
   wire signed [14:0] m88_70;
   assign m88_70 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_71 = W*in
   wire signed [14:0] m88_71;
   assign m88_71 =15'b0;

   // m88_72 = W*in
   wire signed [14:0] m88_72;
   assign m88_72 ={ {3{in88[14]}} , in88[14:3] };

   // m88_73 = W*in
   wire signed [14:0] m88_73;
   assign m88_73 =15'b0;

   // m88_74 = W*in
   wire signed [14:0] m88_74;
   assign m88_74 =15'b0;

   // m88_75 = W*in
   wire signed [14:0] m88_75;
   assign m88_75 =15'b0;

   // m88_76 = W*in
   wire signed [14:0] m88_76;
   assign m88_76 =15'b0;

   // m88_77 = W*in
   wire signed [14:0] m88_77;
   assign m88_77 =15'b0;

   // m88_78 = W*in
   wire signed [14:0] m88_78;
   assign m88_78 ={ {3{in88[14]}} , in88[14:3] };

   // m88_79 = W*in
   wire signed [14:0] m88_79;
   assign m88_79 =15'b0;

   // m88_80 = W*in
   wire signed [14:0] m88_80;
   assign m88_80 =15'b0;

   // m88_81 = W*in
   wire signed [14:0] m88_81;
   assign m88_81 =15'b0;

   // m88_82 = W*in
   wire signed [14:0] m88_82;
   assign m88_82 =15'b0;

   // m88_83 = W*in
   wire signed [14:0] m88_83;
   assign m88_83 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_84 = W*in
   wire signed [14:0] m88_84;
   assign m88_84 =15'b0;

   // m88_85 = W*in
   wire signed [14:0] m88_85;
   assign m88_85 =15'b0;

   // m88_86 = W*in
   wire signed [14:0] m88_86;
   assign m88_86 =15'b0;

   // m88_87 = W*in
   wire signed [14:0] m88_87;
   assign m88_87 =15'b0;

   // m88_88 = W*in
   wire signed [14:0] m88_88;
   assign m88_88 =15'b0;

   // m88_89 = W*in
   wire signed [14:0] m88_89;
   assign m88_89 =15'b0;

   // m88_90 = W*in
   wire signed [14:0] m88_90;
   assign m88_90 =15'b0;

   // m88_91 = W*in
   wire signed [14:0] m88_91;
   assign m88_91 =15'b0;

   // m88_92 = W*in
   wire signed [14:0] m88_92;
   assign m88_92 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_93 = W*in
   wire signed [14:0] m88_93;
   assign m88_93 =15'b0;

   // m88_94 = W*in
   wire signed [14:0] m88_94;
   assign m88_94 ={ {3{neg88[14]}} , neg88[14:3] };

   // m88_95 = W*in
   wire signed [14:0] m88_95;
   assign m88_95 =15'b0;

   // m88_96 = W*in
   wire signed [14:0] m88_96;
   assign m88_96 ={ {3{in88[14]}} , in88[14:3] };

   // m88_97 = W*in
   wire signed [14:0] m88_97;
   assign m88_97 =15'b0;

   // m88_98 = W*in
   wire signed [14:0] m88_98;
   assign m88_98 =15'b0;

   // m88_99 = W*in
   wire signed [14:0] m88_99;
   assign m88_99 ={ {3{in88[14]}} , in88[14:3] };

   // m88_100 = W*in
   wire signed [14:0] m88_100;
   assign m88_100 ={ {3{neg88[14]}} , neg88[14:3] };

   // m89_1 = W*in
   wire signed [14:0] m89_1;
   assign m89_1 ={ {3{in89[14]}} , in89[14:3] };

   // m89_2 = W*in
   wire signed [14:0] m89_2;
   assign m89_2 ={ {3{in89[14]}} , in89[14:3] };

   // m89_3 = W*in
   wire signed [14:0] m89_3;
   assign m89_3 =15'b0;

   // m89_4 = W*in
   wire signed [14:0] m89_4;
   assign m89_4 =15'b0;

   // m89_5 = W*in
   wire signed [14:0] m89_5;
   assign m89_5 =15'b0;

   // m89_6 = W*in
   wire signed [14:0] m89_6;
   assign m89_6 =15'b0;

   // m89_7 = W*in
   wire signed [14:0] m89_7;
   assign m89_7 ={ {3{in89[14]}} , in89[14:3] };

   // m89_8 = W*in
   wire signed [14:0] m89_8;
   assign m89_8 =15'b0;

   // m89_9 = W*in
   wire signed [14:0] m89_9;
   assign m89_9 =15'b0;

   // m89_10 = W*in
   wire signed [14:0] m89_10;
   assign m89_10 =15'b0;

   // m89_11 = W*in
   wire signed [14:0] m89_11;
   assign m89_11 =15'b0;

   // m89_12 = W*in
   wire signed [14:0] m89_12;
   assign m89_12 =15'b0;

   // m89_13 = W*in
   wire signed [14:0] m89_13;
   assign m89_13 ={ {3{in89[14]}} , in89[14:3] };

   // m89_14 = W*in
   wire signed [14:0] m89_14;
   assign m89_14 =15'b0;

   // m89_15 = W*in
   wire signed [14:0] m89_15;
   assign m89_15 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_16 = W*in
   wire signed [14:0] m89_16;
   assign m89_16 =15'b0;

   // m89_17 = W*in
   wire signed [14:0] m89_17;
   assign m89_17 =15'b0;

   // m89_18 = W*in
   wire signed [14:0] m89_18;
   assign m89_18 =15'b0;

   // m89_19 = W*in
   wire signed [14:0] m89_19;
   assign m89_19 =15'b0;

   // m89_20 = W*in
   wire signed [14:0] m89_20;
   assign m89_20 =15'b0;

   // m89_21 = W*in
   wire signed [14:0] m89_21;
   assign m89_21 ={ {4{in89[14]}} , in89[14:4] };

   // m89_22 = W*in
   wire signed [14:0] m89_22;
   assign m89_22 =15'b0;

   // m89_23 = W*in
   wire signed [14:0] m89_23;
   assign m89_23 =15'b0;

   // m89_24 = W*in
   wire signed [14:0] m89_24;
   assign m89_24 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_25 = W*in
   wire signed [14:0] m89_25;
   assign m89_25 =15'b0;

   // m89_26 = W*in
   wire signed [14:0] m89_26;
   assign m89_26 =15'b0;

   // m89_27 = W*in
   wire signed [14:0] m89_27;
   assign m89_27 ={ {3{in89[14]}} , in89[14:3] };

   // m89_28 = W*in
   wire signed [14:0] m89_28;
   assign m89_28 ={ {4{neg89[14]}} , neg89[14:4] };

   // m89_29 = W*in
   wire signed [14:0] m89_29;
   assign m89_29 ={ {3{in89[14]}} , in89[14:3] };

   // m89_30 = W*in
   wire signed [14:0] m89_30;
   assign m89_30 =15'b0;

   // m89_31 = W*in
   wire signed [14:0] m89_31;
   assign m89_31 =15'b0;

   // m89_32 = W*in
   wire signed [14:0] m89_32;
   assign m89_32 ={ {3{in89[14]}} , in89[14:3] };

   // m89_33 = W*in
   wire signed [14:0] m89_33;
   assign m89_33 ={ {3{in89[14]}} , in89[14:3] };

   // m89_34 = W*in
   wire signed [14:0] m89_34;
   assign m89_34 =15'b0;

   // m89_35 = W*in
   wire signed [14:0] m89_35;
   assign m89_35 =15'b0;

   // m89_36 = W*in
   wire signed [14:0] m89_36;
   assign m89_36 =15'b0;

   // m89_37 = W*in
   wire signed [14:0] m89_37;
   assign m89_37 ={ {2{neg89[14]}} , neg89[14:2] };

   // m89_38 = W*in
   wire signed [14:0] m89_38;
   assign m89_38 ={ {3{in89[14]}} , in89[14:3] };

   // m89_39 = W*in
   wire signed [14:0] m89_39;
   assign m89_39 =15'b0;

   // m89_40 = W*in
   wire signed [14:0] m89_40;
   assign m89_40 =15'b0;

   // m89_41 = W*in
   wire signed [14:0] m89_41;
   assign m89_41 ={ {4{neg89[14]}} , neg89[14:4] };

   // m89_42 = W*in
   wire signed [14:0] m89_42;
   assign m89_42 =15'b0;

   // m89_43 = W*in
   wire signed [14:0] m89_43;
   assign m89_43 ={ {3{in89[14]}} , in89[14:3] };

   // m89_44 = W*in
   wire signed [14:0] m89_44;
   assign m89_44 =15'b0;

   // m89_45 = W*in
   wire signed [14:0] m89_45;
   assign m89_45 =15'b0;

   // m89_46 = W*in
   wire signed [14:0] m89_46;
   assign m89_46 =15'b0;

   // m89_47 = W*in
   wire signed [14:0] m89_47;
   assign m89_47 =15'b0;

   // m89_48 = W*in
   wire signed [14:0] m89_48;
   assign m89_48 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_49 = W*in
   wire signed [14:0] m89_49;
   assign m89_49 =15'b0;

   // m89_50 = W*in
   wire signed [14:0] m89_50;
   assign m89_50 =15'b0;

   // m89_51 = W*in
   wire signed [14:0] m89_51;
   assign m89_51 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_52 = W*in
   wire signed [14:0] m89_52;
   assign m89_52 =15'b0;

   // m89_53 = W*in
   wire signed [14:0] m89_53;
   assign m89_53 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_54 = W*in
   wire signed [14:0] m89_54;
   assign m89_54 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_55 = W*in
   wire signed [14:0] m89_55;
   assign m89_55 =15'b0;

   // m89_56 = W*in
   wire signed [14:0] m89_56;
   assign m89_56 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_57 = W*in
   wire signed [14:0] m89_57;
   assign m89_57 =15'b0;

   // m89_58 = W*in
   wire signed [14:0] m89_58;
   assign m89_58 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_59 = W*in
   wire signed [14:0] m89_59;
   assign m89_59 =15'b0;

   // m89_60 = W*in
   wire signed [14:0] m89_60;
   assign m89_60 ={ {4{neg89[14]}} , neg89[14:4] };

   // m89_61 = W*in
   wire signed [14:0] m89_61;
   assign m89_61 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_62 = W*in
   wire signed [14:0] m89_62;
   assign m89_62 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_63 = W*in
   wire signed [14:0] m89_63;
   assign m89_63 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_64 = W*in
   wire signed [14:0] m89_64;
   assign m89_64 ={ {4{neg89[14]}} , neg89[14:4] };

   // m89_65 = W*in
   wire signed [14:0] m89_65;
   assign m89_65 =15'b0;

   // m89_66 = W*in
   wire signed [14:0] m89_66;
   assign m89_66 =15'b0;

   // m89_67 = W*in
   wire signed [14:0] m89_67;
   assign m89_67 =15'b0;

   // m89_68 = W*in
   wire signed [14:0] m89_68;
   assign m89_68 =15'b0;

   // m89_69 = W*in
   wire signed [14:0] m89_69;
   assign m89_69 =15'b0;

   // m89_70 = W*in
   wire signed [14:0] m89_70;
   assign m89_70 =15'b0;

   // m89_71 = W*in
   wire signed [14:0] m89_71;
   assign m89_71 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_72 = W*in
   wire signed [14:0] m89_72;
   assign m89_72 =15'b0;

   // m89_73 = W*in
   wire signed [14:0] m89_73;
   assign m89_73 =15'b0;

   // m89_74 = W*in
   wire signed [14:0] m89_74;
   assign m89_74 =15'b0;

   // m89_75 = W*in
   wire signed [14:0] m89_75;
   assign m89_75 =15'b0;

   // m89_76 = W*in
   wire signed [14:0] m89_76;
   assign m89_76 =15'b0;

   // m89_77 = W*in
   wire signed [14:0] m89_77;
   assign m89_77 ={ {4{neg89[14]}} , neg89[14:4] };

   // m89_78 = W*in
   wire signed [14:0] m89_78;
   assign m89_78 =15'b0;

   // m89_79 = W*in
   wire signed [14:0] m89_79;
   assign m89_79 =15'b0;

   // m89_80 = W*in
   wire signed [14:0] m89_80;
   assign m89_80 =15'b0;

   // m89_81 = W*in
   wire signed [14:0] m89_81;
   assign m89_81 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_82 = W*in
   wire signed [14:0] m89_82;
   assign m89_82 =15'b0;

   // m89_83 = W*in
   wire signed [14:0] m89_83;
   assign m89_83 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_84 = W*in
   wire signed [14:0] m89_84;
   assign m89_84 ={ {3{in89[14]}} , in89[14:3] };

   // m89_85 = W*in
   wire signed [14:0] m89_85;
   assign m89_85 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_86 = W*in
   wire signed [14:0] m89_86;
   assign m89_86 =15'b0;

   // m89_87 = W*in
   wire signed [14:0] m89_87;
   assign m89_87 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_88 = W*in
   wire signed [14:0] m89_88;
   assign m89_88 =15'b0;

   // m89_89 = W*in
   wire signed [14:0] m89_89;
   assign m89_89 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_90 = W*in
   wire signed [14:0] m89_90;
   assign m89_90 ={ {2{in89[14]}} , in89[14:2] };

   // m89_91 = W*in
   wire signed [14:0] m89_91;
   assign m89_91 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_92 = W*in
   wire signed [14:0] m89_92;
   assign m89_92 =15'b0;

   // m89_93 = W*in
   wire signed [14:0] m89_93;
   assign m89_93 ={ {3{neg89[14]}} , neg89[14:3] };

   // m89_94 = W*in
   wire signed [14:0] m89_94;
   assign m89_94 ={ {3{in89[14]}} , in89[14:3] };

   // m89_95 = W*in
   wire signed [14:0] m89_95;
   assign m89_95 ={ {3{in89[14]}} , in89[14:3] };

   // m89_96 = W*in
   wire signed [14:0] m89_96;
   assign m89_96 ={ {4{neg89[14]}} , neg89[14:4] };

   // m89_97 = W*in
   wire signed [14:0] m89_97;
   assign m89_97 ={ {3{in89[14]}} , in89[14:3] };

   // m89_98 = W*in
   wire signed [14:0] m89_98;
   assign m89_98 =15'b0;

   // m89_99 = W*in
   wire signed [14:0] m89_99;
   assign m89_99 =15'b0;

   // m89_100 = W*in
   wire signed [14:0] m89_100;
   assign m89_100 ={ {3{neg89[14]}} , neg89[14:3] };

   // m90_1 = W*in
   wire signed [14:0] m90_1;
   assign m90_1 ={ {4{neg90[14]}} , neg90[14:4] };

   // m90_2 = W*in
   wire signed [14:0] m90_2;
   assign m90_2 =15'b0;

   // m90_3 = W*in
   wire signed [14:0] m90_3;
   assign m90_3 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_4 = W*in
   wire signed [14:0] m90_4;
   assign m90_4 =15'b0;

   // m90_5 = W*in
   wire signed [14:0] m90_5;
   assign m90_5 =15'b0;

   // m90_6 = W*in
   wire signed [14:0] m90_6;
   assign m90_6 =15'b0;

   // m90_7 = W*in
   wire signed [14:0] m90_7;
   assign m90_7 =15'b0;

   // m90_8 = W*in
   wire signed [14:0] m90_8;
   assign m90_8 =15'b0;

   // m90_9 = W*in
   wire signed [14:0] m90_9;
   assign m90_9 =15'b0;

   // m90_10 = W*in
   wire signed [14:0] m90_10;
   assign m90_10 =15'b0;

   // m90_11 = W*in
   wire signed [14:0] m90_11;
   assign m90_11 =15'b0;

   // m90_12 = W*in
   wire signed [14:0] m90_12;
   assign m90_12 =15'b0;

   // m90_13 = W*in
   wire signed [14:0] m90_13;
   assign m90_13 =15'b0;

   // m90_14 = W*in
   wire signed [14:0] m90_14;
   assign m90_14 =15'b0;

   // m90_15 = W*in
   wire signed [14:0] m90_15;
   assign m90_15 =15'b0;

   // m90_16 = W*in
   wire signed [14:0] m90_16;
   assign m90_16 =15'b0;

   // m90_17 = W*in
   wire signed [14:0] m90_17;
   assign m90_17 =15'b0;

   // m90_18 = W*in
   wire signed [14:0] m90_18;
   assign m90_18 ={ {3{in90[14]}} , in90[14:3] };

   // m90_19 = W*in
   wire signed [14:0] m90_19;
   assign m90_19 =15'b0;

   // m90_20 = W*in
   wire signed [14:0] m90_20;
   assign m90_20 =15'b0;

   // m90_21 = W*in
   wire signed [14:0] m90_21;
   assign m90_21 =15'b0;

   // m90_22 = W*in
   wire signed [14:0] m90_22;
   assign m90_22 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_23 = W*in
   wire signed [14:0] m90_23;
   assign m90_23 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_24 = W*in
   wire signed [14:0] m90_24;
   assign m90_24 =15'b0;

   // m90_25 = W*in
   wire signed [14:0] m90_25;
   assign m90_25 =15'b0;

   // m90_26 = W*in
   wire signed [14:0] m90_26;
   assign m90_26 =15'b0;

   // m90_27 = W*in
   wire signed [14:0] m90_27;
   assign m90_27 ={ {4{neg90[14]}} , neg90[14:4] };

   // m90_28 = W*in
   wire signed [14:0] m90_28;
   assign m90_28 ={ {3{in90[14]}} , in90[14:3] };

   // m90_29 = W*in
   wire signed [14:0] m90_29;
   assign m90_29 =15'b0;

   // m90_30 = W*in
   wire signed [14:0] m90_30;
   assign m90_30 =15'b0;

   // m90_31 = W*in
   wire signed [14:0] m90_31;
   assign m90_31 ={ {3{in90[14]}} , in90[14:3] };

   // m90_32 = W*in
   wire signed [14:0] m90_32;
   assign m90_32 =15'b0;

   // m90_33 = W*in
   wire signed [14:0] m90_33;
   assign m90_33 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_34 = W*in
   wire signed [14:0] m90_34;
   assign m90_34 =15'b0;

   // m90_35 = W*in
   wire signed [14:0] m90_35;
   assign m90_35 =15'b0;

   // m90_36 = W*in
   wire signed [14:0] m90_36;
   assign m90_36 =15'b0;

   // m90_37 = W*in
   wire signed [14:0] m90_37;
   assign m90_37 =15'b0;

   // m90_38 = W*in
   wire signed [14:0] m90_38;
   assign m90_38 =15'b0;

   // m90_39 = W*in
   wire signed [14:0] m90_39;
   assign m90_39 =15'b0;

   // m90_40 = W*in
   wire signed [14:0] m90_40;
   assign m90_40 =15'b0;

   // m90_41 = W*in
   wire signed [14:0] m90_41;
   assign m90_41 ={ {3{in90[14]}} , in90[14:3] };

   // m90_42 = W*in
   wire signed [14:0] m90_42;
   assign m90_42 =15'b0;

   // m90_43 = W*in
   wire signed [14:0] m90_43;
   assign m90_43 =15'b0;

   // m90_44 = W*in
   wire signed [14:0] m90_44;
   assign m90_44 =15'b0;

   // m90_45 = W*in
   wire signed [14:0] m90_45;
   assign m90_45 =15'b0;

   // m90_46 = W*in
   wire signed [14:0] m90_46;
   assign m90_46 =15'b0;

   // m90_47 = W*in
   wire signed [14:0] m90_47;
   assign m90_47 =15'b0;

   // m90_48 = W*in
   wire signed [14:0] m90_48;
   assign m90_48 =15'b0;

   // m90_49 = W*in
   wire signed [14:0] m90_49;
   assign m90_49 =15'b0;

   // m90_50 = W*in
   wire signed [14:0] m90_50;
   assign m90_50 =15'b0;

   // m90_51 = W*in
   wire signed [14:0] m90_51;
   assign m90_51 =15'b0;

   // m90_52 = W*in
   wire signed [14:0] m90_52;
   assign m90_52 =15'b0;

   // m90_53 = W*in
   wire signed [14:0] m90_53;
   assign m90_53 =15'b0;

   // m90_54 = W*in
   wire signed [14:0] m90_54;
   assign m90_54 =15'b0;

   // m90_55 = W*in
   wire signed [14:0] m90_55;
   assign m90_55 =15'b0;

   // m90_56 = W*in
   wire signed [14:0] m90_56;
   assign m90_56 =15'b0;

   // m90_57 = W*in
   wire signed [14:0] m90_57;
   assign m90_57 =15'b0;

   // m90_58 = W*in
   wire signed [14:0] m90_58;
   assign m90_58 =15'b0;

   // m90_59 = W*in
   wire signed [14:0] m90_59;
   assign m90_59 =15'b0;

   // m90_60 = W*in
   wire signed [14:0] m90_60;
   assign m90_60 =15'b0;

   // m90_61 = W*in
   wire signed [14:0] m90_61;
   assign m90_61 =15'b0;

   // m90_62 = W*in
   wire signed [14:0] m90_62;
   assign m90_62 =15'b0;

   // m90_63 = W*in
   wire signed [14:0] m90_63;
   assign m90_63 =15'b0;

   // m90_64 = W*in
   wire signed [14:0] m90_64;
   assign m90_64 =15'b0;

   // m90_65 = W*in
   wire signed [14:0] m90_65;
   assign m90_65 =15'b0;

   // m90_66 = W*in
   wire signed [14:0] m90_66;
   assign m90_66 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_67 = W*in
   wire signed [14:0] m90_67;
   assign m90_67 =15'b0;

   // m90_68 = W*in
   wire signed [14:0] m90_68;
   assign m90_68 =15'b0;

   // m90_69 = W*in
   wire signed [14:0] m90_69;
   assign m90_69 =15'b0;

   // m90_70 = W*in
   wire signed [14:0] m90_70;
   assign m90_70 =15'b0;

   // m90_71 = W*in
   wire signed [14:0] m90_71;
   assign m90_71 =15'b0;

   // m90_72 = W*in
   wire signed [14:0] m90_72;
   assign m90_72 =15'b0;

   // m90_73 = W*in
   wire signed [14:0] m90_73;
   assign m90_73 =15'b0;

   // m90_74 = W*in
   wire signed [14:0] m90_74;
   assign m90_74 =15'b0;

   // m90_75 = W*in
   wire signed [14:0] m90_75;
   assign m90_75 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_76 = W*in
   wire signed [14:0] m90_76;
   assign m90_76 =15'b0;

   // m90_77 = W*in
   wire signed [14:0] m90_77;
   assign m90_77 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_78 = W*in
   wire signed [14:0] m90_78;
   assign m90_78 ={ {2{in90[14]}} , in90[14:2] };

   // m90_79 = W*in
   wire signed [14:0] m90_79;
   assign m90_79 =15'b0;

   // m90_80 = W*in
   wire signed [14:0] m90_80;
   assign m90_80 =15'b0;

   // m90_81 = W*in
   wire signed [14:0] m90_81;
   assign m90_81 =15'b0;

   // m90_82 = W*in
   wire signed [14:0] m90_82;
   assign m90_82 =15'b0;

   // m90_83 = W*in
   wire signed [14:0] m90_83;
   assign m90_83 =15'b0;

   // m90_84 = W*in
   wire signed [14:0] m90_84;
   assign m90_84 =15'b0;

   // m90_85 = W*in
   wire signed [14:0] m90_85;
   assign m90_85 =15'b0;

   // m90_86 = W*in
   wire signed [14:0] m90_86;
   assign m90_86 =15'b0;

   // m90_87 = W*in
   wire signed [14:0] m90_87;
   assign m90_87 =15'b0;

   // m90_88 = W*in
   wire signed [14:0] m90_88;
   assign m90_88 =15'b0;

   // m90_89 = W*in
   wire signed [14:0] m90_89;
   assign m90_89 ={ {3{in90[14]}} , in90[14:3] };

   // m90_90 = W*in
   wire signed [14:0] m90_90;
   assign m90_90 =15'b0;

   // m90_91 = W*in
   wire signed [14:0] m90_91;
   assign m90_91 =15'b0;

   // m90_92 = W*in
   wire signed [14:0] m90_92;
   assign m90_92 =15'b0;

   // m90_93 = W*in
   wire signed [14:0] m90_93;
   assign m90_93 ={ {3{neg90[14]}} , neg90[14:3] };

   // m90_94 = W*in
   wire signed [14:0] m90_94;
   assign m90_94 =15'b0;

   // m90_95 = W*in
   wire signed [14:0] m90_95;
   assign m90_95 =15'b0;

   // m90_96 = W*in
   wire signed [14:0] m90_96;
   assign m90_96 =15'b0;

   // m90_97 = W*in
   wire signed [14:0] m90_97;
   assign m90_97 =15'b0;

   // m90_98 = W*in
   wire signed [14:0] m90_98;
   assign m90_98 =15'b0;

   // m90_99 = W*in
   wire signed [14:0] m90_99;
   assign m90_99 =15'b0;

   // m90_100 = W*in
   wire signed [14:0] m90_100;
   assign m90_100 =15'b0;

   // m91_1 = W*in
   wire signed [14:0] m91_1;
   assign m91_1 =15'b0;

   // m91_2 = W*in
   wire signed [14:0] m91_2;
   assign m91_2 =15'b0;

   // m91_3 = W*in
   wire signed [14:0] m91_3;
   assign m91_3 =15'b0;

   // m91_4 = W*in
   wire signed [14:0] m91_4;
   assign m91_4 ={ {3{in91[14]}} , in91[14:3] };

   // m91_5 = W*in
   wire signed [14:0] m91_5;
   assign m91_5 =15'b0;

   // m91_6 = W*in
   wire signed [14:0] m91_6;
   assign m91_6 =15'b0;

   // m91_7 = W*in
   wire signed [14:0] m91_7;
   assign m91_7 =15'b0;

   // m91_8 = W*in
   wire signed [14:0] m91_8;
   assign m91_8 =15'b0;

   // m91_9 = W*in
   wire signed [14:0] m91_9;
   assign m91_9 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_10 = W*in
   wire signed [14:0] m91_10;
   assign m91_10 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_11 = W*in
   wire signed [14:0] m91_11;
   assign m91_11 =15'b0;

   // m91_12 = W*in
   wire signed [14:0] m91_12;
   assign m91_12 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_13 = W*in
   wire signed [14:0] m91_13;
   assign m91_13 =15'b0;

   // m91_14 = W*in
   wire signed [14:0] m91_14;
   assign m91_14 =15'b0;

   // m91_15 = W*in
   wire signed [14:0] m91_15;
   assign m91_15 =15'b0;

   // m91_16 = W*in
   wire signed [14:0] m91_16;
   assign m91_16 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_17 = W*in
   wire signed [14:0] m91_17;
   assign m91_17 ={ {3{in91[14]}} , in91[14:3] };

   // m91_18 = W*in
   wire signed [14:0] m91_18;
   assign m91_18 ={ {3{in91[14]}} , in91[14:3] };

   // m91_19 = W*in
   wire signed [14:0] m91_19;
   assign m91_19 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_20 = W*in
   wire signed [14:0] m91_20;
   assign m91_20 =15'b0;

   // m91_21 = W*in
   wire signed [14:0] m91_21;
   assign m91_21 =15'b0;

   // m91_22 = W*in
   wire signed [14:0] m91_22;
   assign m91_22 =15'b0;

   // m91_23 = W*in
   wire signed [14:0] m91_23;
   assign m91_23 =15'b0;

   // m91_24 = W*in
   wire signed [14:0] m91_24;
   assign m91_24 =15'b0;

   // m91_25 = W*in
   wire signed [14:0] m91_25;
   assign m91_25 =15'b0;

   // m91_26 = W*in
   wire signed [14:0] m91_26;
   assign m91_26 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_27 = W*in
   wire signed [14:0] m91_27;
   assign m91_27 ={ {3{in91[14]}} , in91[14:3] };

   // m91_28 = W*in
   wire signed [14:0] m91_28;
   assign m91_28 ={ {4{in91[14]}} , in91[14:4] };

   // m91_29 = W*in
   wire signed [14:0] m91_29;
   assign m91_29 ={ {4{neg91[14]}} , neg91[14:4] };

   // m91_30 = W*in
   wire signed [14:0] m91_30;
   assign m91_30 =15'b0;

   // m91_31 = W*in
   wire signed [14:0] m91_31;
   assign m91_31 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_32 = W*in
   wire signed [14:0] m91_32;
   assign m91_32 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_33 = W*in
   wire signed [14:0] m91_33;
   assign m91_33 =15'b0;

   // m91_34 = W*in
   wire signed [14:0] m91_34;
   assign m91_34 =15'b0;

   // m91_35 = W*in
   wire signed [14:0] m91_35;
   assign m91_35 =15'b0;

   // m91_36 = W*in
   wire signed [14:0] m91_36;
   assign m91_36 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_37 = W*in
   wire signed [14:0] m91_37;
   assign m91_37 =15'b0;

   // m91_38 = W*in
   wire signed [14:0] m91_38;
   assign m91_38 ={ {3{in91[14]}} , in91[14:3] };

   // m91_39 = W*in
   wire signed [14:0] m91_39;
   assign m91_39 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_40 = W*in
   wire signed [14:0] m91_40;
   assign m91_40 =15'b0;

   // m91_41 = W*in
   wire signed [14:0] m91_41;
   assign m91_41 =15'b0;

   // m91_42 = W*in
   wire signed [14:0] m91_42;
   assign m91_42 =15'b0;

   // m91_43 = W*in
   wire signed [14:0] m91_43;
   assign m91_43 =15'b0;

   // m91_44 = W*in
   wire signed [14:0] m91_44;
   assign m91_44 =15'b0;

   // m91_45 = W*in
   wire signed [14:0] m91_45;
   assign m91_45 =15'b0;

   // m91_46 = W*in
   wire signed [14:0] m91_46;
   assign m91_46 =15'b0;

   // m91_47 = W*in
   wire signed [14:0] m91_47;
   assign m91_47 =15'b0;

   // m91_48 = W*in
   wire signed [14:0] m91_48;
   assign m91_48 =15'b0;

   // m91_49 = W*in
   wire signed [14:0] m91_49;
   assign m91_49 =15'b0;

   // m91_50 = W*in
   wire signed [14:0] m91_50;
   assign m91_50 ={ {3{in91[14]}} , in91[14:3] };

   // m91_51 = W*in
   wire signed [14:0] m91_51;
   assign m91_51 =15'b0;

   // m91_52 = W*in
   wire signed [14:0] m91_52;
   assign m91_52 =15'b0;

   // m91_53 = W*in
   wire signed [14:0] m91_53;
   assign m91_53 =15'b0;

   // m91_54 = W*in
   wire signed [14:0] m91_54;
   assign m91_54 =15'b0;

   // m91_55 = W*in
   wire signed [14:0] m91_55;
   assign m91_55 =15'b0;

   // m91_56 = W*in
   wire signed [14:0] m91_56;
   assign m91_56 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_57 = W*in
   wire signed [14:0] m91_57;
   assign m91_57 ={ {3{neg91[14]}} , neg91[14:3] };

   // m91_58 = W*in
   wire signed [14:0] m91_58;
   assign m91_58 =15'b0;

   // m91_59 = W*in
   wire signed [14:0] m91_59;
   assign m91_59 =15'b0;

   // m91_60 = W*in
   wire signed [14:0] m91_60;
   assign m91_60 =15'b0;

   // m91_61 = W*in
   wire signed [14:0] m91_61;
   assign m91_61 =15'b0;

   // m91_62 = W*in
   wire signed [14:0] m91_62;
   assign m91_62 =15'b0;

   // m91_63 = W*in
   wire signed [14:0] m91_63;
   assign m91_63 =15'b0;

   // m91_64 = W*in
   wire signed [14:0] m91_64;
   assign m91_64 =15'b0;

   // m91_65 = W*in
   wire signed [14:0] m91_65;
   assign m91_65 =15'b0;

   // m91_66 = W*in
   wire signed [14:0] m91_66;
   assign m91_66 =15'b0;

   // m91_67 = W*in
   wire signed [14:0] m91_67;
   assign m91_67 =15'b0;

   // m91_68 = W*in
   wire signed [14:0] m91_68;
   assign m91_68 =15'b0;

   // m91_69 = W*in
   wire signed [14:0] m91_69;
   assign m91_69 ={ {4{neg91[14]}} , neg91[14:4] };

   // m91_70 = W*in
   wire signed [14:0] m91_70;
   assign m91_70 =15'b0;

   // m91_71 = W*in
   wire signed [14:0] m91_71;
   assign m91_71 =15'b0;

   // m91_72 = W*in
   wire signed [14:0] m91_72;
   assign m91_72 =15'b0;

   // m91_73 = W*in
   wire signed [14:0] m91_73;
   assign m91_73 =15'b0;

   // m91_74 = W*in
   wire signed [14:0] m91_74;
   assign m91_74 =15'b0;

   // m91_75 = W*in
   wire signed [14:0] m91_75;
   assign m91_75 =15'b0;

   // m91_76 = W*in
   wire signed [14:0] m91_76;
   assign m91_76 =15'b0;

   // m91_77 = W*in
   wire signed [14:0] m91_77;
   assign m91_77 =15'b0;

   // m91_78 = W*in
   wire signed [14:0] m91_78;
   assign m91_78 =15'b0;

   // m91_79 = W*in
   wire signed [14:0] m91_79;
   assign m91_79 =15'b0;

   // m91_80 = W*in
   wire signed [14:0] m91_80;
   assign m91_80 =15'b0;

   // m91_81 = W*in
   wire signed [14:0] m91_81;
   assign m91_81 =15'b0;

   // m91_82 = W*in
   wire signed [14:0] m91_82;
   assign m91_82 =15'b0;

   // m91_83 = W*in
   wire signed [14:0] m91_83;
   assign m91_83 =15'b0;

   // m91_84 = W*in
   wire signed [14:0] m91_84;
   assign m91_84 ={ {3{in91[14]}} , in91[14:3] };

   // m91_85 = W*in
   wire signed [14:0] m91_85;
   assign m91_85 =15'b0;

   // m91_86 = W*in
   wire signed [14:0] m91_86;
   assign m91_86 =15'b0;

   // m91_87 = W*in
   wire signed [14:0] m91_87;
   assign m91_87 =15'b0;

   // m91_88 = W*in
   wire signed [14:0] m91_88;
   assign m91_88 =15'b0;

   // m91_89 = W*in
   wire signed [14:0] m91_89;
   assign m91_89 =15'b0;

   // m91_90 = W*in
   wire signed [14:0] m91_90;
   assign m91_90 =15'b0;

   // m91_91 = W*in
   wire signed [14:0] m91_91;
   assign m91_91 =15'b0;

   // m91_92 = W*in
   wire signed [14:0] m91_92;
   assign m91_92 =15'b0;

   // m91_93 = W*in
   wire signed [14:0] m91_93;
   assign m91_93 =15'b0;

   // m91_94 = W*in
   wire signed [14:0] m91_94;
   assign m91_94 =15'b0;

   // m91_95 = W*in
   wire signed [14:0] m91_95;
   assign m91_95 =15'b0;

   // m91_96 = W*in
   wire signed [14:0] m91_96;
   assign m91_96 =15'b0;

   // m91_97 = W*in
   wire signed [14:0] m91_97;
   assign m91_97 =15'b0;

   // m91_98 = W*in
   wire signed [14:0] m91_98;
   assign m91_98 =15'b0;

   // m91_99 = W*in
   wire signed [14:0] m91_99;
   assign m91_99 =15'b0;

   // m91_100 = W*in
   wire signed [14:0] m91_100;
   assign m91_100 =15'b0;

   // m92_1 = W*in
   wire signed [14:0] m92_1;
   assign m92_1 =15'b0;

   // m92_2 = W*in
   wire signed [14:0] m92_2;
   assign m92_2 =15'b0;

   // m92_3 = W*in
   wire signed [14:0] m92_3;
   assign m92_3 =15'b0;

   // m92_4 = W*in
   wire signed [14:0] m92_4;
   assign m92_4 =15'b0;

   // m92_5 = W*in
   wire signed [14:0] m92_5;
   assign m92_5 =15'b0;

   // m92_6 = W*in
   wire signed [14:0] m92_6;
   assign m92_6 =15'b0;

   // m92_7 = W*in
   wire signed [14:0] m92_7;
   assign m92_7 =15'b0;

   // m92_8 = W*in
   wire signed [14:0] m92_8;
   assign m92_8 =15'b0;

   // m92_9 = W*in
   wire signed [14:0] m92_9;
   assign m92_9 =15'b0;

   // m92_10 = W*in
   wire signed [14:0] m92_10;
   assign m92_10 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_11 = W*in
   wire signed [14:0] m92_11;
   assign m92_11 =15'b0;

   // m92_12 = W*in
   wire signed [14:0] m92_12;
   assign m92_12 =15'b0;

   // m92_13 = W*in
   wire signed [14:0] m92_13;
   assign m92_13 =15'b0;

   // m92_14 = W*in
   wire signed [14:0] m92_14;
   assign m92_14 =15'b0;

   // m92_15 = W*in
   wire signed [14:0] m92_15;
   assign m92_15 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_16 = W*in
   wire signed [14:0] m92_16;
   assign m92_16 =15'b0;

   // m92_17 = W*in
   wire signed [14:0] m92_17;
   assign m92_17 ={ {3{in92[14]}} , in92[14:3] };

   // m92_18 = W*in
   wire signed [14:0] m92_18;
   assign m92_18 =15'b0;

   // m92_19 = W*in
   wire signed [14:0] m92_19;
   assign m92_19 =15'b0;

   // m92_20 = W*in
   wire signed [14:0] m92_20;
   assign m92_20 =15'b0;

   // m92_21 = W*in
   wire signed [14:0] m92_21;
   assign m92_21 =15'b0;

   // m92_22 = W*in
   wire signed [14:0] m92_22;
   assign m92_22 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_23 = W*in
   wire signed [14:0] m92_23;
   assign m92_23 =15'b0;

   // m92_24 = W*in
   wire signed [14:0] m92_24;
   assign m92_24 =15'b0;

   // m92_25 = W*in
   wire signed [14:0] m92_25;
   assign m92_25 =15'b0;

   // m92_26 = W*in
   wire signed [14:0] m92_26;
   assign m92_26 =15'b0;

   // m92_27 = W*in
   wire signed [14:0] m92_27;
   assign m92_27 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_28 = W*in
   wire signed [14:0] m92_28;
   assign m92_28 =15'b0;

   // m92_29 = W*in
   wire signed [14:0] m92_29;
   assign m92_29 ={ {4{neg92[14]}} , neg92[14:4] };

   // m92_30 = W*in
   wire signed [14:0] m92_30;
   assign m92_30 =15'b0;

   // m92_31 = W*in
   wire signed [14:0] m92_31;
   assign m92_31 =15'b0;

   // m92_32 = W*in
   wire signed [14:0] m92_32;
   assign m92_32 =15'b0;

   // m92_33 = W*in
   wire signed [14:0] m92_33;
   assign m92_33 =15'b0;

   // m92_34 = W*in
   wire signed [14:0] m92_34;
   assign m92_34 =15'b0;

   // m92_35 = W*in
   wire signed [14:0] m92_35;
   assign m92_35 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_36 = W*in
   wire signed [14:0] m92_36;
   assign m92_36 =15'b0;

   // m92_37 = W*in
   wire signed [14:0] m92_37;
   assign m92_37 =15'b0;

   // m92_38 = W*in
   wire signed [14:0] m92_38;
   assign m92_38 =15'b0;

   // m92_39 = W*in
   wire signed [14:0] m92_39;
   assign m92_39 =15'b0;

   // m92_40 = W*in
   wire signed [14:0] m92_40;
   assign m92_40 =15'b0;

   // m92_41 = W*in
   wire signed [14:0] m92_41;
   assign m92_41 =15'b0;

   // m92_42 = W*in
   wire signed [14:0] m92_42;
   assign m92_42 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_43 = W*in
   wire signed [14:0] m92_43;
   assign m92_43 =15'b0;

   // m92_44 = W*in
   wire signed [14:0] m92_44;
   assign m92_44 =15'b0;

   // m92_45 = W*in
   wire signed [14:0] m92_45;
   assign m92_45 =15'b0;

   // m92_46 = W*in
   wire signed [14:0] m92_46;
   assign m92_46 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_47 = W*in
   wire signed [14:0] m92_47;
   assign m92_47 ={ {3{in92[14]}} , in92[14:3] };

   // m92_48 = W*in
   wire signed [14:0] m92_48;
   assign m92_48 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_49 = W*in
   wire signed [14:0] m92_49;
   assign m92_49 =15'b0;

   // m92_50 = W*in
   wire signed [14:0] m92_50;
   assign m92_50 =15'b0;

   // m92_51 = W*in
   wire signed [14:0] m92_51;
   assign m92_51 =15'b0;

   // m92_52 = W*in
   wire signed [14:0] m92_52;
   assign m92_52 ={ {3{in92[14]}} , in92[14:3] };

   // m92_53 = W*in
   wire signed [14:0] m92_53;
   assign m92_53 =15'b0;

   // m92_54 = W*in
   wire signed [14:0] m92_54;
   assign m92_54 =15'b0;

   // m92_55 = W*in
   wire signed [14:0] m92_55;
   assign m92_55 =15'b0;

   // m92_56 = W*in
   wire signed [14:0] m92_56;
   assign m92_56 ={ {3{in92[14]}} , in92[14:3] };

   // m92_57 = W*in
   wire signed [14:0] m92_57;
   assign m92_57 =15'b0;

   // m92_58 = W*in
   wire signed [14:0] m92_58;
   assign m92_58 =15'b0;

   // m92_59 = W*in
   wire signed [14:0] m92_59;
   assign m92_59 ={ {3{in92[14]}} , in92[14:3] };

   // m92_60 = W*in
   wire signed [14:0] m92_60;
   assign m92_60 =15'b0;

   // m92_61 = W*in
   wire signed [14:0] m92_61;
   assign m92_61 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_62 = W*in
   wire signed [14:0] m92_62;
   assign m92_62 =15'b0;

   // m92_63 = W*in
   wire signed [14:0] m92_63;
   assign m92_63 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_64 = W*in
   wire signed [14:0] m92_64;
   assign m92_64 ={ {4{in92[14]}} , in92[14:4] };

   // m92_65 = W*in
   wire signed [14:0] m92_65;
   assign m92_65 =15'b0;

   // m92_66 = W*in
   wire signed [14:0] m92_66;
   assign m92_66 ={ {4{neg92[14]}} , neg92[14:4] };

   // m92_67 = W*in
   wire signed [14:0] m92_67;
   assign m92_67 ={ {4{neg92[14]}} , neg92[14:4] };

   // m92_68 = W*in
   wire signed [14:0] m92_68;
   assign m92_68 =15'b0;

   // m92_69 = W*in
   wire signed [14:0] m92_69;
   assign m92_69 =15'b0;

   // m92_70 = W*in
   wire signed [14:0] m92_70;
   assign m92_70 ={ {3{in92[14]}} , in92[14:3] };

   // m92_71 = W*in
   wire signed [14:0] m92_71;
   assign m92_71 =15'b0;

   // m92_72 = W*in
   wire signed [14:0] m92_72;
   assign m92_72 =15'b0;

   // m92_73 = W*in
   wire signed [14:0] m92_73;
   assign m92_73 =15'b0;

   // m92_74 = W*in
   wire signed [14:0] m92_74;
   assign m92_74 =15'b0;

   // m92_75 = W*in
   wire signed [14:0] m92_75;
   assign m92_75 ={ {3{in92[14]}} , in92[14:3] };

   // m92_76 = W*in
   wire signed [14:0] m92_76;
   assign m92_76 =15'b0;

   // m92_77 = W*in
   wire signed [14:0] m92_77;
   assign m92_77 =15'b0;

   // m92_78 = W*in
   wire signed [14:0] m92_78;
   assign m92_78 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_79 = W*in
   wire signed [14:0] m92_79;
   assign m92_79 ={ {3{in92[14]}} , in92[14:3] };

   // m92_80 = W*in
   wire signed [14:0] m92_80;
   assign m92_80 =15'b0;

   // m92_81 = W*in
   wire signed [14:0] m92_81;
   assign m92_81 =15'b0;

   // m92_82 = W*in
   wire signed [14:0] m92_82;
   assign m92_82 =15'b0;

   // m92_83 = W*in
   wire signed [14:0] m92_83;
   assign m92_83 =15'b0;

   // m92_84 = W*in
   wire signed [14:0] m92_84;
   assign m92_84 =15'b0;

   // m92_85 = W*in
   wire signed [14:0] m92_85;
   assign m92_85 =15'b0;

   // m92_86 = W*in
   wire signed [14:0] m92_86;
   assign m92_86 ={ {3{in92[14]}} , in92[14:3] };

   // m92_87 = W*in
   wire signed [14:0] m92_87;
   assign m92_87 =15'b0;

   // m92_88 = W*in
   wire signed [14:0] m92_88;
   assign m92_88 ={ {3{in92[14]}} , in92[14:3] };

   // m92_89 = W*in
   wire signed [14:0] m92_89;
   assign m92_89 =15'b0;

   // m92_90 = W*in
   wire signed [14:0] m92_90;
   assign m92_90 =15'b0;

   // m92_91 = W*in
   wire signed [14:0] m92_91;
   assign m92_91 =15'b0;

   // m92_92 = W*in
   wire signed [14:0] m92_92;
   assign m92_92 =15'b0;

   // m92_93 = W*in
   wire signed [14:0] m92_93;
   assign m92_93 =15'b0;

   // m92_94 = W*in
   wire signed [14:0] m92_94;
   assign m92_94 =15'b0;

   // m92_95 = W*in
   wire signed [14:0] m92_95;
   assign m92_95 =15'b0;

   // m92_96 = W*in
   wire signed [14:0] m92_96;
   assign m92_96 =15'b0;

   // m92_97 = W*in
   wire signed [14:0] m92_97;
   assign m92_97 ={ {3{neg92[14]}} , neg92[14:3] };

   // m92_98 = W*in
   wire signed [14:0] m92_98;
   assign m92_98 =15'b0;

   // m92_99 = W*in
   wire signed [14:0] m92_99;
   assign m92_99 ={ {3{in92[14]}} , in92[14:3] };

   // m92_100 = W*in
   wire signed [14:0] m92_100;
   assign m92_100 =15'b0;

   // m93_1 = W*in
   wire signed [14:0] m93_1;
   assign m93_1 =15'b0;

   // m93_2 = W*in
   wire signed [14:0] m93_2;
   assign m93_2 =15'b0;

   // m93_3 = W*in
   wire signed [14:0] m93_3;
   assign m93_3 =15'b0;

   // m93_4 = W*in
   wire signed [14:0] m93_4;
   assign m93_4 =15'b0;

   // m93_5 = W*in
   wire signed [14:0] m93_5;
   assign m93_5 =15'b0;

   // m93_6 = W*in
   wire signed [14:0] m93_6;
   assign m93_6 =15'b0;

   // m93_7 = W*in
   wire signed [14:0] m93_7;
   assign m93_7 =15'b0;

   // m93_8 = W*in
   wire signed [14:0] m93_8;
   assign m93_8 =15'b0;

   // m93_9 = W*in
   wire signed [14:0] m93_9;
   assign m93_9 =15'b0;

   // m93_10 = W*in
   wire signed [14:0] m93_10;
   assign m93_10 ={ {3{in93[14]}} , in93[14:3] };

   // m93_11 = W*in
   wire signed [14:0] m93_11;
   assign m93_11 =15'b0;

   // m93_12 = W*in
   wire signed [14:0] m93_12;
   assign m93_12 ={ {3{in93[14]}} , in93[14:3] };

   // m93_13 = W*in
   wire signed [14:0] m93_13;
   assign m93_13 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_14 = W*in
   wire signed [14:0] m93_14;
   assign m93_14 =15'b0;

   // m93_15 = W*in
   wire signed [14:0] m93_15;
   assign m93_15 ={ {3{in93[14]}} , in93[14:3] };

   // m93_16 = W*in
   wire signed [14:0] m93_16;
   assign m93_16 ={ {2{in93[14]}} , in93[14:2] };

   // m93_17 = W*in
   wire signed [14:0] m93_17;
   assign m93_17 ={ {4{neg93[14]}} , neg93[14:4] };

   // m93_18 = W*in
   wire signed [14:0] m93_18;
   assign m93_18 =15'b0;

   // m93_19 = W*in
   wire signed [14:0] m93_19;
   assign m93_19 =15'b0;

   // m93_20 = W*in
   wire signed [14:0] m93_20;
   assign m93_20 ={ {4{neg93[14]}} , neg93[14:4] };

   // m93_21 = W*in
   wire signed [14:0] m93_21;
   assign m93_21 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_22 = W*in
   wire signed [14:0] m93_22;
   assign m93_22 ={ {3{in93[14]}} , in93[14:3] };

   // m93_23 = W*in
   wire signed [14:0] m93_23;
   assign m93_23 =15'b0;

   // m93_24 = W*in
   wire signed [14:0] m93_24;
   assign m93_24 =15'b0;

   // m93_25 = W*in
   wire signed [14:0] m93_25;
   assign m93_25 =15'b0;

   // m93_26 = W*in
   wire signed [14:0] m93_26;
   assign m93_26 ={ {2{in93[14]}} , in93[14:2] };

   // m93_27 = W*in
   wire signed [14:0] m93_27;
   assign m93_27 =15'b0;

   // m93_28 = W*in
   wire signed [14:0] m93_28;
   assign m93_28 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_29 = W*in
   wire signed [14:0] m93_29;
   assign m93_29 =15'b0;

   // m93_30 = W*in
   wire signed [14:0] m93_30;
   assign m93_30 =15'b0;

   // m93_31 = W*in
   wire signed [14:0] m93_31;
   assign m93_31 ={ {3{in93[14]}} , in93[14:3] };

   // m93_32 = W*in
   wire signed [14:0] m93_32;
   assign m93_32 =15'b0;

   // m93_33 = W*in
   wire signed [14:0] m93_33;
   assign m93_33 =15'b0;

   // m93_34 = W*in
   wire signed [14:0] m93_34;
   assign m93_34 =15'b0;

   // m93_35 = W*in
   wire signed [14:0] m93_35;
   assign m93_35 =15'b0;

   // m93_36 = W*in
   wire signed [14:0] m93_36;
   assign m93_36 =15'b0;

   // m93_37 = W*in
   wire signed [14:0] m93_37;
   assign m93_37 =15'b0;

   // m93_38 = W*in
   wire signed [14:0] m93_38;
   assign m93_38 =15'b0;

   // m93_39 = W*in
   wire signed [14:0] m93_39;
   assign m93_39 =15'b0;

   // m93_40 = W*in
   wire signed [14:0] m93_40;
   assign m93_40 =15'b0;

   // m93_41 = W*in
   wire signed [14:0] m93_41;
   assign m93_41 =15'b0;

   // m93_42 = W*in
   wire signed [14:0] m93_42;
   assign m93_42 =15'b0;

   // m93_43 = W*in
   wire signed [14:0] m93_43;
   assign m93_43 =15'b0;

   // m93_44 = W*in
   wire signed [14:0] m93_44;
   assign m93_44 =15'b0;

   // m93_45 = W*in
   wire signed [14:0] m93_45;
   assign m93_45 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_46 = W*in
   wire signed [14:0] m93_46;
   assign m93_46 =15'b0;

   // m93_47 = W*in
   wire signed [14:0] m93_47;
   assign m93_47 ={ {3{in93[14]}} , in93[14:3] };

   // m93_48 = W*in
   wire signed [14:0] m93_48;
   assign m93_48 =15'b0;

   // m93_49 = W*in
   wire signed [14:0] m93_49;
   assign m93_49 =15'b0;

   // m93_50 = W*in
   wire signed [14:0] m93_50;
   assign m93_50 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_51 = W*in
   wire signed [14:0] m93_51;
   assign m93_51 =15'b0;

   // m93_52 = W*in
   wire signed [14:0] m93_52;
   assign m93_52 =15'b0;

   // m93_53 = W*in
   wire signed [14:0] m93_53;
   assign m93_53 =15'b0;

   // m93_54 = W*in
   wire signed [14:0] m93_54;
   assign m93_54 =15'b0;

   // m93_55 = W*in
   wire signed [14:0] m93_55;
   assign m93_55 =15'b0;

   // m93_56 = W*in
   wire signed [14:0] m93_56;
   assign m93_56 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_57 = W*in
   wire signed [14:0] m93_57;
   assign m93_57 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_58 = W*in
   wire signed [14:0] m93_58;
   assign m93_58 =15'b0;

   // m93_59 = W*in
   wire signed [14:0] m93_59;
   assign m93_59 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_60 = W*in
   wire signed [14:0] m93_60;
   assign m93_60 =15'b0;

   // m93_61 = W*in
   wire signed [14:0] m93_61;
   assign m93_61 =15'b0;

   // m93_62 = W*in
   wire signed [14:0] m93_62;
   assign m93_62 =15'b0;

   // m93_63 = W*in
   wire signed [14:0] m93_63;
   assign m93_63 =15'b0;

   // m93_64 = W*in
   wire signed [14:0] m93_64;
   assign m93_64 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_65 = W*in
   wire signed [14:0] m93_65;
   assign m93_65 ={ {2{in93[14]}} , in93[14:2] };

   // m93_66 = W*in
   wire signed [14:0] m93_66;
   assign m93_66 ={ {3{in93[14]}} , in93[14:3] };

   // m93_67 = W*in
   wire signed [14:0] m93_67;
   assign m93_67 =15'b0;

   // m93_68 = W*in
   wire signed [14:0] m93_68;
   assign m93_68 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_69 = W*in
   wire signed [14:0] m93_69;
   assign m93_69 =15'b0;

   // m93_70 = W*in
   wire signed [14:0] m93_70;
   assign m93_70 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_71 = W*in
   wire signed [14:0] m93_71;
   assign m93_71 =15'b0;

   // m93_72 = W*in
   wire signed [14:0] m93_72;
   assign m93_72 =15'b0;

   // m93_73 = W*in
   wire signed [14:0] m93_73;
   assign m93_73 =15'b0;

   // m93_74 = W*in
   wire signed [14:0] m93_74;
   assign m93_74 ={ {4{neg93[14]}} , neg93[14:4] };

   // m93_75 = W*in
   wire signed [14:0] m93_75;
   assign m93_75 =15'b0;

   // m93_76 = W*in
   wire signed [14:0] m93_76;
   assign m93_76 =15'b0;

   // m93_77 = W*in
   wire signed [14:0] m93_77;
   assign m93_77 ={ {4{neg93[14]}} , neg93[14:4] };

   // m93_78 = W*in
   wire signed [14:0] m93_78;
   assign m93_78 =15'b0;

   // m93_79 = W*in
   wire signed [14:0] m93_79;
   assign m93_79 =15'b0;

   // m93_80 = W*in
   wire signed [14:0] m93_80;
   assign m93_80 =15'b0;

   // m93_81 = W*in
   wire signed [14:0] m93_81;
   assign m93_81 =15'b0;

   // m93_82 = W*in
   wire signed [14:0] m93_82;
   assign m93_82 =15'b0;

   // m93_83 = W*in
   wire signed [14:0] m93_83;
   assign m93_83 ={ {3{in93[14]}} , in93[14:3] };

   // m93_84 = W*in
   wire signed [14:0] m93_84;
   assign m93_84 =15'b0;

   // m93_85 = W*in
   wire signed [14:0] m93_85;
   assign m93_85 =15'b0;

   // m93_86 = W*in
   wire signed [14:0] m93_86;
   assign m93_86 =15'b0;

   // m93_87 = W*in
   wire signed [14:0] m93_87;
   assign m93_87 =15'b0;

   // m93_88 = W*in
   wire signed [14:0] m93_88;
   assign m93_88 =15'b0;

   // m93_89 = W*in
   wire signed [14:0] m93_89;
   assign m93_89 =15'b0;

   // m93_90 = W*in
   wire signed [14:0] m93_90;
   assign m93_90 =15'b0;

   // m93_91 = W*in
   wire signed [14:0] m93_91;
   assign m93_91 =15'b0;

   // m93_92 = W*in
   wire signed [14:0] m93_92;
   assign m93_92 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_93 = W*in
   wire signed [14:0] m93_93;
   assign m93_93 =15'b0;

   // m93_94 = W*in
   wire signed [14:0] m93_94;
   assign m93_94 =15'b0;

   // m93_95 = W*in
   wire signed [14:0] m93_95;
   assign m93_95 =15'b0;

   // m93_96 = W*in
   wire signed [14:0] m93_96;
   assign m93_96 =15'b0;

   // m93_97 = W*in
   wire signed [14:0] m93_97;
   assign m93_97 =15'b0;

   // m93_98 = W*in
   wire signed [14:0] m93_98;
   assign m93_98 =15'b0;

   // m93_99 = W*in
   wire signed [14:0] m93_99;
   assign m93_99 ={ {3{neg93[14]}} , neg93[14:3] };

   // m93_100 = W*in
   wire signed [14:0] m93_100;
   assign m93_100 =15'b0;

   // m94_1 = W*in
   wire signed [14:0] m94_1;
   assign m94_1 =15'b0;

   // m94_2 = W*in
   wire signed [14:0] m94_2;
   assign m94_2 =15'b0;

   // m94_3 = W*in
   wire signed [14:0] m94_3;
   assign m94_3 ={ {3{in94[14]}} , in94[14:3] };

   // m94_4 = W*in
   wire signed [14:0] m94_4;
   assign m94_4 =15'b0;

   // m94_5 = W*in
   wire signed [14:0] m94_5;
   assign m94_5 =15'b0;

   // m94_6 = W*in
   wire signed [14:0] m94_6;
   assign m94_6 =15'b0;

   // m94_7 = W*in
   wire signed [14:0] m94_7;
   assign m94_7 =15'b0;

   // m94_8 = W*in
   wire signed [14:0] m94_8;
   assign m94_8 =15'b0;

   // m94_9 = W*in
   wire signed [14:0] m94_9;
   assign m94_9 =15'b0;

   // m94_10 = W*in
   wire signed [14:0] m94_10;
   assign m94_10 =15'b0;

   // m94_11 = W*in
   wire signed [14:0] m94_11;
   assign m94_11 =15'b0;

   // m94_12 = W*in
   wire signed [14:0] m94_12;
   assign m94_12 =15'b0;

   // m94_13 = W*in
   wire signed [14:0] m94_13;
   assign m94_13 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_14 = W*in
   wire signed [14:0] m94_14;
   assign m94_14 =15'b0;

   // m94_15 = W*in
   wire signed [14:0] m94_15;
   assign m94_15 =15'b0;

   // m94_16 = W*in
   wire signed [14:0] m94_16;
   assign m94_16 =15'b0;

   // m94_17 = W*in
   wire signed [14:0] m94_17;
   assign m94_17 =15'b0;

   // m94_18 = W*in
   wire signed [14:0] m94_18;
   assign m94_18 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_19 = W*in
   wire signed [14:0] m94_19;
   assign m94_19 =15'b0;

   // m94_20 = W*in
   wire signed [14:0] m94_20;
   assign m94_20 =15'b0;

   // m94_21 = W*in
   wire signed [14:0] m94_21;
   assign m94_21 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_22 = W*in
   wire signed [14:0] m94_22;
   assign m94_22 =15'b0;

   // m94_23 = W*in
   wire signed [14:0] m94_23;
   assign m94_23 =15'b0;

   // m94_24 = W*in
   wire signed [14:0] m94_24;
   assign m94_24 ={ {3{in94[14]}} , in94[14:3] };

   // m94_25 = W*in
   wire signed [14:0] m94_25;
   assign m94_25 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_26 = W*in
   wire signed [14:0] m94_26;
   assign m94_26 ={ {3{in94[14]}} , in94[14:3] };

   // m94_27 = W*in
   wire signed [14:0] m94_27;
   assign m94_27 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_28 = W*in
   wire signed [14:0] m94_28;
   assign m94_28 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_29 = W*in
   wire signed [14:0] m94_29;
   assign m94_29 ={ {3{in94[14]}} , in94[14:3] };

   // m94_30 = W*in
   wire signed [14:0] m94_30;
   assign m94_30 =15'b0;

   // m94_31 = W*in
   wire signed [14:0] m94_31;
   assign m94_31 ={ {4{in94[14]}} , in94[14:4] };

   // m94_32 = W*in
   wire signed [14:0] m94_32;
   assign m94_32 =15'b0;

   // m94_33 = W*in
   wire signed [14:0] m94_33;
   assign m94_33 =15'b0;

   // m94_34 = W*in
   wire signed [14:0] m94_34;
   assign m94_34 =15'b0;

   // m94_35 = W*in
   wire signed [14:0] m94_35;
   assign m94_35 =15'b0;

   // m94_36 = W*in
   wire signed [14:0] m94_36;
   assign m94_36 =15'b0;

   // m94_37 = W*in
   wire signed [14:0] m94_37;
   assign m94_37 =15'b0;

   // m94_38 = W*in
   wire signed [14:0] m94_38;
   assign m94_38 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_39 = W*in
   wire signed [14:0] m94_39;
   assign m94_39 =15'b0;

   // m94_40 = W*in
   wire signed [14:0] m94_40;
   assign m94_40 ={ {4{neg94[14]}} , neg94[14:4] };

   // m94_41 = W*in
   wire signed [14:0] m94_41;
   assign m94_41 ={ {4{neg94[14]}} , neg94[14:4] };

   // m94_42 = W*in
   wire signed [14:0] m94_42;
   assign m94_42 =15'b0;

   // m94_43 = W*in
   wire signed [14:0] m94_43;
   assign m94_43 =15'b0;

   // m94_44 = W*in
   wire signed [14:0] m94_44;
   assign m94_44 =15'b0;

   // m94_45 = W*in
   wire signed [14:0] m94_45;
   assign m94_45 =15'b0;

   // m94_46 = W*in
   wire signed [14:0] m94_46;
   assign m94_46 =15'b0;

   // m94_47 = W*in
   wire signed [14:0] m94_47;
   assign m94_47 ={ {3{in94[14]}} , in94[14:3] };

   // m94_48 = W*in
   wire signed [14:0] m94_48;
   assign m94_48 =15'b0;

   // m94_49 = W*in
   wire signed [14:0] m94_49;
   assign m94_49 =15'b0;

   // m94_50 = W*in
   wire signed [14:0] m94_50;
   assign m94_50 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_51 = W*in
   wire signed [14:0] m94_51;
   assign m94_51 =15'b0;

   // m94_52 = W*in
   wire signed [14:0] m94_52;
   assign m94_52 =15'b0;

   // m94_53 = W*in
   wire signed [14:0] m94_53;
   assign m94_53 =15'b0;

   // m94_54 = W*in
   wire signed [14:0] m94_54;
   assign m94_54 =15'b0;

   // m94_55 = W*in
   wire signed [14:0] m94_55;
   assign m94_55 =15'b0;

   // m94_56 = W*in
   wire signed [14:0] m94_56;
   assign m94_56 =15'b0;

   // m94_57 = W*in
   wire signed [14:0] m94_57;
   assign m94_57 ={ {3{in94[14]}} , in94[14:3] };

   // m94_58 = W*in
   wire signed [14:0] m94_58;
   assign m94_58 =15'b0;

   // m94_59 = W*in
   wire signed [14:0] m94_59;
   assign m94_59 =15'b0;

   // m94_60 = W*in
   wire signed [14:0] m94_60;
   assign m94_60 =15'b0;

   // m94_61 = W*in
   wire signed [14:0] m94_61;
   assign m94_61 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_62 = W*in
   wire signed [14:0] m94_62;
   assign m94_62 =15'b0;

   // m94_63 = W*in
   wire signed [14:0] m94_63;
   assign m94_63 =15'b0;

   // m94_64 = W*in
   wire signed [14:0] m94_64;
   assign m94_64 =15'b0;

   // m94_65 = W*in
   wire signed [14:0] m94_65;
   assign m94_65 ={ {3{in94[14]}} , in94[14:3] };

   // m94_66 = W*in
   wire signed [14:0] m94_66;
   assign m94_66 =15'b0;

   // m94_67 = W*in
   wire signed [14:0] m94_67;
   assign m94_67 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_68 = W*in
   wire signed [14:0] m94_68;
   assign m94_68 ={ {4{neg94[14]}} , neg94[14:4] };

   // m94_69 = W*in
   wire signed [14:0] m94_69;
   assign m94_69 ={ {4{in94[14]}} , in94[14:4] };

   // m94_70 = W*in
   wire signed [14:0] m94_70;
   assign m94_70 ={ {3{in94[14]}} , in94[14:3] };

   // m94_71 = W*in
   wire signed [14:0] m94_71;
   assign m94_71 =15'b0;

   // m94_72 = W*in
   wire signed [14:0] m94_72;
   assign m94_72 =15'b0;

   // m94_73 = W*in
   wire signed [14:0] m94_73;
   assign m94_73 =15'b0;

   // m94_74 = W*in
   wire signed [14:0] m94_74;
   assign m94_74 =15'b0;

   // m94_75 = W*in
   wire signed [14:0] m94_75;
   assign m94_75 =15'b0;

   // m94_76 = W*in
   wire signed [14:0] m94_76;
   assign m94_76 =15'b0;

   // m94_77 = W*in
   wire signed [14:0] m94_77;
   assign m94_77 =15'b0;

   // m94_78 = W*in
   wire signed [14:0] m94_78;
   assign m94_78 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_79 = W*in
   wire signed [14:0] m94_79;
   assign m94_79 =15'b0;

   // m94_80 = W*in
   wire signed [14:0] m94_80;
   assign m94_80 =15'b0;

   // m94_81 = W*in
   wire signed [14:0] m94_81;
   assign m94_81 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_82 = W*in
   wire signed [14:0] m94_82;
   assign m94_82 =15'b0;

   // m94_83 = W*in
   wire signed [14:0] m94_83;
   assign m94_83 =15'b0;

   // m94_84 = W*in
   wire signed [14:0] m94_84;
   assign m94_84 =15'b0;

   // m94_85 = W*in
   wire signed [14:0] m94_85;
   assign m94_85 =15'b0;

   // m94_86 = W*in
   wire signed [14:0] m94_86;
   assign m94_86 =15'b0;

   // m94_87 = W*in
   wire signed [14:0] m94_87;
   assign m94_87 =15'b0;

   // m94_88 = W*in
   wire signed [14:0] m94_88;
   assign m94_88 =15'b0;

   // m94_89 = W*in
   wire signed [14:0] m94_89;
   assign m94_89 =15'b0;

   // m94_90 = W*in
   wire signed [14:0] m94_90;
   assign m94_90 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_91 = W*in
   wire signed [14:0] m94_91;
   assign m94_91 ={ {3{in94[14]}} , in94[14:3] };

   // m94_92 = W*in
   wire signed [14:0] m94_92;
   assign m94_92 =15'b0;

   // m94_93 = W*in
   wire signed [14:0] m94_93;
   assign m94_93 ={ {3{in94[14]}} , in94[14:3] };

   // m94_94 = W*in
   wire signed [14:0] m94_94;
   assign m94_94 =15'b0;

   // m94_95 = W*in
   wire signed [14:0] m94_95;
   assign m94_95 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_96 = W*in
   wire signed [14:0] m94_96;
   assign m94_96 =15'b0;

   // m94_97 = W*in
   wire signed [14:0] m94_97;
   assign m94_97 ={ {3{neg94[14]}} , neg94[14:3] };

   // m94_98 = W*in
   wire signed [14:0] m94_98;
   assign m94_98 =15'b0;

   // m94_99 = W*in
   wire signed [14:0] m94_99;
   assign m94_99 =15'b0;

   // m94_100 = W*in
   wire signed [14:0] m94_100;
   assign m94_100 =15'b0;

   // m95_1 = W*in
   wire signed [14:0] m95_1;
   assign m95_1 =15'b0;

   // m95_2 = W*in
   wire signed [14:0] m95_2;
   assign m95_2 =15'b0;

   // m95_3 = W*in
   wire signed [14:0] m95_3;
   assign m95_3 =15'b0;

   // m95_4 = W*in
   wire signed [14:0] m95_4;
   assign m95_4 =15'b0;

   // m95_5 = W*in
   wire signed [14:0] m95_5;
   assign m95_5 =15'b0;

   // m95_6 = W*in
   wire signed [14:0] m95_6;
   assign m95_6 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_7 = W*in
   wire signed [14:0] m95_7;
   assign m95_7 =15'b0;

   // m95_8 = W*in
   wire signed [14:0] m95_8;
   assign m95_8 =15'b0;

   // m95_9 = W*in
   wire signed [14:0] m95_9;
   assign m95_9 =15'b0;

   // m95_10 = W*in
   wire signed [14:0] m95_10;
   assign m95_10 ={ {3{in95[14]}} , in95[14:3] };

   // m95_11 = W*in
   wire signed [14:0] m95_11;
   assign m95_11 =15'b0;

   // m95_12 = W*in
   wire signed [14:0] m95_12;
   assign m95_12 =15'b0;

   // m95_13 = W*in
   wire signed [14:0] m95_13;
   assign m95_13 =15'b0;

   // m95_14 = W*in
   wire signed [14:0] m95_14;
   assign m95_14 =15'b0;

   // m95_15 = W*in
   wire signed [14:0] m95_15;
   assign m95_15 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_16 = W*in
   wire signed [14:0] m95_16;
   assign m95_16 =15'b0;

   // m95_17 = W*in
   wire signed [14:0] m95_17;
   assign m95_17 ={ {4{in95[14]}} , in95[14:4] };

   // m95_18 = W*in
   wire signed [14:0] m95_18;
   assign m95_18 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_19 = W*in
   wire signed [14:0] m95_19;
   assign m95_19 ={ {3{in95[14]}} , in95[14:3] };

   // m95_20 = W*in
   wire signed [14:0] m95_20;
   assign m95_20 =15'b0;

   // m95_21 = W*in
   wire signed [14:0] m95_21;
   assign m95_21 =15'b0;

   // m95_22 = W*in
   wire signed [14:0] m95_22;
   assign m95_22 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_23 = W*in
   wire signed [14:0] m95_23;
   assign m95_23 =15'b0;

   // m95_24 = W*in
   wire signed [14:0] m95_24;
   assign m95_24 =15'b0;

   // m95_25 = W*in
   wire signed [14:0] m95_25;
   assign m95_25 ={ {3{in95[14]}} , in95[14:3] };

   // m95_26 = W*in
   wire signed [14:0] m95_26;
   assign m95_26 =15'b0;

   // m95_27 = W*in
   wire signed [14:0] m95_27;
   assign m95_27 =15'b0;

   // m95_28 = W*in
   wire signed [14:0] m95_28;
   assign m95_28 =15'b0;

   // m95_29 = W*in
   wire signed [14:0] m95_29;
   assign m95_29 =15'b0;

   // m95_30 = W*in
   wire signed [14:0] m95_30;
   assign m95_30 =15'b0;

   // m95_31 = W*in
   wire signed [14:0] m95_31;
   assign m95_31 =15'b0;

   // m95_32 = W*in
   wire signed [14:0] m95_32;
   assign m95_32 ={ {3{in95[14]}} , in95[14:3] };

   // m95_33 = W*in
   wire signed [14:0] m95_33;
   assign m95_33 ={ {3{in95[14]}} , in95[14:3] };

   // m95_34 = W*in
   wire signed [14:0] m95_34;
   assign m95_34 =15'b0;

   // m95_35 = W*in
   wire signed [14:0] m95_35;
   assign m95_35 =15'b0;

   // m95_36 = W*in
   wire signed [14:0] m95_36;
   assign m95_36 =15'b0;

   // m95_37 = W*in
   wire signed [14:0] m95_37;
   assign m95_37 =15'b0;

   // m95_38 = W*in
   wire signed [14:0] m95_38;
   assign m95_38 =15'b0;

   // m95_39 = W*in
   wire signed [14:0] m95_39;
   assign m95_39 =15'b0;

   // m95_40 = W*in
   wire signed [14:0] m95_40;
   assign m95_40 =15'b0;

   // m95_41 = W*in
   wire signed [14:0] m95_41;
   assign m95_41 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_42 = W*in
   wire signed [14:0] m95_42;
   assign m95_42 =15'b0;

   // m95_43 = W*in
   wire signed [14:0] m95_43;
   assign m95_43 =15'b0;

   // m95_44 = W*in
   wire signed [14:0] m95_44;
   assign m95_44 ={ {3{in95[14]}} , in95[14:3] };

   // m95_45 = W*in
   wire signed [14:0] m95_45;
   assign m95_45 =15'b0;

   // m95_46 = W*in
   wire signed [14:0] m95_46;
   assign m95_46 =15'b0;

   // m95_47 = W*in
   wire signed [14:0] m95_47;
   assign m95_47 ={ {3{in95[14]}} , in95[14:3] };

   // m95_48 = W*in
   wire signed [14:0] m95_48;
   assign m95_48 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_49 = W*in
   wire signed [14:0] m95_49;
   assign m95_49 =15'b0;

   // m95_50 = W*in
   wire signed [14:0] m95_50;
   assign m95_50 =15'b0;

   // m95_51 = W*in
   wire signed [14:0] m95_51;
   assign m95_51 =15'b0;

   // m95_52 = W*in
   wire signed [14:0] m95_52;
   assign m95_52 =15'b0;

   // m95_53 = W*in
   wire signed [14:0] m95_53;
   assign m95_53 =15'b0;

   // m95_54 = W*in
   wire signed [14:0] m95_54;
   assign m95_54 =15'b0;

   // m95_55 = W*in
   wire signed [14:0] m95_55;
   assign m95_55 =15'b0;

   // m95_56 = W*in
   wire signed [14:0] m95_56;
   assign m95_56 =15'b0;

   // m95_57 = W*in
   wire signed [14:0] m95_57;
   assign m95_57 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_58 = W*in
   wire signed [14:0] m95_58;
   assign m95_58 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_59 = W*in
   wire signed [14:0] m95_59;
   assign m95_59 ={ {3{in95[14]}} , in95[14:3] };

   // m95_60 = W*in
   wire signed [14:0] m95_60;
   assign m95_60 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_61 = W*in
   wire signed [14:0] m95_61;
   assign m95_61 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_62 = W*in
   wire signed [14:0] m95_62;
   assign m95_62 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_63 = W*in
   wire signed [14:0] m95_63;
   assign m95_63 =15'b0;

   // m95_64 = W*in
   wire signed [14:0] m95_64;
   assign m95_64 =15'b0;

   // m95_65 = W*in
   wire signed [14:0] m95_65;
   assign m95_65 =15'b0;

   // m95_66 = W*in
   wire signed [14:0] m95_66;
   assign m95_66 =15'b0;

   // m95_67 = W*in
   wire signed [14:0] m95_67;
   assign m95_67 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_68 = W*in
   wire signed [14:0] m95_68;
   assign m95_68 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_69 = W*in
   wire signed [14:0] m95_69;
   assign m95_69 =15'b0;

   // m95_70 = W*in
   wire signed [14:0] m95_70;
   assign m95_70 ={ {4{in95[14]}} , in95[14:4] };

   // m95_71 = W*in
   wire signed [14:0] m95_71;
   assign m95_71 =15'b0;

   // m95_72 = W*in
   wire signed [14:0] m95_72;
   assign m95_72 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_73 = W*in
   wire signed [14:0] m95_73;
   assign m95_73 =15'b0;

   // m95_74 = W*in
   wire signed [14:0] m95_74;
   assign m95_74 =15'b0;

   // m95_75 = W*in
   wire signed [14:0] m95_75;
   assign m95_75 ={ {3{in95[14]}} , in95[14:3] };

   // m95_76 = W*in
   wire signed [14:0] m95_76;
   assign m95_76 =15'b0;

   // m95_77 = W*in
   wire signed [14:0] m95_77;
   assign m95_77 ={ {4{neg95[14]}} , neg95[14:4] };

   // m95_78 = W*in
   wire signed [14:0] m95_78;
   assign m95_78 =15'b0;

   // m95_79 = W*in
   wire signed [14:0] m95_79;
   assign m95_79 =15'b0;

   // m95_80 = W*in
   wire signed [14:0] m95_80;
   assign m95_80 =15'b0;

   // m95_81 = W*in
   wire signed [14:0] m95_81;
   assign m95_81 =15'b0;

   // m95_82 = W*in
   wire signed [14:0] m95_82;
   assign m95_82 =15'b0;

   // m95_83 = W*in
   wire signed [14:0] m95_83;
   assign m95_83 =15'b0;

   // m95_84 = W*in
   wire signed [14:0] m95_84;
   assign m95_84 =15'b0;

   // m95_85 = W*in
   wire signed [14:0] m95_85;
   assign m95_85 =15'b0;

   // m95_86 = W*in
   wire signed [14:0] m95_86;
   assign m95_86 =15'b0;

   // m95_87 = W*in
   wire signed [14:0] m95_87;
   assign m95_87 =15'b0;

   // m95_88 = W*in
   wire signed [14:0] m95_88;
   assign m95_88 =15'b0;

   // m95_89 = W*in
   wire signed [14:0] m95_89;
   assign m95_89 =15'b0;

   // m95_90 = W*in
   wire signed [14:0] m95_90;
   assign m95_90 ={ {3{in95[14]}} , in95[14:3] };

   // m95_91 = W*in
   wire signed [14:0] m95_91;
   assign m95_91 =15'b0;

   // m95_92 = W*in
   wire signed [14:0] m95_92;
   assign m95_92 =15'b0;

   // m95_93 = W*in
   wire signed [14:0] m95_93;
   assign m95_93 =15'b0;

   // m95_94 = W*in
   wire signed [14:0] m95_94;
   assign m95_94 ={ {3{in95[14]}} , in95[14:3] };

   // m95_95 = W*in
   wire signed [14:0] m95_95;
   assign m95_95 =15'b0;

   // m95_96 = W*in
   wire signed [14:0] m95_96;
   assign m95_96 ={ {3{neg95[14]}} , neg95[14:3] };

   // m95_97 = W*in
   wire signed [14:0] m95_97;
   assign m95_97 =15'b0;

   // m95_98 = W*in
   wire signed [14:0] m95_98;
   assign m95_98 =15'b0;

   // m95_99 = W*in
   wire signed [14:0] m95_99;
   assign m95_99 =15'b0;

   // m95_100 = W*in
   wire signed [14:0] m95_100;
   assign m95_100 =15'b0;

   // m96_1 = W*in
   wire signed [14:0] m96_1;
   assign m96_1 =15'b0;

   // m96_2 = W*in
   wire signed [14:0] m96_2;
   assign m96_2 =15'b0;

   // m96_3 = W*in
   wire signed [14:0] m96_3;
   assign m96_3 =15'b0;

   // m96_4 = W*in
   wire signed [14:0] m96_4;
   assign m96_4 =15'b0;

   // m96_5 = W*in
   wire signed [14:0] m96_5;
   assign m96_5 =15'b0;

   // m96_6 = W*in
   wire signed [14:0] m96_6;
   assign m96_6 =15'b0;

   // m96_7 = W*in
   wire signed [14:0] m96_7;
   assign m96_7 =15'b0;

   // m96_8 = W*in
   wire signed [14:0] m96_8;
   assign m96_8 =15'b0;

   // m96_9 = W*in
   wire signed [14:0] m96_9;
   assign m96_9 =15'b0;

   // m96_10 = W*in
   wire signed [14:0] m96_10;
   assign m96_10 =15'b0;

   // m96_11 = W*in
   wire signed [14:0] m96_11;
   assign m96_11 =15'b0;

   // m96_12 = W*in
   wire signed [14:0] m96_12;
   assign m96_12 =15'b0;

   // m96_13 = W*in
   wire signed [14:0] m96_13;
   assign m96_13 =15'b0;

   // m96_14 = W*in
   wire signed [14:0] m96_14;
   assign m96_14 =15'b0;

   // m96_15 = W*in
   wire signed [14:0] m96_15;
   assign m96_15 =15'b0;

   // m96_16 = W*in
   wire signed [14:0] m96_16;
   assign m96_16 =15'b0;

   // m96_17 = W*in
   wire signed [14:0] m96_17;
   assign m96_17 =15'b0;

   // m96_18 = W*in
   wire signed [14:0] m96_18;
   assign m96_18 =15'b0;

   // m96_19 = W*in
   wire signed [14:0] m96_19;
   assign m96_19 =15'b0;

   // m96_20 = W*in
   wire signed [14:0] m96_20;
   assign m96_20 =15'b0;

   // m96_21 = W*in
   wire signed [14:0] m96_21;
   assign m96_21 =15'b0;

   // m96_22 = W*in
   wire signed [14:0] m96_22;
   assign m96_22 =15'b0;

   // m96_23 = W*in
   wire signed [14:0] m96_23;
   assign m96_23 =15'b0;

   // m96_24 = W*in
   wire signed [14:0] m96_24;
   assign m96_24 ={ {3{in96[14]}} , in96[14:3] };

   // m96_25 = W*in
   wire signed [14:0] m96_25;
   assign m96_25 =15'b0;

   // m96_26 = W*in
   wire signed [14:0] m96_26;
   assign m96_26 =15'b0;

   // m96_27 = W*in
   wire signed [14:0] m96_27;
   assign m96_27 =15'b0;

   // m96_28 = W*in
   wire signed [14:0] m96_28;
   assign m96_28 =15'b0;

   // m96_29 = W*in
   wire signed [14:0] m96_29;
   assign m96_29 =15'b0;

   // m96_30 = W*in
   wire signed [14:0] m96_30;
   assign m96_30 =15'b0;

   // m96_31 = W*in
   wire signed [14:0] m96_31;
   assign m96_31 =15'b0;

   // m96_32 = W*in
   wire signed [14:0] m96_32;
   assign m96_32 =15'b0;

   // m96_33 = W*in
   wire signed [14:0] m96_33;
   assign m96_33 =15'b0;

   // m96_34 = W*in
   wire signed [14:0] m96_34;
   assign m96_34 =15'b0;

   // m96_35 = W*in
   wire signed [14:0] m96_35;
   assign m96_35 ={ {3{in96[14]}} , in96[14:3] };

   // m96_36 = W*in
   wire signed [14:0] m96_36;
   assign m96_36 =15'b0;

   // m96_37 = W*in
   wire signed [14:0] m96_37;
   assign m96_37 =15'b0;

   // m96_38 = W*in
   wire signed [14:0] m96_38;
   assign m96_38 =15'b0;

   // m96_39 = W*in
   wire signed [14:0] m96_39;
   assign m96_39 ={ {3{neg96[14]}} , neg96[14:3] };

   // m96_40 = W*in
   wire signed [14:0] m96_40;
   assign m96_40 =15'b0;

   // m96_41 = W*in
   wire signed [14:0] m96_41;
   assign m96_41 =15'b0;

   // m96_42 = W*in
   wire signed [14:0] m96_42;
   assign m96_42 =15'b0;

   // m96_43 = W*in
   wire signed [14:0] m96_43;
   assign m96_43 =15'b0;

   // m96_44 = W*in
   wire signed [14:0] m96_44;
   assign m96_44 ={ {4{neg96[14]}} , neg96[14:4] };

   // m96_45 = W*in
   wire signed [14:0] m96_45;
   assign m96_45 =15'b0;

   // m96_46 = W*in
   wire signed [14:0] m96_46;
   assign m96_46 =15'b0;

   // m96_47 = W*in
   wire signed [14:0] m96_47;
   assign m96_47 =15'b0;

   // m96_48 = W*in
   wire signed [14:0] m96_48;
   assign m96_48 =15'b0;

   // m96_49 = W*in
   wire signed [14:0] m96_49;
   assign m96_49 =15'b0;

   // m96_50 = W*in
   wire signed [14:0] m96_50;
   assign m96_50 =15'b0;

   // m96_51 = W*in
   wire signed [14:0] m96_51;
   assign m96_51 =15'b0;

   // m96_52 = W*in
   wire signed [14:0] m96_52;
   assign m96_52 =15'b0;

   // m96_53 = W*in
   wire signed [14:0] m96_53;
   assign m96_53 =15'b0;

   // m96_54 = W*in
   wire signed [14:0] m96_54;
   assign m96_54 =15'b0;

   // m96_55 = W*in
   wire signed [14:0] m96_55;
   assign m96_55 =15'b0;

   // m96_56 = W*in
   wire signed [14:0] m96_56;
   assign m96_56 =15'b0;

   // m96_57 = W*in
   wire signed [14:0] m96_57;
   assign m96_57 =15'b0;

   // m96_58 = W*in
   wire signed [14:0] m96_58;
   assign m96_58 =15'b0;

   // m96_59 = W*in
   wire signed [14:0] m96_59;
   assign m96_59 =15'b0;

   // m96_60 = W*in
   wire signed [14:0] m96_60;
   assign m96_60 =15'b0;

   // m96_61 = W*in
   wire signed [14:0] m96_61;
   assign m96_61 =15'b0;

   // m96_62 = W*in
   wire signed [14:0] m96_62;
   assign m96_62 =15'b0;

   // m96_63 = W*in
   wire signed [14:0] m96_63;
   assign m96_63 =15'b0;

   // m96_64 = W*in
   wire signed [14:0] m96_64;
   assign m96_64 =15'b0;

   // m96_65 = W*in
   wire signed [14:0] m96_65;
   assign m96_65 =15'b0;

   // m96_66 = W*in
   wire signed [14:0] m96_66;
   assign m96_66 =15'b0;

   // m96_67 = W*in
   wire signed [14:0] m96_67;
   assign m96_67 ={ {4{in96[14]}} , in96[14:4] };

   // m96_68 = W*in
   wire signed [14:0] m96_68;
   assign m96_68 ={ {4{neg96[14]}} , neg96[14:4] };

   // m96_69 = W*in
   wire signed [14:0] m96_69;
   assign m96_69 ={ {3{neg96[14]}} , neg96[14:3] };

   // m96_70 = W*in
   wire signed [14:0] m96_70;
   assign m96_70 =15'b0;

   // m96_71 = W*in
   wire signed [14:0] m96_71;
   assign m96_71 =15'b0;

   // m96_72 = W*in
   wire signed [14:0] m96_72;
   assign m96_72 =15'b0;

   // m96_73 = W*in
   wire signed [14:0] m96_73;
   assign m96_73 =15'b0;

   // m96_74 = W*in
   wire signed [14:0] m96_74;
   assign m96_74 =15'b0;

   // m96_75 = W*in
   wire signed [14:0] m96_75;
   assign m96_75 =15'b0;

   // m96_76 = W*in
   wire signed [14:0] m96_76;
   assign m96_76 =15'b0;

   // m96_77 = W*in
   wire signed [14:0] m96_77;
   assign m96_77 =15'b0;

   // m96_78 = W*in
   wire signed [14:0] m96_78;
   assign m96_78 =15'b0;

   // m96_79 = W*in
   wire signed [14:0] m96_79;
   assign m96_79 =15'b0;

   // m96_80 = W*in
   wire signed [14:0] m96_80;
   assign m96_80 =15'b0;

   // m96_81 = W*in
   wire signed [14:0] m96_81;
   assign m96_81 =15'b0;

   // m96_82 = W*in
   wire signed [14:0] m96_82;
   assign m96_82 =15'b0;

   // m96_83 = W*in
   wire signed [14:0] m96_83;
   assign m96_83 =15'b0;

   // m96_84 = W*in
   wire signed [14:0] m96_84;
   assign m96_84 ={ {3{in96[14]}} , in96[14:3] };

   // m96_85 = W*in
   wire signed [14:0] m96_85;
   assign m96_85 =15'b0;

   // m96_86 = W*in
   wire signed [14:0] m96_86;
   assign m96_86 =15'b0;

   // m96_87 = W*in
   wire signed [14:0] m96_87;
   assign m96_87 =15'b0;

   // m96_88 = W*in
   wire signed [14:0] m96_88;
   assign m96_88 =15'b0;

   // m96_89 = W*in
   wire signed [14:0] m96_89;
   assign m96_89 =15'b0;

   // m96_90 = W*in
   wire signed [14:0] m96_90;
   assign m96_90 =15'b0;

   // m96_91 = W*in
   wire signed [14:0] m96_91;
   assign m96_91 =15'b0;

   // m96_92 = W*in
   wire signed [14:0] m96_92;
   assign m96_92 =15'b0;

   // m96_93 = W*in
   wire signed [14:0] m96_93;
   assign m96_93 =15'b0;

   // m96_94 = W*in
   wire signed [14:0] m96_94;
   assign m96_94 ={ {3{neg96[14]}} , neg96[14:3] };

   // m96_95 = W*in
   wire signed [14:0] m96_95;
   assign m96_95 =15'b0;

   // m96_96 = W*in
   wire signed [14:0] m96_96;
   assign m96_96 =15'b0;

   // m96_97 = W*in
   wire signed [14:0] m96_97;
   assign m96_97 =15'b0;

   // m96_98 = W*in
   wire signed [14:0] m96_98;
   assign m96_98 =15'b0;

   // m96_99 = W*in
   wire signed [14:0] m96_99;
   assign m96_99 =15'b0;

   // m96_100 = W*in
   wire signed [14:0] m96_100;
   assign m96_100 =15'b0;

   // m97_1 = W*in
   wire signed [14:0] m97_1;
   assign m97_1 =15'b0;

   // m97_2 = W*in
   wire signed [14:0] m97_2;
   assign m97_2 =15'b0;

   // m97_3 = W*in
   wire signed [14:0] m97_3;
   assign m97_3 =15'b0;

   // m97_4 = W*in
   wire signed [14:0] m97_4;
   assign m97_4 =15'b0;

   // m97_5 = W*in
   wire signed [14:0] m97_5;
   assign m97_5 =15'b0;

   // m97_6 = W*in
   wire signed [14:0] m97_6;
   assign m97_6 ={ {4{neg97[14]}} , neg97[14:4] };

   // m97_7 = W*in
   wire signed [14:0] m97_7;
   assign m97_7 =15'b0;

   // m97_8 = W*in
   wire signed [14:0] m97_8;
   assign m97_8 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_9 = W*in
   wire signed [14:0] m97_9;
   assign m97_9 =15'b0;

   // m97_10 = W*in
   wire signed [14:0] m97_10;
   assign m97_10 =15'b0;

   // m97_11 = W*in
   wire signed [14:0] m97_11;
   assign m97_11 ={ {3{in97[14]}} , in97[14:3] };

   // m97_12 = W*in
   wire signed [14:0] m97_12;
   assign m97_12 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_13 = W*in
   wire signed [14:0] m97_13;
   assign m97_13 =15'b0;

   // m97_14 = W*in
   wire signed [14:0] m97_14;
   assign m97_14 =15'b0;

   // m97_15 = W*in
   wire signed [14:0] m97_15;
   assign m97_15 =15'b0;

   // m97_16 = W*in
   wire signed [14:0] m97_16;
   assign m97_16 =15'b0;

   // m97_17 = W*in
   wire signed [14:0] m97_17;
   assign m97_17 =15'b0;

   // m97_18 = W*in
   wire signed [14:0] m97_18;
   assign m97_18 =15'b0;

   // m97_19 = W*in
   wire signed [14:0] m97_19;
   assign m97_19 =15'b0;

   // m97_20 = W*in
   wire signed [14:0] m97_20;
   assign m97_20 =15'b0;

   // m97_21 = W*in
   wire signed [14:0] m97_21;
   assign m97_21 =15'b0;

   // m97_22 = W*in
   wire signed [14:0] m97_22;
   assign m97_22 =15'b0;

   // m97_23 = W*in
   wire signed [14:0] m97_23;
   assign m97_23 =15'b0;

   // m97_24 = W*in
   wire signed [14:0] m97_24;
   assign m97_24 =15'b0;

   // m97_25 = W*in
   wire signed [14:0] m97_25;
   assign m97_25 =15'b0;

   // m97_26 = W*in
   wire signed [14:0] m97_26;
   assign m97_26 ={ {4{neg97[14]}} , neg97[14:4] };

   // m97_27 = W*in
   wire signed [14:0] m97_27;
   assign m97_27 =15'b0;

   // m97_28 = W*in
   wire signed [14:0] m97_28;
   assign m97_28 =15'b0;

   // m97_29 = W*in
   wire signed [14:0] m97_29;
   assign m97_29 =15'b0;

   // m97_30 = W*in
   wire signed [14:0] m97_30;
   assign m97_30 ={ {3{in97[14]}} , in97[14:3] };

   // m97_31 = W*in
   wire signed [14:0] m97_31;
   assign m97_31 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_32 = W*in
   wire signed [14:0] m97_32;
   assign m97_32 =15'b0;

   // m97_33 = W*in
   wire signed [14:0] m97_33;
   assign m97_33 =15'b0;

   // m97_34 = W*in
   wire signed [14:0] m97_34;
   assign m97_34 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_35 = W*in
   wire signed [14:0] m97_35;
   assign m97_35 =15'b0;

   // m97_36 = W*in
   wire signed [14:0] m97_36;
   assign m97_36 =15'b0;

   // m97_37 = W*in
   wire signed [14:0] m97_37;
   assign m97_37 =15'b0;

   // m97_38 = W*in
   wire signed [14:0] m97_38;
   assign m97_38 =15'b0;

   // m97_39 = W*in
   wire signed [14:0] m97_39;
   assign m97_39 =15'b0;

   // m97_40 = W*in
   wire signed [14:0] m97_40;
   assign m97_40 =15'b0;

   // m97_41 = W*in
   wire signed [14:0] m97_41;
   assign m97_41 =15'b0;

   // m97_42 = W*in
   wire signed [14:0] m97_42;
   assign m97_42 =15'b0;

   // m97_43 = W*in
   wire signed [14:0] m97_43;
   assign m97_43 =15'b0;

   // m97_44 = W*in
   wire signed [14:0] m97_44;
   assign m97_44 =15'b0;

   // m97_45 = W*in
   wire signed [14:0] m97_45;
   assign m97_45 =15'b0;

   // m97_46 = W*in
   wire signed [14:0] m97_46;
   assign m97_46 =15'b0;

   // m97_47 = W*in
   wire signed [14:0] m97_47;
   assign m97_47 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_48 = W*in
   wire signed [14:0] m97_48;
   assign m97_48 ={ {4{neg97[14]}} , neg97[14:4] };

   // m97_49 = W*in
   wire signed [14:0] m97_49;
   assign m97_49 =15'b0;

   // m97_50 = W*in
   wire signed [14:0] m97_50;
   assign m97_50 ={ {3{in97[14]}} , in97[14:3] };

   // m97_51 = W*in
   wire signed [14:0] m97_51;
   assign m97_51 =15'b0;

   // m97_52 = W*in
   wire signed [14:0] m97_52;
   assign m97_52 =15'b0;

   // m97_53 = W*in
   wire signed [14:0] m97_53;
   assign m97_53 =15'b0;

   // m97_54 = W*in
   wire signed [14:0] m97_54;
   assign m97_54 =15'b0;

   // m97_55 = W*in
   wire signed [14:0] m97_55;
   assign m97_55 =15'b0;

   // m97_56 = W*in
   wire signed [14:0] m97_56;
   assign m97_56 =15'b0;

   // m97_57 = W*in
   wire signed [14:0] m97_57;
   assign m97_57 =15'b0;

   // m97_58 = W*in
   wire signed [14:0] m97_58;
   assign m97_58 =15'b0;

   // m97_59 = W*in
   wire signed [14:0] m97_59;
   assign m97_59 =15'b0;

   // m97_60 = W*in
   wire signed [14:0] m97_60;
   assign m97_60 =15'b0;

   // m97_61 = W*in
   wire signed [14:0] m97_61;
   assign m97_61 =15'b0;

   // m97_62 = W*in
   wire signed [14:0] m97_62;
   assign m97_62 =15'b0;

   // m97_63 = W*in
   wire signed [14:0] m97_63;
   assign m97_63 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_64 = W*in
   wire signed [14:0] m97_64;
   assign m97_64 =15'b0;

   // m97_65 = W*in
   wire signed [14:0] m97_65;
   assign m97_65 =15'b0;

   // m97_66 = W*in
   wire signed [14:0] m97_66;
   assign m97_66 =15'b0;

   // m97_67 = W*in
   wire signed [14:0] m97_67;
   assign m97_67 ={ {3{in97[14]}} , in97[14:3] };

   // m97_68 = W*in
   wire signed [14:0] m97_68;
   assign m97_68 =15'b0;

   // m97_69 = W*in
   wire signed [14:0] m97_69;
   assign m97_69 =15'b0;

   // m97_70 = W*in
   wire signed [14:0] m97_70;
   assign m97_70 =15'b0;

   // m97_71 = W*in
   wire signed [14:0] m97_71;
   assign m97_71 =15'b0;

   // m97_72 = W*in
   wire signed [14:0] m97_72;
   assign m97_72 =15'b0;

   // m97_73 = W*in
   wire signed [14:0] m97_73;
   assign m97_73 =15'b0;

   // m97_74 = W*in
   wire signed [14:0] m97_74;
   assign m97_74 =15'b0;

   // m97_75 = W*in
   wire signed [14:0] m97_75;
   assign m97_75 =15'b0;

   // m97_76 = W*in
   wire signed [14:0] m97_76;
   assign m97_76 =15'b0;

   // m97_77 = W*in
   wire signed [14:0] m97_77;
   assign m97_77 =15'b0;

   // m97_78 = W*in
   wire signed [14:0] m97_78;
   assign m97_78 =15'b0;

   // m97_79 = W*in
   wire signed [14:0] m97_79;
   assign m97_79 =15'b0;

   // m97_80 = W*in
   wire signed [14:0] m97_80;
   assign m97_80 ={ {3{neg97[14]}} , neg97[14:3] };

   // m97_81 = W*in
   wire signed [14:0] m97_81;
   assign m97_81 =15'b0;

   // m97_82 = W*in
   wire signed [14:0] m97_82;
   assign m97_82 =15'b0;

   // m97_83 = W*in
   wire signed [14:0] m97_83;
   assign m97_83 =15'b0;

   // m97_84 = W*in
   wire signed [14:0] m97_84;
   assign m97_84 =15'b0;

   // m97_85 = W*in
   wire signed [14:0] m97_85;
   assign m97_85 =15'b0;

   // m97_86 = W*in
   wire signed [14:0] m97_86;
   assign m97_86 ={ {3{in97[14]}} , in97[14:3] };

   // m97_87 = W*in
   wire signed [14:0] m97_87;
   assign m97_87 =15'b0;

   // m97_88 = W*in
   wire signed [14:0] m97_88;
   assign m97_88 =15'b0;

   // m97_89 = W*in
   wire signed [14:0] m97_89;
   assign m97_89 =15'b0;

   // m97_90 = W*in
   wire signed [14:0] m97_90;
   assign m97_90 =15'b0;

   // m97_91 = W*in
   wire signed [14:0] m97_91;
   assign m97_91 =15'b0;

   // m97_92 = W*in
   wire signed [14:0] m97_92;
   assign m97_92 =15'b0;

   // m97_93 = W*in
   wire signed [14:0] m97_93;
   assign m97_93 =15'b0;

   // m97_94 = W*in
   wire signed [14:0] m97_94;
   assign m97_94 =15'b0;

   // m97_95 = W*in
   wire signed [14:0] m97_95;
   assign m97_95 =15'b0;

   // m97_96 = W*in
   wire signed [14:0] m97_96;
   assign m97_96 =15'b0;

   // m97_97 = W*in
   wire signed [14:0] m97_97;
   assign m97_97 =15'b0;

   // m97_98 = W*in
   wire signed [14:0] m97_98;
   assign m97_98 =15'b0;

   // m97_99 = W*in
   wire signed [14:0] m97_99;
   assign m97_99 =15'b0;

   // m97_100 = W*in
   wire signed [14:0] m97_100;
   assign m97_100 =15'b0;

   // m98_1 = W*in
   wire signed [14:0] m98_1;
   assign m98_1 =15'b0;

   // m98_2 = W*in
   wire signed [14:0] m98_2;
   assign m98_2 =15'b0;

   // m98_3 = W*in
   wire signed [14:0] m98_3;
   assign m98_3 =15'b0;

   // m98_4 = W*in
   wire signed [14:0] m98_4;
   assign m98_4 =15'b0;

   // m98_5 = W*in
   wire signed [14:0] m98_5;
   assign m98_5 =15'b0;

   // m98_6 = W*in
   wire signed [14:0] m98_6;
   assign m98_6 =15'b0;

   // m98_7 = W*in
   wire signed [14:0] m98_7;
   assign m98_7 =15'b0;

   // m98_8 = W*in
   wire signed [14:0] m98_8;
   assign m98_8 =15'b0;

   // m98_9 = W*in
   wire signed [14:0] m98_9;
   assign m98_9 ={ {4{neg98[14]}} , neg98[14:4] };

   // m98_10 = W*in
   wire signed [14:0] m98_10;
   assign m98_10 =15'b0;

   // m98_11 = W*in
   wire signed [14:0] m98_11;
   assign m98_11 =15'b0;

   // m98_12 = W*in
   wire signed [14:0] m98_12;
   assign m98_12 =15'b0;

   // m98_13 = W*in
   wire signed [14:0] m98_13;
   assign m98_13 =15'b0;

   // m98_14 = W*in
   wire signed [14:0] m98_14;
   assign m98_14 =15'b0;

   // m98_15 = W*in
   wire signed [14:0] m98_15;
   assign m98_15 =15'b0;

   // m98_16 = W*in
   wire signed [14:0] m98_16;
   assign m98_16 =15'b0;

   // m98_17 = W*in
   wire signed [14:0] m98_17;
   assign m98_17 =15'b0;

   // m98_18 = W*in
   wire signed [14:0] m98_18;
   assign m98_18 =15'b0;

   // m98_19 = W*in
   wire signed [14:0] m98_19;
   assign m98_19 =15'b0;

   // m98_20 = W*in
   wire signed [14:0] m98_20;
   assign m98_20 =15'b0;

   // m98_21 = W*in
   wire signed [14:0] m98_21;
   assign m98_21 =15'b0;

   // m98_22 = W*in
   wire signed [14:0] m98_22;
   assign m98_22 =15'b0;

   // m98_23 = W*in
   wire signed [14:0] m98_23;
   assign m98_23 =15'b0;

   // m98_24 = W*in
   wire signed [14:0] m98_24;
   assign m98_24 =15'b0;

   // m98_25 = W*in
   wire signed [14:0] m98_25;
   assign m98_25 =15'b0;

   // m98_26 = W*in
   wire signed [14:0] m98_26;
   assign m98_26 =15'b0;

   // m98_27 = W*in
   wire signed [14:0] m98_27;
   assign m98_27 =15'b0;

   // m98_28 = W*in
   wire signed [14:0] m98_28;
   assign m98_28 =15'b0;

   // m98_29 = W*in
   wire signed [14:0] m98_29;
   assign m98_29 =15'b0;

   // m98_30 = W*in
   wire signed [14:0] m98_30;
   assign m98_30 =15'b0;

   // m98_31 = W*in
   wire signed [14:0] m98_31;
   assign m98_31 =15'b0;

   // m98_32 = W*in
   wire signed [14:0] m98_32;
   assign m98_32 =15'b0;

   // m98_33 = W*in
   wire signed [14:0] m98_33;
   assign m98_33 =15'b0;

   // m98_34 = W*in
   wire signed [14:0] m98_34;
   assign m98_34 =15'b0;

   // m98_35 = W*in
   wire signed [14:0] m98_35;
   assign m98_35 =15'b0;

   // m98_36 = W*in
   wire signed [14:0] m98_36;
   assign m98_36 =15'b0;

   // m98_37 = W*in
   wire signed [14:0] m98_37;
   assign m98_37 =15'b0;

   // m98_38 = W*in
   wire signed [14:0] m98_38;
   assign m98_38 =15'b0;

   // m98_39 = W*in
   wire signed [14:0] m98_39;
   assign m98_39 =15'b0;

   // m98_40 = W*in
   wire signed [14:0] m98_40;
   assign m98_40 ={ {4{neg98[14]}} , neg98[14:4] };

   // m98_41 = W*in
   wire signed [14:0] m98_41;
   assign m98_41 =15'b0;

   // m98_42 = W*in
   wire signed [14:0] m98_42;
   assign m98_42 =15'b0;

   // m98_43 = W*in
   wire signed [14:0] m98_43;
   assign m98_43 =15'b0;

   // m98_44 = W*in
   wire signed [14:0] m98_44;
   assign m98_44 ={ {3{neg98[14]}} , neg98[14:3] };

   // m98_45 = W*in
   wire signed [14:0] m98_45;
   assign m98_45 =15'b0;

   // m98_46 = W*in
   wire signed [14:0] m98_46;
   assign m98_46 =15'b0;

   // m98_47 = W*in
   wire signed [14:0] m98_47;
   assign m98_47 =15'b0;

   // m98_48 = W*in
   wire signed [14:0] m98_48;
   assign m98_48 =15'b0;

   // m98_49 = W*in
   wire signed [14:0] m98_49;
   assign m98_49 =15'b0;

   // m98_50 = W*in
   wire signed [14:0] m98_50;
   assign m98_50 =15'b0;

   // m98_51 = W*in
   wire signed [14:0] m98_51;
   assign m98_51 =15'b0;

   // m98_52 = W*in
   wire signed [14:0] m98_52;
   assign m98_52 =15'b0;

   // m98_53 = W*in
   wire signed [14:0] m98_53;
   assign m98_53 ={ {3{in98[14]}} , in98[14:3] };

   // m98_54 = W*in
   wire signed [14:0] m98_54;
   assign m98_54 =15'b0;

   // m98_55 = W*in
   wire signed [14:0] m98_55;
   assign m98_55 =15'b0;

   // m98_56 = W*in
   wire signed [14:0] m98_56;
   assign m98_56 =15'b0;

   // m98_57 = W*in
   wire signed [14:0] m98_57;
   assign m98_57 ={ {3{neg98[14]}} , neg98[14:3] };

   // m98_58 = W*in
   wire signed [14:0] m98_58;
   assign m98_58 =15'b0;

   // m98_59 = W*in
   wire signed [14:0] m98_59;
   assign m98_59 =15'b0;

   // m98_60 = W*in
   wire signed [14:0] m98_60;
   assign m98_60 =15'b0;

   // m98_61 = W*in
   wire signed [14:0] m98_61;
   assign m98_61 =15'b0;

   // m98_62 = W*in
   wire signed [14:0] m98_62;
   assign m98_62 =15'b0;

   // m98_63 = W*in
   wire signed [14:0] m98_63;
   assign m98_63 =15'b0;

   // m98_64 = W*in
   wire signed [14:0] m98_64;
   assign m98_64 =15'b0;

   // m98_65 = W*in
   wire signed [14:0] m98_65;
   assign m98_65 =15'b0;

   // m98_66 = W*in
   wire signed [14:0] m98_66;
   assign m98_66 ={ {2{in98[14]}} , in98[14:2] };

   // m98_67 = W*in
   wire signed [14:0] m98_67;
   assign m98_67 =15'b0;

   // m98_68 = W*in
   wire signed [14:0] m98_68;
   assign m98_68 =15'b0;

   // m98_69 = W*in
   wire signed [14:0] m98_69;
   assign m98_69 =15'b0;

   // m98_70 = W*in
   wire signed [14:0] m98_70;
   assign m98_70 =15'b0;

   // m98_71 = W*in
   wire signed [14:0] m98_71;
   assign m98_71 =15'b0;

   // m98_72 = W*in
   wire signed [14:0] m98_72;
   assign m98_72 =15'b0;

   // m98_73 = W*in
   wire signed [14:0] m98_73;
   assign m98_73 =15'b0;

   // m98_74 = W*in
   wire signed [14:0] m98_74;
   assign m98_74 =15'b0;

   // m98_75 = W*in
   wire signed [14:0] m98_75;
   assign m98_75 =15'b0;

   // m98_76 = W*in
   wire signed [14:0] m98_76;
   assign m98_76 =15'b0;

   // m98_77 = W*in
   wire signed [14:0] m98_77;
   assign m98_77 =15'b0;

   // m98_78 = W*in
   wire signed [14:0] m98_78;
   assign m98_78 =15'b0;

   // m98_79 = W*in
   wire signed [14:0] m98_79;
   assign m98_79 ={ {3{in98[14]}} , in98[14:3] };

   // m98_80 = W*in
   wire signed [14:0] m98_80;
   assign m98_80 =15'b0;

   // m98_81 = W*in
   wire signed [14:0] m98_81;
   assign m98_81 =15'b0;

   // m98_82 = W*in
   wire signed [14:0] m98_82;
   assign m98_82 =15'b0;

   // m98_83 = W*in
   wire signed [14:0] m98_83;
   assign m98_83 =15'b0;

   // m98_84 = W*in
   wire signed [14:0] m98_84;
   assign m98_84 =15'b0;

   // m98_85 = W*in
   wire signed [14:0] m98_85;
   assign m98_85 =15'b0;

   // m98_86 = W*in
   wire signed [14:0] m98_86;
   assign m98_86 =15'b0;

   // m98_87 = W*in
   wire signed [14:0] m98_87;
   assign m98_87 =15'b0;

   // m98_88 = W*in
   wire signed [14:0] m98_88;
   assign m98_88 =15'b0;

   // m98_89 = W*in
   wire signed [14:0] m98_89;
   assign m98_89 =15'b0;

   // m98_90 = W*in
   wire signed [14:0] m98_90;
   assign m98_90 =15'b0;

   // m98_91 = W*in
   wire signed [14:0] m98_91;
   assign m98_91 ={ {3{neg98[14]}} , neg98[14:3] };

   // m98_92 = W*in
   wire signed [14:0] m98_92;
   assign m98_92 =15'b0;

   // m98_93 = W*in
   wire signed [14:0] m98_93;
   assign m98_93 =15'b0;

   // m98_94 = W*in
   wire signed [14:0] m98_94;
   assign m98_94 ={ {4{neg98[14]}} , neg98[14:4] };

   // m98_95 = W*in
   wire signed [14:0] m98_95;
   assign m98_95 =15'b0;

   // m98_96 = W*in
   wire signed [14:0] m98_96;
   assign m98_96 =15'b0;

   // m98_97 = W*in
   wire signed [14:0] m98_97;
   assign m98_97 =15'b0;

   // m98_98 = W*in
   wire signed [14:0] m98_98;
   assign m98_98 =15'b0;

   // m98_99 = W*in
   wire signed [14:0] m98_99;
   assign m98_99 =15'b0;

   // m98_100 = W*in
   wire signed [14:0] m98_100;
   assign m98_100 =15'b0;

   // m99_1 = W*in
   wire signed [14:0] m99_1;
   assign m99_1 =15'b0;

   // m99_2 = W*in
   wire signed [14:0] m99_2;
   assign m99_2 =15'b0;

   // m99_3 = W*in
   wire signed [14:0] m99_3;
   assign m99_3 =15'b0;

   // m99_4 = W*in
   wire signed [14:0] m99_4;
   assign m99_4 =15'b0;

   // m99_5 = W*in
   wire signed [14:0] m99_5;
   assign m99_5 =15'b0;

   // m99_6 = W*in
   wire signed [14:0] m99_6;
   assign m99_6 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_7 = W*in
   wire signed [14:0] m99_7;
   assign m99_7 =15'b0;

   // m99_8 = W*in
   wire signed [14:0] m99_8;
   assign m99_8 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_9 = W*in
   wire signed [14:0] m99_9;
   assign m99_9 =15'b0;

   // m99_10 = W*in
   wire signed [14:0] m99_10;
   assign m99_10 =15'b0;

   // m99_11 = W*in
   wire signed [14:0] m99_11;
   assign m99_11 =15'b0;

   // m99_12 = W*in
   wire signed [14:0] m99_12;
   assign m99_12 =15'b0;

   // m99_13 = W*in
   wire signed [14:0] m99_13;
   assign m99_13 =15'b0;

   // m99_14 = W*in
   wire signed [14:0] m99_14;
   assign m99_14 =15'b0;

   // m99_15 = W*in
   wire signed [14:0] m99_15;
   assign m99_15 =15'b0;

   // m99_16 = W*in
   wire signed [14:0] m99_16;
   assign m99_16 =15'b0;

   // m99_17 = W*in
   wire signed [14:0] m99_17;
   assign m99_17 =15'b0;

   // m99_18 = W*in
   wire signed [14:0] m99_18;
   assign m99_18 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_19 = W*in
   wire signed [14:0] m99_19;
   assign m99_19 ={ {4{in99[14]}} , in99[14:4] };

   // m99_20 = W*in
   wire signed [14:0] m99_20;
   assign m99_20 =15'b0;

   // m99_21 = W*in
   wire signed [14:0] m99_21;
   assign m99_21 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_22 = W*in
   wire signed [14:0] m99_22;
   assign m99_22 =15'b0;

   // m99_23 = W*in
   wire signed [14:0] m99_23;
   assign m99_23 =15'b0;

   // m99_24 = W*in
   wire signed [14:0] m99_24;
   assign m99_24 =15'b0;

   // m99_25 = W*in
   wire signed [14:0] m99_25;
   assign m99_25 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_26 = W*in
   wire signed [14:0] m99_26;
   assign m99_26 =15'b0;

   // m99_27 = W*in
   wire signed [14:0] m99_27;
   assign m99_27 ={ {3{in99[14]}} , in99[14:3] };

   // m99_28 = W*in
   wire signed [14:0] m99_28;
   assign m99_28 =15'b0;

   // m99_29 = W*in
   wire signed [14:0] m99_29;
   assign m99_29 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_30 = W*in
   wire signed [14:0] m99_30;
   assign m99_30 =15'b0;

   // m99_31 = W*in
   wire signed [14:0] m99_31;
   assign m99_31 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_32 = W*in
   wire signed [14:0] m99_32;
   assign m99_32 ={ {4{in99[14]}} , in99[14:4] };

   // m99_33 = W*in
   wire signed [14:0] m99_33;
   assign m99_33 ={ {3{in99[14]}} , in99[14:3] };

   // m99_34 = W*in
   wire signed [14:0] m99_34;
   assign m99_34 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_35 = W*in
   wire signed [14:0] m99_35;
   assign m99_35 ={ {3{in99[14]}} , in99[14:3] };

   // m99_36 = W*in
   wire signed [14:0] m99_36;
   assign m99_36 =15'b0;

   // m99_37 = W*in
   wire signed [14:0] m99_37;
   assign m99_37 =15'b0;

   // m99_38 = W*in
   wire signed [14:0] m99_38;
   assign m99_38 =15'b0;

   // m99_39 = W*in
   wire signed [14:0] m99_39;
   assign m99_39 =15'b0;

   // m99_40 = W*in
   wire signed [14:0] m99_40;
   assign m99_40 ={ {3{in99[14]}} , in99[14:3] };

   // m99_41 = W*in
   wire signed [14:0] m99_41;
   assign m99_41 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_42 = W*in
   wire signed [14:0] m99_42;
   assign m99_42 ={ {3{in99[14]}} , in99[14:3] };

   // m99_43 = W*in
   wire signed [14:0] m99_43;
   assign m99_43 =15'b0;

   // m99_44 = W*in
   wire signed [14:0] m99_44;
   assign m99_44 =15'b0;

   // m99_45 = W*in
   wire signed [14:0] m99_45;
   assign m99_45 =15'b0;

   // m99_46 = W*in
   wire signed [14:0] m99_46;
   assign m99_46 =15'b0;

   // m99_47 = W*in
   wire signed [14:0] m99_47;
   assign m99_47 =15'b0;

   // m99_48 = W*in
   wire signed [14:0] m99_48;
   assign m99_48 ={ {4{in99[14]}} , in99[14:4] };

   // m99_49 = W*in
   wire signed [14:0] m99_49;
   assign m99_49 =15'b0;

   // m99_50 = W*in
   wire signed [14:0] m99_50;
   assign m99_50 =15'b0;

   // m99_51 = W*in
   wire signed [14:0] m99_51;
   assign m99_51 =15'b0;

   // m99_52 = W*in
   wire signed [14:0] m99_52;
   assign m99_52 =15'b0;

   // m99_53 = W*in
   wire signed [14:0] m99_53;
   assign m99_53 =15'b0;

   // m99_54 = W*in
   wire signed [14:0] m99_54;
   assign m99_54 =15'b0;

   // m99_55 = W*in
   wire signed [14:0] m99_55;
   assign m99_55 =15'b0;

   // m99_56 = W*in
   wire signed [14:0] m99_56;
   assign m99_56 =15'b0;

   // m99_57 = W*in
   wire signed [14:0] m99_57;
   assign m99_57 ={ {4{in99[14]}} , in99[14:4] };

   // m99_58 = W*in
   wire signed [14:0] m99_58;
   assign m99_58 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_59 = W*in
   wire signed [14:0] m99_59;
   assign m99_59 =15'b0;

   // m99_60 = W*in
   wire signed [14:0] m99_60;
   assign m99_60 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_61 = W*in
   wire signed [14:0] m99_61;
   assign m99_61 =15'b0;

   // m99_62 = W*in
   wire signed [14:0] m99_62;
   assign m99_62 =15'b0;

   // m99_63 = W*in
   wire signed [14:0] m99_63;
   assign m99_63 =15'b0;

   // m99_64 = W*in
   wire signed [14:0] m99_64;
   assign m99_64 =15'b0;

   // m99_65 = W*in
   wire signed [14:0] m99_65;
   assign m99_65 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_66 = W*in
   wire signed [14:0] m99_66;
   assign m99_66 =15'b0;

   // m99_67 = W*in
   wire signed [14:0] m99_67;
   assign m99_67 =15'b0;

   // m99_68 = W*in
   wire signed [14:0] m99_68;
   assign m99_68 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_69 = W*in
   wire signed [14:0] m99_69;
   assign m99_69 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_70 = W*in
   wire signed [14:0] m99_70;
   assign m99_70 ={ {4{in99[14]}} , in99[14:4] };

   // m99_71 = W*in
   wire signed [14:0] m99_71;
   assign m99_71 =15'b0;

   // m99_72 = W*in
   wire signed [14:0] m99_72;
   assign m99_72 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_73 = W*in
   wire signed [14:0] m99_73;
   assign m99_73 =15'b0;

   // m99_74 = W*in
   wire signed [14:0] m99_74;
   assign m99_74 =15'b0;

   // m99_75 = W*in
   wire signed [14:0] m99_75;
   assign m99_75 =15'b0;

   // m99_76 = W*in
   wire signed [14:0] m99_76;
   assign m99_76 =15'b0;

   // m99_77 = W*in
   wire signed [14:0] m99_77;
   assign m99_77 ={ {4{neg99[14]}} , neg99[14:4] };

   // m99_78 = W*in
   wire signed [14:0] m99_78;
   assign m99_78 =15'b0;

   // m99_79 = W*in
   wire signed [14:0] m99_79;
   assign m99_79 =15'b0;

   // m99_80 = W*in
   wire signed [14:0] m99_80;
   assign m99_80 =15'b0;

   // m99_81 = W*in
   wire signed [14:0] m99_81;
   assign m99_81 =15'b0;

   // m99_82 = W*in
   wire signed [14:0] m99_82;
   assign m99_82 =15'b0;

   // m99_83 = W*in
   wire signed [14:0] m99_83;
   assign m99_83 =15'b0;

   // m99_84 = W*in
   wire signed [14:0] m99_84;
   assign m99_84 =15'b0;

   // m99_85 = W*in
   wire signed [14:0] m99_85;
   assign m99_85 =15'b0;

   // m99_86 = W*in
   wire signed [14:0] m99_86;
   assign m99_86 =15'b0;

   // m99_87 = W*in
   wire signed [14:0] m99_87;
   assign m99_87 =15'b0;

   // m99_88 = W*in
   wire signed [14:0] m99_88;
   assign m99_88 =15'b0;

   // m99_89 = W*in
   wire signed [14:0] m99_89;
   assign m99_89 =15'b0;

   // m99_90 = W*in
   wire signed [14:0] m99_90;
   assign m99_90 =15'b0;

   // m99_91 = W*in
   wire signed [14:0] m99_91;
   assign m99_91 =15'b0;

   // m99_92 = W*in
   wire signed [14:0] m99_92;
   assign m99_92 =15'b0;

   // m99_93 = W*in
   wire signed [14:0] m99_93;
   assign m99_93 =15'b0;

   // m99_94 = W*in
   wire signed [14:0] m99_94;
   assign m99_94 =15'b0;

   // m99_95 = W*in
   wire signed [14:0] m99_95;
   assign m99_95 =15'b0;

   // m99_96 = W*in
   wire signed [14:0] m99_96;
   assign m99_96 ={ {3{neg99[14]}} , neg99[14:3] };

   // m99_97 = W*in
   wire signed [14:0] m99_97;
   assign m99_97 =15'b0;

   // m99_98 = W*in
   wire signed [14:0] m99_98;
   assign m99_98 =15'b0;

   // m99_99 = W*in
   wire signed [14:0] m99_99;
   assign m99_99 =15'b0;

   // m99_100 = W*in
   wire signed [14:0] m99_100;
   assign m99_100 =15'b0;

   // m100_1 = W*in
   wire signed [14:0] m100_1;
   assign m100_1 =15'b0;

   // m100_2 = W*in
   wire signed [14:0] m100_2;
   assign m100_2 =15'b0;

   // m100_3 = W*in
   wire signed [14:0] m100_3;
   assign m100_3 ={ {3{in100[14]}} , in100[14:3] };

   // m100_4 = W*in
   wire signed [14:0] m100_4;
   assign m100_4 ={ {3{in100[14]}} , in100[14:3] };

   // m100_5 = W*in
   wire signed [14:0] m100_5;
   assign m100_5 =15'b0;

   // m100_6 = W*in
   wire signed [14:0] m100_6;
   assign m100_6 ={ {4{neg100[14]}} , neg100[14:4] };

   // m100_7 = W*in
   wire signed [14:0] m100_7;
   assign m100_7 ={ {4{neg100[14]}} , neg100[14:4] };

   // m100_8 = W*in
   wire signed [14:0] m100_8;
   assign m100_8 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_9 = W*in
   wire signed [14:0] m100_9;
   assign m100_9 =15'b0;

   // m100_10 = W*in
   wire signed [14:0] m100_10;
   assign m100_10 =15'b0;

   // m100_11 = W*in
   wire signed [14:0] m100_11;
   assign m100_11 =15'b0;

   // m100_12 = W*in
   wire signed [14:0] m100_12;
   assign m100_12 =15'b0;

   // m100_13 = W*in
   wire signed [14:0] m100_13;
   assign m100_13 ={ {3{in100[14]}} , in100[14:3] };

   // m100_14 = W*in
   wire signed [14:0] m100_14;
   assign m100_14 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_15 = W*in
   wire signed [14:0] m100_15;
   assign m100_15 =15'b0;

   // m100_16 = W*in
   wire signed [14:0] m100_16;
   assign m100_16 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_17 = W*in
   wire signed [14:0] m100_17;
   assign m100_17 =15'b0;

   // m100_18 = W*in
   wire signed [14:0] m100_18;
   assign m100_18 =15'b0;

   // m100_19 = W*in
   wire signed [14:0] m100_19;
   assign m100_19 =15'b0;

   // m100_20 = W*in
   wire signed [14:0] m100_20;
   assign m100_20 =15'b0;

   // m100_21 = W*in
   wire signed [14:0] m100_21;
   assign m100_21 =15'b0;

   // m100_22 = W*in
   wire signed [14:0] m100_22;
   assign m100_22 =15'b0;

   // m100_23 = W*in
   wire signed [14:0] m100_23;
   assign m100_23 =15'b0;

   // m100_24 = W*in
   wire signed [14:0] m100_24;
   assign m100_24 =15'b0;

   // m100_25 = W*in
   wire signed [14:0] m100_25;
   assign m100_25 =15'b0;

   // m100_26 = W*in
   wire signed [14:0] m100_26;
   assign m100_26 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_27 = W*in
   wire signed [14:0] m100_27;
   assign m100_27 =15'b0;

   // m100_28 = W*in
   wire signed [14:0] m100_28;
   assign m100_28 =15'b0;

   // m100_29 = W*in
   wire signed [14:0] m100_29;
   assign m100_29 =15'b0;

   // m100_30 = W*in
   wire signed [14:0] m100_30;
   assign m100_30 =15'b0;

   // m100_31 = W*in
   wire signed [14:0] m100_31;
   assign m100_31 =15'b0;

   // m100_32 = W*in
   wire signed [14:0] m100_32;
   assign m100_32 =15'b0;

   // m100_33 = W*in
   wire signed [14:0] m100_33;
   assign m100_33 ={ {4{neg100[14]}} , neg100[14:4] };

   // m100_34 = W*in
   wire signed [14:0] m100_34;
   assign m100_34 =15'b0;

   // m100_35 = W*in
   wire signed [14:0] m100_35;
   assign m100_35 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_36 = W*in
   wire signed [14:0] m100_36;
   assign m100_36 =15'b0;

   // m100_37 = W*in
   wire signed [14:0] m100_37;
   assign m100_37 =15'b0;

   // m100_38 = W*in
   wire signed [14:0] m100_38;
   assign m100_38 =15'b0;

   // m100_39 = W*in
   wire signed [14:0] m100_39;
   assign m100_39 =15'b0;

   // m100_40 = W*in
   wire signed [14:0] m100_40;
   assign m100_40 =15'b0;

   // m100_41 = W*in
   wire signed [14:0] m100_41;
   assign m100_41 ={ {4{in100[14]}} , in100[14:4] };

   // m100_42 = W*in
   wire signed [14:0] m100_42;
   assign m100_42 =15'b0;

   // m100_43 = W*in
   wire signed [14:0] m100_43;
   assign m100_43 =15'b0;

   // m100_44 = W*in
   wire signed [14:0] m100_44;
   assign m100_44 =15'b0;

   // m100_45 = W*in
   wire signed [14:0] m100_45;
   assign m100_45 =15'b0;

   // m100_46 = W*in
   wire signed [14:0] m100_46;
   assign m100_46 ={ {4{neg100[14]}} , neg100[14:4] };

   // m100_47 = W*in
   wire signed [14:0] m100_47;
   assign m100_47 =15'b0;

   // m100_48 = W*in
   wire signed [14:0] m100_48;
   assign m100_48 =15'b0;

   // m100_49 = W*in
   wire signed [14:0] m100_49;
   assign m100_49 =15'b0;

   // m100_50 = W*in
   wire signed [14:0] m100_50;
   assign m100_50 =15'b0;

   // m100_51 = W*in
   wire signed [14:0] m100_51;
   assign m100_51 =15'b0;

   // m100_52 = W*in
   wire signed [14:0] m100_52;
   assign m100_52 =15'b0;

   // m100_53 = W*in
   wire signed [14:0] m100_53;
   assign m100_53 =15'b0;

   // m100_54 = W*in
   wire signed [14:0] m100_54;
   assign m100_54 =15'b0;

   // m100_55 = W*in
   wire signed [14:0] m100_55;
   assign m100_55 =15'b0;

   // m100_56 = W*in
   wire signed [14:0] m100_56;
   assign m100_56 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_57 = W*in
   wire signed [14:0] m100_57;
   assign m100_57 =15'b0;

   // m100_58 = W*in
   wire signed [14:0] m100_58;
   assign m100_58 =15'b0;

   // m100_59 = W*in
   wire signed [14:0] m100_59;
   assign m100_59 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_60 = W*in
   wire signed [14:0] m100_60;
   assign m100_60 =15'b0;

   // m100_61 = W*in
   wire signed [14:0] m100_61;
   assign m100_61 =15'b0;

   // m100_62 = W*in
   wire signed [14:0] m100_62;
   assign m100_62 =15'b0;

   // m100_63 = W*in
   wire signed [14:0] m100_63;
   assign m100_63 =15'b0;

   // m100_64 = W*in
   wire signed [14:0] m100_64;
   assign m100_64 =15'b0;

   // m100_65 = W*in
   wire signed [14:0] m100_65;
   assign m100_65 =15'b0;

   // m100_66 = W*in
   wire signed [14:0] m100_66;
   assign m100_66 =15'b0;

   // m100_67 = W*in
   wire signed [14:0] m100_67;
   assign m100_67 =15'b0;

   // m100_68 = W*in
   wire signed [14:0] m100_68;
   assign m100_68 ={ {3{in100[14]}} , in100[14:3] };

   // m100_69 = W*in
   wire signed [14:0] m100_69;
   assign m100_69 =15'b0;

   // m100_70 = W*in
   wire signed [14:0] m100_70;
   assign m100_70 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_71 = W*in
   wire signed [14:0] m100_71;
   assign m100_71 =15'b0;

   // m100_72 = W*in
   wire signed [14:0] m100_72;
   assign m100_72 ={ {3{in100[14]}} , in100[14:3] };

   // m100_73 = W*in
   wire signed [14:0] m100_73;
   assign m100_73 =15'b0;

   // m100_74 = W*in
   wire signed [14:0] m100_74;
   assign m100_74 =15'b0;

   // m100_75 = W*in
   wire signed [14:0] m100_75;
   assign m100_75 ={ {4{in100[14]}} , in100[14:4] };

   // m100_76 = W*in
   wire signed [14:0] m100_76;
   assign m100_76 =15'b0;

   // m100_77 = W*in
   wire signed [14:0] m100_77;
   assign m100_77 ={ {3{in100[14]}} , in100[14:3] };

   // m100_78 = W*in
   wire signed [14:0] m100_78;
   assign m100_78 =15'b0;

   // m100_79 = W*in
   wire signed [14:0] m100_79;
   assign m100_79 =15'b0;

   // m100_80 = W*in
   wire signed [14:0] m100_80;
   assign m100_80 =15'b0;

   // m100_81 = W*in
   wire signed [14:0] m100_81;
   assign m100_81 =15'b0;

   // m100_82 = W*in
   wire signed [14:0] m100_82;
   assign m100_82 =15'b0;

   // m100_83 = W*in
   wire signed [14:0] m100_83;
   assign m100_83 =15'b0;

   // m100_84 = W*in
   wire signed [14:0] m100_84;
   assign m100_84 =15'b0;

   // m100_85 = W*in
   wire signed [14:0] m100_85;
   assign m100_85 ={ {3{in100[14]}} , in100[14:3] };

   // m100_86 = W*in
   wire signed [14:0] m100_86;
   assign m100_86 =15'b0;

   // m100_87 = W*in
   wire signed [14:0] m100_87;
   assign m100_87 =15'b0;

   // m100_88 = W*in
   wire signed [14:0] m100_88;
   assign m100_88 =15'b0;

   // m100_89 = W*in
   wire signed [14:0] m100_89;
   assign m100_89 =15'b0;

   // m100_90 = W*in
   wire signed [14:0] m100_90;
   assign m100_90 =15'b0;

   // m100_91 = W*in
   wire signed [14:0] m100_91;
   assign m100_91 =15'b0;

   // m100_92 = W*in
   wire signed [14:0] m100_92;
   assign m100_92 =15'b0;

   // m100_93 = W*in
   wire signed [14:0] m100_93;
   assign m100_93 =15'b0;

   // m100_94 = W*in
   wire signed [14:0] m100_94;
   assign m100_94 ={ {3{neg100[14]}} , neg100[14:3] };

   // m100_95 = W*in
   wire signed [14:0] m100_95;
   assign m100_95 =15'b0;

   // m100_96 = W*in
   wire signed [14:0] m100_96;
   assign m100_96 ={ {4{in100[14]}} , in100[14:4] };

   // m100_97 = W*in
   wire signed [14:0] m100_97;
   assign m100_97 =15'b0;

   // m100_98 = W*in
   wire signed [14:0] m100_98;
   assign m100_98 =15'b0;

   // m100_99 = W*in
   wire signed [14:0] m100_99;
   assign m100_99 =15'b0;

   // m100_100 = W*in
   wire signed [14:0] m100_100;
   assign m100_100 =15'b0;

   // m101_1 = W*in
   wire signed [14:0] m101_1;
   assign m101_1 =15'b0;

   // m101_2 = W*in
   wire signed [14:0] m101_2;
   assign m101_2 =15'b0;

   // m101_3 = W*in
   wire signed [14:0] m101_3;
   assign m101_3 ={ {4{neg101[14]}} , neg101[14:4] };

   // m101_4 = W*in
   wire signed [14:0] m101_4;
   assign m101_4 =15'b0;

   // m101_5 = W*in
   wire signed [14:0] m101_5;
   assign m101_5 =15'b0;

   // m101_6 = W*in
   wire signed [14:0] m101_6;
   assign m101_6 =15'b0;

   // m101_7 = W*in
   wire signed [14:0] m101_7;
   assign m101_7 =15'b0;

   // m101_8 = W*in
   wire signed [14:0] m101_8;
   assign m101_8 =15'b0;

   // m101_9 = W*in
   wire signed [14:0] m101_9;
   assign m101_9 =15'b0;

   // m101_10 = W*in
   wire signed [14:0] m101_10;
   assign m101_10 =15'b0;

   // m101_11 = W*in
   wire signed [14:0] m101_11;
   assign m101_11 =15'b0;

   // m101_12 = W*in
   wire signed [14:0] m101_12;
   assign m101_12 =15'b0;

   // m101_13 = W*in
   wire signed [14:0] m101_13;
   assign m101_13 =15'b0;

   // m101_14 = W*in
   wire signed [14:0] m101_14;
   assign m101_14 =15'b0;

   // m101_15 = W*in
   wire signed [14:0] m101_15;
   assign m101_15 =15'b0;

   // m101_16 = W*in
   wire signed [14:0] m101_16;
   assign m101_16 =15'b0;

   // m101_17 = W*in
   wire signed [14:0] m101_17;
   assign m101_17 ={ {4{neg101[14]}} , neg101[14:4] };

   // m101_18 = W*in
   wire signed [14:0] m101_18;
   assign m101_18 =15'b0;

   // m101_19 = W*in
   wire signed [14:0] m101_19;
   assign m101_19 =15'b0;

   // m101_20 = W*in
   wire signed [14:0] m101_20;
   assign m101_20 ={ {4{in101[14]}} , in101[14:4] };

   // m101_21 = W*in
   wire signed [14:0] m101_21;
   assign m101_21 =15'b0;

   // m101_22 = W*in
   wire signed [14:0] m101_22;
   assign m101_22 ={ {4{in101[14]}} , in101[14:4] };

   // m101_23 = W*in
   wire signed [14:0] m101_23;
   assign m101_23 =15'b0;

   // m101_24 = W*in
   wire signed [14:0] m101_24;
   assign m101_24 ={ {4{in101[14]}} , in101[14:4] };

   // m101_25 = W*in
   wire signed [14:0] m101_25;
   assign m101_25 =15'b0;

   // m101_26 = W*in
   wire signed [14:0] m101_26;
   assign m101_26 =15'b0;

   // m101_27 = W*in
   wire signed [14:0] m101_27;
   assign m101_27 =15'b0;

   // m101_28 = W*in
   wire signed [14:0] m101_28;
   assign m101_28 =15'b0;

   // m101_29 = W*in
   wire signed [14:0] m101_29;
   assign m101_29 =15'b0;

   // m101_30 = W*in
   wire signed [14:0] m101_30;
   assign m101_30 =15'b0;

   // m101_31 = W*in
   wire signed [14:0] m101_31;
   assign m101_31 =15'b0;

   // m101_32 = W*in
   wire signed [14:0] m101_32;
   assign m101_32 =15'b0;

   // m101_33 = W*in
   wire signed [14:0] m101_33;
   assign m101_33 ={ {4{neg101[14]}} , neg101[14:4] };

   // m101_34 = W*in
   wire signed [14:0] m101_34;
   assign m101_34 =15'b0;

   // m101_35 = W*in
   wire signed [14:0] m101_35;
   assign m101_35 =15'b0;

   // m101_36 = W*in
   wire signed [14:0] m101_36;
   assign m101_36 =15'b0;

   // m101_37 = W*in
   wire signed [14:0] m101_37;
   assign m101_37 =15'b0;

   // m101_38 = W*in
   wire signed [14:0] m101_38;
   assign m101_38 =15'b0;

   // m101_39 = W*in
   wire signed [14:0] m101_39;
   assign m101_39 =15'b0;

   // m101_40 = W*in
   wire signed [14:0] m101_40;
   assign m101_40 ={ {4{neg101[14]}} , neg101[14:4] };

   // m101_41 = W*in
   wire signed [14:0] m101_41;
   assign m101_41 =15'b0;

   // m101_42 = W*in
   wire signed [14:0] m101_42;
   assign m101_42 =15'b0;

   // m101_43 = W*in
   wire signed [14:0] m101_43;
   assign m101_43 =15'b0;

   // m101_44 = W*in
   wire signed [14:0] m101_44;
   assign m101_44 =15'b0;

   // m101_45 = W*in
   wire signed [14:0] m101_45;
   assign m101_45 =15'b0;

   // m101_46 = W*in
   wire signed [14:0] m101_46;
   assign m101_46 =15'b0;

   // m101_47 = W*in
   wire signed [14:0] m101_47;
   assign m101_47 ={ {4{in101[14]}} , in101[14:4] };

   // m101_48 = W*in
   wire signed [14:0] m101_48;
   assign m101_48 =15'b0;

   // m101_49 = W*in
   wire signed [14:0] m101_49;
   assign m101_49 =15'b0;

   // m101_50 = W*in
   wire signed [14:0] m101_50;
   assign m101_50 =15'b0;

   // m101_51 = W*in
   wire signed [14:0] m101_51;
   assign m101_51 =15'b0;

   // m101_52 = W*in
   wire signed [14:0] m101_52;
   assign m101_52 =15'b0;

   // m101_53 = W*in
   wire signed [14:0] m101_53;
   assign m101_53 =15'b0;

   // m101_54 = W*in
   wire signed [14:0] m101_54;
   assign m101_54 =15'b0;

   // m101_55 = W*in
   wire signed [14:0] m101_55;
   assign m101_55 =15'b0;

   // m101_56 = W*in
   wire signed [14:0] m101_56;
   assign m101_56 =15'b0;

   // m101_57 = W*in
   wire signed [14:0] m101_57;
   assign m101_57 =15'b0;

   // m101_58 = W*in
   wire signed [14:0] m101_58;
   assign m101_58 ={ {4{in101[14]}} , in101[14:4] };

   // m101_59 = W*in
   wire signed [14:0] m101_59;
   assign m101_59 =15'b0;

   // m101_60 = W*in
   wire signed [14:0] m101_60;
   assign m101_60 =15'b0;

   // m101_61 = W*in
   wire signed [14:0] m101_61;
   assign m101_61 ={ {3{in101[14]}} , in101[14:3] };

   // m101_62 = W*in
   wire signed [14:0] m101_62;
   assign m101_62 ={ {3{in101[14]}} , in101[14:3] };

   // m101_63 = W*in
   wire signed [14:0] m101_63;
   assign m101_63 =15'b0;

   // m101_64 = W*in
   wire signed [14:0] m101_64;
   assign m101_64 =15'b0;

   // m101_65 = W*in
   wire signed [14:0] m101_65;
   assign m101_65 =15'b0;

   // m101_66 = W*in
   wire signed [14:0] m101_66;
   assign m101_66 ={ {3{neg101[14]}} , neg101[14:3] };

   // m101_67 = W*in
   wire signed [14:0] m101_67;
   assign m101_67 =15'b0;

   // m101_68 = W*in
   wire signed [14:0] m101_68;
   assign m101_68 =15'b0;

   // m101_69 = W*in
   wire signed [14:0] m101_69;
   assign m101_69 =15'b0;

   // m101_70 = W*in
   wire signed [14:0] m101_70;
   assign m101_70 =15'b0;

   // m101_71 = W*in
   wire signed [14:0] m101_71;
   assign m101_71 =15'b0;

   // m101_72 = W*in
   wire signed [14:0] m101_72;
   assign m101_72 ={ {3{in101[14]}} , in101[14:3] };

   // m101_73 = W*in
   wire signed [14:0] m101_73;
   assign m101_73 =15'b0;

   // m101_74 = W*in
   wire signed [14:0] m101_74;
   assign m101_74 =15'b0;

   // m101_75 = W*in
   wire signed [14:0] m101_75;
   assign m101_75 =15'b0;

   // m101_76 = W*in
   wire signed [14:0] m101_76;
   assign m101_76 ={ {3{neg101[14]}} , neg101[14:3] };

   // m101_77 = W*in
   wire signed [14:0] m101_77;
   assign m101_77 =15'b0;

   // m101_78 = W*in
   wire signed [14:0] m101_78;
   assign m101_78 =15'b0;

   // m101_79 = W*in
   wire signed [14:0] m101_79;
   assign m101_79 =15'b0;

   // m101_80 = W*in
   wire signed [14:0] m101_80;
   assign m101_80 =15'b0;

   // m101_81 = W*in
   wire signed [14:0] m101_81;
   assign m101_81 =15'b0;

   // m101_82 = W*in
   wire signed [14:0] m101_82;
   assign m101_82 =15'b0;

   // m101_83 = W*in
   wire signed [14:0] m101_83;
   assign m101_83 =15'b0;

   // m101_84 = W*in
   wire signed [14:0] m101_84;
   assign m101_84 =15'b0;

   // m101_85 = W*in
   wire signed [14:0] m101_85;
   assign m101_85 ={ {3{neg101[14]}} , neg101[14:3] };

   // m101_86 = W*in
   wire signed [14:0] m101_86;
   assign m101_86 =15'b0;

   // m101_87 = W*in
   wire signed [14:0] m101_87;
   assign m101_87 =15'b0;

   // m101_88 = W*in
   wire signed [14:0] m101_88;
   assign m101_88 =15'b0;

   // m101_89 = W*in
   wire signed [14:0] m101_89;
   assign m101_89 =15'b0;

   // m101_90 = W*in
   wire signed [14:0] m101_90;
   assign m101_90 =15'b0;

   // m101_91 = W*in
   wire signed [14:0] m101_91;
   assign m101_91 =15'b0;

   // m101_92 = W*in
   wire signed [14:0] m101_92;
   assign m101_92 =15'b0;

   // m101_93 = W*in
   wire signed [14:0] m101_93;
   assign m101_93 =15'b0;

   // m101_94 = W*in
   wire signed [14:0] m101_94;
   assign m101_94 =15'b0;

   // m101_95 = W*in
   wire signed [14:0] m101_95;
   assign m101_95 ={ {3{neg101[14]}} , neg101[14:3] };

   // m101_96 = W*in
   wire signed [14:0] m101_96;
   assign m101_96 =15'b0;

   // m101_97 = W*in
   wire signed [14:0] m101_97;
   assign m101_97 =15'b0;

   // m101_98 = W*in
   wire signed [14:0] m101_98;
   assign m101_98 =15'b0;

   // m101_99 = W*in
   wire signed [14:0] m101_99;
   assign m101_99 =15'b0;

   // m101_100 = W*in
   wire signed [14:0] m101_100;
   assign m101_100 =15'b0;

   // m102_1 = W*in
   wire signed [14:0] m102_1;
   assign m102_1 =15'b0;

   // m102_2 = W*in
   wire signed [14:0] m102_2;
   assign m102_2 =15'b0;

   // m102_3 = W*in
   wire signed [14:0] m102_3;
   assign m102_3 =15'b0;

   // m102_4 = W*in
   wire signed [14:0] m102_4;
   assign m102_4 =15'b0;

   // m102_5 = W*in
   wire signed [14:0] m102_5;
   assign m102_5 =15'b0;

   // m102_6 = W*in
   wire signed [14:0] m102_6;
   assign m102_6 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_7 = W*in
   wire signed [14:0] m102_7;
   assign m102_7 =15'b0;

   // m102_8 = W*in
   wire signed [14:0] m102_8;
   assign m102_8 =15'b0;

   // m102_9 = W*in
   wire signed [14:0] m102_9;
   assign m102_9 =15'b0;

   // m102_10 = W*in
   wire signed [14:0] m102_10;
   assign m102_10 =15'b0;

   // m102_11 = W*in
   wire signed [14:0] m102_11;
   assign m102_11 =15'b0;

   // m102_12 = W*in
   wire signed [14:0] m102_12;
   assign m102_12 =15'b0;

   // m102_13 = W*in
   wire signed [14:0] m102_13;
   assign m102_13 =15'b0;

   // m102_14 = W*in
   wire signed [14:0] m102_14;
   assign m102_14 =15'b0;

   // m102_15 = W*in
   wire signed [14:0] m102_15;
   assign m102_15 =15'b0;

   // m102_16 = W*in
   wire signed [14:0] m102_16;
   assign m102_16 =15'b0;

   // m102_17 = W*in
   wire signed [14:0] m102_17;
   assign m102_17 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_18 = W*in
   wire signed [14:0] m102_18;
   assign m102_18 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_19 = W*in
   wire signed [14:0] m102_19;
   assign m102_19 ={ {4{in102[14]}} , in102[14:4] };

   // m102_20 = W*in
   wire signed [14:0] m102_20;
   assign m102_20 =15'b0;

   // m102_21 = W*in
   wire signed [14:0] m102_21;
   assign m102_21 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_22 = W*in
   wire signed [14:0] m102_22;
   assign m102_22 ={ {4{in102[14]}} , in102[14:4] };

   // m102_23 = W*in
   wire signed [14:0] m102_23;
   assign m102_23 =15'b0;

   // m102_24 = W*in
   wire signed [14:0] m102_24;
   assign m102_24 =15'b0;

   // m102_25 = W*in
   wire signed [14:0] m102_25;
   assign m102_25 =15'b0;

   // m102_26 = W*in
   wire signed [14:0] m102_26;
   assign m102_26 ={ {4{in102[14]}} , in102[14:4] };

   // m102_27 = W*in
   wire signed [14:0] m102_27;
   assign m102_27 ={ {3{in102[14]}} , in102[14:3] };

   // m102_28 = W*in
   wire signed [14:0] m102_28;
   assign m102_28 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_29 = W*in
   wire signed [14:0] m102_29;
   assign m102_29 =15'b0;

   // m102_30 = W*in
   wire signed [14:0] m102_30;
   assign m102_30 =15'b0;

   // m102_31 = W*in
   wire signed [14:0] m102_31;
   assign m102_31 =15'b0;

   // m102_32 = W*in
   wire signed [14:0] m102_32;
   assign m102_32 ={ {4{in102[14]}} , in102[14:4] };

   // m102_33 = W*in
   wire signed [14:0] m102_33;
   assign m102_33 ={ {4{in102[14]}} , in102[14:4] };

   // m102_34 = W*in
   wire signed [14:0] m102_34;
   assign m102_34 =15'b0;

   // m102_35 = W*in
   wire signed [14:0] m102_35;
   assign m102_35 =15'b0;

   // m102_36 = W*in
   wire signed [14:0] m102_36;
   assign m102_36 =15'b0;

   // m102_37 = W*in
   wire signed [14:0] m102_37;
   assign m102_37 =15'b0;

   // m102_38 = W*in
   wire signed [14:0] m102_38;
   assign m102_38 =15'b0;

   // m102_39 = W*in
   wire signed [14:0] m102_39;
   assign m102_39 =15'b0;

   // m102_40 = W*in
   wire signed [14:0] m102_40;
   assign m102_40 =15'b0;

   // m102_41 = W*in
   wire signed [14:0] m102_41;
   assign m102_41 ={ {3{neg102[14]}} , neg102[14:3] };

   // m102_42 = W*in
   wire signed [14:0] m102_42;
   assign m102_42 =15'b0;

   // m102_43 = W*in
   wire signed [14:0] m102_43;
   assign m102_43 ={ {3{in102[14]}} , in102[14:3] };

   // m102_44 = W*in
   wire signed [14:0] m102_44;
   assign m102_44 =15'b0;

   // m102_45 = W*in
   wire signed [14:0] m102_45;
   assign m102_45 =15'b0;

   // m102_46 = W*in
   wire signed [14:0] m102_46;
   assign m102_46 =15'b0;

   // m102_47 = W*in
   wire signed [14:0] m102_47;
   assign m102_47 =15'b0;

   // m102_48 = W*in
   wire signed [14:0] m102_48;
   assign m102_48 =15'b0;

   // m102_49 = W*in
   wire signed [14:0] m102_49;
   assign m102_49 =15'b0;

   // m102_50 = W*in
   wire signed [14:0] m102_50;
   assign m102_50 =15'b0;

   // m102_51 = W*in
   wire signed [14:0] m102_51;
   assign m102_51 =15'b0;

   // m102_52 = W*in
   wire signed [14:0] m102_52;
   assign m102_52 =15'b0;

   // m102_53 = W*in
   wire signed [14:0] m102_53;
   assign m102_53 =15'b0;

   // m102_54 = W*in
   wire signed [14:0] m102_54;
   assign m102_54 =15'b0;

   // m102_55 = W*in
   wire signed [14:0] m102_55;
   assign m102_55 =15'b0;

   // m102_56 = W*in
   wire signed [14:0] m102_56;
   assign m102_56 =15'b0;

   // m102_57 = W*in
   wire signed [14:0] m102_57;
   assign m102_57 ={ {4{in102[14]}} , in102[14:4] };

   // m102_58 = W*in
   wire signed [14:0] m102_58;
   assign m102_58 =15'b0;

   // m102_59 = W*in
   wire signed [14:0] m102_59;
   assign m102_59 ={ {4{in102[14]}} , in102[14:4] };

   // m102_60 = W*in
   wire signed [14:0] m102_60;
   assign m102_60 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_61 = W*in
   wire signed [14:0] m102_61;
   assign m102_61 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_62 = W*in
   wire signed [14:0] m102_62;
   assign m102_62 =15'b0;

   // m102_63 = W*in
   wire signed [14:0] m102_63;
   assign m102_63 =15'b0;

   // m102_64 = W*in
   wire signed [14:0] m102_64;
   assign m102_64 =15'b0;

   // m102_65 = W*in
   wire signed [14:0] m102_65;
   assign m102_65 ={ {4{in102[14]}} , in102[14:4] };

   // m102_66 = W*in
   wire signed [14:0] m102_66;
   assign m102_66 ={ {4{in102[14]}} , in102[14:4] };

   // m102_67 = W*in
   wire signed [14:0] m102_67;
   assign m102_67 =15'b0;

   // m102_68 = W*in
   wire signed [14:0] m102_68;
   assign m102_68 ={ {4{neg102[14]}} , neg102[14:4] };

   // m102_69 = W*in
   wire signed [14:0] m102_69;
   assign m102_69 =15'b0;

   // m102_70 = W*in
   wire signed [14:0] m102_70;
   assign m102_70 =15'b0;

   // m102_71 = W*in
   wire signed [14:0] m102_71;
   assign m102_71 =15'b0;

   // m102_72 = W*in
   wire signed [14:0] m102_72;
   assign m102_72 =15'b0;

   // m102_73 = W*in
   wire signed [14:0] m102_73;
   assign m102_73 =15'b0;

   // m102_74 = W*in
   wire signed [14:0] m102_74;
   assign m102_74 =15'b0;

   // m102_75 = W*in
   wire signed [14:0] m102_75;
   assign m102_75 =15'b0;

   // m102_76 = W*in
   wire signed [14:0] m102_76;
   assign m102_76 =15'b0;

   // m102_77 = W*in
   wire signed [14:0] m102_77;
   assign m102_77 =15'b0;

   // m102_78 = W*in
   wire signed [14:0] m102_78;
   assign m102_78 =15'b0;

   // m102_79 = W*in
   wire signed [14:0] m102_79;
   assign m102_79 =15'b0;

   // m102_80 = W*in
   wire signed [14:0] m102_80;
   assign m102_80 =15'b0;

   // m102_81 = W*in
   wire signed [14:0] m102_81;
   assign m102_81 =15'b0;

   // m102_82 = W*in
   wire signed [14:0] m102_82;
   assign m102_82 =15'b0;

   // m102_83 = W*in
   wire signed [14:0] m102_83;
   assign m102_83 =15'b0;

   // m102_84 = W*in
   wire signed [14:0] m102_84;
   assign m102_84 =15'b0;

   // m102_85 = W*in
   wire signed [14:0] m102_85;
   assign m102_85 =15'b0;

   // m102_86 = W*in
   wire signed [14:0] m102_86;
   assign m102_86 =15'b0;

   // m102_87 = W*in
   wire signed [14:0] m102_87;
   assign m102_87 =15'b0;

   // m102_88 = W*in
   wire signed [14:0] m102_88;
   assign m102_88 =15'b0;

   // m102_89 = W*in
   wire signed [14:0] m102_89;
   assign m102_89 =15'b0;

   // m102_90 = W*in
   wire signed [14:0] m102_90;
   assign m102_90 =15'b0;

   // m102_91 = W*in
   wire signed [14:0] m102_91;
   assign m102_91 =15'b0;

   // m102_92 = W*in
   wire signed [14:0] m102_92;
   assign m102_92 =15'b0;

   // m102_93 = W*in
   wire signed [14:0] m102_93;
   assign m102_93 =15'b0;

   // m102_94 = W*in
   wire signed [14:0] m102_94;
   assign m102_94 =15'b0;

   // m102_95 = W*in
   wire signed [14:0] m102_95;
   assign m102_95 =15'b0;

   // m102_96 = W*in
   wire signed [14:0] m102_96;
   assign m102_96 ={ {3{neg102[14]}} , neg102[14:3] };

   // m102_97 = W*in
   wire signed [14:0] m102_97;
   assign m102_97 ={ {3{in102[14]}} , in102[14:3] };

   // m102_98 = W*in
   wire signed [14:0] m102_98;
   assign m102_98 =15'b0;

   // m102_99 = W*in
   wire signed [14:0] m102_99;
   assign m102_99 =15'b0;

   // m102_100 = W*in
   wire signed [14:0] m102_100;
   assign m102_100 =15'b0;

   // m103_1 = W*in
   wire signed [14:0] m103_1;
   assign m103_1 =15'b0;

   // m103_2 = W*in
   wire signed [14:0] m103_2;
   assign m103_2 =15'b0;

   // m103_3 = W*in
   wire signed [14:0] m103_3;
   assign m103_3 =15'b0;

   // m103_4 = W*in
   wire signed [14:0] m103_4;
   assign m103_4 ={ {3{in103[14]}} , in103[14:3] };

   // m103_5 = W*in
   wire signed [14:0] m103_5;
   assign m103_5 =15'b0;

   // m103_6 = W*in
   wire signed [14:0] m103_6;
   assign m103_6 ={ {4{neg103[14]}} , neg103[14:4] };

   // m103_7 = W*in
   wire signed [14:0] m103_7;
   assign m103_7 =15'b0;

   // m103_8 = W*in
   wire signed [14:0] m103_8;
   assign m103_8 =15'b0;

   // m103_9 = W*in
   wire signed [14:0] m103_9;
   assign m103_9 =15'b0;

   // m103_10 = W*in
   wire signed [14:0] m103_10;
   assign m103_10 =15'b0;

   // m103_11 = W*in
   wire signed [14:0] m103_11;
   assign m103_11 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_12 = W*in
   wire signed [14:0] m103_12;
   assign m103_12 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_13 = W*in
   wire signed [14:0] m103_13;
   assign m103_13 =15'b0;

   // m103_14 = W*in
   wire signed [14:0] m103_14;
   assign m103_14 =15'b0;

   // m103_15 = W*in
   wire signed [14:0] m103_15;
   assign m103_15 =15'b0;

   // m103_16 = W*in
   wire signed [14:0] m103_16;
   assign m103_16 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_17 = W*in
   wire signed [14:0] m103_17;
   assign m103_17 ={ {3{in103[14]}} , in103[14:3] };

   // m103_18 = W*in
   wire signed [14:0] m103_18;
   assign m103_18 =15'b0;

   // m103_19 = W*in
   wire signed [14:0] m103_19;
   assign m103_19 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_20 = W*in
   wire signed [14:0] m103_20;
   assign m103_20 =15'b0;

   // m103_21 = W*in
   wire signed [14:0] m103_21;
   assign m103_21 =15'b0;

   // m103_22 = W*in
   wire signed [14:0] m103_22;
   assign m103_22 ={ {3{in103[14]}} , in103[14:3] };

   // m103_23 = W*in
   wire signed [14:0] m103_23;
   assign m103_23 =15'b0;

   // m103_24 = W*in
   wire signed [14:0] m103_24;
   assign m103_24 =15'b0;

   // m103_25 = W*in
   wire signed [14:0] m103_25;
   assign m103_25 =15'b0;

   // m103_26 = W*in
   wire signed [14:0] m103_26;
   assign m103_26 ={ {4{neg103[14]}} , neg103[14:4] };

   // m103_27 = W*in
   wire signed [14:0] m103_27;
   assign m103_27 ={ {4{neg103[14]}} , neg103[14:4] };

   // m103_28 = W*in
   wire signed [14:0] m103_28;
   assign m103_28 =15'b0;

   // m103_29 = W*in
   wire signed [14:0] m103_29;
   assign m103_29 =15'b0;

   // m103_30 = W*in
   wire signed [14:0] m103_30;
   assign m103_30 =15'b0;

   // m103_31 = W*in
   wire signed [14:0] m103_31;
   assign m103_31 =15'b0;

   // m103_32 = W*in
   wire signed [14:0] m103_32;
   assign m103_32 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_33 = W*in
   wire signed [14:0] m103_33;
   assign m103_33 =15'b0;

   // m103_34 = W*in
   wire signed [14:0] m103_34;
   assign m103_34 =15'b0;

   // m103_35 = W*in
   wire signed [14:0] m103_35;
   assign m103_35 =15'b0;

   // m103_36 = W*in
   wire signed [14:0] m103_36;
   assign m103_36 =15'b0;

   // m103_37 = W*in
   wire signed [14:0] m103_37;
   assign m103_37 =15'b0;

   // m103_38 = W*in
   wire signed [14:0] m103_38;
   assign m103_38 =15'b0;

   // m103_39 = W*in
   wire signed [14:0] m103_39;
   assign m103_39 =15'b0;

   // m103_40 = W*in
   wire signed [14:0] m103_40;
   assign m103_40 =15'b0;

   // m103_41 = W*in
   wire signed [14:0] m103_41;
   assign m103_41 =15'b0;

   // m103_42 = W*in
   wire signed [14:0] m103_42;
   assign m103_42 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_43 = W*in
   wire signed [14:0] m103_43;
   assign m103_43 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_44 = W*in
   wire signed [14:0] m103_44;
   assign m103_44 =15'b0;

   // m103_45 = W*in
   wire signed [14:0] m103_45;
   assign m103_45 ={ {3{in103[14]}} , in103[14:3] };

   // m103_46 = W*in
   wire signed [14:0] m103_46;
   assign m103_46 =15'b0;

   // m103_47 = W*in
   wire signed [14:0] m103_47;
   assign m103_47 =15'b0;

   // m103_48 = W*in
   wire signed [14:0] m103_48;
   assign m103_48 =15'b0;

   // m103_49 = W*in
   wire signed [14:0] m103_49;
   assign m103_49 =15'b0;

   // m103_50 = W*in
   wire signed [14:0] m103_50;
   assign m103_50 =15'b0;

   // m103_51 = W*in
   wire signed [14:0] m103_51;
   assign m103_51 =15'b0;

   // m103_52 = W*in
   wire signed [14:0] m103_52;
   assign m103_52 =15'b0;

   // m103_53 = W*in
   wire signed [14:0] m103_53;
   assign m103_53 =15'b0;

   // m103_54 = W*in
   wire signed [14:0] m103_54;
   assign m103_54 =15'b0;

   // m103_55 = W*in
   wire signed [14:0] m103_55;
   assign m103_55 =15'b0;

   // m103_56 = W*in
   wire signed [14:0] m103_56;
   assign m103_56 =15'b0;

   // m103_57 = W*in
   wire signed [14:0] m103_57;
   assign m103_57 =15'b0;

   // m103_58 = W*in
   wire signed [14:0] m103_58;
   assign m103_58 ={ {3{in103[14]}} , in103[14:3] };

   // m103_59 = W*in
   wire signed [14:0] m103_59;
   assign m103_59 =15'b0;

   // m103_60 = W*in
   wire signed [14:0] m103_60;
   assign m103_60 =15'b0;

   // m103_61 = W*in
   wire signed [14:0] m103_61;
   assign m103_61 =15'b0;

   // m103_62 = W*in
   wire signed [14:0] m103_62;
   assign m103_62 ={ {3{in103[14]}} , in103[14:3] };

   // m103_63 = W*in
   wire signed [14:0] m103_63;
   assign m103_63 =15'b0;

   // m103_64 = W*in
   wire signed [14:0] m103_64;
   assign m103_64 ={ {3{in103[14]}} , in103[14:3] };

   // m103_65 = W*in
   wire signed [14:0] m103_65;
   assign m103_65 =15'b0;

   // m103_66 = W*in
   wire signed [14:0] m103_66;
   assign m103_66 =15'b0;

   // m103_67 = W*in
   wire signed [14:0] m103_67;
   assign m103_67 =15'b0;

   // m103_68 = W*in
   wire signed [14:0] m103_68;
   assign m103_68 ={ {4{in103[14]}} , in103[14:4] };

   // m103_69 = W*in
   wire signed [14:0] m103_69;
   assign m103_69 =15'b0;

   // m103_70 = W*in
   wire signed [14:0] m103_70;
   assign m103_70 ={ {4{in103[14]}} , in103[14:4] };

   // m103_71 = W*in
   wire signed [14:0] m103_71;
   assign m103_71 =15'b0;

   // m103_72 = W*in
   wire signed [14:0] m103_72;
   assign m103_72 =15'b0;

   // m103_73 = W*in
   wire signed [14:0] m103_73;
   assign m103_73 =15'b0;

   // m103_74 = W*in
   wire signed [14:0] m103_74;
   assign m103_74 ={ {4{in103[14]}} , in103[14:4] };

   // m103_75 = W*in
   wire signed [14:0] m103_75;
   assign m103_75 =15'b0;

   // m103_76 = W*in
   wire signed [14:0] m103_76;
   assign m103_76 =15'b0;

   // m103_77 = W*in
   wire signed [14:0] m103_77;
   assign m103_77 ={ {4{neg103[14]}} , neg103[14:4] };

   // m103_78 = W*in
   wire signed [14:0] m103_78;
   assign m103_78 =15'b0;

   // m103_79 = W*in
   wire signed [14:0] m103_79;
   assign m103_79 =15'b0;

   // m103_80 = W*in
   wire signed [14:0] m103_80;
   assign m103_80 =15'b0;

   // m103_81 = W*in
   wire signed [14:0] m103_81;
   assign m103_81 =15'b0;

   // m103_82 = W*in
   wire signed [14:0] m103_82;
   assign m103_82 =15'b0;

   // m103_83 = W*in
   wire signed [14:0] m103_83;
   assign m103_83 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_84 = W*in
   wire signed [14:0] m103_84;
   assign m103_84 =15'b0;

   // m103_85 = W*in
   wire signed [14:0] m103_85;
   assign m103_85 ={ {3{in103[14]}} , in103[14:3] };

   // m103_86 = W*in
   wire signed [14:0] m103_86;
   assign m103_86 =15'b0;

   // m103_87 = W*in
   wire signed [14:0] m103_87;
   assign m103_87 ={ {3{in103[14]}} , in103[14:3] };

   // m103_88 = W*in
   wire signed [14:0] m103_88;
   assign m103_88 =15'b0;

   // m103_89 = W*in
   wire signed [14:0] m103_89;
   assign m103_89 =15'b0;

   // m103_90 = W*in
   wire signed [14:0] m103_90;
   assign m103_90 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_91 = W*in
   wire signed [14:0] m103_91;
   assign m103_91 =15'b0;

   // m103_92 = W*in
   wire signed [14:0] m103_92;
   assign m103_92 ={ {3{in103[14]}} , in103[14:3] };

   // m103_93 = W*in
   wire signed [14:0] m103_93;
   assign m103_93 =15'b0;

   // m103_94 = W*in
   wire signed [14:0] m103_94;
   assign m103_94 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_95 = W*in
   wire signed [14:0] m103_95;
   assign m103_95 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_96 = W*in
   wire signed [14:0] m103_96;
   assign m103_96 =15'b0;

   // m103_97 = W*in
   wire signed [14:0] m103_97;
   assign m103_97 ={ {3{neg103[14]}} , neg103[14:3] };

   // m103_98 = W*in
   wire signed [14:0] m103_98;
   assign m103_98 =15'b0;

   // m103_99 = W*in
   wire signed [14:0] m103_99;
   assign m103_99 ={ {3{in103[14]}} , in103[14:3] };

   // m103_100 = W*in
   wire signed [14:0] m103_100;
   assign m103_100 =15'b0;

   // m104_1 = W*in
   wire signed [14:0] m104_1;
   assign m104_1 =15'b0;

   // m104_2 = W*in
   wire signed [14:0] m104_2;
   assign m104_2 =15'b0;

   // m104_3 = W*in
   wire signed [14:0] m104_3;
   assign m104_3 =15'b0;

   // m104_4 = W*in
   wire signed [14:0] m104_4;
   assign m104_4 =15'b0;

   // m104_5 = W*in
   wire signed [14:0] m104_5;
   assign m104_5 =15'b0;

   // m104_6 = W*in
   wire signed [14:0] m104_6;
   assign m104_6 =15'b0;

   // m104_7 = W*in
   wire signed [14:0] m104_7;
   assign m104_7 =15'b0;

   // m104_8 = W*in
   wire signed [14:0] m104_8;
   assign m104_8 =15'b0;

   // m104_9 = W*in
   wire signed [14:0] m104_9;
   assign m104_9 =15'b0;

   // m104_10 = W*in
   wire signed [14:0] m104_10;
   assign m104_10 =15'b0;

   // m104_11 = W*in
   wire signed [14:0] m104_11;
   assign m104_11 =15'b0;

   // m104_12 = W*in
   wire signed [14:0] m104_12;
   assign m104_12 =15'b0;

   // m104_13 = W*in
   wire signed [14:0] m104_13;
   assign m104_13 =15'b0;

   // m104_14 = W*in
   wire signed [14:0] m104_14;
   assign m104_14 =15'b0;

   // m104_15 = W*in
   wire signed [14:0] m104_15;
   assign m104_15 =15'b0;

   // m104_16 = W*in
   wire signed [14:0] m104_16;
   assign m104_16 =15'b0;

   // m104_17 = W*in
   wire signed [14:0] m104_17;
   assign m104_17 ={ {4{neg104[14]}} , neg104[14:4] };

   // m104_18 = W*in
   wire signed [14:0] m104_18;
   assign m104_18 =15'b0;

   // m104_19 = W*in
   wire signed [14:0] m104_19;
   assign m104_19 =15'b0;

   // m104_20 = W*in
   wire signed [14:0] m104_20;
   assign m104_20 =15'b0;

   // m104_21 = W*in
   wire signed [14:0] m104_21;
   assign m104_21 ={ {3{in104[14]}} , in104[14:3] };

   // m104_22 = W*in
   wire signed [14:0] m104_22;
   assign m104_22 =15'b0;

   // m104_23 = W*in
   wire signed [14:0] m104_23;
   assign m104_23 =15'b0;

   // m104_24 = W*in
   wire signed [14:0] m104_24;
   assign m104_24 =15'b0;

   // m104_25 = W*in
   wire signed [14:0] m104_25;
   assign m104_25 =15'b0;

   // m104_26 = W*in
   wire signed [14:0] m104_26;
   assign m104_26 =15'b0;

   // m104_27 = W*in
   wire signed [14:0] m104_27;
   assign m104_27 ={ {3{in104[14]}} , in104[14:3] };

   // m104_28 = W*in
   wire signed [14:0] m104_28;
   assign m104_28 =15'b0;

   // m104_29 = W*in
   wire signed [14:0] m104_29;
   assign m104_29 =15'b0;

   // m104_30 = W*in
   wire signed [14:0] m104_30;
   assign m104_30 =15'b0;

   // m104_31 = W*in
   wire signed [14:0] m104_31;
   assign m104_31 =15'b0;

   // m104_32 = W*in
   wire signed [14:0] m104_32;
   assign m104_32 =15'b0;

   // m104_33 = W*in
   wire signed [14:0] m104_33;
   assign m104_33 =15'b0;

   // m104_34 = W*in
   wire signed [14:0] m104_34;
   assign m104_34 =15'b0;

   // m104_35 = W*in
   wire signed [14:0] m104_35;
   assign m104_35 =15'b0;

   // m104_36 = W*in
   wire signed [14:0] m104_36;
   assign m104_36 =15'b0;

   // m104_37 = W*in
   wire signed [14:0] m104_37;
   assign m104_37 =15'b0;

   // m104_38 = W*in
   wire signed [14:0] m104_38;
   assign m104_38 =15'b0;

   // m104_39 = W*in
   wire signed [14:0] m104_39;
   assign m104_39 =15'b0;

   // m104_40 = W*in
   wire signed [14:0] m104_40;
   assign m104_40 =15'b0;

   // m104_41 = W*in
   wire signed [14:0] m104_41;
   assign m104_41 =15'b0;

   // m104_42 = W*in
   wire signed [14:0] m104_42;
   assign m104_42 =15'b0;

   // m104_43 = W*in
   wire signed [14:0] m104_43;
   assign m104_43 =15'b0;

   // m104_44 = W*in
   wire signed [14:0] m104_44;
   assign m104_44 =15'b0;

   // m104_45 = W*in
   wire signed [14:0] m104_45;
   assign m104_45 =15'b0;

   // m104_46 = W*in
   wire signed [14:0] m104_46;
   assign m104_46 =15'b0;

   // m104_47 = W*in
   wire signed [14:0] m104_47;
   assign m104_47 =15'b0;

   // m104_48 = W*in
   wire signed [14:0] m104_48;
   assign m104_48 =15'b0;

   // m104_49 = W*in
   wire signed [14:0] m104_49;
   assign m104_49 =15'b0;

   // m104_50 = W*in
   wire signed [14:0] m104_50;
   assign m104_50 =15'b0;

   // m104_51 = W*in
   wire signed [14:0] m104_51;
   assign m104_51 =15'b0;

   // m104_52 = W*in
   wire signed [14:0] m104_52;
   assign m104_52 =15'b0;

   // m104_53 = W*in
   wire signed [14:0] m104_53;
   assign m104_53 =15'b0;

   // m104_54 = W*in
   wire signed [14:0] m104_54;
   assign m104_54 =15'b0;

   // m104_55 = W*in
   wire signed [14:0] m104_55;
   assign m104_55 =15'b0;

   // m104_56 = W*in
   wire signed [14:0] m104_56;
   assign m104_56 =15'b0;

   // m104_57 = W*in
   wire signed [14:0] m104_57;
   assign m104_57 =15'b0;

   // m104_58 = W*in
   wire signed [14:0] m104_58;
   assign m104_58 =15'b0;

   // m104_59 = W*in
   wire signed [14:0] m104_59;
   assign m104_59 =15'b0;

   // m104_60 = W*in
   wire signed [14:0] m104_60;
   assign m104_60 ={ {4{in104[14]}} , in104[14:4] };

   // m104_61 = W*in
   wire signed [14:0] m104_61;
   assign m104_61 =15'b0;

   // m104_62 = W*in
   wire signed [14:0] m104_62;
   assign m104_62 =15'b0;

   // m104_63 = W*in
   wire signed [14:0] m104_63;
   assign m104_63 =15'b0;

   // m104_64 = W*in
   wire signed [14:0] m104_64;
   assign m104_64 =15'b0;

   // m104_65 = W*in
   wire signed [14:0] m104_65;
   assign m104_65 =15'b0;

   // m104_66 = W*in
   wire signed [14:0] m104_66;
   assign m104_66 =15'b0;

   // m104_67 = W*in
   wire signed [14:0] m104_67;
   assign m104_67 =15'b0;

   // m104_68 = W*in
   wire signed [14:0] m104_68;
   assign m104_68 =15'b0;

   // m104_69 = W*in
   wire signed [14:0] m104_69;
   assign m104_69 =15'b0;

   // m104_70 = W*in
   wire signed [14:0] m104_70;
   assign m104_70 =15'b0;

   // m104_71 = W*in
   wire signed [14:0] m104_71;
   assign m104_71 =15'b0;

   // m104_72 = W*in
   wire signed [14:0] m104_72;
   assign m104_72 =15'b0;

   // m104_73 = W*in
   wire signed [14:0] m104_73;
   assign m104_73 =15'b0;

   // m104_74 = W*in
   wire signed [14:0] m104_74;
   assign m104_74 =15'b0;

   // m104_75 = W*in
   wire signed [14:0] m104_75;
   assign m104_75 =15'b0;

   // m104_76 = W*in
   wire signed [14:0] m104_76;
   assign m104_76 =15'b0;

   // m104_77 = W*in
   wire signed [14:0] m104_77;
   assign m104_77 ={ {4{in104[14]}} , in104[14:4] };

   // m104_78 = W*in
   wire signed [14:0] m104_78;
   assign m104_78 =15'b0;

   // m104_79 = W*in
   wire signed [14:0] m104_79;
   assign m104_79 =15'b0;

   // m104_80 = W*in
   wire signed [14:0] m104_80;
   assign m104_80 =15'b0;

   // m104_81 = W*in
   wire signed [14:0] m104_81;
   assign m104_81 =15'b0;

   // m104_82 = W*in
   wire signed [14:0] m104_82;
   assign m104_82 =15'b0;

   // m104_83 = W*in
   wire signed [14:0] m104_83;
   assign m104_83 =15'b0;

   // m104_84 = W*in
   wire signed [14:0] m104_84;
   assign m104_84 ={ {3{in104[14]}} , in104[14:3] };

   // m104_85 = W*in
   wire signed [14:0] m104_85;
   assign m104_85 =15'b0;

   // m104_86 = W*in
   wire signed [14:0] m104_86;
   assign m104_86 =15'b0;

   // m104_87 = W*in
   wire signed [14:0] m104_87;
   assign m104_87 =15'b0;

   // m104_88 = W*in
   wire signed [14:0] m104_88;
   assign m104_88 =15'b0;

   // m104_89 = W*in
   wire signed [14:0] m104_89;
   assign m104_89 =15'b0;

   // m104_90 = W*in
   wire signed [14:0] m104_90;
   assign m104_90 =15'b0;

   // m104_91 = W*in
   wire signed [14:0] m104_91;
   assign m104_91 =15'b0;

   // m104_92 = W*in
   wire signed [14:0] m104_92;
   assign m104_92 =15'b0;

   // m104_93 = W*in
   wire signed [14:0] m104_93;
   assign m104_93 =15'b0;

   // m104_94 = W*in
   wire signed [14:0] m104_94;
   assign m104_94 =15'b0;

   // m104_95 = W*in
   wire signed [14:0] m104_95;
   assign m104_95 =15'b0;

   // m104_96 = W*in
   wire signed [14:0] m104_96;
   assign m104_96 =15'b0;

   // m104_97 = W*in
   wire signed [14:0] m104_97;
   assign m104_97 =15'b0;

   // m104_98 = W*in
   wire signed [14:0] m104_98;
   assign m104_98 ={ {4{in104[14]}} , in104[14:4] };

   // m104_99 = W*in
   wire signed [14:0] m104_99;
   assign m104_99 =15'b0;

   // m104_100 = W*in
   wire signed [14:0] m104_100;
   assign m104_100 ={ {4{neg104[14]}} , neg104[14:4] };

   // m105_1 = W*in
   wire signed [14:0] m105_1;
   assign m105_1 =15'b0;

   // m105_2 = W*in
   wire signed [14:0] m105_2;
   assign m105_2 =15'b0;

   // m105_3 = W*in
   wire signed [14:0] m105_3;
   assign m105_3 ={ {4{neg105[14]}} , neg105[14:4] };

   // m105_4 = W*in
   wire signed [14:0] m105_4;
   assign m105_4 =15'b0;

   // m105_5 = W*in
   wire signed [14:0] m105_5;
   assign m105_5 =15'b0;

   // m105_6 = W*in
   wire signed [14:0] m105_6;
   assign m105_6 =15'b0;

   // m105_7 = W*in
   wire signed [14:0] m105_7;
   assign m105_7 =15'b0;

   // m105_8 = W*in
   wire signed [14:0] m105_8;
   assign m105_8 =15'b0;

   // m105_9 = W*in
   wire signed [14:0] m105_9;
   assign m105_9 =15'b0;

   // m105_10 = W*in
   wire signed [14:0] m105_10;
   assign m105_10 ={ {4{in105[14]}} , in105[14:4] };

   // m105_11 = W*in
   wire signed [14:0] m105_11;
   assign m105_11 =15'b0;

   // m105_12 = W*in
   wire signed [14:0] m105_12;
   assign m105_12 =15'b0;

   // m105_13 = W*in
   wire signed [14:0] m105_13;
   assign m105_13 =15'b0;

   // m105_14 = W*in
   wire signed [14:0] m105_14;
   assign m105_14 =15'b0;

   // m105_15 = W*in
   wire signed [14:0] m105_15;
   assign m105_15 =15'b0;

   // m105_16 = W*in
   wire signed [14:0] m105_16;
   assign m105_16 ={ {3{in105[14]}} , in105[14:3] };

   // m105_17 = W*in
   wire signed [14:0] m105_17;
   assign m105_17 =15'b0;

   // m105_18 = W*in
   wire signed [14:0] m105_18;
   assign m105_18 =15'b0;

   // m105_19 = W*in
   wire signed [14:0] m105_19;
   assign m105_19 =15'b0;

   // m105_20 = W*in
   wire signed [14:0] m105_20;
   assign m105_20 =15'b0;

   // m105_21 = W*in
   wire signed [14:0] m105_21;
   assign m105_21 =15'b0;

   // m105_22 = W*in
   wire signed [14:0] m105_22;
   assign m105_22 =15'b0;

   // m105_23 = W*in
   wire signed [14:0] m105_23;
   assign m105_23 =15'b0;

   // m105_24 = W*in
   wire signed [14:0] m105_24;
   assign m105_24 =15'b0;

   // m105_25 = W*in
   wire signed [14:0] m105_25;
   assign m105_25 ={ {3{in105[14]}} , in105[14:3] };

   // m105_26 = W*in
   wire signed [14:0] m105_26;
   assign m105_26 =15'b0;

   // m105_27 = W*in
   wire signed [14:0] m105_27;
   assign m105_27 =15'b0;

   // m105_28 = W*in
   wire signed [14:0] m105_28;
   assign m105_28 =15'b0;

   // m105_29 = W*in
   wire signed [14:0] m105_29;
   assign m105_29 =15'b0;

   // m105_30 = W*in
   wire signed [14:0] m105_30;
   assign m105_30 =15'b0;

   // m105_31 = W*in
   wire signed [14:0] m105_31;
   assign m105_31 ={ {4{neg105[14]}} , neg105[14:4] };

   // m105_32 = W*in
   wire signed [14:0] m105_32;
   assign m105_32 =15'b0;

   // m105_33 = W*in
   wire signed [14:0] m105_33;
   assign m105_33 =15'b0;

   // m105_34 = W*in
   wire signed [14:0] m105_34;
   assign m105_34 =15'b0;

   // m105_35 = W*in
   wire signed [14:0] m105_35;
   assign m105_35 =15'b0;

   // m105_36 = W*in
   wire signed [14:0] m105_36;
   assign m105_36 =15'b0;

   // m105_37 = W*in
   wire signed [14:0] m105_37;
   assign m105_37 =15'b0;

   // m105_38 = W*in
   wire signed [14:0] m105_38;
   assign m105_38 =15'b0;

   // m105_39 = W*in
   wire signed [14:0] m105_39;
   assign m105_39 =15'b0;

   // m105_40 = W*in
   wire signed [14:0] m105_40;
   assign m105_40 =15'b0;

   // m105_41 = W*in
   wire signed [14:0] m105_41;
   assign m105_41 =15'b0;

   // m105_42 = W*in
   wire signed [14:0] m105_42;
   assign m105_42 =15'b0;

   // m105_43 = W*in
   wire signed [14:0] m105_43;
   assign m105_43 =15'b0;

   // m105_44 = W*in
   wire signed [14:0] m105_44;
   assign m105_44 =15'b0;

   // m105_45 = W*in
   wire signed [14:0] m105_45;
   assign m105_45 =15'b0;

   // m105_46 = W*in
   wire signed [14:0] m105_46;
   assign m105_46 ={ {4{in105[14]}} , in105[14:4] };

   // m105_47 = W*in
   wire signed [14:0] m105_47;
   assign m105_47 ={ {4{neg105[14]}} , neg105[14:4] };

   // m105_48 = W*in
   wire signed [14:0] m105_48;
   assign m105_48 =15'b0;

   // m105_49 = W*in
   wire signed [14:0] m105_49;
   assign m105_49 ={ {3{in105[14]}} , in105[14:3] };

   // m105_50 = W*in
   wire signed [14:0] m105_50;
   assign m105_50 =15'b0;

   // m105_51 = W*in
   wire signed [14:0] m105_51;
   assign m105_51 =15'b0;

   // m105_52 = W*in
   wire signed [14:0] m105_52;
   assign m105_52 =15'b0;

   // m105_53 = W*in
   wire signed [14:0] m105_53;
   assign m105_53 =15'b0;

   // m105_54 = W*in
   wire signed [14:0] m105_54;
   assign m105_54 =15'b0;

   // m105_55 = W*in
   wire signed [14:0] m105_55;
   assign m105_55 =15'b0;

   // m105_56 = W*in
   wire signed [14:0] m105_56;
   assign m105_56 =15'b0;

   // m105_57 = W*in
   wire signed [14:0] m105_57;
   assign m105_57 =15'b0;

   // m105_58 = W*in
   wire signed [14:0] m105_58;
   assign m105_58 =15'b0;

   // m105_59 = W*in
   wire signed [14:0] m105_59;
   assign m105_59 ={ {3{in105[14]}} , in105[14:3] };

   // m105_60 = W*in
   wire signed [14:0] m105_60;
   assign m105_60 ={ {4{neg105[14]}} , neg105[14:4] };

   // m105_61 = W*in
   wire signed [14:0] m105_61;
   assign m105_61 =15'b0;

   // m105_62 = W*in
   wire signed [14:0] m105_62;
   assign m105_62 =15'b0;

   // m105_63 = W*in
   wire signed [14:0] m105_63;
   assign m105_63 =15'b0;

   // m105_64 = W*in
   wire signed [14:0] m105_64;
   assign m105_64 =15'b0;

   // m105_65 = W*in
   wire signed [14:0] m105_65;
   assign m105_65 =15'b0;

   // m105_66 = W*in
   wire signed [14:0] m105_66;
   assign m105_66 =15'b0;

   // m105_67 = W*in
   wire signed [14:0] m105_67;
   assign m105_67 =15'b0;

   // m105_68 = W*in
   wire signed [14:0] m105_68;
   assign m105_68 =15'b0;

   // m105_69 = W*in
   wire signed [14:0] m105_69;
   assign m105_69 =15'b0;

   // m105_70 = W*in
   wire signed [14:0] m105_70;
   assign m105_70 =15'b0;

   // m105_71 = W*in
   wire signed [14:0] m105_71;
   assign m105_71 =15'b0;

   // m105_72 = W*in
   wire signed [14:0] m105_72;
   assign m105_72 ={ {3{in105[14]}} , in105[14:3] };

   // m105_73 = W*in
   wire signed [14:0] m105_73;
   assign m105_73 =15'b0;

   // m105_74 = W*in
   wire signed [14:0] m105_74;
   assign m105_74 ={ {4{neg105[14]}} , neg105[14:4] };

   // m105_75 = W*in
   wire signed [14:0] m105_75;
   assign m105_75 =15'b0;

   // m105_76 = W*in
   wire signed [14:0] m105_76;
   assign m105_76 =15'b0;

   // m105_77 = W*in
   wire signed [14:0] m105_77;
   assign m105_77 ={ {3{neg105[14]}} , neg105[14:3] };

   // m105_78 = W*in
   wire signed [14:0] m105_78;
   assign m105_78 =15'b0;

   // m105_79 = W*in
   wire signed [14:0] m105_79;
   assign m105_79 =15'b0;

   // m105_80 = W*in
   wire signed [14:0] m105_80;
   assign m105_80 =15'b0;

   // m105_81 = W*in
   wire signed [14:0] m105_81;
   assign m105_81 ={ {4{in105[14]}} , in105[14:4] };

   // m105_82 = W*in
   wire signed [14:0] m105_82;
   assign m105_82 =15'b0;

   // m105_83 = W*in
   wire signed [14:0] m105_83;
   assign m105_83 =15'b0;

   // m105_84 = W*in
   wire signed [14:0] m105_84;
   assign m105_84 =15'b0;

   // m105_85 = W*in
   wire signed [14:0] m105_85;
   assign m105_85 =15'b0;

   // m105_86 = W*in
   wire signed [14:0] m105_86;
   assign m105_86 =15'b0;

   // m105_87 = W*in
   wire signed [14:0] m105_87;
   assign m105_87 =15'b0;

   // m105_88 = W*in
   wire signed [14:0] m105_88;
   assign m105_88 =15'b0;

   // m105_89 = W*in
   wire signed [14:0] m105_89;
   assign m105_89 =15'b0;

   // m105_90 = W*in
   wire signed [14:0] m105_90;
   assign m105_90 =15'b0;

   // m105_91 = W*in
   wire signed [14:0] m105_91;
   assign m105_91 =15'b0;

   // m105_92 = W*in
   wire signed [14:0] m105_92;
   assign m105_92 =15'b0;

   // m105_93 = W*in
   wire signed [14:0] m105_93;
   assign m105_93 =15'b0;

   // m105_94 = W*in
   wire signed [14:0] m105_94;
   assign m105_94 =15'b0;

   // m105_95 = W*in
   wire signed [14:0] m105_95;
   assign m105_95 =15'b0;

   // m105_96 = W*in
   wire signed [14:0] m105_96;
   assign m105_96 ={ {4{in105[14]}} , in105[14:4] };

   // m105_97 = W*in
   wire signed [14:0] m105_97;
   assign m105_97 =15'b0;

   // m105_98 = W*in
   wire signed [14:0] m105_98;
   assign m105_98 ={ {4{neg105[14]}} , neg105[14:4] };

   // m105_99 = W*in
   wire signed [14:0] m105_99;
   assign m105_99 ={ {3{neg105[14]}} , neg105[14:3] };

   // m105_100 = W*in
   wire signed [14:0] m105_100;
   assign m105_100 =15'b0;

   // m106_1 = W*in
   wire signed [14:0] m106_1;
   assign m106_1 =15'b0;

   // m106_2 = W*in
   wire signed [14:0] m106_2;
   assign m106_2 =15'b0;

   // m106_3 = W*in
   wire signed [14:0] m106_3;
   assign m106_3 =15'b0;

   // m106_4 = W*in
   wire signed [14:0] m106_4;
   assign m106_4 =15'b0;

   // m106_5 = W*in
   wire signed [14:0] m106_5;
   assign m106_5 =15'b0;

   // m106_6 = W*in
   wire signed [14:0] m106_6;
   assign m106_6 =15'b0;

   // m106_7 = W*in
   wire signed [14:0] m106_7;
   assign m106_7 =15'b0;

   // m106_8 = W*in
   wire signed [14:0] m106_8;
   assign m106_8 =15'b0;

   // m106_9 = W*in
   wire signed [14:0] m106_9;
   assign m106_9 =15'b0;

   // m106_10 = W*in
   wire signed [14:0] m106_10;
   assign m106_10 =15'b0;

   // m106_11 = W*in
   wire signed [14:0] m106_11;
   assign m106_11 =15'b0;

   // m106_12 = W*in
   wire signed [14:0] m106_12;
   assign m106_12 =15'b0;

   // m106_13 = W*in
   wire signed [14:0] m106_13;
   assign m106_13 =15'b0;

   // m106_14 = W*in
   wire signed [14:0] m106_14;
   assign m106_14 =15'b0;

   // m106_15 = W*in
   wire signed [14:0] m106_15;
   assign m106_15 =15'b0;

   // m106_16 = W*in
   wire signed [14:0] m106_16;
   assign m106_16 ={ {3{neg106[14]}} , neg106[14:3] };

   // m106_17 = W*in
   wire signed [14:0] m106_17;
   assign m106_17 =15'b0;

   // m106_18 = W*in
   wire signed [14:0] m106_18;
   assign m106_18 =15'b0;

   // m106_19 = W*in
   wire signed [14:0] m106_19;
   assign m106_19 =15'b0;

   // m106_20 = W*in
   wire signed [14:0] m106_20;
   assign m106_20 =15'b0;

   // m106_21 = W*in
   wire signed [14:0] m106_21;
   assign m106_21 =15'b0;

   // m106_22 = W*in
   wire signed [14:0] m106_22;
   assign m106_22 =15'b0;

   // m106_23 = W*in
   wire signed [14:0] m106_23;
   assign m106_23 ={ {3{in106[14]}} , in106[14:3] };

   // m106_24 = W*in
   wire signed [14:0] m106_24;
   assign m106_24 =15'b0;

   // m106_25 = W*in
   wire signed [14:0] m106_25;
   assign m106_25 =15'b0;

   // m106_26 = W*in
   wire signed [14:0] m106_26;
   assign m106_26 =15'b0;

   // m106_27 = W*in
   wire signed [14:0] m106_27;
   assign m106_27 =15'b0;

   // m106_28 = W*in
   wire signed [14:0] m106_28;
   assign m106_28 ={ {3{in106[14]}} , in106[14:3] };

   // m106_29 = W*in
   wire signed [14:0] m106_29;
   assign m106_29 ={ {3{in106[14]}} , in106[14:3] };

   // m106_30 = W*in
   wire signed [14:0] m106_30;
   assign m106_30 =15'b0;

   // m106_31 = W*in
   wire signed [14:0] m106_31;
   assign m106_31 =15'b0;

   // m106_32 = W*in
   wire signed [14:0] m106_32;
   assign m106_32 ={ {3{neg106[14]}} , neg106[14:3] };

   // m106_33 = W*in
   wire signed [14:0] m106_33;
   assign m106_33 =15'b0;

   // m106_34 = W*in
   wire signed [14:0] m106_34;
   assign m106_34 =15'b0;

   // m106_35 = W*in
   wire signed [14:0] m106_35;
   assign m106_35 =15'b0;

   // m106_36 = W*in
   wire signed [14:0] m106_36;
   assign m106_36 =15'b0;

   // m106_37 = W*in
   wire signed [14:0] m106_37;
   assign m106_37 =15'b0;

   // m106_38 = W*in
   wire signed [14:0] m106_38;
   assign m106_38 =15'b0;

   // m106_39 = W*in
   wire signed [14:0] m106_39;
   assign m106_39 =15'b0;

   // m106_40 = W*in
   wire signed [14:0] m106_40;
   assign m106_40 =15'b0;

   // m106_41 = W*in
   wire signed [14:0] m106_41;
   assign m106_41 =15'b0;

   // m106_42 = W*in
   wire signed [14:0] m106_42;
   assign m106_42 =15'b0;

   // m106_43 = W*in
   wire signed [14:0] m106_43;
   assign m106_43 =15'b0;

   // m106_44 = W*in
   wire signed [14:0] m106_44;
   assign m106_44 =15'b0;

   // m106_45 = W*in
   wire signed [14:0] m106_45;
   assign m106_45 =15'b0;

   // m106_46 = W*in
   wire signed [14:0] m106_46;
   assign m106_46 =15'b0;

   // m106_47 = W*in
   wire signed [14:0] m106_47;
   assign m106_47 =15'b0;

   // m106_48 = W*in
   wire signed [14:0] m106_48;
   assign m106_48 ={ {4{neg106[14]}} , neg106[14:4] };

   // m106_49 = W*in
   wire signed [14:0] m106_49;
   assign m106_49 ={ {4{in106[14]}} , in106[14:4] };

   // m106_50 = W*in
   wire signed [14:0] m106_50;
   assign m106_50 ={ {3{in106[14]}} , in106[14:3] };

   // m106_51 = W*in
   wire signed [14:0] m106_51;
   assign m106_51 ={ {3{neg106[14]}} , neg106[14:3] };

   // m106_52 = W*in
   wire signed [14:0] m106_52;
   assign m106_52 =15'b0;

   // m106_53 = W*in
   wire signed [14:0] m106_53;
   assign m106_53 =15'b0;

   // m106_54 = W*in
   wire signed [14:0] m106_54;
   assign m106_54 =15'b0;

   // m106_55 = W*in
   wire signed [14:0] m106_55;
   assign m106_55 =15'b0;

   // m106_56 = W*in
   wire signed [14:0] m106_56;
   assign m106_56 =15'b0;

   // m106_57 = W*in
   wire signed [14:0] m106_57;
   assign m106_57 =15'b0;

   // m106_58 = W*in
   wire signed [14:0] m106_58;
   assign m106_58 =15'b0;

   // m106_59 = W*in
   wire signed [14:0] m106_59;
   assign m106_59 =15'b0;

   // m106_60 = W*in
   wire signed [14:0] m106_60;
   assign m106_60 =15'b0;

   // m106_61 = W*in
   wire signed [14:0] m106_61;
   assign m106_61 =15'b0;

   // m106_62 = W*in
   wire signed [14:0] m106_62;
   assign m106_62 =15'b0;

   // m106_63 = W*in
   wire signed [14:0] m106_63;
   assign m106_63 =15'b0;

   // m106_64 = W*in
   wire signed [14:0] m106_64;
   assign m106_64 ={ {2{in106[14]}} , in106[14:2] };

   // m106_65 = W*in
   wire signed [14:0] m106_65;
   assign m106_65 =15'b0;

   // m106_66 = W*in
   wire signed [14:0] m106_66;
   assign m106_66 =15'b0;

   // m106_67 = W*in
   wire signed [14:0] m106_67;
   assign m106_67 =15'b0;

   // m106_68 = W*in
   wire signed [14:0] m106_68;
   assign m106_68 =15'b0;

   // m106_69 = W*in
   wire signed [14:0] m106_69;
   assign m106_69 =15'b0;

   // m106_70 = W*in
   wire signed [14:0] m106_70;
   assign m106_70 =15'b0;

   // m106_71 = W*in
   wire signed [14:0] m106_71;
   assign m106_71 =15'b0;

   // m106_72 = W*in
   wire signed [14:0] m106_72;
   assign m106_72 =15'b0;

   // m106_73 = W*in
   wire signed [14:0] m106_73;
   assign m106_73 =15'b0;

   // m106_74 = W*in
   wire signed [14:0] m106_74;
   assign m106_74 =15'b0;

   // m106_75 = W*in
   wire signed [14:0] m106_75;
   assign m106_75 =15'b0;

   // m106_76 = W*in
   wire signed [14:0] m106_76;
   assign m106_76 =15'b0;

   // m106_77 = W*in
   wire signed [14:0] m106_77;
   assign m106_77 =15'b0;

   // m106_78 = W*in
   wire signed [14:0] m106_78;
   assign m106_78 ={ {4{neg106[14]}} , neg106[14:4] };

   // m106_79 = W*in
   wire signed [14:0] m106_79;
   assign m106_79 =15'b0;

   // m106_80 = W*in
   wire signed [14:0] m106_80;
   assign m106_80 =15'b0;

   // m106_81 = W*in
   wire signed [14:0] m106_81;
   assign m106_81 =15'b0;

   // m106_82 = W*in
   wire signed [14:0] m106_82;
   assign m106_82 =15'b0;

   // m106_83 = W*in
   wire signed [14:0] m106_83;
   assign m106_83 =15'b0;

   // m106_84 = W*in
   wire signed [14:0] m106_84;
   assign m106_84 =15'b0;

   // m106_85 = W*in
   wire signed [14:0] m106_85;
   assign m106_85 ={ {3{in106[14]}} , in106[14:3] };

   // m106_86 = W*in
   wire signed [14:0] m106_86;
   assign m106_86 =15'b0;

   // m106_87 = W*in
   wire signed [14:0] m106_87;
   assign m106_87 ={ {3{in106[14]}} , in106[14:3] };

   // m106_88 = W*in
   wire signed [14:0] m106_88;
   assign m106_88 =15'b0;

   // m106_89 = W*in
   wire signed [14:0] m106_89;
   assign m106_89 =15'b0;

   // m106_90 = W*in
   wire signed [14:0] m106_90;
   assign m106_90 =15'b0;

   // m106_91 = W*in
   wire signed [14:0] m106_91;
   assign m106_91 =15'b0;

   // m106_92 = W*in
   wire signed [14:0] m106_92;
   assign m106_92 =15'b0;

   // m106_93 = W*in
   wire signed [14:0] m106_93;
   assign m106_93 =15'b0;

   // m106_94 = W*in
   wire signed [14:0] m106_94;
   assign m106_94 =15'b0;

   // m106_95 = W*in
   wire signed [14:0] m106_95;
   assign m106_95 =15'b0;

   // m106_96 = W*in
   wire signed [14:0] m106_96;
   assign m106_96 =15'b0;

   // m106_97 = W*in
   wire signed [14:0] m106_97;
   assign m106_97 =15'b0;

   // m106_98 = W*in
   wire signed [14:0] m106_98;
   assign m106_98 =15'b0;

   // m106_99 = W*in
   wire signed [14:0] m106_99;
   assign m106_99 =15'b0;

   // m106_100 = W*in
   wire signed [14:0] m106_100;
   assign m106_100 =15'b0;

   // m107_1 = W*in
   wire signed [14:0] m107_1;
   assign m107_1 =15'b0;

   // m107_2 = W*in
   wire signed [14:0] m107_2;
   assign m107_2 =15'b0;

   // m107_3 = W*in
   wire signed [14:0] m107_3;
   assign m107_3 ={ {3{neg107[14]}} , neg107[14:3] };

   // m107_4 = W*in
   wire signed [14:0] m107_4;
   assign m107_4 =15'b0;

   // m107_5 = W*in
   wire signed [14:0] m107_5;
   assign m107_5 =15'b0;

   // m107_6 = W*in
   wire signed [14:0] m107_6;
   assign m107_6 ={ {3{neg107[14]}} , neg107[14:3] };

   // m107_7 = W*in
   wire signed [14:0] m107_7;
   assign m107_7 =15'b0;

   // m107_8 = W*in
   wire signed [14:0] m107_8;
   assign m107_8 =15'b0;

   // m107_9 = W*in
   wire signed [14:0] m107_9;
   assign m107_9 =15'b0;

   // m107_10 = W*in
   wire signed [14:0] m107_10;
   assign m107_10 =15'b0;

   // m107_11 = W*in
   wire signed [14:0] m107_11;
   assign m107_11 =15'b0;

   // m107_12 = W*in
   wire signed [14:0] m107_12;
   assign m107_12 =15'b0;

   // m107_13 = W*in
   wire signed [14:0] m107_13;
   assign m107_13 =15'b0;

   // m107_14 = W*in
   wire signed [14:0] m107_14;
   assign m107_14 =15'b0;

   // m107_15 = W*in
   wire signed [14:0] m107_15;
   assign m107_15 =15'b0;

   // m107_16 = W*in
   wire signed [14:0] m107_16;
   assign m107_16 =15'b0;

   // m107_17 = W*in
   wire signed [14:0] m107_17;
   assign m107_17 =15'b0;

   // m107_18 = W*in
   wire signed [14:0] m107_18;
   assign m107_18 =15'b0;

   // m107_19 = W*in
   wire signed [14:0] m107_19;
   assign m107_19 ={ {3{in107[14]}} , in107[14:3] };

   // m107_20 = W*in
   wire signed [14:0] m107_20;
   assign m107_20 =15'b0;

   // m107_21 = W*in
   wire signed [14:0] m107_21;
   assign m107_21 =15'b0;

   // m107_22 = W*in
   wire signed [14:0] m107_22;
   assign m107_22 =15'b0;

   // m107_23 = W*in
   wire signed [14:0] m107_23;
   assign m107_23 =15'b0;

   // m107_24 = W*in
   wire signed [14:0] m107_24;
   assign m107_24 =15'b0;

   // m107_25 = W*in
   wire signed [14:0] m107_25;
   assign m107_25 =15'b0;

   // m107_26 = W*in
   wire signed [14:0] m107_26;
   assign m107_26 =15'b0;

   // m107_27 = W*in
   wire signed [14:0] m107_27;
   assign m107_27 =15'b0;

   // m107_28 = W*in
   wire signed [14:0] m107_28;
   assign m107_28 =15'b0;

   // m107_29 = W*in
   wire signed [14:0] m107_29;
   assign m107_29 ={ {3{neg107[14]}} , neg107[14:3] };

   // m107_30 = W*in
   wire signed [14:0] m107_30;
   assign m107_30 =15'b0;

   // m107_31 = W*in
   wire signed [14:0] m107_31;
   assign m107_31 =15'b0;

   // m107_32 = W*in
   wire signed [14:0] m107_32;
   assign m107_32 =15'b0;

   // m107_33 = W*in
   wire signed [14:0] m107_33;
   assign m107_33 =15'b0;

   // m107_34 = W*in
   wire signed [14:0] m107_34;
   assign m107_34 =15'b0;

   // m107_35 = W*in
   wire signed [14:0] m107_35;
   assign m107_35 =15'b0;

   // m107_36 = W*in
   wire signed [14:0] m107_36;
   assign m107_36 =15'b0;

   // m107_37 = W*in
   wire signed [14:0] m107_37;
   assign m107_37 =15'b0;

   // m107_38 = W*in
   wire signed [14:0] m107_38;
   assign m107_38 =15'b0;

   // m107_39 = W*in
   wire signed [14:0] m107_39;
   assign m107_39 =15'b0;

   // m107_40 = W*in
   wire signed [14:0] m107_40;
   assign m107_40 ={ {3{in107[14]}} , in107[14:3] };

   // m107_41 = W*in
   wire signed [14:0] m107_41;
   assign m107_41 =15'b0;

   // m107_42 = W*in
   wire signed [14:0] m107_42;
   assign m107_42 =15'b0;

   // m107_43 = W*in
   wire signed [14:0] m107_43;
   assign m107_43 =15'b0;

   // m107_44 = W*in
   wire signed [14:0] m107_44;
   assign m107_44 =15'b0;

   // m107_45 = W*in
   wire signed [14:0] m107_45;
   assign m107_45 =15'b0;

   // m107_46 = W*in
   wire signed [14:0] m107_46;
   assign m107_46 =15'b0;

   // m107_47 = W*in
   wire signed [14:0] m107_47;
   assign m107_47 =15'b0;

   // m107_48 = W*in
   wire signed [14:0] m107_48;
   assign m107_48 =15'b0;

   // m107_49 = W*in
   wire signed [14:0] m107_49;
   assign m107_49 =15'b0;

   // m107_50 = W*in
   wire signed [14:0] m107_50;
   assign m107_50 =15'b0;

   // m107_51 = W*in
   wire signed [14:0] m107_51;
   assign m107_51 =15'b0;

   // m107_52 = W*in
   wire signed [14:0] m107_52;
   assign m107_52 =15'b0;

   // m107_53 = W*in
   wire signed [14:0] m107_53;
   assign m107_53 =15'b0;

   // m107_54 = W*in
   wire signed [14:0] m107_54;
   assign m107_54 ={ {3{neg107[14]}} , neg107[14:3] };

   // m107_55 = W*in
   wire signed [14:0] m107_55;
   assign m107_55 =15'b0;

   // m107_56 = W*in
   wire signed [14:0] m107_56;
   assign m107_56 =15'b0;

   // m107_57 = W*in
   wire signed [14:0] m107_57;
   assign m107_57 =15'b0;

   // m107_58 = W*in
   wire signed [14:0] m107_58;
   assign m107_58 =15'b0;

   // m107_59 = W*in
   wire signed [14:0] m107_59;
   assign m107_59 =15'b0;

   // m107_60 = W*in
   wire signed [14:0] m107_60;
   assign m107_60 ={ {2{neg107[14]}} , neg107[14:2] };

   // m107_61 = W*in
   wire signed [14:0] m107_61;
   assign m107_61 =15'b0;

   // m107_62 = W*in
   wire signed [14:0] m107_62;
   assign m107_62 =15'b0;

   // m107_63 = W*in
   wire signed [14:0] m107_63;
   assign m107_63 =15'b0;

   // m107_64 = W*in
   wire signed [14:0] m107_64;
   assign m107_64 ={ {3{in107[14]}} , in107[14:3] };

   // m107_65 = W*in
   wire signed [14:0] m107_65;
   assign m107_65 =15'b0;

   // m107_66 = W*in
   wire signed [14:0] m107_66;
   assign m107_66 =15'b0;

   // m107_67 = W*in
   wire signed [14:0] m107_67;
   assign m107_67 =15'b0;

   // m107_68 = W*in
   wire signed [14:0] m107_68;
   assign m107_68 =15'b0;

   // m107_69 = W*in
   wire signed [14:0] m107_69;
   assign m107_69 =15'b0;

   // m107_70 = W*in
   wire signed [14:0] m107_70;
   assign m107_70 ={ {3{in107[14]}} , in107[14:3] };

   // m107_71 = W*in
   wire signed [14:0] m107_71;
   assign m107_71 =15'b0;

   // m107_72 = W*in
   wire signed [14:0] m107_72;
   assign m107_72 ={ {2{neg107[14]}} , neg107[14:2] };

   // m107_73 = W*in
   wire signed [14:0] m107_73;
   assign m107_73 =15'b0;

   // m107_74 = W*in
   wire signed [14:0] m107_74;
   assign m107_74 ={ {4{in107[14]}} , in107[14:4] };

   // m107_75 = W*in
   wire signed [14:0] m107_75;
   assign m107_75 ={ {3{in107[14]}} , in107[14:3] };

   // m107_76 = W*in
   wire signed [14:0] m107_76;
   assign m107_76 =15'b0;

   // m107_77 = W*in
   wire signed [14:0] m107_77;
   assign m107_77 =15'b0;

   // m107_78 = W*in
   wire signed [14:0] m107_78;
   assign m107_78 =15'b0;

   // m107_79 = W*in
   wire signed [14:0] m107_79;
   assign m107_79 =15'b0;

   // m107_80 = W*in
   wire signed [14:0] m107_80;
   assign m107_80 ={ {3{neg107[14]}} , neg107[14:3] };

   // m107_81 = W*in
   wire signed [14:0] m107_81;
   assign m107_81 =15'b0;

   // m107_82 = W*in
   wire signed [14:0] m107_82;
   assign m107_82 =15'b0;

   // m107_83 = W*in
   wire signed [14:0] m107_83;
   assign m107_83 =15'b0;

   // m107_84 = W*in
   wire signed [14:0] m107_84;
   assign m107_84 =15'b0;

   // m107_85 = W*in
   wire signed [14:0] m107_85;
   assign m107_85 =15'b0;

   // m107_86 = W*in
   wire signed [14:0] m107_86;
   assign m107_86 =15'b0;

   // m107_87 = W*in
   wire signed [14:0] m107_87;
   assign m107_87 =15'b0;

   // m107_88 = W*in
   wire signed [14:0] m107_88;
   assign m107_88 =15'b0;

   // m107_89 = W*in
   wire signed [14:0] m107_89;
   assign m107_89 =15'b0;

   // m107_90 = W*in
   wire signed [14:0] m107_90;
   assign m107_90 ={ {3{in107[14]}} , in107[14:3] };

   // m107_91 = W*in
   wire signed [14:0] m107_91;
   assign m107_91 =15'b0;

   // m107_92 = W*in
   wire signed [14:0] m107_92;
   assign m107_92 ={ {3{in107[14]}} , in107[14:3] };

   // m107_93 = W*in
   wire signed [14:0] m107_93;
   assign m107_93 =15'b0;

   // m107_94 = W*in
   wire signed [14:0] m107_94;
   assign m107_94 ={ {3{in107[14]}} , in107[14:3] };

   // m107_95 = W*in
   wire signed [14:0] m107_95;
   assign m107_95 =15'b0;

   // m107_96 = W*in
   wire signed [14:0] m107_96;
   assign m107_96 ={ {3{neg107[14]}} , neg107[14:3] };

   // m107_97 = W*in
   wire signed [14:0] m107_97;
   assign m107_97 ={ {3{in107[14]}} , in107[14:3] };

   // m107_98 = W*in
   wire signed [14:0] m107_98;
   assign m107_98 =15'b0;

   // m107_99 = W*in
   wire signed [14:0] m107_99;
   assign m107_99 =15'b0;

   // m107_100 = W*in
   wire signed [14:0] m107_100;
   assign m107_100 =15'b0;

   // m108_1 = W*in
   wire signed [14:0] m108_1;
   assign m108_1 =15'b0;

   // m108_2 = W*in
   wire signed [14:0] m108_2;
   assign m108_2 =15'b0;

   // m108_3 = W*in
   wire signed [14:0] m108_3;
   assign m108_3 =15'b0;

   // m108_4 = W*in
   wire signed [14:0] m108_4;
   assign m108_4 =15'b0;

   // m108_5 = W*in
   wire signed [14:0] m108_5;
   assign m108_5 =15'b0;

   // m108_6 = W*in
   wire signed [14:0] m108_6;
   assign m108_6 =15'b0;

   // m108_7 = W*in
   wire signed [14:0] m108_7;
   assign m108_7 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_8 = W*in
   wire signed [14:0] m108_8;
   assign m108_8 =15'b0;

   // m108_9 = W*in
   wire signed [14:0] m108_9;
   assign m108_9 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_10 = W*in
   wire signed [14:0] m108_10;
   assign m108_10 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_11 = W*in
   wire signed [14:0] m108_11;
   assign m108_11 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_12 = W*in
   wire signed [14:0] m108_12;
   assign m108_12 =15'b0;

   // m108_13 = W*in
   wire signed [14:0] m108_13;
   assign m108_13 =15'b0;

   // m108_14 = W*in
   wire signed [14:0] m108_14;
   assign m108_14 =15'b0;

   // m108_15 = W*in
   wire signed [14:0] m108_15;
   assign m108_15 =15'b0;

   // m108_16 = W*in
   wire signed [14:0] m108_16;
   assign m108_16 =15'b0;

   // m108_17 = W*in
   wire signed [14:0] m108_17;
   assign m108_17 =15'b0;

   // m108_18 = W*in
   wire signed [14:0] m108_18;
   assign m108_18 =15'b0;

   // m108_19 = W*in
   wire signed [14:0] m108_19;
   assign m108_19 ={ {4{neg108[14]}} , neg108[14:4] };

   // m108_20 = W*in
   wire signed [14:0] m108_20;
   assign m108_20 ={ {3{in108[14]}} , in108[14:3] };

   // m108_21 = W*in
   wire signed [14:0] m108_21;
   assign m108_21 =15'b0;

   // m108_22 = W*in
   wire signed [14:0] m108_22;
   assign m108_22 =15'b0;

   // m108_23 = W*in
   wire signed [14:0] m108_23;
   assign m108_23 ={ {3{in108[14]}} , in108[14:3] };

   // m108_24 = W*in
   wire signed [14:0] m108_24;
   assign m108_24 =15'b0;

   // m108_25 = W*in
   wire signed [14:0] m108_25;
   assign m108_25 =15'b0;

   // m108_26 = W*in
   wire signed [14:0] m108_26;
   assign m108_26 =15'b0;

   // m108_27 = W*in
   wire signed [14:0] m108_27;
   assign m108_27 =15'b0;

   // m108_28 = W*in
   wire signed [14:0] m108_28;
   assign m108_28 =15'b0;

   // m108_29 = W*in
   wire signed [14:0] m108_29;
   assign m108_29 =15'b0;

   // m108_30 = W*in
   wire signed [14:0] m108_30;
   assign m108_30 =15'b0;

   // m108_31 = W*in
   wire signed [14:0] m108_31;
   assign m108_31 =15'b0;

   // m108_32 = W*in
   wire signed [14:0] m108_32;
   assign m108_32 =15'b0;

   // m108_33 = W*in
   wire signed [14:0] m108_33;
   assign m108_33 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_34 = W*in
   wire signed [14:0] m108_34;
   assign m108_34 =15'b0;

   // m108_35 = W*in
   wire signed [14:0] m108_35;
   assign m108_35 =15'b0;

   // m108_36 = W*in
   wire signed [14:0] m108_36;
   assign m108_36 =15'b0;

   // m108_37 = W*in
   wire signed [14:0] m108_37;
   assign m108_37 =15'b0;

   // m108_38 = W*in
   wire signed [14:0] m108_38;
   assign m108_38 =15'b0;

   // m108_39 = W*in
   wire signed [14:0] m108_39;
   assign m108_39 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_40 = W*in
   wire signed [14:0] m108_40;
   assign m108_40 ={ {3{in108[14]}} , in108[14:3] };

   // m108_41 = W*in
   wire signed [14:0] m108_41;
   assign m108_41 =15'b0;

   // m108_42 = W*in
   wire signed [14:0] m108_42;
   assign m108_42 =15'b0;

   // m108_43 = W*in
   wire signed [14:0] m108_43;
   assign m108_43 =15'b0;

   // m108_44 = W*in
   wire signed [14:0] m108_44;
   assign m108_44 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_45 = W*in
   wire signed [14:0] m108_45;
   assign m108_45 ={ {3{in108[14]}} , in108[14:3] };

   // m108_46 = W*in
   wire signed [14:0] m108_46;
   assign m108_46 =15'b0;

   // m108_47 = W*in
   wire signed [14:0] m108_47;
   assign m108_47 =15'b0;

   // m108_48 = W*in
   wire signed [14:0] m108_48;
   assign m108_48 =15'b0;

   // m108_49 = W*in
   wire signed [14:0] m108_49;
   assign m108_49 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_50 = W*in
   wire signed [14:0] m108_50;
   assign m108_50 =15'b0;

   // m108_51 = W*in
   wire signed [14:0] m108_51;
   assign m108_51 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_52 = W*in
   wire signed [14:0] m108_52;
   assign m108_52 =15'b0;

   // m108_53 = W*in
   wire signed [14:0] m108_53;
   assign m108_53 =15'b0;

   // m108_54 = W*in
   wire signed [14:0] m108_54;
   assign m108_54 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_55 = W*in
   wire signed [14:0] m108_55;
   assign m108_55 =15'b0;

   // m108_56 = W*in
   wire signed [14:0] m108_56;
   assign m108_56 =15'b0;

   // m108_57 = W*in
   wire signed [14:0] m108_57;
   assign m108_57 =15'b0;

   // m108_58 = W*in
   wire signed [14:0] m108_58;
   assign m108_58 =15'b0;

   // m108_59 = W*in
   wire signed [14:0] m108_59;
   assign m108_59 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_60 = W*in
   wire signed [14:0] m108_60;
   assign m108_60 =15'b0;

   // m108_61 = W*in
   wire signed [14:0] m108_61;
   assign m108_61 =15'b0;

   // m108_62 = W*in
   wire signed [14:0] m108_62;
   assign m108_62 ={ {3{in108[14]}} , in108[14:3] };

   // m108_63 = W*in
   wire signed [14:0] m108_63;
   assign m108_63 =15'b0;

   // m108_64 = W*in
   wire signed [14:0] m108_64;
   assign m108_64 ={ {3{in108[14]}} , in108[14:3] };

   // m108_65 = W*in
   wire signed [14:0] m108_65;
   assign m108_65 =15'b0;

   // m108_66 = W*in
   wire signed [14:0] m108_66;
   assign m108_66 =15'b0;

   // m108_67 = W*in
   wire signed [14:0] m108_67;
   assign m108_67 =15'b0;

   // m108_68 = W*in
   wire signed [14:0] m108_68;
   assign m108_68 =15'b0;

   // m108_69 = W*in
   wire signed [14:0] m108_69;
   assign m108_69 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_70 = W*in
   wire signed [14:0] m108_70;
   assign m108_70 =15'b0;

   // m108_71 = W*in
   wire signed [14:0] m108_71;
   assign m108_71 =15'b0;

   // m108_72 = W*in
   wire signed [14:0] m108_72;
   assign m108_72 =15'b0;

   // m108_73 = W*in
   wire signed [14:0] m108_73;
   assign m108_73 =15'b0;

   // m108_74 = W*in
   wire signed [14:0] m108_74;
   assign m108_74 ={ {4{in108[14]}} , in108[14:4] };

   // m108_75 = W*in
   wire signed [14:0] m108_75;
   assign m108_75 =15'b0;

   // m108_76 = W*in
   wire signed [14:0] m108_76;
   assign m108_76 =15'b0;

   // m108_77 = W*in
   wire signed [14:0] m108_77;
   assign m108_77 =15'b0;

   // m108_78 = W*in
   wire signed [14:0] m108_78;
   assign m108_78 =15'b0;

   // m108_79 = W*in
   wire signed [14:0] m108_79;
   assign m108_79 =15'b0;

   // m108_80 = W*in
   wire signed [14:0] m108_80;
   assign m108_80 =15'b0;

   // m108_81 = W*in
   wire signed [14:0] m108_81;
   assign m108_81 =15'b0;

   // m108_82 = W*in
   wire signed [14:0] m108_82;
   assign m108_82 =15'b0;

   // m108_83 = W*in
   wire signed [14:0] m108_83;
   assign m108_83 =15'b0;

   // m108_84 = W*in
   wire signed [14:0] m108_84;
   assign m108_84 =15'b0;

   // m108_85 = W*in
   wire signed [14:0] m108_85;
   assign m108_85 =15'b0;

   // m108_86 = W*in
   wire signed [14:0] m108_86;
   assign m108_86 =15'b0;

   // m108_87 = W*in
   wire signed [14:0] m108_87;
   assign m108_87 ={ {3{in108[14]}} , in108[14:3] };

   // m108_88 = W*in
   wire signed [14:0] m108_88;
   assign m108_88 =15'b0;

   // m108_89 = W*in
   wire signed [14:0] m108_89;
   assign m108_89 =15'b0;

   // m108_90 = W*in
   wire signed [14:0] m108_90;
   assign m108_90 =15'b0;

   // m108_91 = W*in
   wire signed [14:0] m108_91;
   assign m108_91 =15'b0;

   // m108_92 = W*in
   wire signed [14:0] m108_92;
   assign m108_92 =15'b0;

   // m108_93 = W*in
   wire signed [14:0] m108_93;
   assign m108_93 =15'b0;

   // m108_94 = W*in
   wire signed [14:0] m108_94;
   assign m108_94 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_95 = W*in
   wire signed [14:0] m108_95;
   assign m108_95 ={ {3{neg108[14]}} , neg108[14:3] };

   // m108_96 = W*in
   wire signed [14:0] m108_96;
   assign m108_96 =15'b0;

   // m108_97 = W*in
   wire signed [14:0] m108_97;
   assign m108_97 =15'b0;

   // m108_98 = W*in
   wire signed [14:0] m108_98;
   assign m108_98 =15'b0;

   // m108_99 = W*in
   wire signed [14:0] m108_99;
   assign m108_99 =15'b0;

   // m108_100 = W*in
   wire signed [14:0] m108_100;
   assign m108_100 =15'b0;

   // m109_1 = W*in
   wire signed [14:0] m109_1;
   assign m109_1 =15'b0;

   // m109_2 = W*in
   wire signed [14:0] m109_2;
   assign m109_2 =15'b0;

   // m109_3 = W*in
   wire signed [14:0] m109_3;
   assign m109_3 =15'b0;

   // m109_4 = W*in
   wire signed [14:0] m109_4;
   assign m109_4 =15'b0;

   // m109_5 = W*in
   wire signed [14:0] m109_5;
   assign m109_5 =15'b0;

   // m109_6 = W*in
   wire signed [14:0] m109_6;
   assign m109_6 =15'b0;

   // m109_7 = W*in
   wire signed [14:0] m109_7;
   assign m109_7 =15'b0;

   // m109_8 = W*in
   wire signed [14:0] m109_8;
   assign m109_8 =15'b0;

   // m109_9 = W*in
   wire signed [14:0] m109_9;
   assign m109_9 =15'b0;

   // m109_10 = W*in
   wire signed [14:0] m109_10;
   assign m109_10 ={ {3{in109[14]}} , in109[14:3] };

   // m109_11 = W*in
   wire signed [14:0] m109_11;
   assign m109_11 =15'b0;

   // m109_12 = W*in
   wire signed [14:0] m109_12;
   assign m109_12 =15'b0;

   // m109_13 = W*in
   wire signed [14:0] m109_13;
   assign m109_13 =15'b0;

   // m109_14 = W*in
   wire signed [14:0] m109_14;
   assign m109_14 =15'b0;

   // m109_15 = W*in
   wire signed [14:0] m109_15;
   assign m109_15 =15'b0;

   // m109_16 = W*in
   wire signed [14:0] m109_16;
   assign m109_16 =15'b0;

   // m109_17 = W*in
   wire signed [14:0] m109_17;
   assign m109_17 =15'b0;

   // m109_18 = W*in
   wire signed [14:0] m109_18;
   assign m109_18 =15'b0;

   // m109_19 = W*in
   wire signed [14:0] m109_19;
   assign m109_19 =15'b0;

   // m109_20 = W*in
   wire signed [14:0] m109_20;
   assign m109_20 =15'b0;

   // m109_21 = W*in
   wire signed [14:0] m109_21;
   assign m109_21 =15'b0;

   // m109_22 = W*in
   wire signed [14:0] m109_22;
   assign m109_22 =15'b0;

   // m109_23 = W*in
   wire signed [14:0] m109_23;
   assign m109_23 =15'b0;

   // m109_24 = W*in
   wire signed [14:0] m109_24;
   assign m109_24 =15'b0;

   // m109_25 = W*in
   wire signed [14:0] m109_25;
   assign m109_25 =15'b0;

   // m109_26 = W*in
   wire signed [14:0] m109_26;
   assign m109_26 =15'b0;

   // m109_27 = W*in
   wire signed [14:0] m109_27;
   assign m109_27 =15'b0;

   // m109_28 = W*in
   wire signed [14:0] m109_28;
   assign m109_28 =15'b0;

   // m109_29 = W*in
   wire signed [14:0] m109_29;
   assign m109_29 =15'b0;

   // m109_30 = W*in
   wire signed [14:0] m109_30;
   assign m109_30 ={ {3{neg109[14]}} , neg109[14:3] };

   // m109_31 = W*in
   wire signed [14:0] m109_31;
   assign m109_31 =15'b0;

   // m109_32 = W*in
   wire signed [14:0] m109_32;
   assign m109_32 =15'b0;

   // m109_33 = W*in
   wire signed [14:0] m109_33;
   assign m109_33 =15'b0;

   // m109_34 = W*in
   wire signed [14:0] m109_34;
   assign m109_34 =15'b0;

   // m109_35 = W*in
   wire signed [14:0] m109_35;
   assign m109_35 =15'b0;

   // m109_36 = W*in
   wire signed [14:0] m109_36;
   assign m109_36 =15'b0;

   // m109_37 = W*in
   wire signed [14:0] m109_37;
   assign m109_37 ={ {3{in109[14]}} , in109[14:3] };

   // m109_38 = W*in
   wire signed [14:0] m109_38;
   assign m109_38 =15'b0;

   // m109_39 = W*in
   wire signed [14:0] m109_39;
   assign m109_39 =15'b0;

   // m109_40 = W*in
   wire signed [14:0] m109_40;
   assign m109_40 =15'b0;

   // m109_41 = W*in
   wire signed [14:0] m109_41;
   assign m109_41 =15'b0;

   // m109_42 = W*in
   wire signed [14:0] m109_42;
   assign m109_42 =15'b0;

   // m109_43 = W*in
   wire signed [14:0] m109_43;
   assign m109_43 =15'b0;

   // m109_44 = W*in
   wire signed [14:0] m109_44;
   assign m109_44 =15'b0;

   // m109_45 = W*in
   wire signed [14:0] m109_45;
   assign m109_45 ={ {4{in109[14]}} , in109[14:4] };

   // m109_46 = W*in
   wire signed [14:0] m109_46;
   assign m109_46 =15'b0;

   // m109_47 = W*in
   wire signed [14:0] m109_47;
   assign m109_47 =15'b0;

   // m109_48 = W*in
   wire signed [14:0] m109_48;
   assign m109_48 =15'b0;

   // m109_49 = W*in
   wire signed [14:0] m109_49;
   assign m109_49 =15'b0;

   // m109_50 = W*in
   wire signed [14:0] m109_50;
   assign m109_50 =15'b0;

   // m109_51 = W*in
   wire signed [14:0] m109_51;
   assign m109_51 =15'b0;

   // m109_52 = W*in
   wire signed [14:0] m109_52;
   assign m109_52 =15'b0;

   // m109_53 = W*in
   wire signed [14:0] m109_53;
   assign m109_53 =15'b0;

   // m109_54 = W*in
   wire signed [14:0] m109_54;
   assign m109_54 =15'b0;

   // m109_55 = W*in
   wire signed [14:0] m109_55;
   assign m109_55 =15'b0;

   // m109_56 = W*in
   wire signed [14:0] m109_56;
   assign m109_56 =15'b0;

   // m109_57 = W*in
   wire signed [14:0] m109_57;
   assign m109_57 =15'b0;

   // m109_58 = W*in
   wire signed [14:0] m109_58;
   assign m109_58 =15'b0;

   // m109_59 = W*in
   wire signed [14:0] m109_59;
   assign m109_59 =15'b0;

   // m109_60 = W*in
   wire signed [14:0] m109_60;
   assign m109_60 =15'b0;

   // m109_61 = W*in
   wire signed [14:0] m109_61;
   assign m109_61 ={ {3{in109[14]}} , in109[14:3] };

   // m109_62 = W*in
   wire signed [14:0] m109_62;
   assign m109_62 =15'b0;

   // m109_63 = W*in
   wire signed [14:0] m109_63;
   assign m109_63 ={ {3{in109[14]}} , in109[14:3] };

   // m109_64 = W*in
   wire signed [14:0] m109_64;
   assign m109_64 =15'b0;

   // m109_65 = W*in
   wire signed [14:0] m109_65;
   assign m109_65 =15'b0;

   // m109_66 = W*in
   wire signed [14:0] m109_66;
   assign m109_66 =15'b0;

   // m109_67 = W*in
   wire signed [14:0] m109_67;
   assign m109_67 =15'b0;

   // m109_68 = W*in
   wire signed [14:0] m109_68;
   assign m109_68 =15'b0;

   // m109_69 = W*in
   wire signed [14:0] m109_69;
   assign m109_69 =15'b0;

   // m109_70 = W*in
   wire signed [14:0] m109_70;
   assign m109_70 =15'b0;

   // m109_71 = W*in
   wire signed [14:0] m109_71;
   assign m109_71 ={ {3{in109[14]}} , in109[14:3] };

   // m109_72 = W*in
   wire signed [14:0] m109_72;
   assign m109_72 =15'b0;

   // m109_73 = W*in
   wire signed [14:0] m109_73;
   assign m109_73 =15'b0;

   // m109_74 = W*in
   wire signed [14:0] m109_74;
   assign m109_74 =15'b0;

   // m109_75 = W*in
   wire signed [14:0] m109_75;
   assign m109_75 =15'b0;

   // m109_76 = W*in
   wire signed [14:0] m109_76;
   assign m109_76 =15'b0;

   // m109_77 = W*in
   wire signed [14:0] m109_77;
   assign m109_77 =15'b0;

   // m109_78 = W*in
   wire signed [14:0] m109_78;
   assign m109_78 =15'b0;

   // m109_79 = W*in
   wire signed [14:0] m109_79;
   assign m109_79 =15'b0;

   // m109_80 = W*in
   wire signed [14:0] m109_80;
   assign m109_80 =15'b0;

   // m109_81 = W*in
   wire signed [14:0] m109_81;
   assign m109_81 =15'b0;

   // m109_82 = W*in
   wire signed [14:0] m109_82;
   assign m109_82 ={ {4{neg109[14]}} , neg109[14:4] };

   // m109_83 = W*in
   wire signed [14:0] m109_83;
   assign m109_83 =15'b0;

   // m109_84 = W*in
   wire signed [14:0] m109_84;
   assign m109_84 =15'b0;

   // m109_85 = W*in
   wire signed [14:0] m109_85;
   assign m109_85 =15'b0;

   // m109_86 = W*in
   wire signed [14:0] m109_86;
   assign m109_86 ={ {3{neg109[14]}} , neg109[14:3] };

   // m109_87 = W*in
   wire signed [14:0] m109_87;
   assign m109_87 =15'b0;

   // m109_88 = W*in
   wire signed [14:0] m109_88;
   assign m109_88 ={ {3{neg109[14]}} , neg109[14:3] };

   // m109_89 = W*in
   wire signed [14:0] m109_89;
   assign m109_89 =15'b0;

   // m109_90 = W*in
   wire signed [14:0] m109_90;
   assign m109_90 =15'b0;

   // m109_91 = W*in
   wire signed [14:0] m109_91;
   assign m109_91 =15'b0;

   // m109_92 = W*in
   wire signed [14:0] m109_92;
   assign m109_92 =15'b0;

   // m109_93 = W*in
   wire signed [14:0] m109_93;
   assign m109_93 =15'b0;

   // m109_94 = W*in
   wire signed [14:0] m109_94;
   assign m109_94 =15'b0;

   // m109_95 = W*in
   wire signed [14:0] m109_95;
   assign m109_95 =15'b0;

   // m109_96 = W*in
   wire signed [14:0] m109_96;
   assign m109_96 =15'b0;

   // m109_97 = W*in
   wire signed [14:0] m109_97;
   assign m109_97 =15'b0;

   // m109_98 = W*in
   wire signed [14:0] m109_98;
   assign m109_98 =15'b0;

   // m109_99 = W*in
   wire signed [14:0] m109_99;
   assign m109_99 =15'b0;

   // m109_100 = W*in
   wire signed [14:0] m109_100;
   assign m109_100 =15'b0;

   // m110_1 = W*in
   wire signed [14:0] m110_1;
   assign m110_1 =15'b0;

   // m110_2 = W*in
   wire signed [14:0] m110_2;
   assign m110_2 =15'b0;

   // m110_3 = W*in
   wire signed [14:0] m110_3;
   assign m110_3 =15'b0;

   // m110_4 = W*in
   wire signed [14:0] m110_4;
   assign m110_4 =15'b0;

   // m110_5 = W*in
   wire signed [14:0] m110_5;
   assign m110_5 ={ {4{neg110[14]}} , neg110[14:4] };

   // m110_6 = W*in
   wire signed [14:0] m110_6;
   assign m110_6 ={ {4{in110[14]}} , in110[14:4] };

   // m110_7 = W*in
   wire signed [14:0] m110_7;
   assign m110_7 =15'b0;

   // m110_8 = W*in
   wire signed [14:0] m110_8;
   assign m110_8 =15'b0;

   // m110_9 = W*in
   wire signed [14:0] m110_9;
   assign m110_9 =15'b0;

   // m110_10 = W*in
   wire signed [14:0] m110_10;
   assign m110_10 =15'b0;

   // m110_11 = W*in
   wire signed [14:0] m110_11;
   assign m110_11 =15'b0;

   // m110_12 = W*in
   wire signed [14:0] m110_12;
   assign m110_12 =15'b0;

   // m110_13 = W*in
   wire signed [14:0] m110_13;
   assign m110_13 =15'b0;

   // m110_14 = W*in
   wire signed [14:0] m110_14;
   assign m110_14 =15'b0;

   // m110_15 = W*in
   wire signed [14:0] m110_15;
   assign m110_15 =15'b0;

   // m110_16 = W*in
   wire signed [14:0] m110_16;
   assign m110_16 =15'b0;

   // m110_17 = W*in
   wire signed [14:0] m110_17;
   assign m110_17 =15'b0;

   // m110_18 = W*in
   wire signed [14:0] m110_18;
   assign m110_18 =15'b0;

   // m110_19 = W*in
   wire signed [14:0] m110_19;
   assign m110_19 =15'b0;

   // m110_20 = W*in
   wire signed [14:0] m110_20;
   assign m110_20 =15'b0;

   // m110_21 = W*in
   wire signed [14:0] m110_21;
   assign m110_21 ={ {4{in110[14]}} , in110[14:4] };

   // m110_22 = W*in
   wire signed [14:0] m110_22;
   assign m110_22 =15'b0;

   // m110_23 = W*in
   wire signed [14:0] m110_23;
   assign m110_23 =15'b0;

   // m110_24 = W*in
   wire signed [14:0] m110_24;
   assign m110_24 =15'b0;

   // m110_25 = W*in
   wire signed [14:0] m110_25;
   assign m110_25 ={ {4{in110[14]}} , in110[14:4] };

   // m110_26 = W*in
   wire signed [14:0] m110_26;
   assign m110_26 =15'b0;

   // m110_27 = W*in
   wire signed [14:0] m110_27;
   assign m110_27 ={ {4{neg110[14]}} , neg110[14:4] };

   // m110_28 = W*in
   wire signed [14:0] m110_28;
   assign m110_28 =15'b0;

   // m110_29 = W*in
   wire signed [14:0] m110_29;
   assign m110_29 =15'b0;

   // m110_30 = W*in
   wire signed [14:0] m110_30;
   assign m110_30 =15'b0;

   // m110_31 = W*in
   wire signed [14:0] m110_31;
   assign m110_31 =15'b0;

   // m110_32 = W*in
   wire signed [14:0] m110_32;
   assign m110_32 =15'b0;

   // m110_33 = W*in
   wire signed [14:0] m110_33;
   assign m110_33 ={ {4{neg110[14]}} , neg110[14:4] };

   // m110_34 = W*in
   wire signed [14:0] m110_34;
   assign m110_34 =15'b0;

   // m110_35 = W*in
   wire signed [14:0] m110_35;
   assign m110_35 =15'b0;

   // m110_36 = W*in
   wire signed [14:0] m110_36;
   assign m110_36 =15'b0;

   // m110_37 = W*in
   wire signed [14:0] m110_37;
   assign m110_37 =15'b0;

   // m110_38 = W*in
   wire signed [14:0] m110_38;
   assign m110_38 =15'b0;

   // m110_39 = W*in
   wire signed [14:0] m110_39;
   assign m110_39 =15'b0;

   // m110_40 = W*in
   wire signed [14:0] m110_40;
   assign m110_40 =15'b0;

   // m110_41 = W*in
   wire signed [14:0] m110_41;
   assign m110_41 =15'b0;

   // m110_42 = W*in
   wire signed [14:0] m110_42;
   assign m110_42 =15'b0;

   // m110_43 = W*in
   wire signed [14:0] m110_43;
   assign m110_43 =15'b0;

   // m110_44 = W*in
   wire signed [14:0] m110_44;
   assign m110_44 =15'b0;

   // m110_45 = W*in
   wire signed [14:0] m110_45;
   assign m110_45 =15'b0;

   // m110_46 = W*in
   wire signed [14:0] m110_46;
   assign m110_46 =15'b0;

   // m110_47 = W*in
   wire signed [14:0] m110_47;
   assign m110_47 =15'b0;

   // m110_48 = W*in
   wire signed [14:0] m110_48;
   assign m110_48 =15'b0;

   // m110_49 = W*in
   wire signed [14:0] m110_49;
   assign m110_49 =15'b0;

   // m110_50 = W*in
   wire signed [14:0] m110_50;
   assign m110_50 =15'b0;

   // m110_51 = W*in
   wire signed [14:0] m110_51;
   assign m110_51 =15'b0;

   // m110_52 = W*in
   wire signed [14:0] m110_52;
   assign m110_52 =15'b0;

   // m110_53 = W*in
   wire signed [14:0] m110_53;
   assign m110_53 =15'b0;

   // m110_54 = W*in
   wire signed [14:0] m110_54;
   assign m110_54 =15'b0;

   // m110_55 = W*in
   wire signed [14:0] m110_55;
   assign m110_55 =15'b0;

   // m110_56 = W*in
   wire signed [14:0] m110_56;
   assign m110_56 =15'b0;

   // m110_57 = W*in
   wire signed [14:0] m110_57;
   assign m110_57 ={ {4{neg110[14]}} , neg110[14:4] };

   // m110_58 = W*in
   wire signed [14:0] m110_58;
   assign m110_58 =15'b0;

   // m110_59 = W*in
   wire signed [14:0] m110_59;
   assign m110_59 =15'b0;

   // m110_60 = W*in
   wire signed [14:0] m110_60;
   assign m110_60 ={ {4{in110[14]}} , in110[14:4] };

   // m110_61 = W*in
   wire signed [14:0] m110_61;
   assign m110_61 =15'b0;

   // m110_62 = W*in
   wire signed [14:0] m110_62;
   assign m110_62 =15'b0;

   // m110_63 = W*in
   wire signed [14:0] m110_63;
   assign m110_63 =15'b0;

   // m110_64 = W*in
   wire signed [14:0] m110_64;
   assign m110_64 ={ {4{in110[14]}} , in110[14:4] };

   // m110_65 = W*in
   wire signed [14:0] m110_65;
   assign m110_65 ={ {4{neg110[14]}} , neg110[14:4] };

   // m110_66 = W*in
   wire signed [14:0] m110_66;
   assign m110_66 =15'b0;

   // m110_67 = W*in
   wire signed [14:0] m110_67;
   assign m110_67 =15'b0;

   // m110_68 = W*in
   wire signed [14:0] m110_68;
   assign m110_68 ={ {4{neg110[14]}} , neg110[14:4] };

   // m110_69 = W*in
   wire signed [14:0] m110_69;
   assign m110_69 ={ {4{in110[14]}} , in110[14:4] };

   // m110_70 = W*in
   wire signed [14:0] m110_70;
   assign m110_70 =15'b0;

   // m110_71 = W*in
   wire signed [14:0] m110_71;
   assign m110_71 =15'b0;

   // m110_72 = W*in
   wire signed [14:0] m110_72;
   assign m110_72 =15'b0;

   // m110_73 = W*in
   wire signed [14:0] m110_73;
   assign m110_73 =15'b0;

   // m110_74 = W*in
   wire signed [14:0] m110_74;
   assign m110_74 =15'b0;

   // m110_75 = W*in
   wire signed [14:0] m110_75;
   assign m110_75 =15'b0;

   // m110_76 = W*in
   wire signed [14:0] m110_76;
   assign m110_76 =15'b0;

   // m110_77 = W*in
   wire signed [14:0] m110_77;
   assign m110_77 ={ {4{in110[14]}} , in110[14:4] };

   // m110_78 = W*in
   wire signed [14:0] m110_78;
   assign m110_78 =15'b0;

   // m110_79 = W*in
   wire signed [14:0] m110_79;
   assign m110_79 =15'b0;

   // m110_80 = W*in
   wire signed [14:0] m110_80;
   assign m110_80 =15'b0;

   // m110_81 = W*in
   wire signed [14:0] m110_81;
   assign m110_81 =15'b0;

   // m110_82 = W*in
   wire signed [14:0] m110_82;
   assign m110_82 =15'b0;

   // m110_83 = W*in
   wire signed [14:0] m110_83;
   assign m110_83 =15'b0;

   // m110_84 = W*in
   wire signed [14:0] m110_84;
   assign m110_84 =15'b0;

   // m110_85 = W*in
   wire signed [14:0] m110_85;
   assign m110_85 =15'b0;

   // m110_86 = W*in
   wire signed [14:0] m110_86;
   assign m110_86 =15'b0;

   // m110_87 = W*in
   wire signed [14:0] m110_87;
   assign m110_87 =15'b0;

   // m110_88 = W*in
   wire signed [14:0] m110_88;
   assign m110_88 =15'b0;

   // m110_89 = W*in
   wire signed [14:0] m110_89;
   assign m110_89 =15'b0;

   // m110_90 = W*in
   wire signed [14:0] m110_90;
   assign m110_90 =15'b0;

   // m110_91 = W*in
   wire signed [14:0] m110_91;
   assign m110_91 =15'b0;

   // m110_92 = W*in
   wire signed [14:0] m110_92;
   assign m110_92 =15'b0;

   // m110_93 = W*in
   wire signed [14:0] m110_93;
   assign m110_93 =15'b0;

   // m110_94 = W*in
   wire signed [14:0] m110_94;
   assign m110_94 =15'b0;

   // m110_95 = W*in
   wire signed [14:0] m110_95;
   assign m110_95 =15'b0;

   // m110_96 = W*in
   wire signed [14:0] m110_96;
   assign m110_96 =15'b0;

   // m110_97 = W*in
   wire signed [14:0] m110_97;
   assign m110_97 =15'b0;

   // m110_98 = W*in
   wire signed [14:0] m110_98;
   assign m110_98 =15'b0;

   // m110_99 = W*in
   wire signed [14:0] m110_99;
   assign m110_99 =15'b0;

   // m110_100 = W*in
   wire signed [14:0] m110_100;
   assign m110_100 =15'b0;

   // m111_1 = W*in
   wire signed [14:0] m111_1;
   assign m111_1 =15'b0;

   // m111_2 = W*in
   wire signed [14:0] m111_2;
   assign m111_2 ={ {3{in111[14]}} , in111[14:3] };

   // m111_3 = W*in
   wire signed [14:0] m111_3;
   assign m111_3 =15'b0;

   // m111_4 = W*in
   wire signed [14:0] m111_4;
   assign m111_4 =15'b0;

   // m111_5 = W*in
   wire signed [14:0] m111_5;
   assign m111_5 =15'b0;

   // m111_6 = W*in
   wire signed [14:0] m111_6;
   assign m111_6 =15'b0;

   // m111_7 = W*in
   wire signed [14:0] m111_7;
   assign m111_7 ={ {3{in111[14]}} , in111[14:3] };

   // m111_8 = W*in
   wire signed [14:0] m111_8;
   assign m111_8 =15'b0;

   // m111_9 = W*in
   wire signed [14:0] m111_9;
   assign m111_9 =15'b0;

   // m111_10 = W*in
   wire signed [14:0] m111_10;
   assign m111_10 ={ {3{in111[14]}} , in111[14:3] };

   // m111_11 = W*in
   wire signed [14:0] m111_11;
   assign m111_11 =15'b0;

   // m111_12 = W*in
   wire signed [14:0] m111_12;
   assign m111_12 ={ {3{in111[14]}} , in111[14:3] };

   // m111_13 = W*in
   wire signed [14:0] m111_13;
   assign m111_13 =15'b0;

   // m111_14 = W*in
   wire signed [14:0] m111_14;
   assign m111_14 =15'b0;

   // m111_15 = W*in
   wire signed [14:0] m111_15;
   assign m111_15 =15'b0;

   // m111_16 = W*in
   wire signed [14:0] m111_16;
   assign m111_16 =15'b0;

   // m111_17 = W*in
   wire signed [14:0] m111_17;
   assign m111_17 =15'b0;

   // m111_18 = W*in
   wire signed [14:0] m111_18;
   assign m111_18 =15'b0;

   // m111_19 = W*in
   wire signed [14:0] m111_19;
   assign m111_19 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_20 = W*in
   wire signed [14:0] m111_20;
   assign m111_20 =15'b0;

   // m111_21 = W*in
   wire signed [14:0] m111_21;
   assign m111_21 =15'b0;

   // m111_22 = W*in
   wire signed [14:0] m111_22;
   assign m111_22 =15'b0;

   // m111_23 = W*in
   wire signed [14:0] m111_23;
   assign m111_23 =15'b0;

   // m111_24 = W*in
   wire signed [14:0] m111_24;
   assign m111_24 =15'b0;

   // m111_25 = W*in
   wire signed [14:0] m111_25;
   assign m111_25 ={ {4{in111[14]}} , in111[14:4] };

   // m111_26 = W*in
   wire signed [14:0] m111_26;
   assign m111_26 ={ {4{neg111[14]}} , neg111[14:4] };

   // m111_27 = W*in
   wire signed [14:0] m111_27;
   assign m111_27 ={ {3{in111[14]}} , in111[14:3] };

   // m111_28 = W*in
   wire signed [14:0] m111_28;
   assign m111_28 =15'b0;

   // m111_29 = W*in
   wire signed [14:0] m111_29;
   assign m111_29 =15'b0;

   // m111_30 = W*in
   wire signed [14:0] m111_30;
   assign m111_30 =15'b0;

   // m111_31 = W*in
   wire signed [14:0] m111_31;
   assign m111_31 =15'b0;

   // m111_32 = W*in
   wire signed [14:0] m111_32;
   assign m111_32 =15'b0;

   // m111_33 = W*in
   wire signed [14:0] m111_33;
   assign m111_33 ={ {4{in111[14]}} , in111[14:4] };

   // m111_34 = W*in
   wire signed [14:0] m111_34;
   assign m111_34 ={ {3{in111[14]}} , in111[14:3] };

   // m111_35 = W*in
   wire signed [14:0] m111_35;
   assign m111_35 =15'b0;

   // m111_36 = W*in
   wire signed [14:0] m111_36;
   assign m111_36 =15'b0;

   // m111_37 = W*in
   wire signed [14:0] m111_37;
   assign m111_37 =15'b0;

   // m111_38 = W*in
   wire signed [14:0] m111_38;
   assign m111_38 ={ {3{in111[14]}} , in111[14:3] };

   // m111_39 = W*in
   wire signed [14:0] m111_39;
   assign m111_39 ={ {3{in111[14]}} , in111[14:3] };

   // m111_40 = W*in
   wire signed [14:0] m111_40;
   assign m111_40 =15'b0;

   // m111_41 = W*in
   wire signed [14:0] m111_41;
   assign m111_41 =15'b0;

   // m111_42 = W*in
   wire signed [14:0] m111_42;
   assign m111_42 =15'b0;

   // m111_43 = W*in
   wire signed [14:0] m111_43;
   assign m111_43 =15'b0;

   // m111_44 = W*in
   wire signed [14:0] m111_44;
   assign m111_44 ={ {3{in111[14]}} , in111[14:3] };

   // m111_45 = W*in
   wire signed [14:0] m111_45;
   assign m111_45 =15'b0;

   // m111_46 = W*in
   wire signed [14:0] m111_46;
   assign m111_46 =15'b0;

   // m111_47 = W*in
   wire signed [14:0] m111_47;
   assign m111_47 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_48 = W*in
   wire signed [14:0] m111_48;
   assign m111_48 =15'b0;

   // m111_49 = W*in
   wire signed [14:0] m111_49;
   assign m111_49 =15'b0;

   // m111_50 = W*in
   wire signed [14:0] m111_50;
   assign m111_50 =15'b0;

   // m111_51 = W*in
   wire signed [14:0] m111_51;
   assign m111_51 =15'b0;

   // m111_52 = W*in
   wire signed [14:0] m111_52;
   assign m111_52 ={ {3{in111[14]}} , in111[14:3] };

   // m111_53 = W*in
   wire signed [14:0] m111_53;
   assign m111_53 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_54 = W*in
   wire signed [14:0] m111_54;
   assign m111_54 =15'b0;

   // m111_55 = W*in
   wire signed [14:0] m111_55;
   assign m111_55 =15'b0;

   // m111_56 = W*in
   wire signed [14:0] m111_56;
   assign m111_56 =15'b0;

   // m111_57 = W*in
   wire signed [14:0] m111_57;
   assign m111_57 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_58 = W*in
   wire signed [14:0] m111_58;
   assign m111_58 ={ {4{neg111[14]}} , neg111[14:4] };

   // m111_59 = W*in
   wire signed [14:0] m111_59;
   assign m111_59 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_60 = W*in
   wire signed [14:0] m111_60;
   assign m111_60 =15'b0;

   // m111_61 = W*in
   wire signed [14:0] m111_61;
   assign m111_61 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_62 = W*in
   wire signed [14:0] m111_62;
   assign m111_62 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_63 = W*in
   wire signed [14:0] m111_63;
   assign m111_63 =15'b0;

   // m111_64 = W*in
   wire signed [14:0] m111_64;
   assign m111_64 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_65 = W*in
   wire signed [14:0] m111_65;
   assign m111_65 ={ {3{in111[14]}} , in111[14:3] };

   // m111_66 = W*in
   wire signed [14:0] m111_66;
   assign m111_66 ={ {3{in111[14]}} , in111[14:3] };

   // m111_67 = W*in
   wire signed [14:0] m111_67;
   assign m111_67 =15'b0;

   // m111_68 = W*in
   wire signed [14:0] m111_68;
   assign m111_68 =15'b0;

   // m111_69 = W*in
   wire signed [14:0] m111_69;
   assign m111_69 =15'b0;

   // m111_70 = W*in
   wire signed [14:0] m111_70;
   assign m111_70 =15'b0;

   // m111_71 = W*in
   wire signed [14:0] m111_71;
   assign m111_71 =15'b0;

   // m111_72 = W*in
   wire signed [14:0] m111_72;
   assign m111_72 =15'b0;

   // m111_73 = W*in
   wire signed [14:0] m111_73;
   assign m111_73 =15'b0;

   // m111_74 = W*in
   wire signed [14:0] m111_74;
   assign m111_74 =15'b0;

   // m111_75 = W*in
   wire signed [14:0] m111_75;
   assign m111_75 =15'b0;

   // m111_76 = W*in
   wire signed [14:0] m111_76;
   assign m111_76 =15'b0;

   // m111_77 = W*in
   wire signed [14:0] m111_77;
   assign m111_77 =15'b0;

   // m111_78 = W*in
   wire signed [14:0] m111_78;
   assign m111_78 =15'b0;

   // m111_79 = W*in
   wire signed [14:0] m111_79;
   assign m111_79 =15'b0;

   // m111_80 = W*in
   wire signed [14:0] m111_80;
   assign m111_80 ={ {3{in111[14]}} , in111[14:3] };

   // m111_81 = W*in
   wire signed [14:0] m111_81;
   assign m111_81 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_82 = W*in
   wire signed [14:0] m111_82;
   assign m111_82 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_83 = W*in
   wire signed [14:0] m111_83;
   assign m111_83 =15'b0;

   // m111_84 = W*in
   wire signed [14:0] m111_84;
   assign m111_84 ={ {3{in111[14]}} , in111[14:3] };

   // m111_85 = W*in
   wire signed [14:0] m111_85;
   assign m111_85 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_86 = W*in
   wire signed [14:0] m111_86;
   assign m111_86 =15'b0;

   // m111_87 = W*in
   wire signed [14:0] m111_87;
   assign m111_87 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_88 = W*in
   wire signed [14:0] m111_88;
   assign m111_88 =15'b0;

   // m111_89 = W*in
   wire signed [14:0] m111_89;
   assign m111_89 =15'b0;

   // m111_90 = W*in
   wire signed [14:0] m111_90;
   assign m111_90 ={ {3{in111[14]}} , in111[14:3] };

   // m111_91 = W*in
   wire signed [14:0] m111_91;
   assign m111_91 =15'b0;

   // m111_92 = W*in
   wire signed [14:0] m111_92;
   assign m111_92 ={ {3{neg111[14]}} , neg111[14:3] };

   // m111_93 = W*in
   wire signed [14:0] m111_93;
   assign m111_93 =15'b0;

   // m111_94 = W*in
   wire signed [14:0] m111_94;
   assign m111_94 =15'b0;

   // m111_95 = W*in
   wire signed [14:0] m111_95;
   assign m111_95 =15'b0;

   // m111_96 = W*in
   wire signed [14:0] m111_96;
   assign m111_96 =15'b0;

   // m111_97 = W*in
   wire signed [14:0] m111_97;
   assign m111_97 =15'b0;

   // m111_98 = W*in
   wire signed [14:0] m111_98;
   assign m111_98 =15'b0;

   // m111_99 = W*in
   wire signed [14:0] m111_99;
   assign m111_99 =15'b0;

   // m111_100 = W*in
   wire signed [14:0] m111_100;
   assign m111_100 =15'b0;

   // m112_1 = W*in
   wire signed [14:0] m112_1;
   assign m112_1 =15'b0;

   // m112_2 = W*in
   wire signed [14:0] m112_2;
   assign m112_2 =15'b0;

   // m112_3 = W*in
   wire signed [14:0] m112_3;
   assign m112_3 =15'b0;

   // m112_4 = W*in
   wire signed [14:0] m112_4;
   assign m112_4 =15'b0;

   // m112_5 = W*in
   wire signed [14:0] m112_5;
   assign m112_5 =15'b0;

   // m112_6 = W*in
   wire signed [14:0] m112_6;
   assign m112_6 =15'b0;

   // m112_7 = W*in
   wire signed [14:0] m112_7;
   assign m112_7 =15'b0;

   // m112_8 = W*in
   wire signed [14:0] m112_8;
   assign m112_8 =15'b0;

   // m112_9 = W*in
   wire signed [14:0] m112_9;
   assign m112_9 =15'b0;

   // m112_10 = W*in
   wire signed [14:0] m112_10;
   assign m112_10 ={ {3{in112[14]}} , in112[14:3] };

   // m112_11 = W*in
   wire signed [14:0] m112_11;
   assign m112_11 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_12 = W*in
   wire signed [14:0] m112_12;
   assign m112_12 =15'b0;

   // m112_13 = W*in
   wire signed [14:0] m112_13;
   assign m112_13 ={ {3{in112[14]}} , in112[14:3] };

   // m112_14 = W*in
   wire signed [14:0] m112_14;
   assign m112_14 =15'b0;

   // m112_15 = W*in
   wire signed [14:0] m112_15;
   assign m112_15 =15'b0;

   // m112_16 = W*in
   wire signed [14:0] m112_16;
   assign m112_16 =15'b0;

   // m112_17 = W*in
   wire signed [14:0] m112_17;
   assign m112_17 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_18 = W*in
   wire signed [14:0] m112_18;
   assign m112_18 =15'b0;

   // m112_19 = W*in
   wire signed [14:0] m112_19;
   assign m112_19 ={ {4{neg112[14]}} , neg112[14:4] };

   // m112_20 = W*in
   wire signed [14:0] m112_20;
   assign m112_20 ={ {4{neg112[14]}} , neg112[14:4] };

   // m112_21 = W*in
   wire signed [14:0] m112_21;
   assign m112_21 ={ {4{neg112[14]}} , neg112[14:4] };

   // m112_22 = W*in
   wire signed [14:0] m112_22;
   assign m112_22 =15'b0;

   // m112_23 = W*in
   wire signed [14:0] m112_23;
   assign m112_23 =15'b0;

   // m112_24 = W*in
   wire signed [14:0] m112_24;
   assign m112_24 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_25 = W*in
   wire signed [14:0] m112_25;
   assign m112_25 =15'b0;

   // m112_26 = W*in
   wire signed [14:0] m112_26;
   assign m112_26 =15'b0;

   // m112_27 = W*in
   wire signed [14:0] m112_27;
   assign m112_27 ={ {4{in112[14]}} , in112[14:4] };

   // m112_28 = W*in
   wire signed [14:0] m112_28;
   assign m112_28 ={ {4{neg112[14]}} , neg112[14:4] };

   // m112_29 = W*in
   wire signed [14:0] m112_29;
   assign m112_29 ={ {3{in112[14]}} , in112[14:3] };

   // m112_30 = W*in
   wire signed [14:0] m112_30;
   assign m112_30 =15'b0;

   // m112_31 = W*in
   wire signed [14:0] m112_31;
   assign m112_31 =15'b0;

   // m112_32 = W*in
   wire signed [14:0] m112_32;
   assign m112_32 =15'b0;

   // m112_33 = W*in
   wire signed [14:0] m112_33;
   assign m112_33 =15'b0;

   // m112_34 = W*in
   wire signed [14:0] m112_34;
   assign m112_34 =15'b0;

   // m112_35 = W*in
   wire signed [14:0] m112_35;
   assign m112_35 =15'b0;

   // m112_36 = W*in
   wire signed [14:0] m112_36;
   assign m112_36 =15'b0;

   // m112_37 = W*in
   wire signed [14:0] m112_37;
   assign m112_37 =15'b0;

   // m112_38 = W*in
   wire signed [14:0] m112_38;
   assign m112_38 ={ {3{in112[14]}} , in112[14:3] };

   // m112_39 = W*in
   wire signed [14:0] m112_39;
   assign m112_39 =15'b0;

   // m112_40 = W*in
   wire signed [14:0] m112_40;
   assign m112_40 =15'b0;

   // m112_41 = W*in
   wire signed [14:0] m112_41;
   assign m112_41 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_42 = W*in
   wire signed [14:0] m112_42;
   assign m112_42 =15'b0;

   // m112_43 = W*in
   wire signed [14:0] m112_43;
   assign m112_43 =15'b0;

   // m112_44 = W*in
   wire signed [14:0] m112_44;
   assign m112_44 =15'b0;

   // m112_45 = W*in
   wire signed [14:0] m112_45;
   assign m112_45 =15'b0;

   // m112_46 = W*in
   wire signed [14:0] m112_46;
   assign m112_46 =15'b0;

   // m112_47 = W*in
   wire signed [14:0] m112_47;
   assign m112_47 =15'b0;

   // m112_48 = W*in
   wire signed [14:0] m112_48;
   assign m112_48 =15'b0;

   // m112_49 = W*in
   wire signed [14:0] m112_49;
   assign m112_49 =15'b0;

   // m112_50 = W*in
   wire signed [14:0] m112_50;
   assign m112_50 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_51 = W*in
   wire signed [14:0] m112_51;
   assign m112_51 =15'b0;

   // m112_52 = W*in
   wire signed [14:0] m112_52;
   assign m112_52 =15'b0;

   // m112_53 = W*in
   wire signed [14:0] m112_53;
   assign m112_53 =15'b0;

   // m112_54 = W*in
   wire signed [14:0] m112_54;
   assign m112_54 =15'b0;

   // m112_55 = W*in
   wire signed [14:0] m112_55;
   assign m112_55 =15'b0;

   // m112_56 = W*in
   wire signed [14:0] m112_56;
   assign m112_56 =15'b0;

   // m112_57 = W*in
   wire signed [14:0] m112_57;
   assign m112_57 =15'b0;

   // m112_58 = W*in
   wire signed [14:0] m112_58;
   assign m112_58 =15'b0;

   // m112_59 = W*in
   wire signed [14:0] m112_59;
   assign m112_59 =15'b0;

   // m112_60 = W*in
   wire signed [14:0] m112_60;
   assign m112_60 =15'b0;

   // m112_61 = W*in
   wire signed [14:0] m112_61;
   assign m112_61 =15'b0;

   // m112_62 = W*in
   wire signed [14:0] m112_62;
   assign m112_62 =15'b0;

   // m112_63 = W*in
   wire signed [14:0] m112_63;
   assign m112_63 =15'b0;

   // m112_64 = W*in
   wire signed [14:0] m112_64;
   assign m112_64 =15'b0;

   // m112_65 = W*in
   wire signed [14:0] m112_65;
   assign m112_65 =15'b0;

   // m112_66 = W*in
   wire signed [14:0] m112_66;
   assign m112_66 ={ {3{in112[14]}} , in112[14:3] };

   // m112_67 = W*in
   wire signed [14:0] m112_67;
   assign m112_67 =15'b0;

   // m112_68 = W*in
   wire signed [14:0] m112_68;
   assign m112_68 =15'b0;

   // m112_69 = W*in
   wire signed [14:0] m112_69;
   assign m112_69 =15'b0;

   // m112_70 = W*in
   wire signed [14:0] m112_70;
   assign m112_70 =15'b0;

   // m112_71 = W*in
   wire signed [14:0] m112_71;
   assign m112_71 =15'b0;

   // m112_72 = W*in
   wire signed [14:0] m112_72;
   assign m112_72 =15'b0;

   // m112_73 = W*in
   wire signed [14:0] m112_73;
   assign m112_73 =15'b0;

   // m112_74 = W*in
   wire signed [14:0] m112_74;
   assign m112_74 =15'b0;

   // m112_75 = W*in
   wire signed [14:0] m112_75;
   assign m112_75 =15'b0;

   // m112_76 = W*in
   wire signed [14:0] m112_76;
   assign m112_76 =15'b0;

   // m112_77 = W*in
   wire signed [14:0] m112_77;
   assign m112_77 =15'b0;

   // m112_78 = W*in
   wire signed [14:0] m112_78;
   assign m112_78 =15'b0;

   // m112_79 = W*in
   wire signed [14:0] m112_79;
   assign m112_79 =15'b0;

   // m112_80 = W*in
   wire signed [14:0] m112_80;
   assign m112_80 =15'b0;

   // m112_81 = W*in
   wire signed [14:0] m112_81;
   assign m112_81 =15'b0;

   // m112_82 = W*in
   wire signed [14:0] m112_82;
   assign m112_82 =15'b0;

   // m112_83 = W*in
   wire signed [14:0] m112_83;
   assign m112_83 ={ {3{in112[14]}} , in112[14:3] };

   // m112_84 = W*in
   wire signed [14:0] m112_84;
   assign m112_84 =15'b0;

   // m112_85 = W*in
   wire signed [14:0] m112_85;
   assign m112_85 =15'b0;

   // m112_86 = W*in
   wire signed [14:0] m112_86;
   assign m112_86 =15'b0;

   // m112_87 = W*in
   wire signed [14:0] m112_87;
   assign m112_87 =15'b0;

   // m112_88 = W*in
   wire signed [14:0] m112_88;
   assign m112_88 =15'b0;

   // m112_89 = W*in
   wire signed [14:0] m112_89;
   assign m112_89 =15'b0;

   // m112_90 = W*in
   wire signed [14:0] m112_90;
   assign m112_90 =15'b0;

   // m112_91 = W*in
   wire signed [14:0] m112_91;
   assign m112_91 =15'b0;

   // m112_92 = W*in
   wire signed [14:0] m112_92;
   assign m112_92 =15'b0;

   // m112_93 = W*in
   wire signed [14:0] m112_93;
   assign m112_93 =15'b0;

   // m112_94 = W*in
   wire signed [14:0] m112_94;
   assign m112_94 =15'b0;

   // m112_95 = W*in
   wire signed [14:0] m112_95;
   assign m112_95 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_96 = W*in
   wire signed [14:0] m112_96;
   assign m112_96 =15'b0;

   // m112_97 = W*in
   wire signed [14:0] m112_97;
   assign m112_97 ={ {3{in112[14]}} , in112[14:3] };

   // m112_98 = W*in
   wire signed [14:0] m112_98;
   assign m112_98 ={ {3{neg112[14]}} , neg112[14:3] };

   // m112_99 = W*in
   wire signed [14:0] m112_99;
   assign m112_99 =15'b0;

   // m112_100 = W*in
   wire signed [14:0] m112_100;
   assign m112_100 ={ {3{in112[14]}} , in112[14:3] };

   // m113_1 = W*in
   wire signed [14:0] m113_1;
   assign m113_1 =15'b0;

   // m113_2 = W*in
   wire signed [14:0] m113_2;
   assign m113_2 =15'b0;

   // m113_3 = W*in
   wire signed [14:0] m113_3;
   assign m113_3 =15'b0;

   // m113_4 = W*in
   wire signed [14:0] m113_4;
   assign m113_4 ={ {3{in113[14]}} , in113[14:3] };

   // m113_5 = W*in
   wire signed [14:0] m113_5;
   assign m113_5 =15'b0;

   // m113_6 = W*in
   wire signed [14:0] m113_6;
   assign m113_6 ={ {4{neg113[14]}} , neg113[14:4] };

   // m113_7 = W*in
   wire signed [14:0] m113_7;
   assign m113_7 =15'b0;

   // m113_8 = W*in
   wire signed [14:0] m113_8;
   assign m113_8 =15'b0;

   // m113_9 = W*in
   wire signed [14:0] m113_9;
   assign m113_9 =15'b0;

   // m113_10 = W*in
   wire signed [14:0] m113_10;
   assign m113_10 ={ {3{in113[14]}} , in113[14:3] };

   // m113_11 = W*in
   wire signed [14:0] m113_11;
   assign m113_11 =15'b0;

   // m113_12 = W*in
   wire signed [14:0] m113_12;
   assign m113_12 =15'b0;

   // m113_13 = W*in
   wire signed [14:0] m113_13;
   assign m113_13 =15'b0;

   // m113_14 = W*in
   wire signed [14:0] m113_14;
   assign m113_14 =15'b0;

   // m113_15 = W*in
   wire signed [14:0] m113_15;
   assign m113_15 =15'b0;

   // m113_16 = W*in
   wire signed [14:0] m113_16;
   assign m113_16 =15'b0;

   // m113_17 = W*in
   wire signed [14:0] m113_17;
   assign m113_17 =15'b0;

   // m113_18 = W*in
   wire signed [14:0] m113_18;
   assign m113_18 =15'b0;

   // m113_19 = W*in
   wire signed [14:0] m113_19;
   assign m113_19 ={ {4{in113[14]}} , in113[14:4] };

   // m113_20 = W*in
   wire signed [14:0] m113_20;
   assign m113_20 =15'b0;

   // m113_21 = W*in
   wire signed [14:0] m113_21;
   assign m113_21 ={ {4{neg113[14]}} , neg113[14:4] };

   // m113_22 = W*in
   wire signed [14:0] m113_22;
   assign m113_22 ={ {4{neg113[14]}} , neg113[14:4] };

   // m113_23 = W*in
   wire signed [14:0] m113_23;
   assign m113_23 =15'b0;

   // m113_24 = W*in
   wire signed [14:0] m113_24;
   assign m113_24 =15'b0;

   // m113_25 = W*in
   wire signed [14:0] m113_25;
   assign m113_25 ={ {3{in113[14]}} , in113[14:3] };

   // m113_26 = W*in
   wire signed [14:0] m113_26;
   assign m113_26 =15'b0;

   // m113_27 = W*in
   wire signed [14:0] m113_27;
   assign m113_27 =15'b0;

   // m113_28 = W*in
   wire signed [14:0] m113_28;
   assign m113_28 =15'b0;

   // m113_29 = W*in
   wire signed [14:0] m113_29;
   assign m113_29 ={ {4{in113[14]}} , in113[14:4] };

   // m113_30 = W*in
   wire signed [14:0] m113_30;
   assign m113_30 ={ {3{in113[14]}} , in113[14:3] };

   // m113_31 = W*in
   wire signed [14:0] m113_31;
   assign m113_31 ={ {4{in113[14]}} , in113[14:4] };

   // m113_32 = W*in
   wire signed [14:0] m113_32;
   assign m113_32 ={ {3{in113[14]}} , in113[14:3] };

   // m113_33 = W*in
   wire signed [14:0] m113_33;
   assign m113_33 ={ {4{in113[14]}} , in113[14:4] };

   // m113_34 = W*in
   wire signed [14:0] m113_34;
   assign m113_34 =15'b0;

   // m113_35 = W*in
   wire signed [14:0] m113_35;
   assign m113_35 =15'b0;

   // m113_36 = W*in
   wire signed [14:0] m113_36;
   assign m113_36 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_37 = W*in
   wire signed [14:0] m113_37;
   assign m113_37 =15'b0;

   // m113_38 = W*in
   wire signed [14:0] m113_38;
   assign m113_38 =15'b0;

   // m113_39 = W*in
   wire signed [14:0] m113_39;
   assign m113_39 ={ {3{in113[14]}} , in113[14:3] };

   // m113_40 = W*in
   wire signed [14:0] m113_40;
   assign m113_40 =15'b0;

   // m113_41 = W*in
   wire signed [14:0] m113_41;
   assign m113_41 =15'b0;

   // m113_42 = W*in
   wire signed [14:0] m113_42;
   assign m113_42 =15'b0;

   // m113_43 = W*in
   wire signed [14:0] m113_43;
   assign m113_43 =15'b0;

   // m113_44 = W*in
   wire signed [14:0] m113_44;
   assign m113_44 ={ {3{in113[14]}} , in113[14:3] };

   // m113_45 = W*in
   wire signed [14:0] m113_45;
   assign m113_45 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_46 = W*in
   wire signed [14:0] m113_46;
   assign m113_46 =15'b0;

   // m113_47 = W*in
   wire signed [14:0] m113_47;
   assign m113_47 =15'b0;

   // m113_48 = W*in
   wire signed [14:0] m113_48;
   assign m113_48 =15'b0;

   // m113_49 = W*in
   wire signed [14:0] m113_49;
   assign m113_49 =15'b0;

   // m113_50 = W*in
   wire signed [14:0] m113_50;
   assign m113_50 =15'b0;

   // m113_51 = W*in
   wire signed [14:0] m113_51;
   assign m113_51 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_52 = W*in
   wire signed [14:0] m113_52;
   assign m113_52 =15'b0;

   // m113_53 = W*in
   wire signed [14:0] m113_53;
   assign m113_53 =15'b0;

   // m113_54 = W*in
   wire signed [14:0] m113_54;
   assign m113_54 =15'b0;

   // m113_55 = W*in
   wire signed [14:0] m113_55;
   assign m113_55 =15'b0;

   // m113_56 = W*in
   wire signed [14:0] m113_56;
   assign m113_56 =15'b0;

   // m113_57 = W*in
   wire signed [14:0] m113_57;
   assign m113_57 =15'b0;

   // m113_58 = W*in
   wire signed [14:0] m113_58;
   assign m113_58 ={ {4{neg113[14]}} , neg113[14:4] };

   // m113_59 = W*in
   wire signed [14:0] m113_59;
   assign m113_59 ={ {4{in113[14]}} , in113[14:4] };

   // m113_60 = W*in
   wire signed [14:0] m113_60;
   assign m113_60 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_61 = W*in
   wire signed [14:0] m113_61;
   assign m113_61 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_62 = W*in
   wire signed [14:0] m113_62;
   assign m113_62 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_63 = W*in
   wire signed [14:0] m113_63;
   assign m113_63 =15'b0;

   // m113_64 = W*in
   wire signed [14:0] m113_64;
   assign m113_64 ={ {4{neg113[14]}} , neg113[14:4] };

   // m113_65 = W*in
   wire signed [14:0] m113_65;
   assign m113_65 ={ {4{in113[14]}} , in113[14:4] };

   // m113_66 = W*in
   wire signed [14:0] m113_66;
   assign m113_66 =15'b0;

   // m113_67 = W*in
   wire signed [14:0] m113_67;
   assign m113_67 ={ {4{in113[14]}} , in113[14:4] };

   // m113_68 = W*in
   wire signed [14:0] m113_68;
   assign m113_68 =15'b0;

   // m113_69 = W*in
   wire signed [14:0] m113_69;
   assign m113_69 =15'b0;

   // m113_70 = W*in
   wire signed [14:0] m113_70;
   assign m113_70 =15'b0;

   // m113_71 = W*in
   wire signed [14:0] m113_71;
   assign m113_71 =15'b0;

   // m113_72 = W*in
   wire signed [14:0] m113_72;
   assign m113_72 =15'b0;

   // m113_73 = W*in
   wire signed [14:0] m113_73;
   assign m113_73 =15'b0;

   // m113_74 = W*in
   wire signed [14:0] m113_74;
   assign m113_74 ={ {4{neg113[14]}} , neg113[14:4] };

   // m113_75 = W*in
   wire signed [14:0] m113_75;
   assign m113_75 =15'b0;

   // m113_76 = W*in
   wire signed [14:0] m113_76;
   assign m113_76 =15'b0;

   // m113_77 = W*in
   wire signed [14:0] m113_77;
   assign m113_77 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_78 = W*in
   wire signed [14:0] m113_78;
   assign m113_78 =15'b0;

   // m113_79 = W*in
   wire signed [14:0] m113_79;
   assign m113_79 =15'b0;

   // m113_80 = W*in
   wire signed [14:0] m113_80;
   assign m113_80 =15'b0;

   // m113_81 = W*in
   wire signed [14:0] m113_81;
   assign m113_81 =15'b0;

   // m113_82 = W*in
   wire signed [14:0] m113_82;
   assign m113_82 =15'b0;

   // m113_83 = W*in
   wire signed [14:0] m113_83;
   assign m113_83 =15'b0;

   // m113_84 = W*in
   wire signed [14:0] m113_84;
   assign m113_84 =15'b0;

   // m113_85 = W*in
   wire signed [14:0] m113_85;
   assign m113_85 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_86 = W*in
   wire signed [14:0] m113_86;
   assign m113_86 =15'b0;

   // m113_87 = W*in
   wire signed [14:0] m113_87;
   assign m113_87 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_88 = W*in
   wire signed [14:0] m113_88;
   assign m113_88 =15'b0;

   // m113_89 = W*in
   wire signed [14:0] m113_89;
   assign m113_89 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_90 = W*in
   wire signed [14:0] m113_90;
   assign m113_90 ={ {3{in113[14]}} , in113[14:3] };

   // m113_91 = W*in
   wire signed [14:0] m113_91;
   assign m113_91 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_92 = W*in
   wire signed [14:0] m113_92;
   assign m113_92 =15'b0;

   // m113_93 = W*in
   wire signed [14:0] m113_93;
   assign m113_93 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_94 = W*in
   wire signed [14:0] m113_94;
   assign m113_94 =15'b0;

   // m113_95 = W*in
   wire signed [14:0] m113_95;
   assign m113_95 ={ {3{in113[14]}} , in113[14:3] };

   // m113_96 = W*in
   wire signed [14:0] m113_96;
   assign m113_96 ={ {3{neg113[14]}} , neg113[14:3] };

   // m113_97 = W*in
   wire signed [14:0] m113_97;
   assign m113_97 =15'b0;

   // m113_98 = W*in
   wire signed [14:0] m113_98;
   assign m113_98 =15'b0;

   // m113_99 = W*in
   wire signed [14:0] m113_99;
   assign m113_99 =15'b0;

   // m113_100 = W*in
   wire signed [14:0] m113_100;
   assign m113_100 =15'b0;

   // m114_1 = W*in
   wire signed [14:0] m114_1;
   assign m114_1 =15'b0;

   // m114_2 = W*in
   wire signed [14:0] m114_2;
   assign m114_2 ={ {3{in114[14]}} , in114[14:3] };

   // m114_3 = W*in
   wire signed [14:0] m114_3;
   assign m114_3 =15'b0;

   // m114_4 = W*in
   wire signed [14:0] m114_4;
   assign m114_4 =15'b0;

   // m114_5 = W*in
   wire signed [14:0] m114_5;
   assign m114_5 ={ {4{neg114[14]}} , neg114[14:4] };

   // m114_6 = W*in
   wire signed [14:0] m114_6;
   assign m114_6 =15'b0;

   // m114_7 = W*in
   wire signed [14:0] m114_7;
   assign m114_7 =15'b0;

   // m114_8 = W*in
   wire signed [14:0] m114_8;
   assign m114_8 =15'b0;

   // m114_9 = W*in
   wire signed [14:0] m114_9;
   assign m114_9 =15'b0;

   // m114_10 = W*in
   wire signed [14:0] m114_10;
   assign m114_10 =15'b0;

   // m114_11 = W*in
   wire signed [14:0] m114_11;
   assign m114_11 =15'b0;

   // m114_12 = W*in
   wire signed [14:0] m114_12;
   assign m114_12 =15'b0;

   // m114_13 = W*in
   wire signed [14:0] m114_13;
   assign m114_13 ={ {3{in114[14]}} , in114[14:3] };

   // m114_14 = W*in
   wire signed [14:0] m114_14;
   assign m114_14 =15'b0;

   // m114_15 = W*in
   wire signed [14:0] m114_15;
   assign m114_15 =15'b0;

   // m114_16 = W*in
   wire signed [14:0] m114_16;
   assign m114_16 =15'b0;

   // m114_17 = W*in
   wire signed [14:0] m114_17;
   assign m114_17 =15'b0;

   // m114_18 = W*in
   wire signed [14:0] m114_18;
   assign m114_18 =15'b0;

   // m114_19 = W*in
   wire signed [14:0] m114_19;
   assign m114_19 ={ {4{neg114[14]}} , neg114[14:4] };

   // m114_20 = W*in
   wire signed [14:0] m114_20;
   assign m114_20 ={ {3{in114[14]}} , in114[14:3] };

   // m114_21 = W*in
   wire signed [14:0] m114_21;
   assign m114_21 =15'b0;

   // m114_22 = W*in
   wire signed [14:0] m114_22;
   assign m114_22 =15'b0;

   // m114_23 = W*in
   wire signed [14:0] m114_23;
   assign m114_23 =15'b0;

   // m114_24 = W*in
   wire signed [14:0] m114_24;
   assign m114_24 =15'b0;

   // m114_25 = W*in
   wire signed [14:0] m114_25;
   assign m114_25 =15'b0;

   // m114_26 = W*in
   wire signed [14:0] m114_26;
   assign m114_26 =15'b0;

   // m114_27 = W*in
   wire signed [14:0] m114_27;
   assign m114_27 =15'b0;

   // m114_28 = W*in
   wire signed [14:0] m114_28;
   assign m114_28 =15'b0;

   // m114_29 = W*in
   wire signed [14:0] m114_29;
   assign m114_29 ={ {3{in114[14]}} , in114[14:3] };

   // m114_30 = W*in
   wire signed [14:0] m114_30;
   assign m114_30 =15'b0;

   // m114_31 = W*in
   wire signed [14:0] m114_31;
   assign m114_31 =15'b0;

   // m114_32 = W*in
   wire signed [14:0] m114_32;
   assign m114_32 ={ {4{in114[14]}} , in114[14:4] };

   // m114_33 = W*in
   wire signed [14:0] m114_33;
   assign m114_33 ={ {3{in114[14]}} , in114[14:3] };

   // m114_34 = W*in
   wire signed [14:0] m114_34;
   assign m114_34 ={ {3{in114[14]}} , in114[14:3] };

   // m114_35 = W*in
   wire signed [14:0] m114_35;
   assign m114_35 =15'b0;

   // m114_36 = W*in
   wire signed [14:0] m114_36;
   assign m114_36 =15'b0;

   // m114_37 = W*in
   wire signed [14:0] m114_37;
   assign m114_37 =15'b0;

   // m114_38 = W*in
   wire signed [14:0] m114_38;
   assign m114_38 =15'b0;

   // m114_39 = W*in
   wire signed [14:0] m114_39;
   assign m114_39 =15'b0;

   // m114_40 = W*in
   wire signed [14:0] m114_40;
   assign m114_40 =15'b0;

   // m114_41 = W*in
   wire signed [14:0] m114_41;
   assign m114_41 =15'b0;

   // m114_42 = W*in
   wire signed [14:0] m114_42;
   assign m114_42 =15'b0;

   // m114_43 = W*in
   wire signed [14:0] m114_43;
   assign m114_43 =15'b0;

   // m114_44 = W*in
   wire signed [14:0] m114_44;
   assign m114_44 ={ {3{in114[14]}} , in114[14:3] };

   // m114_45 = W*in
   wire signed [14:0] m114_45;
   assign m114_45 =15'b0;

   // m114_46 = W*in
   wire signed [14:0] m114_46;
   assign m114_46 =15'b0;

   // m114_47 = W*in
   wire signed [14:0] m114_47;
   assign m114_47 ={ {3{neg114[14]}} , neg114[14:3] };

   // m114_48 = W*in
   wire signed [14:0] m114_48;
   assign m114_48 ={ {4{neg114[14]}} , neg114[14:4] };

   // m114_49 = W*in
   wire signed [14:0] m114_49;
   assign m114_49 =15'b0;

   // m114_50 = W*in
   wire signed [14:0] m114_50;
   assign m114_50 =15'b0;

   // m114_51 = W*in
   wire signed [14:0] m114_51;
   assign m114_51 ={ {3{neg114[14]}} , neg114[14:3] };

   // m114_52 = W*in
   wire signed [14:0] m114_52;
   assign m114_52 =15'b0;

   // m114_53 = W*in
   wire signed [14:0] m114_53;
   assign m114_53 =15'b0;

   // m114_54 = W*in
   wire signed [14:0] m114_54;
   assign m114_54 =15'b0;

   // m114_55 = W*in
   wire signed [14:0] m114_55;
   assign m114_55 =15'b0;

   // m114_56 = W*in
   wire signed [14:0] m114_56;
   assign m114_56 =15'b0;

   // m114_57 = W*in
   wire signed [14:0] m114_57;
   assign m114_57 =15'b0;

   // m114_58 = W*in
   wire signed [14:0] m114_58;
   assign m114_58 ={ {3{neg114[14]}} , neg114[14:3] };

   // m114_59 = W*in
   wire signed [14:0] m114_59;
   assign m114_59 ={ {4{neg114[14]}} , neg114[14:4] };

   // m114_60 = W*in
   wire signed [14:0] m114_60;
   assign m114_60 ={ {4{in114[14]}} , in114[14:4] };

   // m114_61 = W*in
   wire signed [14:0] m114_61;
   assign m114_61 ={ {3{neg114[14]}} , neg114[14:3] };

   // m114_62 = W*in
   wire signed [14:0] m114_62;
   assign m114_62 =15'b0;

   // m114_63 = W*in
   wire signed [14:0] m114_63;
   assign m114_63 =15'b0;

   // m114_64 = W*in
   wire signed [14:0] m114_64;
   assign m114_64 =15'b0;

   // m114_65 = W*in
   wire signed [14:0] m114_65;
   assign m114_65 =15'b0;

   // m114_66 = W*in
   wire signed [14:0] m114_66;
   assign m114_66 =15'b0;

   // m114_67 = W*in
   wire signed [14:0] m114_67;
   assign m114_67 =15'b0;

   // m114_68 = W*in
   wire signed [14:0] m114_68;
   assign m114_68 =15'b0;

   // m114_69 = W*in
   wire signed [14:0] m114_69;
   assign m114_69 =15'b0;

   // m114_70 = W*in
   wire signed [14:0] m114_70;
   assign m114_70 =15'b0;

   // m114_71 = W*in
   wire signed [14:0] m114_71;
   assign m114_71 =15'b0;

   // m114_72 = W*in
   wire signed [14:0] m114_72;
   assign m114_72 =15'b0;

   // m114_73 = W*in
   wire signed [14:0] m114_73;
   assign m114_73 =15'b0;

   // m114_74 = W*in
   wire signed [14:0] m114_74;
   assign m114_74 =15'b0;

   // m114_75 = W*in
   wire signed [14:0] m114_75;
   assign m114_75 =15'b0;

   // m114_76 = W*in
   wire signed [14:0] m114_76;
   assign m114_76 =15'b0;

   // m114_77 = W*in
   wire signed [14:0] m114_77;
   assign m114_77 ={ {4{neg114[14]}} , neg114[14:4] };

   // m114_78 = W*in
   wire signed [14:0] m114_78;
   assign m114_78 =15'b0;

   // m114_79 = W*in
   wire signed [14:0] m114_79;
   assign m114_79 =15'b0;

   // m114_80 = W*in
   wire signed [14:0] m114_80;
   assign m114_80 =15'b0;

   // m114_81 = W*in
   wire signed [14:0] m114_81;
   assign m114_81 =15'b0;

   // m114_82 = W*in
   wire signed [14:0] m114_82;
   assign m114_82 =15'b0;

   // m114_83 = W*in
   wire signed [14:0] m114_83;
   assign m114_83 =15'b0;

   // m114_84 = W*in
   wire signed [14:0] m114_84;
   assign m114_84 =15'b0;

   // m114_85 = W*in
   wire signed [14:0] m114_85;
   assign m114_85 =15'b0;

   // m114_86 = W*in
   wire signed [14:0] m114_86;
   assign m114_86 =15'b0;

   // m114_87 = W*in
   wire signed [14:0] m114_87;
   assign m114_87 =15'b0;

   // m114_88 = W*in
   wire signed [14:0] m114_88;
   assign m114_88 =15'b0;

   // m114_89 = W*in
   wire signed [14:0] m114_89;
   assign m114_89 ={ {3{neg114[14]}} , neg114[14:3] };

   // m114_90 = W*in
   wire signed [14:0] m114_90;
   assign m114_90 ={ {3{in114[14]}} , in114[14:3] };

   // m114_91 = W*in
   wire signed [14:0] m114_91;
   assign m114_91 ={ {3{neg114[14]}} , neg114[14:3] };

   // m114_92 = W*in
   wire signed [14:0] m114_92;
   assign m114_92 =15'b0;

   // m114_93 = W*in
   wire signed [14:0] m114_93;
   assign m114_93 =15'b0;

   // m114_94 = W*in
   wire signed [14:0] m114_94;
   assign m114_94 ={ {3{in114[14]}} , in114[14:3] };

   // m114_95 = W*in
   wire signed [14:0] m114_95;
   assign m114_95 ={ {3{in114[14]}} , in114[14:3] };

   // m114_96 = W*in
   wire signed [14:0] m114_96;
   assign m114_96 =15'b0;

   // m114_97 = W*in
   wire signed [14:0] m114_97;
   assign m114_97 =15'b0;

   // m114_98 = W*in
   wire signed [14:0] m114_98;
   assign m114_98 =15'b0;

   // m114_99 = W*in
   wire signed [14:0] m114_99;
   assign m114_99 =15'b0;

   // m114_100 = W*in
   wire signed [14:0] m114_100;
   assign m114_100 =15'b0;

   // m115_1 = W*in
   wire signed [14:0] m115_1;
   assign m115_1 ={ {3{in115[14]}} , in115[14:3] };

   // m115_2 = W*in
   wire signed [14:0] m115_2;
   assign m115_2 =15'b0;

   // m115_3 = W*in
   wire signed [14:0] m115_3;
   assign m115_3 =15'b0;

   // m115_4 = W*in
   wire signed [14:0] m115_4;
   assign m115_4 =15'b0;

   // m115_5 = W*in
   wire signed [14:0] m115_5;
   assign m115_5 =15'b0;

   // m115_6 = W*in
   wire signed [14:0] m115_6;
   assign m115_6 =15'b0;

   // m115_7 = W*in
   wire signed [14:0] m115_7;
   assign m115_7 =15'b0;

   // m115_8 = W*in
   wire signed [14:0] m115_8;
   assign m115_8 =15'b0;

   // m115_9 = W*in
   wire signed [14:0] m115_9;
   assign m115_9 =15'b0;

   // m115_10 = W*in
   wire signed [14:0] m115_10;
   assign m115_10 ={ {3{in115[14]}} , in115[14:3] };

   // m115_11 = W*in
   wire signed [14:0] m115_11;
   assign m115_11 =15'b0;

   // m115_12 = W*in
   wire signed [14:0] m115_12;
   assign m115_12 ={ {4{in115[14]}} , in115[14:4] };

   // m115_13 = W*in
   wire signed [14:0] m115_13;
   assign m115_13 =15'b0;

   // m115_14 = W*in
   wire signed [14:0] m115_14;
   assign m115_14 ={ {3{neg115[14]}} , neg115[14:3] };

   // m115_15 = W*in
   wire signed [14:0] m115_15;
   assign m115_15 =15'b0;

   // m115_16 = W*in
   wire signed [14:0] m115_16;
   assign m115_16 =15'b0;

   // m115_17 = W*in
   wire signed [14:0] m115_17;
   assign m115_17 ={ {3{neg115[14]}} , neg115[14:3] };

   // m115_18 = W*in
   wire signed [14:0] m115_18;
   assign m115_18 =15'b0;

   // m115_19 = W*in
   wire signed [14:0] m115_19;
   assign m115_19 ={ {4{neg115[14]}} , neg115[14:4] };

   // m115_20 = W*in
   wire signed [14:0] m115_20;
   assign m115_20 =15'b0;

   // m115_21 = W*in
   wire signed [14:0] m115_21;
   assign m115_21 =15'b0;

   // m115_22 = W*in
   wire signed [14:0] m115_22;
   assign m115_22 ={ {4{in115[14]}} , in115[14:4] };

   // m115_23 = W*in
   wire signed [14:0] m115_23;
   assign m115_23 =15'b0;

   // m115_24 = W*in
   wire signed [14:0] m115_24;
   assign m115_24 ={ {3{neg115[14]}} , neg115[14:3] };

   // m115_25 = W*in
   wire signed [14:0] m115_25;
   assign m115_25 =15'b0;

   // m115_26 = W*in
   wire signed [14:0] m115_26;
   assign m115_26 ={ {4{neg115[14]}} , neg115[14:4] };

   // m115_27 = W*in
   wire signed [14:0] m115_27;
   assign m115_27 =15'b0;

   // m115_28 = W*in
   wire signed [14:0] m115_28;
   assign m115_28 ={ {3{neg115[14]}} , neg115[14:3] };

   // m115_29 = W*in
   wire signed [14:0] m115_29;
   assign m115_29 =15'b0;

   // m115_30 = W*in
   wire signed [14:0] m115_30;
   assign m115_30 =15'b0;

   // m115_31 = W*in
   wire signed [14:0] m115_31;
   assign m115_31 =15'b0;

   // m115_32 = W*in
   wire signed [14:0] m115_32;
   assign m115_32 =15'b0;

   // m115_33 = W*in
   wire signed [14:0] m115_33;
   assign m115_33 =15'b0;

   // m115_34 = W*in
   wire signed [14:0] m115_34;
   assign m115_34 ={ {4{in115[14]}} , in115[14:4] };

   // m115_35 = W*in
   wire signed [14:0] m115_35;
   assign m115_35 =15'b0;

   // m115_36 = W*in
   wire signed [14:0] m115_36;
   assign m115_36 ={ {3{in115[14]}} , in115[14:3] };

   // m115_37 = W*in
   wire signed [14:0] m115_37;
   assign m115_37 =15'b0;

   // m115_38 = W*in
   wire signed [14:0] m115_38;
   assign m115_38 =15'b0;

   // m115_39 = W*in
   wire signed [14:0] m115_39;
   assign m115_39 =15'b0;

   // m115_40 = W*in
   wire signed [14:0] m115_40;
   assign m115_40 =15'b0;

   // m115_41 = W*in
   wire signed [14:0] m115_41;
   assign m115_41 =15'b0;

   // m115_42 = W*in
   wire signed [14:0] m115_42;
   assign m115_42 =15'b0;

   // m115_43 = W*in
   wire signed [14:0] m115_43;
   assign m115_43 =15'b0;

   // m115_44 = W*in
   wire signed [14:0] m115_44;
   assign m115_44 =15'b0;

   // m115_45 = W*in
   wire signed [14:0] m115_45;
   assign m115_45 =15'b0;

   // m115_46 = W*in
   wire signed [14:0] m115_46;
   assign m115_46 =15'b0;

   // m115_47 = W*in
   wire signed [14:0] m115_47;
   assign m115_47 =15'b0;

   // m115_48 = W*in
   wire signed [14:0] m115_48;
   assign m115_48 =15'b0;

   // m115_49 = W*in
   wire signed [14:0] m115_49;
   assign m115_49 =15'b0;

   // m115_50 = W*in
   wire signed [14:0] m115_50;
   assign m115_50 =15'b0;

   // m115_51 = W*in
   wire signed [14:0] m115_51;
   assign m115_51 =15'b0;

   // m115_52 = W*in
   wire signed [14:0] m115_52;
   assign m115_52 =15'b0;

   // m115_53 = W*in
   wire signed [14:0] m115_53;
   assign m115_53 =15'b0;

   // m115_54 = W*in
   wire signed [14:0] m115_54;
   assign m115_54 =15'b0;

   // m115_55 = W*in
   wire signed [14:0] m115_55;
   assign m115_55 ={ {3{neg115[14]}} , neg115[14:3] };

   // m115_56 = W*in
   wire signed [14:0] m115_56;
   assign m115_56 =15'b0;

   // m115_57 = W*in
   wire signed [14:0] m115_57;
   assign m115_57 =15'b0;

   // m115_58 = W*in
   wire signed [14:0] m115_58;
   assign m115_58 =15'b0;

   // m115_59 = W*in
   wire signed [14:0] m115_59;
   assign m115_59 =15'b0;

   // m115_60 = W*in
   wire signed [14:0] m115_60;
   assign m115_60 =15'b0;

   // m115_61 = W*in
   wire signed [14:0] m115_61;
   assign m115_61 =15'b0;

   // m115_62 = W*in
   wire signed [14:0] m115_62;
   assign m115_62 =15'b0;

   // m115_63 = W*in
   wire signed [14:0] m115_63;
   assign m115_63 =15'b0;

   // m115_64 = W*in
   wire signed [14:0] m115_64;
   assign m115_64 =15'b0;

   // m115_65 = W*in
   wire signed [14:0] m115_65;
   assign m115_65 ={ {3{in115[14]}} , in115[14:3] };

   // m115_66 = W*in
   wire signed [14:0] m115_66;
   assign m115_66 =15'b0;

   // m115_67 = W*in
   wire signed [14:0] m115_67;
   assign m115_67 ={ {4{neg115[14]}} , neg115[14:4] };

   // m115_68 = W*in
   wire signed [14:0] m115_68;
   assign m115_68 =15'b0;

   // m115_69 = W*in
   wire signed [14:0] m115_69;
   assign m115_69 =15'b0;

   // m115_70 = W*in
   wire signed [14:0] m115_70;
   assign m115_70 =15'b0;

   // m115_71 = W*in
   wire signed [14:0] m115_71;
   assign m115_71 =15'b0;

   // m115_72 = W*in
   wire signed [14:0] m115_72;
   assign m115_72 =15'b0;

   // m115_73 = W*in
   wire signed [14:0] m115_73;
   assign m115_73 ={ {4{in115[14]}} , in115[14:4] };

   // m115_74 = W*in
   wire signed [14:0] m115_74;
   assign m115_74 ={ {3{neg115[14]}} , neg115[14:3] };

   // m115_75 = W*in
   wire signed [14:0] m115_75;
   assign m115_75 =15'b0;

   // m115_76 = W*in
   wire signed [14:0] m115_76;
   assign m115_76 =15'b0;

   // m115_77 = W*in
   wire signed [14:0] m115_77;
   assign m115_77 =15'b0;

   // m115_78 = W*in
   wire signed [14:0] m115_78;
   assign m115_78 =15'b0;

   // m115_79 = W*in
   wire signed [14:0] m115_79;
   assign m115_79 =15'b0;

   // m115_80 = W*in
   wire signed [14:0] m115_80;
   assign m115_80 =15'b0;

   // m115_81 = W*in
   wire signed [14:0] m115_81;
   assign m115_81 =15'b0;

   // m115_82 = W*in
   wire signed [14:0] m115_82;
   assign m115_82 =15'b0;

   // m115_83 = W*in
   wire signed [14:0] m115_83;
   assign m115_83 =15'b0;

   // m115_84 = W*in
   wire signed [14:0] m115_84;
   assign m115_84 =15'b0;

   // m115_85 = W*in
   wire signed [14:0] m115_85;
   assign m115_85 =15'b0;

   // m115_86 = W*in
   wire signed [14:0] m115_86;
   assign m115_86 =15'b0;

   // m115_87 = W*in
   wire signed [14:0] m115_87;
   assign m115_87 =15'b0;

   // m115_88 = W*in
   wire signed [14:0] m115_88;
   assign m115_88 =15'b0;

   // m115_89 = W*in
   wire signed [14:0] m115_89;
   assign m115_89 =15'b0;

   // m115_90 = W*in
   wire signed [14:0] m115_90;
   assign m115_90 =15'b0;

   // m115_91 = W*in
   wire signed [14:0] m115_91;
   assign m115_91 =15'b0;

   // m115_92 = W*in
   wire signed [14:0] m115_92;
   assign m115_92 ={ {4{neg115[14]}} , neg115[14:4] };

   // m115_93 = W*in
   wire signed [14:0] m115_93;
   assign m115_93 =15'b0;

   // m115_94 = W*in
   wire signed [14:0] m115_94;
   assign m115_94 =15'b0;

   // m115_95 = W*in
   wire signed [14:0] m115_95;
   assign m115_95 =15'b0;

   // m115_96 = W*in
   wire signed [14:0] m115_96;
   assign m115_96 =15'b0;

   // m115_97 = W*in
   wire signed [14:0] m115_97;
   assign m115_97 =15'b0;

   // m115_98 = W*in
   wire signed [14:0] m115_98;
   assign m115_98 =15'b0;

   // m115_99 = W*in
   wire signed [14:0] m115_99;
   assign m115_99 =15'b0;

   // m115_100 = W*in
   wire signed [14:0] m115_100;
   assign m115_100 =15'b0;

   // m116_1 = W*in
   wire signed [14:0] m116_1;
   assign m116_1 =15'b0;

   // m116_2 = W*in
   wire signed [14:0] m116_2;
   assign m116_2 =15'b0;

   // m116_3 = W*in
   wire signed [14:0] m116_3;
   assign m116_3 =15'b0;

   // m116_4 = W*in
   wire signed [14:0] m116_4;
   assign m116_4 ={ {3{neg116[14]}} , neg116[14:3] };

   // m116_5 = W*in
   wire signed [14:0] m116_5;
   assign m116_5 =15'b0;

   // m116_6 = W*in
   wire signed [14:0] m116_6;
   assign m116_6 =15'b0;

   // m116_7 = W*in
   wire signed [14:0] m116_7;
   assign m116_7 =15'b0;

   // m116_8 = W*in
   wire signed [14:0] m116_8;
   assign m116_8 =15'b0;

   // m116_9 = W*in
   wire signed [14:0] m116_9;
   assign m116_9 =15'b0;

   // m116_10 = W*in
   wire signed [14:0] m116_10;
   assign m116_10 =15'b0;

   // m116_11 = W*in
   wire signed [14:0] m116_11;
   assign m116_11 =15'b0;

   // m116_12 = W*in
   wire signed [14:0] m116_12;
   assign m116_12 =15'b0;

   // m116_13 = W*in
   wire signed [14:0] m116_13;
   assign m116_13 =15'b0;

   // m116_14 = W*in
   wire signed [14:0] m116_14;
   assign m116_14 =15'b0;

   // m116_15 = W*in
   wire signed [14:0] m116_15;
   assign m116_15 =15'b0;

   // m116_16 = W*in
   wire signed [14:0] m116_16;
   assign m116_16 =15'b0;

   // m116_17 = W*in
   wire signed [14:0] m116_17;
   assign m116_17 =15'b0;

   // m116_18 = W*in
   wire signed [14:0] m116_18;
   assign m116_18 =15'b0;

   // m116_19 = W*in
   wire signed [14:0] m116_19;
   assign m116_19 ={ {3{in116[14]}} , in116[14:3] };

   // m116_20 = W*in
   wire signed [14:0] m116_20;
   assign m116_20 =15'b0;

   // m116_21 = W*in
   wire signed [14:0] m116_21;
   assign m116_21 =15'b0;

   // m116_22 = W*in
   wire signed [14:0] m116_22;
   assign m116_22 =15'b0;

   // m116_23 = W*in
   wire signed [14:0] m116_23;
   assign m116_23 =15'b0;

   // m116_24 = W*in
   wire signed [14:0] m116_24;
   assign m116_24 =15'b0;

   // m116_25 = W*in
   wire signed [14:0] m116_25;
   assign m116_25 =15'b0;

   // m116_26 = W*in
   wire signed [14:0] m116_26;
   assign m116_26 =15'b0;

   // m116_27 = W*in
   wire signed [14:0] m116_27;
   assign m116_27 =15'b0;

   // m116_28 = W*in
   wire signed [14:0] m116_28;
   assign m116_28 ={ {3{in116[14]}} , in116[14:3] };

   // m116_29 = W*in
   wire signed [14:0] m116_29;
   assign m116_29 ={ {4{neg116[14]}} , neg116[14:4] };

   // m116_30 = W*in
   wire signed [14:0] m116_30;
   assign m116_30 =15'b0;

   // m116_31 = W*in
   wire signed [14:0] m116_31;
   assign m116_31 =15'b0;

   // m116_32 = W*in
   wire signed [14:0] m116_32;
   assign m116_32 =15'b0;

   // m116_33 = W*in
   wire signed [14:0] m116_33;
   assign m116_33 ={ {3{in116[14]}} , in116[14:3] };

   // m116_34 = W*in
   wire signed [14:0] m116_34;
   assign m116_34 =15'b0;

   // m116_35 = W*in
   wire signed [14:0] m116_35;
   assign m116_35 =15'b0;

   // m116_36 = W*in
   wire signed [14:0] m116_36;
   assign m116_36 =15'b0;

   // m116_37 = W*in
   wire signed [14:0] m116_37;
   assign m116_37 =15'b0;

   // m116_38 = W*in
   wire signed [14:0] m116_38;
   assign m116_38 =15'b0;

   // m116_39 = W*in
   wire signed [14:0] m116_39;
   assign m116_39 =15'b0;

   // m116_40 = W*in
   wire signed [14:0] m116_40;
   assign m116_40 =15'b0;

   // m116_41 = W*in
   wire signed [14:0] m116_41;
   assign m116_41 =15'b0;

   // m116_42 = W*in
   wire signed [14:0] m116_42;
   assign m116_42 =15'b0;

   // m116_43 = W*in
   wire signed [14:0] m116_43;
   assign m116_43 =15'b0;

   // m116_44 = W*in
   wire signed [14:0] m116_44;
   assign m116_44 =15'b0;

   // m116_45 = W*in
   wire signed [14:0] m116_45;
   assign m116_45 =15'b0;

   // m116_46 = W*in
   wire signed [14:0] m116_46;
   assign m116_46 ={ {4{in116[14]}} , in116[14:4] };

   // m116_47 = W*in
   wire signed [14:0] m116_47;
   assign m116_47 =15'b0;

   // m116_48 = W*in
   wire signed [14:0] m116_48;
   assign m116_48 =15'b0;

   // m116_49 = W*in
   wire signed [14:0] m116_49;
   assign m116_49 =15'b0;

   // m116_50 = W*in
   wire signed [14:0] m116_50;
   assign m116_50 =15'b0;

   // m116_51 = W*in
   wire signed [14:0] m116_51;
   assign m116_51 =15'b0;

   // m116_52 = W*in
   wire signed [14:0] m116_52;
   assign m116_52 =15'b0;

   // m116_53 = W*in
   wire signed [14:0] m116_53;
   assign m116_53 =15'b0;

   // m116_54 = W*in
   wire signed [14:0] m116_54;
   assign m116_54 =15'b0;

   // m116_55 = W*in
   wire signed [14:0] m116_55;
   assign m116_55 =15'b0;

   // m116_56 = W*in
   wire signed [14:0] m116_56;
   assign m116_56 =15'b0;

   // m116_57 = W*in
   wire signed [14:0] m116_57;
   assign m116_57 ={ {4{neg116[14]}} , neg116[14:4] };

   // m116_58 = W*in
   wire signed [14:0] m116_58;
   assign m116_58 =15'b0;

   // m116_59 = W*in
   wire signed [14:0] m116_59;
   assign m116_59 =15'b0;

   // m116_60 = W*in
   wire signed [14:0] m116_60;
   assign m116_60 =15'b0;

   // m116_61 = W*in
   wire signed [14:0] m116_61;
   assign m116_61 =15'b0;

   // m116_62 = W*in
   wire signed [14:0] m116_62;
   assign m116_62 =15'b0;

   // m116_63 = W*in
   wire signed [14:0] m116_63;
   assign m116_63 =15'b0;

   // m116_64 = W*in
   wire signed [14:0] m116_64;
   assign m116_64 ={ {4{in116[14]}} , in116[14:4] };

   // m116_65 = W*in
   wire signed [14:0] m116_65;
   assign m116_65 ={ {4{neg116[14]}} , neg116[14:4] };

   // m116_66 = W*in
   wire signed [14:0] m116_66;
   assign m116_66 ={ {3{neg116[14]}} , neg116[14:3] };

   // m116_67 = W*in
   wire signed [14:0] m116_67;
   assign m116_67 =15'b0;

   // m116_68 = W*in
   wire signed [14:0] m116_68;
   assign m116_68 =15'b0;

   // m116_69 = W*in
   wire signed [14:0] m116_69;
   assign m116_69 =15'b0;

   // m116_70 = W*in
   wire signed [14:0] m116_70;
   assign m116_70 =15'b0;

   // m116_71 = W*in
   wire signed [14:0] m116_71;
   assign m116_71 =15'b0;

   // m116_72 = W*in
   wire signed [14:0] m116_72;
   assign m116_72 =15'b0;

   // m116_73 = W*in
   wire signed [14:0] m116_73;
   assign m116_73 =15'b0;

   // m116_74 = W*in
   wire signed [14:0] m116_74;
   assign m116_74 ={ {3{in116[14]}} , in116[14:3] };

   // m116_75 = W*in
   wire signed [14:0] m116_75;
   assign m116_75 ={ {3{in116[14]}} , in116[14:3] };

   // m116_76 = W*in
   wire signed [14:0] m116_76;
   assign m116_76 =15'b0;

   // m116_77 = W*in
   wire signed [14:0] m116_77;
   assign m116_77 =15'b0;

   // m116_78 = W*in
   wire signed [14:0] m116_78;
   assign m116_78 =15'b0;

   // m116_79 = W*in
   wire signed [14:0] m116_79;
   assign m116_79 =15'b0;

   // m116_80 = W*in
   wire signed [14:0] m116_80;
   assign m116_80 ={ {4{neg116[14]}} , neg116[14:4] };

   // m116_81 = W*in
   wire signed [14:0] m116_81;
   assign m116_81 =15'b0;

   // m116_82 = W*in
   wire signed [14:0] m116_82;
   assign m116_82 =15'b0;

   // m116_83 = W*in
   wire signed [14:0] m116_83;
   assign m116_83 =15'b0;

   // m116_84 = W*in
   wire signed [14:0] m116_84;
   assign m116_84 =15'b0;

   // m116_85 = W*in
   wire signed [14:0] m116_85;
   assign m116_85 ={ {3{neg116[14]}} , neg116[14:3] };

   // m116_86 = W*in
   wire signed [14:0] m116_86;
   assign m116_86 =15'b0;

   // m116_87 = W*in
   wire signed [14:0] m116_87;
   assign m116_87 =15'b0;

   // m116_88 = W*in
   wire signed [14:0] m116_88;
   assign m116_88 =15'b0;

   // m116_89 = W*in
   wire signed [14:0] m116_89;
   assign m116_89 =15'b0;

   // m116_90 = W*in
   wire signed [14:0] m116_90;
   assign m116_90 ={ {4{in116[14]}} , in116[14:4] };

   // m116_91 = W*in
   wire signed [14:0] m116_91;
   assign m116_91 =15'b0;

   // m116_92 = W*in
   wire signed [14:0] m116_92;
   assign m116_92 =15'b0;

   // m116_93 = W*in
   wire signed [14:0] m116_93;
   assign m116_93 =15'b0;

   // m116_94 = W*in
   wire signed [14:0] m116_94;
   assign m116_94 ={ {3{in116[14]}} , in116[14:3] };

   // m116_95 = W*in
   wire signed [14:0] m116_95;
   assign m116_95 =15'b0;

   // m116_96 = W*in
   wire signed [14:0] m116_96;
   assign m116_96 =15'b0;

   // m116_97 = W*in
   wire signed [14:0] m116_97;
   assign m116_97 =15'b0;

   // m116_98 = W*in
   wire signed [14:0] m116_98;
   assign m116_98 =15'b0;

   // m116_99 = W*in
   wire signed [14:0] m116_99;
   assign m116_99 =15'b0;

   // m116_100 = W*in
   wire signed [14:0] m116_100;
   assign m116_100 =15'b0;

   // m117_1 = W*in
   wire signed [14:0] m117_1;
   assign m117_1 =15'b0;

   // m117_2 = W*in
   wire signed [14:0] m117_2;
   assign m117_2 =15'b0;

   // m117_3 = W*in
   wire signed [14:0] m117_3;
   assign m117_3 =15'b0;

   // m117_4 = W*in
   wire signed [14:0] m117_4;
   assign m117_4 =15'b0;

   // m117_5 = W*in
   wire signed [14:0] m117_5;
   assign m117_5 =15'b0;

   // m117_6 = W*in
   wire signed [14:0] m117_6;
   assign m117_6 =15'b0;

   // m117_7 = W*in
   wire signed [14:0] m117_7;
   assign m117_7 =15'b0;

   // m117_8 = W*in
   wire signed [14:0] m117_8;
   assign m117_8 =15'b0;

   // m117_9 = W*in
   wire signed [14:0] m117_9;
   assign m117_9 =15'b0;

   // m117_10 = W*in
   wire signed [14:0] m117_10;
   assign m117_10 =15'b0;

   // m117_11 = W*in
   wire signed [14:0] m117_11;
   assign m117_11 =15'b0;

   // m117_12 = W*in
   wire signed [14:0] m117_12;
   assign m117_12 =15'b0;

   // m117_13 = W*in
   wire signed [14:0] m117_13;
   assign m117_13 =15'b0;

   // m117_14 = W*in
   wire signed [14:0] m117_14;
   assign m117_14 ={ {3{in117[14]}} , in117[14:3] };

   // m117_15 = W*in
   wire signed [14:0] m117_15;
   assign m117_15 =15'b0;

   // m117_16 = W*in
   wire signed [14:0] m117_16;
   assign m117_16 =15'b0;

   // m117_17 = W*in
   wire signed [14:0] m117_17;
   assign m117_17 =15'b0;

   // m117_18 = W*in
   wire signed [14:0] m117_18;
   assign m117_18 =15'b0;

   // m117_19 = W*in
   wire signed [14:0] m117_19;
   assign m117_19 =15'b0;

   // m117_20 = W*in
   wire signed [14:0] m117_20;
   assign m117_20 ={ {4{neg117[14]}} , neg117[14:4] };

   // m117_21 = W*in
   wire signed [14:0] m117_21;
   assign m117_21 =15'b0;

   // m117_22 = W*in
   wire signed [14:0] m117_22;
   assign m117_22 =15'b0;

   // m117_23 = W*in
   wire signed [14:0] m117_23;
   assign m117_23 =15'b0;

   // m117_24 = W*in
   wire signed [14:0] m117_24;
   assign m117_24 ={ {3{in117[14]}} , in117[14:3] };

   // m117_25 = W*in
   wire signed [14:0] m117_25;
   assign m117_25 =15'b0;

   // m117_26 = W*in
   wire signed [14:0] m117_26;
   assign m117_26 =15'b0;

   // m117_27 = W*in
   wire signed [14:0] m117_27;
   assign m117_27 =15'b0;

   // m117_28 = W*in
   wire signed [14:0] m117_28;
   assign m117_28 =15'b0;

   // m117_29 = W*in
   wire signed [14:0] m117_29;
   assign m117_29 =15'b0;

   // m117_30 = W*in
   wire signed [14:0] m117_30;
   assign m117_30 ={ {3{neg117[14]}} , neg117[14:3] };

   // m117_31 = W*in
   wire signed [14:0] m117_31;
   assign m117_31 =15'b0;

   // m117_32 = W*in
   wire signed [14:0] m117_32;
   assign m117_32 =15'b0;

   // m117_33 = W*in
   wire signed [14:0] m117_33;
   assign m117_33 =15'b0;

   // m117_34 = W*in
   wire signed [14:0] m117_34;
   assign m117_34 =15'b0;

   // m117_35 = W*in
   wire signed [14:0] m117_35;
   assign m117_35 =15'b0;

   // m117_36 = W*in
   wire signed [14:0] m117_36;
   assign m117_36 =15'b0;

   // m117_37 = W*in
   wire signed [14:0] m117_37;
   assign m117_37 =15'b0;

   // m117_38 = W*in
   wire signed [14:0] m117_38;
   assign m117_38 =15'b0;

   // m117_39 = W*in
   wire signed [14:0] m117_39;
   assign m117_39 =15'b0;

   // m117_40 = W*in
   wire signed [14:0] m117_40;
   assign m117_40 =15'b0;

   // m117_41 = W*in
   wire signed [14:0] m117_41;
   assign m117_41 =15'b0;

   // m117_42 = W*in
   wire signed [14:0] m117_42;
   assign m117_42 ={ {3{in117[14]}} , in117[14:3] };

   // m117_43 = W*in
   wire signed [14:0] m117_43;
   assign m117_43 =15'b0;

   // m117_44 = W*in
   wire signed [14:0] m117_44;
   assign m117_44 =15'b0;

   // m117_45 = W*in
   wire signed [14:0] m117_45;
   assign m117_45 =15'b0;

   // m117_46 = W*in
   wire signed [14:0] m117_46;
   assign m117_46 =15'b0;

   // m117_47 = W*in
   wire signed [14:0] m117_47;
   assign m117_47 =15'b0;

   // m117_48 = W*in
   wire signed [14:0] m117_48;
   assign m117_48 =15'b0;

   // m117_49 = W*in
   wire signed [14:0] m117_49;
   assign m117_49 =15'b0;

   // m117_50 = W*in
   wire signed [14:0] m117_50;
   assign m117_50 =15'b0;

   // m117_51 = W*in
   wire signed [14:0] m117_51;
   assign m117_51 =15'b0;

   // m117_52 = W*in
   wire signed [14:0] m117_52;
   assign m117_52 =15'b0;

   // m117_53 = W*in
   wire signed [14:0] m117_53;
   assign m117_53 =15'b0;

   // m117_54 = W*in
   wire signed [14:0] m117_54;
   assign m117_54 =15'b0;

   // m117_55 = W*in
   wire signed [14:0] m117_55;
   assign m117_55 =15'b0;

   // m117_56 = W*in
   wire signed [14:0] m117_56;
   assign m117_56 =15'b0;

   // m117_57 = W*in
   wire signed [14:0] m117_57;
   assign m117_57 =15'b0;

   // m117_58 = W*in
   wire signed [14:0] m117_58;
   assign m117_58 =15'b0;

   // m117_59 = W*in
   wire signed [14:0] m117_59;
   assign m117_59 ={ {3{neg117[14]}} , neg117[14:3] };

   // m117_60 = W*in
   wire signed [14:0] m117_60;
   assign m117_60 =15'b0;

   // m117_61 = W*in
   wire signed [14:0] m117_61;
   assign m117_61 =15'b0;

   // m117_62 = W*in
   wire signed [14:0] m117_62;
   assign m117_62 =15'b0;

   // m117_63 = W*in
   wire signed [14:0] m117_63;
   assign m117_63 =15'b0;

   // m117_64 = W*in
   wire signed [14:0] m117_64;
   assign m117_64 =15'b0;

   // m117_65 = W*in
   wire signed [14:0] m117_65;
   assign m117_65 =15'b0;

   // m117_66 = W*in
   wire signed [14:0] m117_66;
   assign m117_66 =15'b0;

   // m117_67 = W*in
   wire signed [14:0] m117_67;
   assign m117_67 =15'b0;

   // m117_68 = W*in
   wire signed [14:0] m117_68;
   assign m117_68 =15'b0;

   // m117_69 = W*in
   wire signed [14:0] m117_69;
   assign m117_69 =15'b0;

   // m117_70 = W*in
   wire signed [14:0] m117_70;
   assign m117_70 =15'b0;

   // m117_71 = W*in
   wire signed [14:0] m117_71;
   assign m117_71 ={ {3{in117[14]}} , in117[14:3] };

   // m117_72 = W*in
   wire signed [14:0] m117_72;
   assign m117_72 =15'b0;

   // m117_73 = W*in
   wire signed [14:0] m117_73;
   assign m117_73 =15'b0;

   // m117_74 = W*in
   wire signed [14:0] m117_74;
   assign m117_74 ={ {3{in117[14]}} , in117[14:3] };

   // m117_75 = W*in
   wire signed [14:0] m117_75;
   assign m117_75 =15'b0;

   // m117_76 = W*in
   wire signed [14:0] m117_76;
   assign m117_76 =15'b0;

   // m117_77 = W*in
   wire signed [14:0] m117_77;
   assign m117_77 =15'b0;

   // m117_78 = W*in
   wire signed [14:0] m117_78;
   assign m117_78 =15'b0;

   // m117_79 = W*in
   wire signed [14:0] m117_79;
   assign m117_79 =15'b0;

   // m117_80 = W*in
   wire signed [14:0] m117_80;
   assign m117_80 =15'b0;

   // m117_81 = W*in
   wire signed [14:0] m117_81;
   assign m117_81 =15'b0;

   // m117_82 = W*in
   wire signed [14:0] m117_82;
   assign m117_82 =15'b0;

   // m117_83 = W*in
   wire signed [14:0] m117_83;
   assign m117_83 =15'b0;

   // m117_84 = W*in
   wire signed [14:0] m117_84;
   assign m117_84 =15'b0;

   // m117_85 = W*in
   wire signed [14:0] m117_85;
   assign m117_85 =15'b0;

   // m117_86 = W*in
   wire signed [14:0] m117_86;
   assign m117_86 =15'b0;

   // m117_87 = W*in
   wire signed [14:0] m117_87;
   assign m117_87 =15'b0;

   // m117_88 = W*in
   wire signed [14:0] m117_88;
   assign m117_88 ={ {3{in117[14]}} , in117[14:3] };

   // m117_89 = W*in
   wire signed [14:0] m117_89;
   assign m117_89 =15'b0;

   // m117_90 = W*in
   wire signed [14:0] m117_90;
   assign m117_90 =15'b0;

   // m117_91 = W*in
   wire signed [14:0] m117_91;
   assign m117_91 ={ {3{in117[14]}} , in117[14:3] };

   // m117_92 = W*in
   wire signed [14:0] m117_92;
   assign m117_92 =15'b0;

   // m117_93 = W*in
   wire signed [14:0] m117_93;
   assign m117_93 =15'b0;

   // m117_94 = W*in
   wire signed [14:0] m117_94;
   assign m117_94 =15'b0;

   // m117_95 = W*in
   wire signed [14:0] m117_95;
   assign m117_95 =15'b0;

   // m117_96 = W*in
   wire signed [14:0] m117_96;
   assign m117_96 =15'b0;

   // m117_97 = W*in
   wire signed [14:0] m117_97;
   assign m117_97 =15'b0;

   // m117_98 = W*in
   wire signed [14:0] m117_98;
   assign m117_98 ={ {3{in117[14]}} , in117[14:3] };

   // m117_99 = W*in
   wire signed [14:0] m117_99;
   assign m117_99 =15'b0;

   // m117_100 = W*in
   wire signed [14:0] m117_100;
   assign m117_100 =15'b0;

   // m118_1 = W*in
   wire signed [14:0] m118_1;
   assign m118_1 =15'b0;

   // m118_2 = W*in
   wire signed [14:0] m118_2;
   assign m118_2 =15'b0;

   // m118_3 = W*in
   wire signed [14:0] m118_3;
   assign m118_3 =15'b0;

   // m118_4 = W*in
   wire signed [14:0] m118_4;
   assign m118_4 =15'b0;

   // m118_5 = W*in
   wire signed [14:0] m118_5;
   assign m118_5 =15'b0;

   // m118_6 = W*in
   wire signed [14:0] m118_6;
   assign m118_6 =15'b0;

   // m118_7 = W*in
   wire signed [14:0] m118_7;
   assign m118_7 =15'b0;

   // m118_8 = W*in
   wire signed [14:0] m118_8;
   assign m118_8 =15'b0;

   // m118_9 = W*in
   wire signed [14:0] m118_9;
   assign m118_9 ={ {3{in118[14]}} , in118[14:3] };

   // m118_10 = W*in
   wire signed [14:0] m118_10;
   assign m118_10 =15'b0;

   // m118_11 = W*in
   wire signed [14:0] m118_11;
   assign m118_11 =15'b0;

   // m118_12 = W*in
   wire signed [14:0] m118_12;
   assign m118_12 =15'b0;

   // m118_13 = W*in
   wire signed [14:0] m118_13;
   assign m118_13 =15'b0;

   // m118_14 = W*in
   wire signed [14:0] m118_14;
   assign m118_14 =15'b0;

   // m118_15 = W*in
   wire signed [14:0] m118_15;
   assign m118_15 =15'b0;

   // m118_16 = W*in
   wire signed [14:0] m118_16;
   assign m118_16 =15'b0;

   // m118_17 = W*in
   wire signed [14:0] m118_17;
   assign m118_17 =15'b0;

   // m118_18 = W*in
   wire signed [14:0] m118_18;
   assign m118_18 =15'b0;

   // m118_19 = W*in
   wire signed [14:0] m118_19;
   assign m118_19 =15'b0;

   // m118_20 = W*in
   wire signed [14:0] m118_20;
   assign m118_20 =15'b0;

   // m118_21 = W*in
   wire signed [14:0] m118_21;
   assign m118_21 =15'b0;

   // m118_22 = W*in
   wire signed [14:0] m118_22;
   assign m118_22 =15'b0;

   // m118_23 = W*in
   wire signed [14:0] m118_23;
   assign m118_23 =15'b0;

   // m118_24 = W*in
   wire signed [14:0] m118_24;
   assign m118_24 =15'b0;

   // m118_25 = W*in
   wire signed [14:0] m118_25;
   assign m118_25 =15'b0;

   // m118_26 = W*in
   wire signed [14:0] m118_26;
   assign m118_26 =15'b0;

   // m118_27 = W*in
   wire signed [14:0] m118_27;
   assign m118_27 =15'b0;

   // m118_28 = W*in
   wire signed [14:0] m118_28;
   assign m118_28 ={ {4{in118[14]}} , in118[14:4] };

   // m118_29 = W*in
   wire signed [14:0] m118_29;
   assign m118_29 =15'b0;

   // m118_30 = W*in
   wire signed [14:0] m118_30;
   assign m118_30 =15'b0;

   // m118_31 = W*in
   wire signed [14:0] m118_31;
   assign m118_31 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_32 = W*in
   wire signed [14:0] m118_32;
   assign m118_32 =15'b0;

   // m118_33 = W*in
   wire signed [14:0] m118_33;
   assign m118_33 =15'b0;

   // m118_34 = W*in
   wire signed [14:0] m118_34;
   assign m118_34 =15'b0;

   // m118_35 = W*in
   wire signed [14:0] m118_35;
   assign m118_35 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_36 = W*in
   wire signed [14:0] m118_36;
   assign m118_36 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_37 = W*in
   wire signed [14:0] m118_37;
   assign m118_37 =15'b0;

   // m118_38 = W*in
   wire signed [14:0] m118_38;
   assign m118_38 =15'b0;

   // m118_39 = W*in
   wire signed [14:0] m118_39;
   assign m118_39 =15'b0;

   // m118_40 = W*in
   wire signed [14:0] m118_40;
   assign m118_40 =15'b0;

   // m118_41 = W*in
   wire signed [14:0] m118_41;
   assign m118_41 =15'b0;

   // m118_42 = W*in
   wire signed [14:0] m118_42;
   assign m118_42 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_43 = W*in
   wire signed [14:0] m118_43;
   assign m118_43 =15'b0;

   // m118_44 = W*in
   wire signed [14:0] m118_44;
   assign m118_44 =15'b0;

   // m118_45 = W*in
   wire signed [14:0] m118_45;
   assign m118_45 ={ {3{in118[14]}} , in118[14:3] };

   // m118_46 = W*in
   wire signed [14:0] m118_46;
   assign m118_46 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_47 = W*in
   wire signed [14:0] m118_47;
   assign m118_47 =15'b0;

   // m118_48 = W*in
   wire signed [14:0] m118_48;
   assign m118_48 =15'b0;

   // m118_49 = W*in
   wire signed [14:0] m118_49;
   assign m118_49 =15'b0;

   // m118_50 = W*in
   wire signed [14:0] m118_50;
   assign m118_50 ={ {3{in118[14]}} , in118[14:3] };

   // m118_51 = W*in
   wire signed [14:0] m118_51;
   assign m118_51 =15'b0;

   // m118_52 = W*in
   wire signed [14:0] m118_52;
   assign m118_52 =15'b0;

   // m118_53 = W*in
   wire signed [14:0] m118_53;
   assign m118_53 =15'b0;

   // m118_54 = W*in
   wire signed [14:0] m118_54;
   assign m118_54 =15'b0;

   // m118_55 = W*in
   wire signed [14:0] m118_55;
   assign m118_55 =15'b0;

   // m118_56 = W*in
   wire signed [14:0] m118_56;
   assign m118_56 ={ {3{in118[14]}} , in118[14:3] };

   // m118_57 = W*in
   wire signed [14:0] m118_57;
   assign m118_57 =15'b0;

   // m118_58 = W*in
   wire signed [14:0] m118_58;
   assign m118_58 =15'b0;

   // m118_59 = W*in
   wire signed [14:0] m118_59;
   assign m118_59 =15'b0;

   // m118_60 = W*in
   wire signed [14:0] m118_60;
   assign m118_60 ={ {4{neg118[14]}} , neg118[14:4] };

   // m118_61 = W*in
   wire signed [14:0] m118_61;
   assign m118_61 =15'b0;

   // m118_62 = W*in
   wire signed [14:0] m118_62;
   assign m118_62 =15'b0;

   // m118_63 = W*in
   wire signed [14:0] m118_63;
   assign m118_63 =15'b0;

   // m118_64 = W*in
   wire signed [14:0] m118_64;
   assign m118_64 =15'b0;

   // m118_65 = W*in
   wire signed [14:0] m118_65;
   assign m118_65 =15'b0;

   // m118_66 = W*in
   wire signed [14:0] m118_66;
   assign m118_66 =15'b0;

   // m118_67 = W*in
   wire signed [14:0] m118_67;
   assign m118_67 =15'b0;

   // m118_68 = W*in
   wire signed [14:0] m118_68;
   assign m118_68 =15'b0;

   // m118_69 = W*in
   wire signed [14:0] m118_69;
   assign m118_69 =15'b0;

   // m118_70 = W*in
   wire signed [14:0] m118_70;
   assign m118_70 =15'b0;

   // m118_71 = W*in
   wire signed [14:0] m118_71;
   assign m118_71 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_72 = W*in
   wire signed [14:0] m118_72;
   assign m118_72 =15'b0;

   // m118_73 = W*in
   wire signed [14:0] m118_73;
   assign m118_73 =15'b0;

   // m118_74 = W*in
   wire signed [14:0] m118_74;
   assign m118_74 ={ {4{in118[14]}} , in118[14:4] };

   // m118_75 = W*in
   wire signed [14:0] m118_75;
   assign m118_75 =15'b0;

   // m118_76 = W*in
   wire signed [14:0] m118_76;
   assign m118_76 =15'b0;

   // m118_77 = W*in
   wire signed [14:0] m118_77;
   assign m118_77 =15'b0;

   // m118_78 = W*in
   wire signed [14:0] m118_78;
   assign m118_78 =15'b0;

   // m118_79 = W*in
   wire signed [14:0] m118_79;
   assign m118_79 =15'b0;

   // m118_80 = W*in
   wire signed [14:0] m118_80;
   assign m118_80 =15'b0;

   // m118_81 = W*in
   wire signed [14:0] m118_81;
   assign m118_81 =15'b0;

   // m118_82 = W*in
   wire signed [14:0] m118_82;
   assign m118_82 ={ {3{neg118[14]}} , neg118[14:3] };

   // m118_83 = W*in
   wire signed [14:0] m118_83;
   assign m118_83 =15'b0;

   // m118_84 = W*in
   wire signed [14:0] m118_84;
   assign m118_84 =15'b0;

   // m118_85 = W*in
   wire signed [14:0] m118_85;
   assign m118_85 =15'b0;

   // m118_86 = W*in
   wire signed [14:0] m118_86;
   assign m118_86 ={ {3{in118[14]}} , in118[14:3] };

   // m118_87 = W*in
   wire signed [14:0] m118_87;
   assign m118_87 ={ {3{in118[14]}} , in118[14:3] };

   // m118_88 = W*in
   wire signed [14:0] m118_88;
   assign m118_88 =15'b0;

   // m118_89 = W*in
   wire signed [14:0] m118_89;
   assign m118_89 =15'b0;

   // m118_90 = W*in
   wire signed [14:0] m118_90;
   assign m118_90 =15'b0;

   // m118_91 = W*in
   wire signed [14:0] m118_91;
   assign m118_91 =15'b0;

   // m118_92 = W*in
   wire signed [14:0] m118_92;
   assign m118_92 =15'b0;

   // m118_93 = W*in
   wire signed [14:0] m118_93;
   assign m118_93 =15'b0;

   // m118_94 = W*in
   wire signed [14:0] m118_94;
   assign m118_94 =15'b0;

   // m118_95 = W*in
   wire signed [14:0] m118_95;
   assign m118_95 =15'b0;

   // m118_96 = W*in
   wire signed [14:0] m118_96;
   assign m118_96 ={ {4{neg118[14]}} , neg118[14:4] };

   // m118_97 = W*in
   wire signed [14:0] m118_97;
   assign m118_97 =15'b0;

   // m118_98 = W*in
   wire signed [14:0] m118_98;
   assign m118_98 =15'b0;

   // m118_99 = W*in
   wire signed [14:0] m118_99;
   assign m118_99 ={ {3{in118[14]}} , in118[14:3] };

   // m118_100 = W*in
   wire signed [14:0] m118_100;
   assign m118_100 =15'b0;

   // m119_1 = W*in
   wire signed [14:0] m119_1;
   assign m119_1 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_2 = W*in
   wire signed [14:0] m119_2;
   assign m119_2 =15'b0;

   // m119_3 = W*in
   wire signed [14:0] m119_3;
   assign m119_3 =15'b0;

   // m119_4 = W*in
   wire signed [14:0] m119_4;
   assign m119_4 =15'b0;

   // m119_5 = W*in
   wire signed [14:0] m119_5;
   assign m119_5 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_6 = W*in
   wire signed [14:0] m119_6;
   assign m119_6 ={ {3{in119[14]}} , in119[14:3] };

   // m119_7 = W*in
   wire signed [14:0] m119_7;
   assign m119_7 ={ {3{in119[14]}} , in119[14:3] };

   // m119_8 = W*in
   wire signed [14:0] m119_8;
   assign m119_8 =15'b0;

   // m119_9 = W*in
   wire signed [14:0] m119_9;
   assign m119_9 =15'b0;

   // m119_10 = W*in
   wire signed [14:0] m119_10;
   assign m119_10 =15'b0;

   // m119_11 = W*in
   wire signed [14:0] m119_11;
   assign m119_11 =15'b0;

   // m119_12 = W*in
   wire signed [14:0] m119_12;
   assign m119_12 =15'b0;

   // m119_13 = W*in
   wire signed [14:0] m119_13;
   assign m119_13 =15'b0;

   // m119_14 = W*in
   wire signed [14:0] m119_14;
   assign m119_14 =15'b0;

   // m119_15 = W*in
   wire signed [14:0] m119_15;
   assign m119_15 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_16 = W*in
   wire signed [14:0] m119_16;
   assign m119_16 =15'b0;

   // m119_17 = W*in
   wire signed [14:0] m119_17;
   assign m119_17 =15'b0;

   // m119_18 = W*in
   wire signed [14:0] m119_18;
   assign m119_18 =15'b0;

   // m119_19 = W*in
   wire signed [14:0] m119_19;
   assign m119_19 =15'b0;

   // m119_20 = W*in
   wire signed [14:0] m119_20;
   assign m119_20 =15'b0;

   // m119_21 = W*in
   wire signed [14:0] m119_21;
   assign m119_21 =15'b0;

   // m119_22 = W*in
   wire signed [14:0] m119_22;
   assign m119_22 =15'b0;

   // m119_23 = W*in
   wire signed [14:0] m119_23;
   assign m119_23 =15'b0;

   // m119_24 = W*in
   wire signed [14:0] m119_24;
   assign m119_24 ={ {3{in119[14]}} , in119[14:3] };

   // m119_25 = W*in
   wire signed [14:0] m119_25;
   assign m119_25 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_26 = W*in
   wire signed [14:0] m119_26;
   assign m119_26 =15'b0;

   // m119_27 = W*in
   wire signed [14:0] m119_27;
   assign m119_27 =15'b0;

   // m119_28 = W*in
   wire signed [14:0] m119_28;
   assign m119_28 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_29 = W*in
   wire signed [14:0] m119_29;
   assign m119_29 =15'b0;

   // m119_30 = W*in
   wire signed [14:0] m119_30;
   assign m119_30 =15'b0;

   // m119_31 = W*in
   wire signed [14:0] m119_31;
   assign m119_31 ={ {2{in119[14]}} , in119[14:2] };

   // m119_32 = W*in
   wire signed [14:0] m119_32;
   assign m119_32 ={ {3{in119[14]}} , in119[14:3] };

   // m119_33 = W*in
   wire signed [14:0] m119_33;
   assign m119_33 =15'b0;

   // m119_34 = W*in
   wire signed [14:0] m119_34;
   assign m119_34 =15'b0;

   // m119_35 = W*in
   wire signed [14:0] m119_35;
   assign m119_35 =15'b0;

   // m119_36 = W*in
   wire signed [14:0] m119_36;
   assign m119_36 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_37 = W*in
   wire signed [14:0] m119_37;
   assign m119_37 ={ {3{in119[14]}} , in119[14:3] };

   // m119_38 = W*in
   wire signed [14:0] m119_38;
   assign m119_38 =15'b0;

   // m119_39 = W*in
   wire signed [14:0] m119_39;
   assign m119_39 =15'b0;

   // m119_40 = W*in
   wire signed [14:0] m119_40;
   assign m119_40 =15'b0;

   // m119_41 = W*in
   wire signed [14:0] m119_41;
   assign m119_41 =15'b0;

   // m119_42 = W*in
   wire signed [14:0] m119_42;
   assign m119_42 =15'b0;

   // m119_43 = W*in
   wire signed [14:0] m119_43;
   assign m119_43 =15'b0;

   // m119_44 = W*in
   wire signed [14:0] m119_44;
   assign m119_44 =15'b0;

   // m119_45 = W*in
   wire signed [14:0] m119_45;
   assign m119_45 =15'b0;

   // m119_46 = W*in
   wire signed [14:0] m119_46;
   assign m119_46 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_47 = W*in
   wire signed [14:0] m119_47;
   assign m119_47 ={ {3{in119[14]}} , in119[14:3] };

   // m119_48 = W*in
   wire signed [14:0] m119_48;
   assign m119_48 =15'b0;

   // m119_49 = W*in
   wire signed [14:0] m119_49;
   assign m119_49 =15'b0;

   // m119_50 = W*in
   wire signed [14:0] m119_50;
   assign m119_50 =15'b0;

   // m119_51 = W*in
   wire signed [14:0] m119_51;
   assign m119_51 =15'b0;

   // m119_52 = W*in
   wire signed [14:0] m119_52;
   assign m119_52 ={ {3{in119[14]}} , in119[14:3] };

   // m119_53 = W*in
   wire signed [14:0] m119_53;
   assign m119_53 =15'b0;

   // m119_54 = W*in
   wire signed [14:0] m119_54;
   assign m119_54 =15'b0;

   // m119_55 = W*in
   wire signed [14:0] m119_55;
   assign m119_55 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_56 = W*in
   wire signed [14:0] m119_56;
   assign m119_56 =15'b0;

   // m119_57 = W*in
   wire signed [14:0] m119_57;
   assign m119_57 =15'b0;

   // m119_58 = W*in
   wire signed [14:0] m119_58;
   assign m119_58 =15'b0;

   // m119_59 = W*in
   wire signed [14:0] m119_59;
   assign m119_59 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_60 = W*in
   wire signed [14:0] m119_60;
   assign m119_60 =15'b0;

   // m119_61 = W*in
   wire signed [14:0] m119_61;
   assign m119_61 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_62 = W*in
   wire signed [14:0] m119_62;
   assign m119_62 =15'b0;

   // m119_63 = W*in
   wire signed [14:0] m119_63;
   assign m119_63 =15'b0;

   // m119_64 = W*in
   wire signed [14:0] m119_64;
   assign m119_64 =15'b0;

   // m119_65 = W*in
   wire signed [14:0] m119_65;
   assign m119_65 =15'b0;

   // m119_66 = W*in
   wire signed [14:0] m119_66;
   assign m119_66 =15'b0;

   // m119_67 = W*in
   wire signed [14:0] m119_67;
   assign m119_67 =15'b0;

   // m119_68 = W*in
   wire signed [14:0] m119_68;
   assign m119_68 =15'b0;

   // m119_69 = W*in
   wire signed [14:0] m119_69;
   assign m119_69 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_70 = W*in
   wire signed [14:0] m119_70;
   assign m119_70 =15'b0;

   // m119_71 = W*in
   wire signed [14:0] m119_71;
   assign m119_71 =15'b0;

   // m119_72 = W*in
   wire signed [14:0] m119_72;
   assign m119_72 =15'b0;

   // m119_73 = W*in
   wire signed [14:0] m119_73;
   assign m119_73 =15'b0;

   // m119_74 = W*in
   wire signed [14:0] m119_74;
   assign m119_74 =15'b0;

   // m119_75 = W*in
   wire signed [14:0] m119_75;
   assign m119_75 =15'b0;

   // m119_76 = W*in
   wire signed [14:0] m119_76;
   assign m119_76 =15'b0;

   // m119_77 = W*in
   wire signed [14:0] m119_77;
   assign m119_77 =15'b0;

   // m119_78 = W*in
   wire signed [14:0] m119_78;
   assign m119_78 =15'b0;

   // m119_79 = W*in
   wire signed [14:0] m119_79;
   assign m119_79 =15'b0;

   // m119_80 = W*in
   wire signed [14:0] m119_80;
   assign m119_80 =15'b0;

   // m119_81 = W*in
   wire signed [14:0] m119_81;
   assign m119_81 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_82 = W*in
   wire signed [14:0] m119_82;
   assign m119_82 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_83 = W*in
   wire signed [14:0] m119_83;
   assign m119_83 =15'b0;

   // m119_84 = W*in
   wire signed [14:0] m119_84;
   assign m119_84 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_85 = W*in
   wire signed [14:0] m119_85;
   assign m119_85 =15'b0;

   // m119_86 = W*in
   wire signed [14:0] m119_86;
   assign m119_86 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_87 = W*in
   wire signed [14:0] m119_87;
   assign m119_87 =15'b0;

   // m119_88 = W*in
   wire signed [14:0] m119_88;
   assign m119_88 =15'b0;

   // m119_89 = W*in
   wire signed [14:0] m119_89;
   assign m119_89 ={ {3{in119[14]}} , in119[14:3] };

   // m119_90 = W*in
   wire signed [14:0] m119_90;
   assign m119_90 =15'b0;

   // m119_91 = W*in
   wire signed [14:0] m119_91;
   assign m119_91 =15'b0;

   // m119_92 = W*in
   wire signed [14:0] m119_92;
   assign m119_92 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_93 = W*in
   wire signed [14:0] m119_93;
   assign m119_93 =15'b0;

   // m119_94 = W*in
   wire signed [14:0] m119_94;
   assign m119_94 =15'b0;

   // m119_95 = W*in
   wire signed [14:0] m119_95;
   assign m119_95 ={ {3{neg119[14]}} , neg119[14:3] };

   // m119_96 = W*in
   wire signed [14:0] m119_96;
   assign m119_96 =15'b0;

   // m119_97 = W*in
   wire signed [14:0] m119_97;
   assign m119_97 =15'b0;

   // m119_98 = W*in
   wire signed [14:0] m119_98;
   assign m119_98 =15'b0;

   // m119_99 = W*in
   wire signed [14:0] m119_99;
   assign m119_99 =15'b0;

   // m119_100 = W*in
   wire signed [14:0] m119_100;
   assign m119_100 =15'b0;

   // m120_1 = W*in
   wire signed [14:0] m120_1;
   assign m120_1 =15'b0;

   // m120_2 = W*in
   wire signed [14:0] m120_2;
   assign m120_2 =15'b0;

   // m120_3 = W*in
   wire signed [14:0] m120_3;
   assign m120_3 =15'b0;

   // m120_4 = W*in
   wire signed [14:0] m120_4;
   assign m120_4 ={ {3{in120[14]}} , in120[14:3] };

   // m120_5 = W*in
   wire signed [14:0] m120_5;
   assign m120_5 =15'b0;

   // m120_6 = W*in
   wire signed [14:0] m120_6;
   assign m120_6 =15'b0;

   // m120_7 = W*in
   wire signed [14:0] m120_7;
   assign m120_7 =15'b0;

   // m120_8 = W*in
   wire signed [14:0] m120_8;
   assign m120_8 ={ {3{in120[14]}} , in120[14:3] };

   // m120_9 = W*in
   wire signed [14:0] m120_9;
   assign m120_9 =15'b0;

   // m120_10 = W*in
   wire signed [14:0] m120_10;
   assign m120_10 =15'b0;

   // m120_11 = W*in
   wire signed [14:0] m120_11;
   assign m120_11 ={ {3{in120[14]}} , in120[14:3] };

   // m120_12 = W*in
   wire signed [14:0] m120_12;
   assign m120_12 =15'b0;

   // m120_13 = W*in
   wire signed [14:0] m120_13;
   assign m120_13 =15'b0;

   // m120_14 = W*in
   wire signed [14:0] m120_14;
   assign m120_14 =15'b0;

   // m120_15 = W*in
   wire signed [14:0] m120_15;
   assign m120_15 =15'b0;

   // m120_16 = W*in
   wire signed [14:0] m120_16;
   assign m120_16 ={ {3{in120[14]}} , in120[14:3] };

   // m120_17 = W*in
   wire signed [14:0] m120_17;
   assign m120_17 ={ {4{neg120[14]}} , neg120[14:4] };

   // m120_18 = W*in
   wire signed [14:0] m120_18;
   assign m120_18 =15'b0;

   // m120_19 = W*in
   wire signed [14:0] m120_19;
   assign m120_19 =15'b0;

   // m120_20 = W*in
   wire signed [14:0] m120_20;
   assign m120_20 =15'b0;

   // m120_21 = W*in
   wire signed [14:0] m120_21;
   assign m120_21 =15'b0;

   // m120_22 = W*in
   wire signed [14:0] m120_22;
   assign m120_22 =15'b0;

   // m120_23 = W*in
   wire signed [14:0] m120_23;
   assign m120_23 =15'b0;

   // m120_24 = W*in
   wire signed [14:0] m120_24;
   assign m120_24 =15'b0;

   // m120_25 = W*in
   wire signed [14:0] m120_25;
   assign m120_25 ={ {3{neg120[14]}} , neg120[14:3] };

   // m120_26 = W*in
   wire signed [14:0] m120_26;
   assign m120_26 ={ {3{in120[14]}} , in120[14:3] };

   // m120_27 = W*in
   wire signed [14:0] m120_27;
   assign m120_27 =15'b0;

   // m120_28 = W*in
   wire signed [14:0] m120_28;
   assign m120_28 =15'b0;

   // m120_29 = W*in
   wire signed [14:0] m120_29;
   assign m120_29 ={ {4{in120[14]}} , in120[14:4] };

   // m120_30 = W*in
   wire signed [14:0] m120_30;
   assign m120_30 =15'b0;

   // m120_31 = W*in
   wire signed [14:0] m120_31;
   assign m120_31 ={ {2{in120[14]}} , in120[14:2] };

   // m120_32 = W*in
   wire signed [14:0] m120_32;
   assign m120_32 =15'b0;

   // m120_33 = W*in
   wire signed [14:0] m120_33;
   assign m120_33 =15'b0;

   // m120_34 = W*in
   wire signed [14:0] m120_34;
   assign m120_34 =15'b0;

   // m120_35 = W*in
   wire signed [14:0] m120_35;
   assign m120_35 =15'b0;

   // m120_36 = W*in
   wire signed [14:0] m120_36;
   assign m120_36 ={ {3{neg120[14]}} , neg120[14:3] };

   // m120_37 = W*in
   wire signed [14:0] m120_37;
   assign m120_37 =15'b0;

   // m120_38 = W*in
   wire signed [14:0] m120_38;
   assign m120_38 =15'b0;

   // m120_39 = W*in
   wire signed [14:0] m120_39;
   assign m120_39 =15'b0;

   // m120_40 = W*in
   wire signed [14:0] m120_40;
   assign m120_40 =15'b0;

   // m120_41 = W*in
   wire signed [14:0] m120_41;
   assign m120_41 =15'b0;

   // m120_42 = W*in
   wire signed [14:0] m120_42;
   assign m120_42 =15'b0;

   // m120_43 = W*in
   wire signed [14:0] m120_43;
   assign m120_43 =15'b0;

   // m120_44 = W*in
   wire signed [14:0] m120_44;
   assign m120_44 =15'b0;

   // m120_45 = W*in
   wire signed [14:0] m120_45;
   assign m120_45 =15'b0;

   // m120_46 = W*in
   wire signed [14:0] m120_46;
   assign m120_46 =15'b0;

   // m120_47 = W*in
   wire signed [14:0] m120_47;
   assign m120_47 =15'b0;

   // m120_48 = W*in
   wire signed [14:0] m120_48;
   assign m120_48 =15'b0;

   // m120_49 = W*in
   wire signed [14:0] m120_49;
   assign m120_49 ={ {3{neg120[14]}} , neg120[14:3] };

   // m120_50 = W*in
   wire signed [14:0] m120_50;
   assign m120_50 =15'b0;

   // m120_51 = W*in
   wire signed [14:0] m120_51;
   assign m120_51 =15'b0;

   // m120_52 = W*in
   wire signed [14:0] m120_52;
   assign m120_52 =15'b0;

   // m120_53 = W*in
   wire signed [14:0] m120_53;
   assign m120_53 =15'b0;

   // m120_54 = W*in
   wire signed [14:0] m120_54;
   assign m120_54 =15'b0;

   // m120_55 = W*in
   wire signed [14:0] m120_55;
   assign m120_55 =15'b0;

   // m120_56 = W*in
   wire signed [14:0] m120_56;
   assign m120_56 =15'b0;

   // m120_57 = W*in
   wire signed [14:0] m120_57;
   assign m120_57 =15'b0;

   // m120_58 = W*in
   wire signed [14:0] m120_58;
   assign m120_58 =15'b0;

   // m120_59 = W*in
   wire signed [14:0] m120_59;
   assign m120_59 =15'b0;

   // m120_60 = W*in
   wire signed [14:0] m120_60;
   assign m120_60 =15'b0;

   // m120_61 = W*in
   wire signed [14:0] m120_61;
   assign m120_61 =15'b0;

   // m120_62 = W*in
   wire signed [14:0] m120_62;
   assign m120_62 =15'b0;

   // m120_63 = W*in
   wire signed [14:0] m120_63;
   assign m120_63 ={ {3{neg120[14]}} , neg120[14:3] };

   // m120_64 = W*in
   wire signed [14:0] m120_64;
   assign m120_64 =15'b0;

   // m120_65 = W*in
   wire signed [14:0] m120_65;
   assign m120_65 =15'b0;

   // m120_66 = W*in
   wire signed [14:0] m120_66;
   assign m120_66 =15'b0;

   // m120_67 = W*in
   wire signed [14:0] m120_67;
   assign m120_67 =15'b0;

   // m120_68 = W*in
   wire signed [14:0] m120_68;
   assign m120_68 =15'b0;

   // m120_69 = W*in
   wire signed [14:0] m120_69;
   assign m120_69 =15'b0;

   // m120_70 = W*in
   wire signed [14:0] m120_70;
   assign m120_70 =15'b0;

   // m120_71 = W*in
   wire signed [14:0] m120_71;
   assign m120_71 =15'b0;

   // m120_72 = W*in
   wire signed [14:0] m120_72;
   assign m120_72 ={ {3{neg120[14]}} , neg120[14:3] };

   // m120_73 = W*in
   wire signed [14:0] m120_73;
   assign m120_73 =15'b0;

   // m120_74 = W*in
   wire signed [14:0] m120_74;
   assign m120_74 =15'b0;

   // m120_75 = W*in
   wire signed [14:0] m120_75;
   assign m120_75 =15'b0;

   // m120_76 = W*in
   wire signed [14:0] m120_76;
   assign m120_76 =15'b0;

   // m120_77 = W*in
   wire signed [14:0] m120_77;
   assign m120_77 =15'b0;

   // m120_78 = W*in
   wire signed [14:0] m120_78;
   assign m120_78 =15'b0;

   // m120_79 = W*in
   wire signed [14:0] m120_79;
   assign m120_79 =15'b0;

   // m120_80 = W*in
   wire signed [14:0] m120_80;
   assign m120_80 =15'b0;

   // m120_81 = W*in
   wire signed [14:0] m120_81;
   assign m120_81 =15'b0;

   // m120_82 = W*in
   wire signed [14:0] m120_82;
   assign m120_82 =15'b0;

   // m120_83 = W*in
   wire signed [14:0] m120_83;
   assign m120_83 =15'b0;

   // m120_84 = W*in
   wire signed [14:0] m120_84;
   assign m120_84 =15'b0;

   // m120_85 = W*in
   wire signed [14:0] m120_85;
   assign m120_85 =15'b0;

   // m120_86 = W*in
   wire signed [14:0] m120_86;
   assign m120_86 ={ {3{neg120[14]}} , neg120[14:3] };

   // m120_87 = W*in
   wire signed [14:0] m120_87;
   assign m120_87 =15'b0;

   // m120_88 = W*in
   wire signed [14:0] m120_88;
   assign m120_88 =15'b0;

   // m120_89 = W*in
   wire signed [14:0] m120_89;
   assign m120_89 =15'b0;

   // m120_90 = W*in
   wire signed [14:0] m120_90;
   assign m120_90 =15'b0;

   // m120_91 = W*in
   wire signed [14:0] m120_91;
   assign m120_91 =15'b0;

   // m120_92 = W*in
   wire signed [14:0] m120_92;
   assign m120_92 =15'b0;

   // m120_93 = W*in
   wire signed [14:0] m120_93;
   assign m120_93 =15'b0;

   // m120_94 = W*in
   wire signed [14:0] m120_94;
   assign m120_94 =15'b0;

   // m120_95 = W*in
   wire signed [14:0] m120_95;
   assign m120_95 =15'b0;

   // m120_96 = W*in
   wire signed [14:0] m120_96;
   assign m120_96 ={ {3{in120[14]}} , in120[14:3] };

   // m120_97 = W*in
   wire signed [14:0] m120_97;
   assign m120_97 =15'b0;

   // m120_98 = W*in
   wire signed [14:0] m120_98;
   assign m120_98 =15'b0;

   // m120_99 = W*in
   wire signed [14:0] m120_99;
   assign m120_99 =15'b0;

   // m120_100 = W*in
   wire signed [14:0] m120_100;
   assign m120_100 =15'b0;

   // m121_1 = W*in
   wire signed [14:0] m121_1;
   assign m121_1 =15'b0;

   // m121_2 = W*in
   wire signed [14:0] m121_2;
   assign m121_2 =15'b0;

   // m121_3 = W*in
   wire signed [14:0] m121_3;
   assign m121_3 =15'b0;

   // m121_4 = W*in
   wire signed [14:0] m121_4;
   assign m121_4 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_5 = W*in
   wire signed [14:0] m121_5;
   assign m121_5 =15'b0;

   // m121_6 = W*in
   wire signed [14:0] m121_6;
   assign m121_6 =15'b0;

   // m121_7 = W*in
   wire signed [14:0] m121_7;
   assign m121_7 =15'b0;

   // m121_8 = W*in
   wire signed [14:0] m121_8;
   assign m121_8 =15'b0;

   // m121_9 = W*in
   wire signed [14:0] m121_9;
   assign m121_9 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_10 = W*in
   wire signed [14:0] m121_10;
   assign m121_10 =15'b0;

   // m121_11 = W*in
   wire signed [14:0] m121_11;
   assign m121_11 =15'b0;

   // m121_12 = W*in
   wire signed [14:0] m121_12;
   assign m121_12 =15'b0;

   // m121_13 = W*in
   wire signed [14:0] m121_13;
   assign m121_13 =15'b0;

   // m121_14 = W*in
   wire signed [14:0] m121_14;
   assign m121_14 =15'b0;

   // m121_15 = W*in
   wire signed [14:0] m121_15;
   assign m121_15 =15'b0;

   // m121_16 = W*in
   wire signed [14:0] m121_16;
   assign m121_16 =15'b0;

   // m121_17 = W*in
   wire signed [14:0] m121_17;
   assign m121_17 =15'b0;

   // m121_18 = W*in
   wire signed [14:0] m121_18;
   assign m121_18 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_19 = W*in
   wire signed [14:0] m121_19;
   assign m121_19 =15'b0;

   // m121_20 = W*in
   wire signed [14:0] m121_20;
   assign m121_20 =15'b0;

   // m121_21 = W*in
   wire signed [14:0] m121_21;
   assign m121_21 =15'b0;

   // m121_22 = W*in
   wire signed [14:0] m121_22;
   assign m121_22 ={ {4{in121[14]}} , in121[14:4] };

   // m121_23 = W*in
   wire signed [14:0] m121_23;
   assign m121_23 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_24 = W*in
   wire signed [14:0] m121_24;
   assign m121_24 =15'b0;

   // m121_25 = W*in
   wire signed [14:0] m121_25;
   assign m121_25 =15'b0;

   // m121_26 = W*in
   wire signed [14:0] m121_26;
   assign m121_26 =15'b0;

   // m121_27 = W*in
   wire signed [14:0] m121_27;
   assign m121_27 =15'b0;

   // m121_28 = W*in
   wire signed [14:0] m121_28;
   assign m121_28 =15'b0;

   // m121_29 = W*in
   wire signed [14:0] m121_29;
   assign m121_29 =15'b0;

   // m121_30 = W*in
   wire signed [14:0] m121_30;
   assign m121_30 =15'b0;

   // m121_31 = W*in
   wire signed [14:0] m121_31;
   assign m121_31 =15'b0;

   // m121_32 = W*in
   wire signed [14:0] m121_32;
   assign m121_32 =15'b0;

   // m121_33 = W*in
   wire signed [14:0] m121_33;
   assign m121_33 =15'b0;

   // m121_34 = W*in
   wire signed [14:0] m121_34;
   assign m121_34 =15'b0;

   // m121_35 = W*in
   wire signed [14:0] m121_35;
   assign m121_35 =15'b0;

   // m121_36 = W*in
   wire signed [14:0] m121_36;
   assign m121_36 =15'b0;

   // m121_37 = W*in
   wire signed [14:0] m121_37;
   assign m121_37 =15'b0;

   // m121_38 = W*in
   wire signed [14:0] m121_38;
   assign m121_38 =15'b0;

   // m121_39 = W*in
   wire signed [14:0] m121_39;
   assign m121_39 =15'b0;

   // m121_40 = W*in
   wire signed [14:0] m121_40;
   assign m121_40 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_41 = W*in
   wire signed [14:0] m121_41;
   assign m121_41 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_42 = W*in
   wire signed [14:0] m121_42;
   assign m121_42 =15'b0;

   // m121_43 = W*in
   wire signed [14:0] m121_43;
   assign m121_43 =15'b0;

   // m121_44 = W*in
   wire signed [14:0] m121_44;
   assign m121_44 ={ {3{in121[14]}} , in121[14:3] };

   // m121_45 = W*in
   wire signed [14:0] m121_45;
   assign m121_45 =15'b0;

   // m121_46 = W*in
   wire signed [14:0] m121_46;
   assign m121_46 ={ {3{in121[14]}} , in121[14:3] };

   // m121_47 = W*in
   wire signed [14:0] m121_47;
   assign m121_47 =15'b0;

   // m121_48 = W*in
   wire signed [14:0] m121_48;
   assign m121_48 =15'b0;

   // m121_49 = W*in
   wire signed [14:0] m121_49;
   assign m121_49 =15'b0;

   // m121_50 = W*in
   wire signed [14:0] m121_50;
   assign m121_50 =15'b0;

   // m121_51 = W*in
   wire signed [14:0] m121_51;
   assign m121_51 =15'b0;

   // m121_52 = W*in
   wire signed [14:0] m121_52;
   assign m121_52 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_53 = W*in
   wire signed [14:0] m121_53;
   assign m121_53 =15'b0;

   // m121_54 = W*in
   wire signed [14:0] m121_54;
   assign m121_54 =15'b0;

   // m121_55 = W*in
   wire signed [14:0] m121_55;
   assign m121_55 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_56 = W*in
   wire signed [14:0] m121_56;
   assign m121_56 =15'b0;

   // m121_57 = W*in
   wire signed [14:0] m121_57;
   assign m121_57 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_58 = W*in
   wire signed [14:0] m121_58;
   assign m121_58 =15'b0;

   // m121_59 = W*in
   wire signed [14:0] m121_59;
   assign m121_59 =15'b0;

   // m121_60 = W*in
   wire signed [14:0] m121_60;
   assign m121_60 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_61 = W*in
   wire signed [14:0] m121_61;
   assign m121_61 =15'b0;

   // m121_62 = W*in
   wire signed [14:0] m121_62;
   assign m121_62 =15'b0;

   // m121_63 = W*in
   wire signed [14:0] m121_63;
   assign m121_63 ={ {3{in121[14]}} , in121[14:3] };

   // m121_64 = W*in
   wire signed [14:0] m121_64;
   assign m121_64 =15'b0;

   // m121_65 = W*in
   wire signed [14:0] m121_65;
   assign m121_65 =15'b0;

   // m121_66 = W*in
   wire signed [14:0] m121_66;
   assign m121_66 =15'b0;

   // m121_67 = W*in
   wire signed [14:0] m121_67;
   assign m121_67 =15'b0;

   // m121_68 = W*in
   wire signed [14:0] m121_68;
   assign m121_68 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_69 = W*in
   wire signed [14:0] m121_69;
   assign m121_69 =15'b0;

   // m121_70 = W*in
   wire signed [14:0] m121_70;
   assign m121_70 =15'b0;

   // m121_71 = W*in
   wire signed [14:0] m121_71;
   assign m121_71 =15'b0;

   // m121_72 = W*in
   wire signed [14:0] m121_72;
   assign m121_72 =15'b0;

   // m121_73 = W*in
   wire signed [14:0] m121_73;
   assign m121_73 =15'b0;

   // m121_74 = W*in
   wire signed [14:0] m121_74;
   assign m121_74 ={ {4{neg121[14]}} , neg121[14:4] };

   // m121_75 = W*in
   wire signed [14:0] m121_75;
   assign m121_75 ={ {3{in121[14]}} , in121[14:3] };

   // m121_76 = W*in
   wire signed [14:0] m121_76;
   assign m121_76 =15'b0;

   // m121_77 = W*in
   wire signed [14:0] m121_77;
   assign m121_77 ={ {4{neg121[14]}} , neg121[14:4] };

   // m121_78 = W*in
   wire signed [14:0] m121_78;
   assign m121_78 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_79 = W*in
   wire signed [14:0] m121_79;
   assign m121_79 =15'b0;

   // m121_80 = W*in
   wire signed [14:0] m121_80;
   assign m121_80 ={ {3{neg121[14]}} , neg121[14:3] };

   // m121_81 = W*in
   wire signed [14:0] m121_81;
   assign m121_81 =15'b0;

   // m121_82 = W*in
   wire signed [14:0] m121_82;
   assign m121_82 =15'b0;

   // m121_83 = W*in
   wire signed [14:0] m121_83;
   assign m121_83 ={ {3{in121[14]}} , in121[14:3] };

   // m121_84 = W*in
   wire signed [14:0] m121_84;
   assign m121_84 =15'b0;

   // m121_85 = W*in
   wire signed [14:0] m121_85;
   assign m121_85 =15'b0;

   // m121_86 = W*in
   wire signed [14:0] m121_86;
   assign m121_86 =15'b0;

   // m121_87 = W*in
   wire signed [14:0] m121_87;
   assign m121_87 =15'b0;

   // m121_88 = W*in
   wire signed [14:0] m121_88;
   assign m121_88 =15'b0;

   // m121_89 = W*in
   wire signed [14:0] m121_89;
   assign m121_89 =15'b0;

   // m121_90 = W*in
   wire signed [14:0] m121_90;
   assign m121_90 =15'b0;

   // m121_91 = W*in
   wire signed [14:0] m121_91;
   assign m121_91 =15'b0;

   // m121_92 = W*in
   wire signed [14:0] m121_92;
   assign m121_92 =15'b0;

   // m121_93 = W*in
   wire signed [14:0] m121_93;
   assign m121_93 =15'b0;

   // m121_94 = W*in
   wire signed [14:0] m121_94;
   assign m121_94 ={ {3{in121[14]}} , in121[14:3] };

   // m121_95 = W*in
   wire signed [14:0] m121_95;
   assign m121_95 =15'b0;

   // m121_96 = W*in
   wire signed [14:0] m121_96;
   assign m121_96 =15'b0;

   // m121_97 = W*in
   wire signed [14:0] m121_97;
   assign m121_97 =15'b0;

   // m121_98 = W*in
   wire signed [14:0] m121_98;
   assign m121_98 =15'b0;

   // m121_99 = W*in
   wire signed [14:0] m121_99;
   assign m121_99 =15'b0;

   // m121_100 = W*in
   wire signed [14:0] m121_100;
   assign m121_100 =15'b0;

   // m122_1 = W*in
   wire signed [14:0] m122_1;
   assign m122_1 =15'b0;

   // m122_2 = W*in
   wire signed [14:0] m122_2;
   assign m122_2 =15'b0;

   // m122_3 = W*in
   wire signed [14:0] m122_3;
   assign m122_3 =15'b0;

   // m122_4 = W*in
   wire signed [14:0] m122_4;
   assign m122_4 =15'b0;

   // m122_5 = W*in
   wire signed [14:0] m122_5;
   assign m122_5 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_6 = W*in
   wire signed [14:0] m122_6;
   assign m122_6 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_7 = W*in
   wire signed [14:0] m122_7;
   assign m122_7 ={ {3{in122[14]}} , in122[14:3] };

   // m122_8 = W*in
   wire signed [14:0] m122_8;
   assign m122_8 =15'b0;

   // m122_9 = W*in
   wire signed [14:0] m122_9;
   assign m122_9 ={ {3{in122[14]}} , in122[14:3] };

   // m122_10 = W*in
   wire signed [14:0] m122_10;
   assign m122_10 =15'b0;

   // m122_11 = W*in
   wire signed [14:0] m122_11;
   assign m122_11 =15'b0;

   // m122_12 = W*in
   wire signed [14:0] m122_12;
   assign m122_12 =15'b0;

   // m122_13 = W*in
   wire signed [14:0] m122_13;
   assign m122_13 =15'b0;

   // m122_14 = W*in
   wire signed [14:0] m122_14;
   assign m122_14 =15'b0;

   // m122_15 = W*in
   wire signed [14:0] m122_15;
   assign m122_15 =15'b0;

   // m122_16 = W*in
   wire signed [14:0] m122_16;
   assign m122_16 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_17 = W*in
   wire signed [14:0] m122_17;
   assign m122_17 ={ {3{in122[14]}} , in122[14:3] };

   // m122_18 = W*in
   wire signed [14:0] m122_18;
   assign m122_18 =15'b0;

   // m122_19 = W*in
   wire signed [14:0] m122_19;
   assign m122_19 =15'b0;

   // m122_20 = W*in
   wire signed [14:0] m122_20;
   assign m122_20 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_21 = W*in
   wire signed [14:0] m122_21;
   assign m122_21 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_22 = W*in
   wire signed [14:0] m122_22;
   assign m122_22 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_23 = W*in
   wire signed [14:0] m122_23;
   assign m122_23 =15'b0;

   // m122_24 = W*in
   wire signed [14:0] m122_24;
   assign m122_24 =15'b0;

   // m122_25 = W*in
   wire signed [14:0] m122_25;
   assign m122_25 =15'b0;

   // m122_26 = W*in
   wire signed [14:0] m122_26;
   assign m122_26 ={ {4{in122[14]}} , in122[14:4] };

   // m122_27 = W*in
   wire signed [14:0] m122_27;
   assign m122_27 =15'b0;

   // m122_28 = W*in
   wire signed [14:0] m122_28;
   assign m122_28 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_29 = W*in
   wire signed [14:0] m122_29;
   assign m122_29 =15'b0;

   // m122_30 = W*in
   wire signed [14:0] m122_30;
   assign m122_30 =15'b0;

   // m122_31 = W*in
   wire signed [14:0] m122_31;
   assign m122_31 ={ {3{in122[14]}} , in122[14:3] };

   // m122_32 = W*in
   wire signed [14:0] m122_32;
   assign m122_32 ={ {4{in122[14]}} , in122[14:4] };

   // m122_33 = W*in
   wire signed [14:0] m122_33;
   assign m122_33 =15'b0;

   // m122_34 = W*in
   wire signed [14:0] m122_34;
   assign m122_34 =15'b0;

   // m122_35 = W*in
   wire signed [14:0] m122_35;
   assign m122_35 ={ {3{in122[14]}} , in122[14:3] };

   // m122_36 = W*in
   wire signed [14:0] m122_36;
   assign m122_36 =15'b0;

   // m122_37 = W*in
   wire signed [14:0] m122_37;
   assign m122_37 =15'b0;

   // m122_38 = W*in
   wire signed [14:0] m122_38;
   assign m122_38 =15'b0;

   // m122_39 = W*in
   wire signed [14:0] m122_39;
   assign m122_39 ={ {3{in122[14]}} , in122[14:3] };

   // m122_40 = W*in
   wire signed [14:0] m122_40;
   assign m122_40 ={ {3{in122[14]}} , in122[14:3] };

   // m122_41 = W*in
   wire signed [14:0] m122_41;
   assign m122_41 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_42 = W*in
   wire signed [14:0] m122_42;
   assign m122_42 ={ {3{in122[14]}} , in122[14:3] };

   // m122_43 = W*in
   wire signed [14:0] m122_43;
   assign m122_43 =15'b0;

   // m122_44 = W*in
   wire signed [14:0] m122_44;
   assign m122_44 ={ {3{in122[14]}} , in122[14:3] };

   // m122_45 = W*in
   wire signed [14:0] m122_45;
   assign m122_45 =15'b0;

   // m122_46 = W*in
   wire signed [14:0] m122_46;
   assign m122_46 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_47 = W*in
   wire signed [14:0] m122_47;
   assign m122_47 =15'b0;

   // m122_48 = W*in
   wire signed [14:0] m122_48;
   assign m122_48 =15'b0;

   // m122_49 = W*in
   wire signed [14:0] m122_49;
   assign m122_49 =15'b0;

   // m122_50 = W*in
   wire signed [14:0] m122_50;
   assign m122_50 =15'b0;

   // m122_51 = W*in
   wire signed [14:0] m122_51;
   assign m122_51 =15'b0;

   // m122_52 = W*in
   wire signed [14:0] m122_52;
   assign m122_52 =15'b0;

   // m122_53 = W*in
   wire signed [14:0] m122_53;
   assign m122_53 =15'b0;

   // m122_54 = W*in
   wire signed [14:0] m122_54;
   assign m122_54 ={ {3{in122[14]}} , in122[14:3] };

   // m122_55 = W*in
   wire signed [14:0] m122_55;
   assign m122_55 =15'b0;

   // m122_56 = W*in
   wire signed [14:0] m122_56;
   assign m122_56 ={ {3{in122[14]}} , in122[14:3] };

   // m122_57 = W*in
   wire signed [14:0] m122_57;
   assign m122_57 =15'b0;

   // m122_58 = W*in
   wire signed [14:0] m122_58;
   assign m122_58 =15'b0;

   // m122_59 = W*in
   wire signed [14:0] m122_59;
   assign m122_59 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_60 = W*in
   wire signed [14:0] m122_60;
   assign m122_60 =15'b0;

   // m122_61 = W*in
   wire signed [14:0] m122_61;
   assign m122_61 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_62 = W*in
   wire signed [14:0] m122_62;
   assign m122_62 =15'b0;

   // m122_63 = W*in
   wire signed [14:0] m122_63;
   assign m122_63 =15'b0;

   // m122_64 = W*in
   wire signed [14:0] m122_64;
   assign m122_64 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_65 = W*in
   wire signed [14:0] m122_65;
   assign m122_65 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_66 = W*in
   wire signed [14:0] m122_66;
   assign m122_66 ={ {3{in122[14]}} , in122[14:3] };

   // m122_67 = W*in
   wire signed [14:0] m122_67;
   assign m122_67 =15'b0;

   // m122_68 = W*in
   wire signed [14:0] m122_68;
   assign m122_68 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_69 = W*in
   wire signed [14:0] m122_69;
   assign m122_69 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_70 = W*in
   wire signed [14:0] m122_70;
   assign m122_70 ={ {4{in122[14]}} , in122[14:4] };

   // m122_71 = W*in
   wire signed [14:0] m122_71;
   assign m122_71 =15'b0;

   // m122_72 = W*in
   wire signed [14:0] m122_72;
   assign m122_72 =15'b0;

   // m122_73 = W*in
   wire signed [14:0] m122_73;
   assign m122_73 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_74 = W*in
   wire signed [14:0] m122_74;
   assign m122_74 =15'b0;

   // m122_75 = W*in
   wire signed [14:0] m122_75;
   assign m122_75 =15'b0;

   // m122_76 = W*in
   wire signed [14:0] m122_76;
   assign m122_76 =15'b0;

   // m122_77 = W*in
   wire signed [14:0] m122_77;
   assign m122_77 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_78 = W*in
   wire signed [14:0] m122_78;
   assign m122_78 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_79 = W*in
   wire signed [14:0] m122_79;
   assign m122_79 =15'b0;

   // m122_80 = W*in
   wire signed [14:0] m122_80;
   assign m122_80 =15'b0;

   // m122_81 = W*in
   wire signed [14:0] m122_81;
   assign m122_81 =15'b0;

   // m122_82 = W*in
   wire signed [14:0] m122_82;
   assign m122_82 =15'b0;

   // m122_83 = W*in
   wire signed [14:0] m122_83;
   assign m122_83 =15'b0;

   // m122_84 = W*in
   wire signed [14:0] m122_84;
   assign m122_84 ={ {3{in122[14]}} , in122[14:3] };

   // m122_85 = W*in
   wire signed [14:0] m122_85;
   assign m122_85 =15'b0;

   // m122_86 = W*in
   wire signed [14:0] m122_86;
   assign m122_86 =15'b0;

   // m122_87 = W*in
   wire signed [14:0] m122_87;
   assign m122_87 =15'b0;

   // m122_88 = W*in
   wire signed [14:0] m122_88;
   assign m122_88 =15'b0;

   // m122_89 = W*in
   wire signed [14:0] m122_89;
   assign m122_89 =15'b0;

   // m122_90 = W*in
   wire signed [14:0] m122_90;
   assign m122_90 =15'b0;

   // m122_91 = W*in
   wire signed [14:0] m122_91;
   assign m122_91 =15'b0;

   // m122_92 = W*in
   wire signed [14:0] m122_92;
   assign m122_92 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_93 = W*in
   wire signed [14:0] m122_93;
   assign m122_93 =15'b0;

   // m122_94 = W*in
   wire signed [14:0] m122_94;
   assign m122_94 ={ {3{in122[14]}} , in122[14:3] };

   // m122_95 = W*in
   wire signed [14:0] m122_95;
   assign m122_95 =15'b0;

   // m122_96 = W*in
   wire signed [14:0] m122_96;
   assign m122_96 ={ {4{neg122[14]}} , neg122[14:4] };

   // m122_97 = W*in
   wire signed [14:0] m122_97;
   assign m122_97 ={ {3{neg122[14]}} , neg122[14:3] };

   // m122_98 = W*in
   wire signed [14:0] m122_98;
   assign m122_98 =15'b0;

   // m122_99 = W*in
   wire signed [14:0] m122_99;
   assign m122_99 =15'b0;

   // m122_100 = W*in
   wire signed [14:0] m122_100;
   assign m122_100 =15'b0;

   // m123_1 = W*in
   wire signed [14:0] m123_1;
   assign m123_1 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_2 = W*in
   wire signed [14:0] m123_2;
   assign m123_2 =15'b0;

   // m123_3 = W*in
   wire signed [14:0] m123_3;
   assign m123_3 ={ {3{in123[14]}} , in123[14:3] };

   // m123_4 = W*in
   wire signed [14:0] m123_4;
   assign m123_4 =15'b0;

   // m123_5 = W*in
   wire signed [14:0] m123_5;
   assign m123_5 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_6 = W*in
   wire signed [14:0] m123_6;
   assign m123_6 ={ {2{in123[14]}} , in123[14:2] };

   // m123_7 = W*in
   wire signed [14:0] m123_7;
   assign m123_7 =15'b0;

   // m123_8 = W*in
   wire signed [14:0] m123_8;
   assign m123_8 =15'b0;

   // m123_9 = W*in
   wire signed [14:0] m123_9;
   assign m123_9 =15'b0;

   // m123_10 = W*in
   wire signed [14:0] m123_10;
   assign m123_10 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_11 = W*in
   wire signed [14:0] m123_11;
   assign m123_11 ={ {3{in123[14]}} , in123[14:3] };

   // m123_12 = W*in
   wire signed [14:0] m123_12;
   assign m123_12 =15'b0;

   // m123_13 = W*in
   wire signed [14:0] m123_13;
   assign m123_13 =15'b0;

   // m123_14 = W*in
   wire signed [14:0] m123_14;
   assign m123_14 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_15 = W*in
   wire signed [14:0] m123_15;
   assign m123_15 =15'b0;

   // m123_16 = W*in
   wire signed [14:0] m123_16;
   assign m123_16 =15'b0;

   // m123_17 = W*in
   wire signed [14:0] m123_17;
   assign m123_17 =15'b0;

   // m123_18 = W*in
   wire signed [14:0] m123_18;
   assign m123_18 =15'b0;

   // m123_19 = W*in
   wire signed [14:0] m123_19;
   assign m123_19 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_20 = W*in
   wire signed [14:0] m123_20;
   assign m123_20 =15'b0;

   // m123_21 = W*in
   wire signed [14:0] m123_21;
   assign m123_21 =15'b0;

   // m123_22 = W*in
   wire signed [14:0] m123_22;
   assign m123_22 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_23 = W*in
   wire signed [14:0] m123_23;
   assign m123_23 =15'b0;

   // m123_24 = W*in
   wire signed [14:0] m123_24;
   assign m123_24 =15'b0;

   // m123_25 = W*in
   wire signed [14:0] m123_25;
   assign m123_25 ={ {4{in123[14]}} , in123[14:4] };

   // m123_26 = W*in
   wire signed [14:0] m123_26;
   assign m123_26 ={ {4{neg123[14]}} , neg123[14:4] };

   // m123_27 = W*in
   wire signed [14:0] m123_27;
   assign m123_27 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_28 = W*in
   wire signed [14:0] m123_28;
   assign m123_28 ={ {4{in123[14]}} , in123[14:4] };

   // m123_29 = W*in
   wire signed [14:0] m123_29;
   assign m123_29 ={ {3{in123[14]}} , in123[14:3] };

   // m123_30 = W*in
   wire signed [14:0] m123_30;
   assign m123_30 =15'b0;

   // m123_31 = W*in
   wire signed [14:0] m123_31;
   assign m123_31 ={ {4{neg123[14]}} , neg123[14:4] };

   // m123_32 = W*in
   wire signed [14:0] m123_32;
   assign m123_32 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_33 = W*in
   wire signed [14:0] m123_33;
   assign m123_33 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_34 = W*in
   wire signed [14:0] m123_34;
   assign m123_34 ={ {3{in123[14]}} , in123[14:3] };

   // m123_35 = W*in
   wire signed [14:0] m123_35;
   assign m123_35 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_36 = W*in
   wire signed [14:0] m123_36;
   assign m123_36 =15'b0;

   // m123_37 = W*in
   wire signed [14:0] m123_37;
   assign m123_37 =15'b0;

   // m123_38 = W*in
   wire signed [14:0] m123_38;
   assign m123_38 =15'b0;

   // m123_39 = W*in
   wire signed [14:0] m123_39;
   assign m123_39 =15'b0;

   // m123_40 = W*in
   wire signed [14:0] m123_40;
   assign m123_40 =15'b0;

   // m123_41 = W*in
   wire signed [14:0] m123_41;
   assign m123_41 ={ {3{in123[14]}} , in123[14:3] };

   // m123_42 = W*in
   wire signed [14:0] m123_42;
   assign m123_42 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_43 = W*in
   wire signed [14:0] m123_43;
   assign m123_43 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_44 = W*in
   wire signed [14:0] m123_44;
   assign m123_44 =15'b0;

   // m123_45 = W*in
   wire signed [14:0] m123_45;
   assign m123_45 ={ {3{in123[14]}} , in123[14:3] };

   // m123_46 = W*in
   wire signed [14:0] m123_46;
   assign m123_46 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_47 = W*in
   wire signed [14:0] m123_47;
   assign m123_47 =15'b0;

   // m123_48 = W*in
   wire signed [14:0] m123_48;
   assign m123_48 ={ {4{neg123[14]}} , neg123[14:4] };

   // m123_49 = W*in
   wire signed [14:0] m123_49;
   assign m123_49 ={ {3{in123[14]}} , in123[14:3] };

   // m123_50 = W*in
   wire signed [14:0] m123_50;
   assign m123_50 =15'b0;

   // m123_51 = W*in
   wire signed [14:0] m123_51;
   assign m123_51 =15'b0;

   // m123_52 = W*in
   wire signed [14:0] m123_52;
   assign m123_52 ={ {3{in123[14]}} , in123[14:3] };

   // m123_53 = W*in
   wire signed [14:0] m123_53;
   assign m123_53 =15'b0;

   // m123_54 = W*in
   wire signed [14:0] m123_54;
   assign m123_54 =15'b0;

   // m123_55 = W*in
   wire signed [14:0] m123_55;
   assign m123_55 =15'b0;

   // m123_56 = W*in
   wire signed [14:0] m123_56;
   assign m123_56 =15'b0;

   // m123_57 = W*in
   wire signed [14:0] m123_57;
   assign m123_57 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_58 = W*in
   wire signed [14:0] m123_58;
   assign m123_58 ={ {3{in123[14]}} , in123[14:3] };

   // m123_59 = W*in
   wire signed [14:0] m123_59;
   assign m123_59 =15'b0;

   // m123_60 = W*in
   wire signed [14:0] m123_60;
   assign m123_60 ={ {3{in123[14]}} , in123[14:3] };

   // m123_61 = W*in
   wire signed [14:0] m123_61;
   assign m123_61 ={ {4{neg123[14]}} , neg123[14:4] };

   // m123_62 = W*in
   wire signed [14:0] m123_62;
   assign m123_62 =15'b0;

   // m123_63 = W*in
   wire signed [14:0] m123_63;
   assign m123_63 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_64 = W*in
   wire signed [14:0] m123_64;
   assign m123_64 =15'b0;

   // m123_65 = W*in
   wire signed [14:0] m123_65;
   assign m123_65 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_66 = W*in
   wire signed [14:0] m123_66;
   assign m123_66 ={ {4{neg123[14]}} , neg123[14:4] };

   // m123_67 = W*in
   wire signed [14:0] m123_67;
   assign m123_67 ={ {4{in123[14]}} , in123[14:4] };

   // m123_68 = W*in
   wire signed [14:0] m123_68;
   assign m123_68 ={ {4{in123[14]}} , in123[14:4] };

   // m123_69 = W*in
   wire signed [14:0] m123_69;
   assign m123_69 =15'b0;

   // m123_70 = W*in
   wire signed [14:0] m123_70;
   assign m123_70 =15'b0;

   // m123_71 = W*in
   wire signed [14:0] m123_71;
   assign m123_71 =15'b0;

   // m123_72 = W*in
   wire signed [14:0] m123_72;
   assign m123_72 =15'b0;

   // m123_73 = W*in
   wire signed [14:0] m123_73;
   assign m123_73 =15'b0;

   // m123_74 = W*in
   wire signed [14:0] m123_74;
   assign m123_74 =15'b0;

   // m123_75 = W*in
   wire signed [14:0] m123_75;
   assign m123_75 =15'b0;

   // m123_76 = W*in
   wire signed [14:0] m123_76;
   assign m123_76 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_77 = W*in
   wire signed [14:0] m123_77;
   assign m123_77 ={ {3{in123[14]}} , in123[14:3] };

   // m123_78 = W*in
   wire signed [14:0] m123_78;
   assign m123_78 =15'b0;

   // m123_79 = W*in
   wire signed [14:0] m123_79;
   assign m123_79 =15'b0;

   // m123_80 = W*in
   wire signed [14:0] m123_80;
   assign m123_80 =15'b0;

   // m123_81 = W*in
   wire signed [14:0] m123_81;
   assign m123_81 =15'b0;

   // m123_82 = W*in
   wire signed [14:0] m123_82;
   assign m123_82 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_83 = W*in
   wire signed [14:0] m123_83;
   assign m123_83 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_84 = W*in
   wire signed [14:0] m123_84;
   assign m123_84 =15'b0;

   // m123_85 = W*in
   wire signed [14:0] m123_85;
   assign m123_85 =15'b0;

   // m123_86 = W*in
   wire signed [14:0] m123_86;
   assign m123_86 =15'b0;

   // m123_87 = W*in
   wire signed [14:0] m123_87;
   assign m123_87 =15'b0;

   // m123_88 = W*in
   wire signed [14:0] m123_88;
   assign m123_88 ={ {3{in123[14]}} , in123[14:3] };

   // m123_89 = W*in
   wire signed [14:0] m123_89;
   assign m123_89 =15'b0;

   // m123_90 = W*in
   wire signed [14:0] m123_90;
   assign m123_90 =15'b0;

   // m123_91 = W*in
   wire signed [14:0] m123_91;
   assign m123_91 =15'b0;

   // m123_92 = W*in
   wire signed [14:0] m123_92;
   assign m123_92 =15'b0;

   // m123_93 = W*in
   wire signed [14:0] m123_93;
   assign m123_93 =15'b0;

   // m123_94 = W*in
   wire signed [14:0] m123_94;
   assign m123_94 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_95 = W*in
   wire signed [14:0] m123_95;
   assign m123_95 ={ {3{in123[14]}} , in123[14:3] };

   // m123_96 = W*in
   wire signed [14:0] m123_96;
   assign m123_96 ={ {2{in123[14]}} , in123[14:2] };

   // m123_97 = W*in
   wire signed [14:0] m123_97;
   assign m123_97 ={ {3{neg123[14]}} , neg123[14:3] };

   // m123_98 = W*in
   wire signed [14:0] m123_98;
   assign m123_98 =15'b0;

   // m123_99 = W*in
   wire signed [14:0] m123_99;
   assign m123_99 =15'b0;

   // m123_100 = W*in
   wire signed [14:0] m123_100;
   assign m123_100 ={ {3{neg123[14]}} , neg123[14:3] };

   // m124_1 = W*in
   wire signed [14:0] m124_1;
   assign m124_1 =15'b0;

   // m124_2 = W*in
   wire signed [14:0] m124_2;
   assign m124_2 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_3 = W*in
   wire signed [14:0] m124_3;
   assign m124_3 =15'b0;

   // m124_4 = W*in
   wire signed [14:0] m124_4;
   assign m124_4 =15'b0;

   // m124_5 = W*in
   wire signed [14:0] m124_5;
   assign m124_5 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_6 = W*in
   wire signed [14:0] m124_6;
   assign m124_6 =15'b0;

   // m124_7 = W*in
   wire signed [14:0] m124_7;
   assign m124_7 =15'b0;

   // m124_8 = W*in
   wire signed [14:0] m124_8;
   assign m124_8 =15'b0;

   // m124_9 = W*in
   wire signed [14:0] m124_9;
   assign m124_9 =15'b0;

   // m124_10 = W*in
   wire signed [14:0] m124_10;
   assign m124_10 =15'b0;

   // m124_11 = W*in
   wire signed [14:0] m124_11;
   assign m124_11 =15'b0;

   // m124_12 = W*in
   wire signed [14:0] m124_12;
   assign m124_12 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_13 = W*in
   wire signed [14:0] m124_13;
   assign m124_13 =15'b0;

   // m124_14 = W*in
   wire signed [14:0] m124_14;
   assign m124_14 =15'b0;

   // m124_15 = W*in
   wire signed [14:0] m124_15;
   assign m124_15 =15'b0;

   // m124_16 = W*in
   wire signed [14:0] m124_16;
   assign m124_16 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_17 = W*in
   wire signed [14:0] m124_17;
   assign m124_17 ={ {3{in124[14]}} , in124[14:3] };

   // m124_18 = W*in
   wire signed [14:0] m124_18;
   assign m124_18 =15'b0;

   // m124_19 = W*in
   wire signed [14:0] m124_19;
   assign m124_19 =15'b0;

   // m124_20 = W*in
   wire signed [14:0] m124_20;
   assign m124_20 =15'b0;

   // m124_21 = W*in
   wire signed [14:0] m124_21;
   assign m124_21 ={ {3{in124[14]}} , in124[14:3] };

   // m124_22 = W*in
   wire signed [14:0] m124_22;
   assign m124_22 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_23 = W*in
   wire signed [14:0] m124_23;
   assign m124_23 =15'b0;

   // m124_24 = W*in
   wire signed [14:0] m124_24;
   assign m124_24 =15'b0;

   // m124_25 = W*in
   wire signed [14:0] m124_25;
   assign m124_25 =15'b0;

   // m124_26 = W*in
   wire signed [14:0] m124_26;
   assign m124_26 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_27 = W*in
   wire signed [14:0] m124_27;
   assign m124_27 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_28 = W*in
   wire signed [14:0] m124_28;
   assign m124_28 ={ {4{in124[14]}} , in124[14:4] };

   // m124_29 = W*in
   wire signed [14:0] m124_29;
   assign m124_29 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_30 = W*in
   wire signed [14:0] m124_30;
   assign m124_30 =15'b0;

   // m124_31 = W*in
   wire signed [14:0] m124_31;
   assign m124_31 =15'b0;

   // m124_32 = W*in
   wire signed [14:0] m124_32;
   assign m124_32 =15'b0;

   // m124_33 = W*in
   wire signed [14:0] m124_33;
   assign m124_33 =15'b0;

   // m124_34 = W*in
   wire signed [14:0] m124_34;
   assign m124_34 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_35 = W*in
   wire signed [14:0] m124_35;
   assign m124_35 =15'b0;

   // m124_36 = W*in
   wire signed [14:0] m124_36;
   assign m124_36 =15'b0;

   // m124_37 = W*in
   wire signed [14:0] m124_37;
   assign m124_37 =15'b0;

   // m124_38 = W*in
   wire signed [14:0] m124_38;
   assign m124_38 =15'b0;

   // m124_39 = W*in
   wire signed [14:0] m124_39;
   assign m124_39 =15'b0;

   // m124_40 = W*in
   wire signed [14:0] m124_40;
   assign m124_40 =15'b0;

   // m124_41 = W*in
   wire signed [14:0] m124_41;
   assign m124_41 =15'b0;

   // m124_42 = W*in
   wire signed [14:0] m124_42;
   assign m124_42 =15'b0;

   // m124_43 = W*in
   wire signed [14:0] m124_43;
   assign m124_43 =15'b0;

   // m124_44 = W*in
   wire signed [14:0] m124_44;
   assign m124_44 ={ {3{in124[14]}} , in124[14:3] };

   // m124_45 = W*in
   wire signed [14:0] m124_45;
   assign m124_45 =15'b0;

   // m124_46 = W*in
   wire signed [14:0] m124_46;
   assign m124_46 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_47 = W*in
   wire signed [14:0] m124_47;
   assign m124_47 ={ {3{in124[14]}} , in124[14:3] };

   // m124_48 = W*in
   wire signed [14:0] m124_48;
   assign m124_48 =15'b0;

   // m124_49 = W*in
   wire signed [14:0] m124_49;
   assign m124_49 =15'b0;

   // m124_50 = W*in
   wire signed [14:0] m124_50;
   assign m124_50 ={ {3{in124[14]}} , in124[14:3] };

   // m124_51 = W*in
   wire signed [14:0] m124_51;
   assign m124_51 =15'b0;

   // m124_52 = W*in
   wire signed [14:0] m124_52;
   assign m124_52 =15'b0;

   // m124_53 = W*in
   wire signed [14:0] m124_53;
   assign m124_53 =15'b0;

   // m124_54 = W*in
   wire signed [14:0] m124_54;
   assign m124_54 =15'b0;

   // m124_55 = W*in
   wire signed [14:0] m124_55;
   assign m124_55 =15'b0;

   // m124_56 = W*in
   wire signed [14:0] m124_56;
   assign m124_56 =15'b0;

   // m124_57 = W*in
   wire signed [14:0] m124_57;
   assign m124_57 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_58 = W*in
   wire signed [14:0] m124_58;
   assign m124_58 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_59 = W*in
   wire signed [14:0] m124_59;
   assign m124_59 ={ {3{in124[14]}} , in124[14:3] };

   // m124_60 = W*in
   wire signed [14:0] m124_60;
   assign m124_60 =15'b0;

   // m124_61 = W*in
   wire signed [14:0] m124_61;
   assign m124_61 ={ {4{neg124[14]}} , neg124[14:4] };

   // m124_62 = W*in
   wire signed [14:0] m124_62;
   assign m124_62 =15'b0;

   // m124_63 = W*in
   wire signed [14:0] m124_63;
   assign m124_63 =15'b0;

   // m124_64 = W*in
   wire signed [14:0] m124_64;
   assign m124_64 =15'b0;

   // m124_65 = W*in
   wire signed [14:0] m124_65;
   assign m124_65 ={ {4{neg124[14]}} , neg124[14:4] };

   // m124_66 = W*in
   wire signed [14:0] m124_66;
   assign m124_66 =15'b0;

   // m124_67 = W*in
   wire signed [14:0] m124_67;
   assign m124_67 =15'b0;

   // m124_68 = W*in
   wire signed [14:0] m124_68;
   assign m124_68 =15'b0;

   // m124_69 = W*in
   wire signed [14:0] m124_69;
   assign m124_69 =15'b0;

   // m124_70 = W*in
   wire signed [14:0] m124_70;
   assign m124_70 =15'b0;

   // m124_71 = W*in
   wire signed [14:0] m124_71;
   assign m124_71 =15'b0;

   // m124_72 = W*in
   wire signed [14:0] m124_72;
   assign m124_72 =15'b0;

   // m124_73 = W*in
   wire signed [14:0] m124_73;
   assign m124_73 ={ {3{in124[14]}} , in124[14:3] };

   // m124_74 = W*in
   wire signed [14:0] m124_74;
   assign m124_74 =15'b0;

   // m124_75 = W*in
   wire signed [14:0] m124_75;
   assign m124_75 ={ {3{in124[14]}} , in124[14:3] };

   // m124_76 = W*in
   wire signed [14:0] m124_76;
   assign m124_76 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_77 = W*in
   wire signed [14:0] m124_77;
   assign m124_77 ={ {3{in124[14]}} , in124[14:3] };

   // m124_78 = W*in
   wire signed [14:0] m124_78;
   assign m124_78 =15'b0;

   // m124_79 = W*in
   wire signed [14:0] m124_79;
   assign m124_79 =15'b0;

   // m124_80 = W*in
   wire signed [14:0] m124_80;
   assign m124_80 =15'b0;

   // m124_81 = W*in
   wire signed [14:0] m124_81;
   assign m124_81 =15'b0;

   // m124_82 = W*in
   wire signed [14:0] m124_82;
   assign m124_82 ={ {3{neg124[14]}} , neg124[14:3] };

   // m124_83 = W*in
   wire signed [14:0] m124_83;
   assign m124_83 =15'b0;

   // m124_84 = W*in
   wire signed [14:0] m124_84;
   assign m124_84 =15'b0;

   // m124_85 = W*in
   wire signed [14:0] m124_85;
   assign m124_85 =15'b0;

   // m124_86 = W*in
   wire signed [14:0] m124_86;
   assign m124_86 ={ {3{in124[14]}} , in124[14:3] };

   // m124_87 = W*in
   wire signed [14:0] m124_87;
   assign m124_87 =15'b0;

   // m124_88 = W*in
   wire signed [14:0] m124_88;
   assign m124_88 =15'b0;

   // m124_89 = W*in
   wire signed [14:0] m124_89;
   assign m124_89 =15'b0;

   // m124_90 = W*in
   wire signed [14:0] m124_90;
   assign m124_90 =15'b0;

   // m124_91 = W*in
   wire signed [14:0] m124_91;
   assign m124_91 =15'b0;

   // m124_92 = W*in
   wire signed [14:0] m124_92;
   assign m124_92 =15'b0;

   // m124_93 = W*in
   wire signed [14:0] m124_93;
   assign m124_93 =15'b0;

   // m124_94 = W*in
   wire signed [14:0] m124_94;
   assign m124_94 ={ {3{in124[14]}} , in124[14:3] };

   // m124_95 = W*in
   wire signed [14:0] m124_95;
   assign m124_95 =15'b0;

   // m124_96 = W*in
   wire signed [14:0] m124_96;
   assign m124_96 =15'b0;

   // m124_97 = W*in
   wire signed [14:0] m124_97;
   assign m124_97 =15'b0;

   // m124_98 = W*in
   wire signed [14:0] m124_98;
   assign m124_98 =15'b0;

   // m124_99 = W*in
   wire signed [14:0] m124_99;
   assign m124_99 ={ {3{in124[14]}} , in124[14:3] };

   // m124_100 = W*in
   wire signed [14:0] m124_100;
   assign m124_100 =15'b0;

   // m125_1 = W*in
   wire signed [14:0] m125_1;
   assign m125_1 =15'b0;

   // m125_2 = W*in
   wire signed [14:0] m125_2;
   assign m125_2 =15'b0;

   // m125_3 = W*in
   wire signed [14:0] m125_3;
   assign m125_3 =15'b0;

   // m125_4 = W*in
   wire signed [14:0] m125_4;
   assign m125_4 =15'b0;

   // m125_5 = W*in
   wire signed [14:0] m125_5;
   assign m125_5 =15'b0;

   // m125_6 = W*in
   wire signed [14:0] m125_6;
   assign m125_6 =15'b0;

   // m125_7 = W*in
   wire signed [14:0] m125_7;
   assign m125_7 =15'b0;

   // m125_8 = W*in
   wire signed [14:0] m125_8;
   assign m125_8 =15'b0;

   // m125_9 = W*in
   wire signed [14:0] m125_9;
   assign m125_9 =15'b0;

   // m125_10 = W*in
   wire signed [14:0] m125_10;
   assign m125_10 ={ {2{in125[14]}} , in125[14:2] };

   // m125_11 = W*in
   wire signed [14:0] m125_11;
   assign m125_11 =15'b0;

   // m125_12 = W*in
   wire signed [14:0] m125_12;
   assign m125_12 =15'b0;

   // m125_13 = W*in
   wire signed [14:0] m125_13;
   assign m125_13 =15'b0;

   // m125_14 = W*in
   wire signed [14:0] m125_14;
   assign m125_14 =15'b0;

   // m125_15 = W*in
   wire signed [14:0] m125_15;
   assign m125_15 =15'b0;

   // m125_16 = W*in
   wire signed [14:0] m125_16;
   assign m125_16 =15'b0;

   // m125_17 = W*in
   wire signed [14:0] m125_17;
   assign m125_17 =15'b0;

   // m125_18 = W*in
   wire signed [14:0] m125_18;
   assign m125_18 =15'b0;

   // m125_19 = W*in
   wire signed [14:0] m125_19;
   assign m125_19 ={ {4{in125[14]}} , in125[14:4] };

   // m125_20 = W*in
   wire signed [14:0] m125_20;
   assign m125_20 =15'b0;

   // m125_21 = W*in
   wire signed [14:0] m125_21;
   assign m125_21 ={ {4{in125[14]}} , in125[14:4] };

   // m125_22 = W*in
   wire signed [14:0] m125_22;
   assign m125_22 ={ {4{neg125[14]}} , neg125[14:4] };

   // m125_23 = W*in
   wire signed [14:0] m125_23;
   assign m125_23 =15'b0;

   // m125_24 = W*in
   wire signed [14:0] m125_24;
   assign m125_24 =15'b0;

   // m125_25 = W*in
   wire signed [14:0] m125_25;
   assign m125_25 =15'b0;

   // m125_26 = W*in
   wire signed [14:0] m125_26;
   assign m125_26 =15'b0;

   // m125_27 = W*in
   wire signed [14:0] m125_27;
   assign m125_27 =15'b0;

   // m125_28 = W*in
   wire signed [14:0] m125_28;
   assign m125_28 ={ {3{neg125[14]}} , neg125[14:3] };

   // m125_29 = W*in
   wire signed [14:0] m125_29;
   assign m125_29 ={ {4{in125[14]}} , in125[14:4] };

   // m125_30 = W*in
   wire signed [14:0] m125_30;
   assign m125_30 =15'b0;

   // m125_31 = W*in
   wire signed [14:0] m125_31;
   assign m125_31 =15'b0;

   // m125_32 = W*in
   wire signed [14:0] m125_32;
   assign m125_32 =15'b0;

   // m125_33 = W*in
   wire signed [14:0] m125_33;
   assign m125_33 =15'b0;

   // m125_34 = W*in
   wire signed [14:0] m125_34;
   assign m125_34 =15'b0;

   // m125_35 = W*in
   wire signed [14:0] m125_35;
   assign m125_35 =15'b0;

   // m125_36 = W*in
   wire signed [14:0] m125_36;
   assign m125_36 =15'b0;

   // m125_37 = W*in
   wire signed [14:0] m125_37;
   assign m125_37 =15'b0;

   // m125_38 = W*in
   wire signed [14:0] m125_38;
   assign m125_38 =15'b0;

   // m125_39 = W*in
   wire signed [14:0] m125_39;
   assign m125_39 =15'b0;

   // m125_40 = W*in
   wire signed [14:0] m125_40;
   assign m125_40 =15'b0;

   // m125_41 = W*in
   wire signed [14:0] m125_41;
   assign m125_41 =15'b0;

   // m125_42 = W*in
   wire signed [14:0] m125_42;
   assign m125_42 =15'b0;

   // m125_43 = W*in
   wire signed [14:0] m125_43;
   assign m125_43 =15'b0;

   // m125_44 = W*in
   wire signed [14:0] m125_44;
   assign m125_44 =15'b0;

   // m125_45 = W*in
   wire signed [14:0] m125_45;
   assign m125_45 ={ {3{neg125[14]}} , neg125[14:3] };

   // m125_46 = W*in
   wire signed [14:0] m125_46;
   assign m125_46 ={ {4{in125[14]}} , in125[14:4] };

   // m125_47 = W*in
   wire signed [14:0] m125_47;
   assign m125_47 ={ {3{in125[14]}} , in125[14:3] };

   // m125_48 = W*in
   wire signed [14:0] m125_48;
   assign m125_48 =15'b0;

   // m125_49 = W*in
   wire signed [14:0] m125_49;
   assign m125_49 =15'b0;

   // m125_50 = W*in
   wire signed [14:0] m125_50;
   assign m125_50 =15'b0;

   // m125_51 = W*in
   wire signed [14:0] m125_51;
   assign m125_51 =15'b0;

   // m125_52 = W*in
   wire signed [14:0] m125_52;
   assign m125_52 =15'b0;

   // m125_53 = W*in
   wire signed [14:0] m125_53;
   assign m125_53 =15'b0;

   // m125_54 = W*in
   wire signed [14:0] m125_54;
   assign m125_54 =15'b0;

   // m125_55 = W*in
   wire signed [14:0] m125_55;
   assign m125_55 ={ {3{neg125[14]}} , neg125[14:3] };

   // m125_56 = W*in
   wire signed [14:0] m125_56;
   assign m125_56 =15'b0;

   // m125_57 = W*in
   wire signed [14:0] m125_57;
   assign m125_57 =15'b0;

   // m125_58 = W*in
   wire signed [14:0] m125_58;
   assign m125_58 ={ {4{neg125[14]}} , neg125[14:4] };

   // m125_59 = W*in
   wire signed [14:0] m125_59;
   assign m125_59 =15'b0;

   // m125_60 = W*in
   wire signed [14:0] m125_60;
   assign m125_60 ={ {4{neg125[14]}} , neg125[14:4] };

   // m125_61 = W*in
   wire signed [14:0] m125_61;
   assign m125_61 ={ {4{neg125[14]}} , neg125[14:4] };

   // m125_62 = W*in
   wire signed [14:0] m125_62;
   assign m125_62 =15'b0;

   // m125_63 = W*in
   wire signed [14:0] m125_63;
   assign m125_63 ={ {3{in125[14]}} , in125[14:3] };

   // m125_64 = W*in
   wire signed [14:0] m125_64;
   assign m125_64 ={ {4{neg125[14]}} , neg125[14:4] };

   // m125_65 = W*in
   wire signed [14:0] m125_65;
   assign m125_65 ={ {4{in125[14]}} , in125[14:4] };

   // m125_66 = W*in
   wire signed [14:0] m125_66;
   assign m125_66 ={ {4{in125[14]}} , in125[14:4] };

   // m125_67 = W*in
   wire signed [14:0] m125_67;
   assign m125_67 =15'b0;

   // m125_68 = W*in
   wire signed [14:0] m125_68;
   assign m125_68 ={ {3{neg125[14]}} , neg125[14:3] };

   // m125_69 = W*in
   wire signed [14:0] m125_69;
   assign m125_69 =15'b0;

   // m125_70 = W*in
   wire signed [14:0] m125_70;
   assign m125_70 =15'b0;

   // m125_71 = W*in
   wire signed [14:0] m125_71;
   assign m125_71 =15'b0;

   // m125_72 = W*in
   wire signed [14:0] m125_72;
   assign m125_72 =15'b0;

   // m125_73 = W*in
   wire signed [14:0] m125_73;
   assign m125_73 =15'b0;

   // m125_74 = W*in
   wire signed [14:0] m125_74;
   assign m125_74 =15'b0;

   // m125_75 = W*in
   wire signed [14:0] m125_75;
   assign m125_75 =15'b0;

   // m125_76 = W*in
   wire signed [14:0] m125_76;
   assign m125_76 =15'b0;

   // m125_77 = W*in
   wire signed [14:0] m125_77;
   assign m125_77 =15'b0;

   // m125_78 = W*in
   wire signed [14:0] m125_78;
   assign m125_78 =15'b0;

   // m125_79 = W*in
   wire signed [14:0] m125_79;
   assign m125_79 ={ {3{in125[14]}} , in125[14:3] };

   // m125_80 = W*in
   wire signed [14:0] m125_80;
   assign m125_80 =15'b0;

   // m125_81 = W*in
   wire signed [14:0] m125_81;
   assign m125_81 =15'b0;

   // m125_82 = W*in
   wire signed [14:0] m125_82;
   assign m125_82 =15'b0;

   // m125_83 = W*in
   wire signed [14:0] m125_83;
   assign m125_83 =15'b0;

   // m125_84 = W*in
   wire signed [14:0] m125_84;
   assign m125_84 =15'b0;

   // m125_85 = W*in
   wire signed [14:0] m125_85;
   assign m125_85 =15'b0;

   // m125_86 = W*in
   wire signed [14:0] m125_86;
   assign m125_86 =15'b0;

   // m125_87 = W*in
   wire signed [14:0] m125_87;
   assign m125_87 =15'b0;

   // m125_88 = W*in
   wire signed [14:0] m125_88;
   assign m125_88 =15'b0;

   // m125_89 = W*in
   wire signed [14:0] m125_89;
   assign m125_89 =15'b0;

   // m125_90 = W*in
   wire signed [14:0] m125_90;
   assign m125_90 =15'b0;

   // m125_91 = W*in
   wire signed [14:0] m125_91;
   assign m125_91 =15'b0;

   // m125_92 = W*in
   wire signed [14:0] m125_92;
   assign m125_92 =15'b0;

   // m125_93 = W*in
   wire signed [14:0] m125_93;
   assign m125_93 =15'b0;

   // m125_94 = W*in
   wire signed [14:0] m125_94;
   assign m125_94 =15'b0;

   // m125_95 = W*in
   wire signed [14:0] m125_95;
   assign m125_95 =15'b0;

   // m125_96 = W*in
   wire signed [14:0] m125_96;
   assign m125_96 =15'b0;

   // m125_97 = W*in
   wire signed [14:0] m125_97;
   assign m125_97 =15'b0;

   // m125_98 = W*in
   wire signed [14:0] m125_98;
   assign m125_98 =15'b0;

   // m125_99 = W*in
   wire signed [14:0] m125_99;
   assign m125_99 =15'b0;

   // m125_100 = W*in
   wire signed [14:0] m125_100;
   assign m125_100 =15'b0;

   // m126_1 = W*in
   wire signed [14:0] m126_1;
   assign m126_1 =15'b0;

   // m126_2 = W*in
   wire signed [14:0] m126_2;
   assign m126_2 =15'b0;

   // m126_3 = W*in
   wire signed [14:0] m126_3;
   assign m126_3 =15'b0;

   // m126_4 = W*in
   wire signed [14:0] m126_4;
   assign m126_4 =15'b0;

   // m126_5 = W*in
   wire signed [14:0] m126_5;
   assign m126_5 ={ {3{neg126[14]}} , neg126[14:3] };

   // m126_6 = W*in
   wire signed [14:0] m126_6;
   assign m126_6 =15'b0;

   // m126_7 = W*in
   wire signed [14:0] m126_7;
   assign m126_7 =15'b0;

   // m126_8 = W*in
   wire signed [14:0] m126_8;
   assign m126_8 =15'b0;

   // m126_9 = W*in
   wire signed [14:0] m126_9;
   assign m126_9 =15'b0;

   // m126_10 = W*in
   wire signed [14:0] m126_10;
   assign m126_10 =15'b0;

   // m126_11 = W*in
   wire signed [14:0] m126_11;
   assign m126_11 ={ {3{neg126[14]}} , neg126[14:3] };

   // m126_12 = W*in
   wire signed [14:0] m126_12;
   assign m126_12 =15'b0;

   // m126_13 = W*in
   wire signed [14:0] m126_13;
   assign m126_13 =15'b0;

   // m126_14 = W*in
   wire signed [14:0] m126_14;
   assign m126_14 ={ {4{neg126[14]}} , neg126[14:4] };

   // m126_15 = W*in
   wire signed [14:0] m126_15;
   assign m126_15 =15'b0;

   // m126_16 = W*in
   wire signed [14:0] m126_16;
   assign m126_16 =15'b0;

   // m126_17 = W*in
   wire signed [14:0] m126_17;
   assign m126_17 =15'b0;

   // m126_18 = W*in
   wire signed [14:0] m126_18;
   assign m126_18 =15'b0;

   // m126_19 = W*in
   wire signed [14:0] m126_19;
   assign m126_19 =15'b0;

   // m126_20 = W*in
   wire signed [14:0] m126_20;
   assign m126_20 =15'b0;

   // m126_21 = W*in
   wire signed [14:0] m126_21;
   assign m126_21 ={ {4{neg126[14]}} , neg126[14:4] };

   // m126_22 = W*in
   wire signed [14:0] m126_22;
   assign m126_22 =15'b0;

   // m126_23 = W*in
   wire signed [14:0] m126_23;
   assign m126_23 ={ {4{in126[14]}} , in126[14:4] };

   // m126_24 = W*in
   wire signed [14:0] m126_24;
   assign m126_24 =15'b0;

   // m126_25 = W*in
   wire signed [14:0] m126_25;
   assign m126_25 =15'b0;

   // m126_26 = W*in
   wire signed [14:0] m126_26;
   assign m126_26 =15'b0;

   // m126_27 = W*in
   wire signed [14:0] m126_27;
   assign m126_27 ={ {4{in126[14]}} , in126[14:4] };

   // m126_28 = W*in
   wire signed [14:0] m126_28;
   assign m126_28 =15'b0;

   // m126_29 = W*in
   wire signed [14:0] m126_29;
   assign m126_29 =15'b0;

   // m126_30 = W*in
   wire signed [14:0] m126_30;
   assign m126_30 =15'b0;

   // m126_31 = W*in
   wire signed [14:0] m126_31;
   assign m126_31 =15'b0;

   // m126_32 = W*in
   wire signed [14:0] m126_32;
   assign m126_32 =15'b0;

   // m126_33 = W*in
   wire signed [14:0] m126_33;
   assign m126_33 =15'b0;

   // m126_34 = W*in
   wire signed [14:0] m126_34;
   assign m126_34 =15'b0;

   // m126_35 = W*in
   wire signed [14:0] m126_35;
   assign m126_35 =15'b0;

   // m126_36 = W*in
   wire signed [14:0] m126_36;
   assign m126_36 =15'b0;

   // m126_37 = W*in
   wire signed [14:0] m126_37;
   assign m126_37 =15'b0;

   // m126_38 = W*in
   wire signed [14:0] m126_38;
   assign m126_38 =15'b0;

   // m126_39 = W*in
   wire signed [14:0] m126_39;
   assign m126_39 =15'b0;

   // m126_40 = W*in
   wire signed [14:0] m126_40;
   assign m126_40 =15'b0;

   // m126_41 = W*in
   wire signed [14:0] m126_41;
   assign m126_41 ={ {4{in126[14]}} , in126[14:4] };

   // m126_42 = W*in
   wire signed [14:0] m126_42;
   assign m126_42 =15'b0;

   // m126_43 = W*in
   wire signed [14:0] m126_43;
   assign m126_43 =15'b0;

   // m126_44 = W*in
   wire signed [14:0] m126_44;
   assign m126_44 =15'b0;

   // m126_45 = W*in
   wire signed [14:0] m126_45;
   assign m126_45 =15'b0;

   // m126_46 = W*in
   wire signed [14:0] m126_46;
   assign m126_46 =15'b0;

   // m126_47 = W*in
   wire signed [14:0] m126_47;
   assign m126_47 ={ {4{in126[14]}} , in126[14:4] };

   // m126_48 = W*in
   wire signed [14:0] m126_48;
   assign m126_48 =15'b0;

   // m126_49 = W*in
   wire signed [14:0] m126_49;
   assign m126_49 =15'b0;

   // m126_50 = W*in
   wire signed [14:0] m126_50;
   assign m126_50 =15'b0;

   // m126_51 = W*in
   wire signed [14:0] m126_51;
   assign m126_51 =15'b0;

   // m126_52 = W*in
   wire signed [14:0] m126_52;
   assign m126_52 =15'b0;

   // m126_53 = W*in
   wire signed [14:0] m126_53;
   assign m126_53 ={ {4{in126[14]}} , in126[14:4] };

   // m126_54 = W*in
   wire signed [14:0] m126_54;
   assign m126_54 =15'b0;

   // m126_55 = W*in
   wire signed [14:0] m126_55;
   assign m126_55 ={ {4{neg126[14]}} , neg126[14:4] };

   // m126_56 = W*in
   wire signed [14:0] m126_56;
   assign m126_56 =15'b0;

   // m126_57 = W*in
   wire signed [14:0] m126_57;
   assign m126_57 ={ {4{in126[14]}} , in126[14:4] };

   // m126_58 = W*in
   wire signed [14:0] m126_58;
   assign m126_58 =15'b0;

   // m126_59 = W*in
   wire signed [14:0] m126_59;
   assign m126_59 =15'b0;

   // m126_60 = W*in
   wire signed [14:0] m126_60;
   assign m126_60 =15'b0;

   // m126_61 = W*in
   wire signed [14:0] m126_61;
   assign m126_61 =15'b0;

   // m126_62 = W*in
   wire signed [14:0] m126_62;
   assign m126_62 =15'b0;

   // m126_63 = W*in
   wire signed [14:0] m126_63;
   assign m126_63 =15'b0;

   // m126_64 = W*in
   wire signed [14:0] m126_64;
   assign m126_64 =15'b0;

   // m126_65 = W*in
   wire signed [14:0] m126_65;
   assign m126_65 ={ {4{neg126[14]}} , neg126[14:4] };

   // m126_66 = W*in
   wire signed [14:0] m126_66;
   assign m126_66 =15'b0;

   // m126_67 = W*in
   wire signed [14:0] m126_67;
   assign m126_67 =15'b0;

   // m126_68 = W*in
   wire signed [14:0] m126_68;
   assign m126_68 =15'b0;

   // m126_69 = W*in
   wire signed [14:0] m126_69;
   assign m126_69 =15'b0;

   // m126_70 = W*in
   wire signed [14:0] m126_70;
   assign m126_70 =15'b0;

   // m126_71 = W*in
   wire signed [14:0] m126_71;
   assign m126_71 =15'b0;

   // m126_72 = W*in
   wire signed [14:0] m126_72;
   assign m126_72 =15'b0;

   // m126_73 = W*in
   wire signed [14:0] m126_73;
   assign m126_73 =15'b0;

   // m126_74 = W*in
   wire signed [14:0] m126_74;
   assign m126_74 ={ {4{neg126[14]}} , neg126[14:4] };

   // m126_75 = W*in
   wire signed [14:0] m126_75;
   assign m126_75 =15'b0;

   // m126_76 = W*in
   wire signed [14:0] m126_76;
   assign m126_76 ={ {3{neg126[14]}} , neg126[14:3] };

   // m126_77 = W*in
   wire signed [14:0] m126_77;
   assign m126_77 ={ {4{neg126[14]}} , neg126[14:4] };

   // m126_78 = W*in
   wire signed [14:0] m126_78;
   assign m126_78 =15'b0;

   // m126_79 = W*in
   wire signed [14:0] m126_79;
   assign m126_79 ={ {3{neg126[14]}} , neg126[14:3] };

   // m126_80 = W*in
   wire signed [14:0] m126_80;
   assign m126_80 =15'b0;

   // m126_81 = W*in
   wire signed [14:0] m126_81;
   assign m126_81 ={ {4{in126[14]}} , in126[14:4] };

   // m126_82 = W*in
   wire signed [14:0] m126_82;
   assign m126_82 =15'b0;

   // m126_83 = W*in
   wire signed [14:0] m126_83;
   assign m126_83 =15'b0;

   // m126_84 = W*in
   wire signed [14:0] m126_84;
   assign m126_84 =15'b0;

   // m126_85 = W*in
   wire signed [14:0] m126_85;
   assign m126_85 =15'b0;

   // m126_86 = W*in
   wire signed [14:0] m126_86;
   assign m126_86 =15'b0;

   // m126_87 = W*in
   wire signed [14:0] m126_87;
   assign m126_87 =15'b0;

   // m126_88 = W*in
   wire signed [14:0] m126_88;
   assign m126_88 ={ {3{neg126[14]}} , neg126[14:3] };

   // m126_89 = W*in
   wire signed [14:0] m126_89;
   assign m126_89 =15'b0;

   // m126_90 = W*in
   wire signed [14:0] m126_90;
   assign m126_90 =15'b0;

   // m126_91 = W*in
   wire signed [14:0] m126_91;
   assign m126_91 =15'b0;

   // m126_92 = W*in
   wire signed [14:0] m126_92;
   assign m126_92 =15'b0;

   // m126_93 = W*in
   wire signed [14:0] m126_93;
   assign m126_93 =15'b0;

   // m126_94 = W*in
   wire signed [14:0] m126_94;
   assign m126_94 =15'b0;

   // m126_95 = W*in
   wire signed [14:0] m126_95;
   assign m126_95 =15'b0;

   // m126_96 = W*in
   wire signed [14:0] m126_96;
   assign m126_96 =15'b0;

   // m126_97 = W*in
   wire signed [14:0] m126_97;
   assign m126_97 =15'b0;

   // m126_98 = W*in
   wire signed [14:0] m126_98;
   assign m126_98 =15'b0;

   // m126_99 = W*in
   wire signed [14:0] m126_99;
   assign m126_99 =15'b0;

   // m126_100 = W*in
   wire signed [14:0] m126_100;
   assign m126_100 =15'b0;

   // m127_1 = W*in
   wire signed [14:0] m127_1;
   assign m127_1 =15'b0;

   // m127_2 = W*in
   wire signed [14:0] m127_2;
   assign m127_2 =15'b0;

   // m127_3 = W*in
   wire signed [14:0] m127_3;
   assign m127_3 =15'b0;

   // m127_4 = W*in
   wire signed [14:0] m127_4;
   assign m127_4 =15'b0;

   // m127_5 = W*in
   wire signed [14:0] m127_5;
   assign m127_5 ={ {4{in127[14]}} , in127[14:4] };

   // m127_6 = W*in
   wire signed [14:0] m127_6;
   assign m127_6 =15'b0;

   // m127_7 = W*in
   wire signed [14:0] m127_7;
   assign m127_7 =15'b0;

   // m127_8 = W*in
   wire signed [14:0] m127_8;
   assign m127_8 =15'b0;

   // m127_9 = W*in
   wire signed [14:0] m127_9;
   assign m127_9 =15'b0;

   // m127_10 = W*in
   wire signed [14:0] m127_10;
   assign m127_10 =15'b0;

   // m127_11 = W*in
   wire signed [14:0] m127_11;
   assign m127_11 =15'b0;

   // m127_12 = W*in
   wire signed [14:0] m127_12;
   assign m127_12 =15'b0;

   // m127_13 = W*in
   wire signed [14:0] m127_13;
   assign m127_13 =15'b0;

   // m127_14 = W*in
   wire signed [14:0] m127_14;
   assign m127_14 =15'b0;

   // m127_15 = W*in
   wire signed [14:0] m127_15;
   assign m127_15 =15'b0;

   // m127_16 = W*in
   wire signed [14:0] m127_16;
   assign m127_16 =15'b0;

   // m127_17 = W*in
   wire signed [14:0] m127_17;
   assign m127_17 =15'b0;

   // m127_18 = W*in
   wire signed [14:0] m127_18;
   assign m127_18 ={ {4{in127[14]}} , in127[14:4] };

   // m127_19 = W*in
   wire signed [14:0] m127_19;
   assign m127_19 =15'b0;

   // m127_20 = W*in
   wire signed [14:0] m127_20;
   assign m127_20 =15'b0;

   // m127_21 = W*in
   wire signed [14:0] m127_21;
   assign m127_21 =15'b0;

   // m127_22 = W*in
   wire signed [14:0] m127_22;
   assign m127_22 =15'b0;

   // m127_23 = W*in
   wire signed [14:0] m127_23;
   assign m127_23 =15'b0;

   // m127_24 = W*in
   wire signed [14:0] m127_24;
   assign m127_24 =15'b0;

   // m127_25 = W*in
   wire signed [14:0] m127_25;
   assign m127_25 =15'b0;

   // m127_26 = W*in
   wire signed [14:0] m127_26;
   assign m127_26 =15'b0;

   // m127_27 = W*in
   wire signed [14:0] m127_27;
   assign m127_27 =15'b0;

   // m127_28 = W*in
   wire signed [14:0] m127_28;
   assign m127_28 =15'b0;

   // m127_29 = W*in
   wire signed [14:0] m127_29;
   assign m127_29 =15'b0;

   // m127_30 = W*in
   wire signed [14:0] m127_30;
   assign m127_30 =15'b0;

   // m127_31 = W*in
   wire signed [14:0] m127_31;
   assign m127_31 =15'b0;

   // m127_32 = W*in
   wire signed [14:0] m127_32;
   assign m127_32 =15'b0;

   // m127_33 = W*in
   wire signed [14:0] m127_33;
   assign m127_33 =15'b0;

   // m127_34 = W*in
   wire signed [14:0] m127_34;
   assign m127_34 =15'b0;

   // m127_35 = W*in
   wire signed [14:0] m127_35;
   assign m127_35 =15'b0;

   // m127_36 = W*in
   wire signed [14:0] m127_36;
   assign m127_36 =15'b0;

   // m127_37 = W*in
   wire signed [14:0] m127_37;
   assign m127_37 =15'b0;

   // m127_38 = W*in
   wire signed [14:0] m127_38;
   assign m127_38 =15'b0;

   // m127_39 = W*in
   wire signed [14:0] m127_39;
   assign m127_39 =15'b0;

   // m127_40 = W*in
   wire signed [14:0] m127_40;
   assign m127_40 =15'b0;

   // m127_41 = W*in
   wire signed [14:0] m127_41;
   assign m127_41 =15'b0;

   // m127_42 = W*in
   wire signed [14:0] m127_42;
   assign m127_42 ={ {4{neg127[14]}} , neg127[14:4] };

   // m127_43 = W*in
   wire signed [14:0] m127_43;
   assign m127_43 =15'b0;

   // m127_44 = W*in
   wire signed [14:0] m127_44;
   assign m127_44 =15'b0;

   // m127_45 = W*in
   wire signed [14:0] m127_45;
   assign m127_45 =15'b0;

   // m127_46 = W*in
   wire signed [14:0] m127_46;
   assign m127_46 =15'b0;

   // m127_47 = W*in
   wire signed [14:0] m127_47;
   assign m127_47 =15'b0;

   // m127_48 = W*in
   wire signed [14:0] m127_48;
   assign m127_48 =15'b0;

   // m127_49 = W*in
   wire signed [14:0] m127_49;
   assign m127_49 =15'b0;

   // m127_50 = W*in
   wire signed [14:0] m127_50;
   assign m127_50 =15'b0;

   // m127_51 = W*in
   wire signed [14:0] m127_51;
   assign m127_51 =15'b0;

   // m127_52 = W*in
   wire signed [14:0] m127_52;
   assign m127_52 =15'b0;

   // m127_53 = W*in
   wire signed [14:0] m127_53;
   assign m127_53 =15'b0;

   // m127_54 = W*in
   wire signed [14:0] m127_54;
   assign m127_54 =15'b0;

   // m127_55 = W*in
   wire signed [14:0] m127_55;
   assign m127_55 =15'b0;

   // m127_56 = W*in
   wire signed [14:0] m127_56;
   assign m127_56 =15'b0;

   // m127_57 = W*in
   wire signed [14:0] m127_57;
   assign m127_57 =15'b0;

   // m127_58 = W*in
   wire signed [14:0] m127_58;
   assign m127_58 =15'b0;

   // m127_59 = W*in
   wire signed [14:0] m127_59;
   assign m127_59 =15'b0;

   // m127_60 = W*in
   wire signed [14:0] m127_60;
   assign m127_60 =15'b0;

   // m127_61 = W*in
   wire signed [14:0] m127_61;
   assign m127_61 =15'b0;

   // m127_62 = W*in
   wire signed [14:0] m127_62;
   assign m127_62 =15'b0;

   // m127_63 = W*in
   wire signed [14:0] m127_63;
   assign m127_63 =15'b0;

   // m127_64 = W*in
   wire signed [14:0] m127_64;
   assign m127_64 =15'b0;

   // m127_65 = W*in
   wire signed [14:0] m127_65;
   assign m127_65 =15'b0;

   // m127_66 = W*in
   wire signed [14:0] m127_66;
   assign m127_66 =15'b0;

   // m127_67 = W*in
   wire signed [14:0] m127_67;
   assign m127_67 =15'b0;

   // m127_68 = W*in
   wire signed [14:0] m127_68;
   assign m127_68 =15'b0;

   // m127_69 = W*in
   wire signed [14:0] m127_69;
   assign m127_69 =15'b0;

   // m127_70 = W*in
   wire signed [14:0] m127_70;
   assign m127_70 =15'b0;

   // m127_71 = W*in
   wire signed [14:0] m127_71;
   assign m127_71 =15'b0;

   // m127_72 = W*in
   wire signed [14:0] m127_72;
   assign m127_72 =15'b0;

   // m127_73 = W*in
   wire signed [14:0] m127_73;
   assign m127_73 =15'b0;

   // m127_74 = W*in
   wire signed [14:0] m127_74;
   assign m127_74 =15'b0;

   // m127_75 = W*in
   wire signed [14:0] m127_75;
   assign m127_75 =15'b0;

   // m127_76 = W*in
   wire signed [14:0] m127_76;
   assign m127_76 =15'b0;

   // m127_77 = W*in
   wire signed [14:0] m127_77;
   assign m127_77 =15'b0;

   // m127_78 = W*in
   wire signed [14:0] m127_78;
   assign m127_78 ={ {3{in127[14]}} , in127[14:3] };

   // m127_79 = W*in
   wire signed [14:0] m127_79;
   assign m127_79 =15'b0;

   // m127_80 = W*in
   wire signed [14:0] m127_80;
   assign m127_80 =15'b0;

   // m127_81 = W*in
   wire signed [14:0] m127_81;
   assign m127_81 =15'b0;

   // m127_82 = W*in
   wire signed [14:0] m127_82;
   assign m127_82 ={ {3{neg127[14]}} , neg127[14:3] };

   // m127_83 = W*in
   wire signed [14:0] m127_83;
   assign m127_83 ={ {4{in127[14]}} , in127[14:4] };

   // m127_84 = W*in
   wire signed [14:0] m127_84;
   assign m127_84 =15'b0;

   // m127_85 = W*in
   wire signed [14:0] m127_85;
   assign m127_85 ={ {4{neg127[14]}} , neg127[14:4] };

   // m127_86 = W*in
   wire signed [14:0] m127_86;
   assign m127_86 =15'b0;

   // m127_87 = W*in
   wire signed [14:0] m127_87;
   assign m127_87 =15'b0;

   // m127_88 = W*in
   wire signed [14:0] m127_88;
   assign m127_88 =15'b0;

   // m127_89 = W*in
   wire signed [14:0] m127_89;
   assign m127_89 =15'b0;

   // m127_90 = W*in
   wire signed [14:0] m127_90;
   assign m127_90 =15'b0;

   // m127_91 = W*in
   wire signed [14:0] m127_91;
   assign m127_91 =15'b0;

   // m127_92 = W*in
   wire signed [14:0] m127_92;
   assign m127_92 =15'b0;

   // m127_93 = W*in
   wire signed [14:0] m127_93;
   assign m127_93 =15'b0;

   // m127_94 = W*in
   wire signed [14:0] m127_94;
   assign m127_94 ={ {3{in127[14]}} , in127[14:3] };

   // m127_95 = W*in
   wire signed [14:0] m127_95;
   assign m127_95 =15'b0;

   // m127_96 = W*in
   wire signed [14:0] m127_96;
   assign m127_96 =15'b0;

   // m127_97 = W*in
   wire signed [14:0] m127_97;
   assign m127_97 =15'b0;

   // m127_98 = W*in
   wire signed [14:0] m127_98;
   assign m127_98 =15'b0;

   // m127_99 = W*in
   wire signed [14:0] m127_99;
   assign m127_99 =15'b0;

   // m127_100 = W*in
   wire signed [14:0] m127_100;
   assign m127_100 =15'b0;

   // m128_1 = W*in
   wire signed [14:0] m128_1;
   assign m128_1 =15'b0;

   // m128_2 = W*in
   wire signed [14:0] m128_2;
   assign m128_2 =15'b0;

   // m128_3 = W*in
   wire signed [14:0] m128_3;
   assign m128_3 =15'b0;

   // m128_4 = W*in
   wire signed [14:0] m128_4;
   assign m128_4 ={ {3{in128[14]}} , in128[14:3] };

   // m128_5 = W*in
   wire signed [14:0] m128_5;
   assign m128_5 ={ {4{in128[14]}} , in128[14:4] };

   // m128_6 = W*in
   wire signed [14:0] m128_6;
   assign m128_6 =15'b0;

   // m128_7 = W*in
   wire signed [14:0] m128_7;
   assign m128_7 =15'b0;

   // m128_8 = W*in
   wire signed [14:0] m128_8;
   assign m128_8 =15'b0;

   // m128_9 = W*in
   wire signed [14:0] m128_9;
   assign m128_9 =15'b0;

   // m128_10 = W*in
   wire signed [14:0] m128_10;
   assign m128_10 =15'b0;

   // m128_11 = W*in
   wire signed [14:0] m128_11;
   assign m128_11 =15'b0;

   // m128_12 = W*in
   wire signed [14:0] m128_12;
   assign m128_12 =15'b0;

   // m128_13 = W*in
   wire signed [14:0] m128_13;
   assign m128_13 ={ {2{in128[14]}} , in128[14:2] };

   // m128_14 = W*in
   wire signed [14:0] m128_14;
   assign m128_14 =15'b0;

   // m128_15 = W*in
   wire signed [14:0] m128_15;
   assign m128_15 =15'b0;

   // m128_16 = W*in
   wire signed [14:0] m128_16;
   assign m128_16 =15'b0;

   // m128_17 = W*in
   wire signed [14:0] m128_17;
   assign m128_17 =15'b0;

   // m128_18 = W*in
   wire signed [14:0] m128_18;
   assign m128_18 ={ {3{in128[14]}} , in128[14:3] };

   // m128_19 = W*in
   wire signed [14:0] m128_19;
   assign m128_19 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_20 = W*in
   wire signed [14:0] m128_20;
   assign m128_20 =15'b0;

   // m128_21 = W*in
   wire signed [14:0] m128_21;
   assign m128_21 =15'b0;

   // m128_22 = W*in
   wire signed [14:0] m128_22;
   assign m128_22 ={ {3{in128[14]}} , in128[14:3] };

   // m128_23 = W*in
   wire signed [14:0] m128_23;
   assign m128_23 =15'b0;

   // m128_24 = W*in
   wire signed [14:0] m128_24;
   assign m128_24 =15'b0;

   // m128_25 = W*in
   wire signed [14:0] m128_25;
   assign m128_25 ={ {4{in128[14]}} , in128[14:4] };

   // m128_26 = W*in
   wire signed [14:0] m128_26;
   assign m128_26 ={ {4{neg128[14]}} , neg128[14:4] };

   // m128_27 = W*in
   wire signed [14:0] m128_27;
   assign m128_27 =15'b0;

   // m128_28 = W*in
   wire signed [14:0] m128_28;
   assign m128_28 ={ {4{in128[14]}} , in128[14:4] };

   // m128_29 = W*in
   wire signed [14:0] m128_29;
   assign m128_29 ={ {4{in128[14]}} , in128[14:4] };

   // m128_30 = W*in
   wire signed [14:0] m128_30;
   assign m128_30 =15'b0;

   // m128_31 = W*in
   wire signed [14:0] m128_31;
   assign m128_31 ={ {4{neg128[14]}} , neg128[14:4] };

   // m128_32 = W*in
   wire signed [14:0] m128_32;
   assign m128_32 =15'b0;

   // m128_33 = W*in
   wire signed [14:0] m128_33;
   assign m128_33 =15'b0;

   // m128_34 = W*in
   wire signed [14:0] m128_34;
   assign m128_34 =15'b0;

   // m128_35 = W*in
   wire signed [14:0] m128_35;
   assign m128_35 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_36 = W*in
   wire signed [14:0] m128_36;
   assign m128_36 =15'b0;

   // m128_37 = W*in
   wire signed [14:0] m128_37;
   assign m128_37 =15'b0;

   // m128_38 = W*in
   wire signed [14:0] m128_38;
   assign m128_38 ={ {3{in128[14]}} , in128[14:3] };

   // m128_39 = W*in
   wire signed [14:0] m128_39;
   assign m128_39 =15'b0;

   // m128_40 = W*in
   wire signed [14:0] m128_40;
   assign m128_40 =15'b0;

   // m128_41 = W*in
   wire signed [14:0] m128_41;
   assign m128_41 =15'b0;

   // m128_42 = W*in
   wire signed [14:0] m128_42;
   assign m128_42 =15'b0;

   // m128_43 = W*in
   wire signed [14:0] m128_43;
   assign m128_43 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_44 = W*in
   wire signed [14:0] m128_44;
   assign m128_44 =15'b0;

   // m128_45 = W*in
   wire signed [14:0] m128_45;
   assign m128_45 =15'b0;

   // m128_46 = W*in
   wire signed [14:0] m128_46;
   assign m128_46 =15'b0;

   // m128_47 = W*in
   wire signed [14:0] m128_47;
   assign m128_47 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_48 = W*in
   wire signed [14:0] m128_48;
   assign m128_48 =15'b0;

   // m128_49 = W*in
   wire signed [14:0] m128_49;
   assign m128_49 =15'b0;

   // m128_50 = W*in
   wire signed [14:0] m128_50;
   assign m128_50 =15'b0;

   // m128_51 = W*in
   wire signed [14:0] m128_51;
   assign m128_51 =15'b0;

   // m128_52 = W*in
   wire signed [14:0] m128_52;
   assign m128_52 =15'b0;

   // m128_53 = W*in
   wire signed [14:0] m128_53;
   assign m128_53 =15'b0;

   // m128_54 = W*in
   wire signed [14:0] m128_54;
   assign m128_54 =15'b0;

   // m128_55 = W*in
   wire signed [14:0] m128_55;
   assign m128_55 ={ {3{in128[14]}} , in128[14:3] };

   // m128_56 = W*in
   wire signed [14:0] m128_56;
   assign m128_56 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_57 = W*in
   wire signed [14:0] m128_57;
   assign m128_57 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_58 = W*in
   wire signed [14:0] m128_58;
   assign m128_58 =15'b0;

   // m128_59 = W*in
   wire signed [14:0] m128_59;
   assign m128_59 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_60 = W*in
   wire signed [14:0] m128_60;
   assign m128_60 ={ {3{in128[14]}} , in128[14:3] };

   // m128_61 = W*in
   wire signed [14:0] m128_61;
   assign m128_61 ={ {4{in128[14]}} , in128[14:4] };

   // m128_62 = W*in
   wire signed [14:0] m128_62;
   assign m128_62 =15'b0;

   // m128_63 = W*in
   wire signed [14:0] m128_63;
   assign m128_63 ={ {3{in128[14]}} , in128[14:3] };

   // m128_64 = W*in
   wire signed [14:0] m128_64;
   assign m128_64 =15'b0;

   // m128_65 = W*in
   wire signed [14:0] m128_65;
   assign m128_65 =15'b0;

   // m128_66 = W*in
   wire signed [14:0] m128_66;
   assign m128_66 =15'b0;

   // m128_67 = W*in
   wire signed [14:0] m128_67;
   assign m128_67 ={ {4{in128[14]}} , in128[14:4] };

   // m128_68 = W*in
   wire signed [14:0] m128_68;
   assign m128_68 ={ {3{in128[14]}} , in128[14:3] };

   // m128_69 = W*in
   wire signed [14:0] m128_69;
   assign m128_69 ={ {4{in128[14]}} , in128[14:4] };

   // m128_70 = W*in
   wire signed [14:0] m128_70;
   assign m128_70 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_71 = W*in
   wire signed [14:0] m128_71;
   assign m128_71 =15'b0;

   // m128_72 = W*in
   wire signed [14:0] m128_72;
   assign m128_72 ={ {3{in128[14]}} , in128[14:3] };

   // m128_73 = W*in
   wire signed [14:0] m128_73;
   assign m128_73 =15'b0;

   // m128_74 = W*in
   wire signed [14:0] m128_74;
   assign m128_74 ={ {4{neg128[14]}} , neg128[14:4] };

   // m128_75 = W*in
   wire signed [14:0] m128_75;
   assign m128_75 =15'b0;

   // m128_76 = W*in
   wire signed [14:0] m128_76;
   assign m128_76 =15'b0;

   // m128_77 = W*in
   wire signed [14:0] m128_77;
   assign m128_77 =15'b0;

   // m128_78 = W*in
   wire signed [14:0] m128_78;
   assign m128_78 ={ {3{in128[14]}} , in128[14:3] };

   // m128_79 = W*in
   wire signed [14:0] m128_79;
   assign m128_79 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_80 = W*in
   wire signed [14:0] m128_80;
   assign m128_80 ={ {3{in128[14]}} , in128[14:3] };

   // m128_81 = W*in
   wire signed [14:0] m128_81;
   assign m128_81 =15'b0;

   // m128_82 = W*in
   wire signed [14:0] m128_82;
   assign m128_82 =15'b0;

   // m128_83 = W*in
   wire signed [14:0] m128_83;
   assign m128_83 =15'b0;

   // m128_84 = W*in
   wire signed [14:0] m128_84;
   assign m128_84 =15'b0;

   // m128_85 = W*in
   wire signed [14:0] m128_85;
   assign m128_85 =15'b0;

   // m128_86 = W*in
   wire signed [14:0] m128_86;
   assign m128_86 =15'b0;

   // m128_87 = W*in
   wire signed [14:0] m128_87;
   assign m128_87 =15'b0;

   // m128_88 = W*in
   wire signed [14:0] m128_88;
   assign m128_88 =15'b0;

   // m128_89 = W*in
   wire signed [14:0] m128_89;
   assign m128_89 =15'b0;

   // m128_90 = W*in
   wire signed [14:0] m128_90;
   assign m128_90 =15'b0;

   // m128_91 = W*in
   wire signed [14:0] m128_91;
   assign m128_91 =15'b0;

   // m128_92 = W*in
   wire signed [14:0] m128_92;
   assign m128_92 =15'b0;

   // m128_93 = W*in
   wire signed [14:0] m128_93;
   assign m128_93 =15'b0;

   // m128_94 = W*in
   wire signed [14:0] m128_94;
   assign m128_94 ={ {3{neg128[14]}} , neg128[14:3] };

   // m128_95 = W*in
   wire signed [14:0] m128_95;
   assign m128_95 ={ {4{neg128[14]}} , neg128[14:4] };

   // m128_96 = W*in
   wire signed [14:0] m128_96;
   assign m128_96 ={ {4{in128[14]}} , in128[14:4] };

   // m128_97 = W*in
   wire signed [14:0] m128_97;
   assign m128_97 ={ {3{in128[14]}} , in128[14:3] };

   // m128_98 = W*in
   wire signed [14:0] m128_98;
   assign m128_98 =15'b0;

   // m128_99 = W*in
   wire signed [14:0] m128_99;
   assign m128_99 =15'b0;

   // m128_100 = W*in
   wire signed [14:0] m128_100;
   assign m128_100 =15'b0;

   // m129_1 = W*in
   wire signed [14:0] m129_1;
   assign m129_1 =15'b0;

   // m129_2 = W*in
   wire signed [14:0] m129_2;
   assign m129_2 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_3 = W*in
   wire signed [14:0] m129_3;
   assign m129_3 =15'b0;

   // m129_4 = W*in
   wire signed [14:0] m129_4;
   assign m129_4 =15'b0;

   // m129_5 = W*in
   wire signed [14:0] m129_5;
   assign m129_5 =15'b0;

   // m129_6 = W*in
   wire signed [14:0] m129_6;
   assign m129_6 =15'b0;

   // m129_7 = W*in
   wire signed [14:0] m129_7;
   assign m129_7 =15'b0;

   // m129_8 = W*in
   wire signed [14:0] m129_8;
   assign m129_8 ={ {3{in129[14]}} , in129[14:3] };

   // m129_9 = W*in
   wire signed [14:0] m129_9;
   assign m129_9 =15'b0;

   // m129_10 = W*in
   wire signed [14:0] m129_10;
   assign m129_10 =15'b0;

   // m129_11 = W*in
   wire signed [14:0] m129_11;
   assign m129_11 =15'b0;

   // m129_12 = W*in
   wire signed [14:0] m129_12;
   assign m129_12 =15'b0;

   // m129_13 = W*in
   wire signed [14:0] m129_13;
   assign m129_13 =15'b0;

   // m129_14 = W*in
   wire signed [14:0] m129_14;
   assign m129_14 ={ {3{in129[14]}} , in129[14:3] };

   // m129_15 = W*in
   wire signed [14:0] m129_15;
   assign m129_15 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_16 = W*in
   wire signed [14:0] m129_16;
   assign m129_16 =15'b0;

   // m129_17 = W*in
   wire signed [14:0] m129_17;
   assign m129_17 =15'b0;

   // m129_18 = W*in
   wire signed [14:0] m129_18;
   assign m129_18 =15'b0;

   // m129_19 = W*in
   wire signed [14:0] m129_19;
   assign m129_19 =15'b0;

   // m129_20 = W*in
   wire signed [14:0] m129_20;
   assign m129_20 =15'b0;

   // m129_21 = W*in
   wire signed [14:0] m129_21;
   assign m129_21 ={ {3{in129[14]}} , in129[14:3] };

   // m129_22 = W*in
   wire signed [14:0] m129_22;
   assign m129_22 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_23 = W*in
   wire signed [14:0] m129_23;
   assign m129_23 =15'b0;

   // m129_24 = W*in
   wire signed [14:0] m129_24;
   assign m129_24 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_25 = W*in
   wire signed [14:0] m129_25;
   assign m129_25 ={ {3{in129[14]}} , in129[14:3] };

   // m129_26 = W*in
   wire signed [14:0] m129_26;
   assign m129_26 ={ {4{in129[14]}} , in129[14:4] };

   // m129_27 = W*in
   wire signed [14:0] m129_27;
   assign m129_27 ={ {4{neg129[14]}} , neg129[14:4] };

   // m129_28 = W*in
   wire signed [14:0] m129_28;
   assign m129_28 =15'b0;

   // m129_29 = W*in
   wire signed [14:0] m129_29;
   assign m129_29 ={ {3{in129[14]}} , in129[14:3] };

   // m129_30 = W*in
   wire signed [14:0] m129_30;
   assign m129_30 =15'b0;

   // m129_31 = W*in
   wire signed [14:0] m129_31;
   assign m129_31 ={ {3{in129[14]}} , in129[14:3] };

   // m129_32 = W*in
   wire signed [14:0] m129_32;
   assign m129_32 ={ {3{in129[14]}} , in129[14:3] };

   // m129_33 = W*in
   wire signed [14:0] m129_33;
   assign m129_33 ={ {4{neg129[14]}} , neg129[14:4] };

   // m129_34 = W*in
   wire signed [14:0] m129_34;
   assign m129_34 =15'b0;

   // m129_35 = W*in
   wire signed [14:0] m129_35;
   assign m129_35 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_36 = W*in
   wire signed [14:0] m129_36;
   assign m129_36 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_37 = W*in
   wire signed [14:0] m129_37;
   assign m129_37 ={ {3{in129[14]}} , in129[14:3] };

   // m129_38 = W*in
   wire signed [14:0] m129_38;
   assign m129_38 =15'b0;

   // m129_39 = W*in
   wire signed [14:0] m129_39;
   assign m129_39 =15'b0;

   // m129_40 = W*in
   wire signed [14:0] m129_40;
   assign m129_40 =15'b0;

   // m129_41 = W*in
   wire signed [14:0] m129_41;
   assign m129_41 =15'b0;

   // m129_42 = W*in
   wire signed [14:0] m129_42;
   assign m129_42 =15'b0;

   // m129_43 = W*in
   wire signed [14:0] m129_43;
   assign m129_43 =15'b0;

   // m129_44 = W*in
   wire signed [14:0] m129_44;
   assign m129_44 ={ {3{in129[14]}} , in129[14:3] };

   // m129_45 = W*in
   wire signed [14:0] m129_45;
   assign m129_45 =15'b0;

   // m129_46 = W*in
   wire signed [14:0] m129_46;
   assign m129_46 =15'b0;

   // m129_47 = W*in
   wire signed [14:0] m129_47;
   assign m129_47 =15'b0;

   // m129_48 = W*in
   wire signed [14:0] m129_48;
   assign m129_48 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_49 = W*in
   wire signed [14:0] m129_49;
   assign m129_49 =15'b0;

   // m129_50 = W*in
   wire signed [14:0] m129_50;
   assign m129_50 =15'b0;

   // m129_51 = W*in
   wire signed [14:0] m129_51;
   assign m129_51 =15'b0;

   // m129_52 = W*in
   wire signed [14:0] m129_52;
   assign m129_52 ={ {3{in129[14]}} , in129[14:3] };

   // m129_53 = W*in
   wire signed [14:0] m129_53;
   assign m129_53 =15'b0;

   // m129_54 = W*in
   wire signed [14:0] m129_54;
   assign m129_54 =15'b0;

   // m129_55 = W*in
   wire signed [14:0] m129_55;
   assign m129_55 =15'b0;

   // m129_56 = W*in
   wire signed [14:0] m129_56;
   assign m129_56 =15'b0;

   // m129_57 = W*in
   wire signed [14:0] m129_57;
   assign m129_57 =15'b0;

   // m129_58 = W*in
   wire signed [14:0] m129_58;
   assign m129_58 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_59 = W*in
   wire signed [14:0] m129_59;
   assign m129_59 =15'b0;

   // m129_60 = W*in
   wire signed [14:0] m129_60;
   assign m129_60 =15'b0;

   // m129_61 = W*in
   wire signed [14:0] m129_61;
   assign m129_61 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_62 = W*in
   wire signed [14:0] m129_62;
   assign m129_62 ={ {2{neg129[14]}} , neg129[14:2] };

   // m129_63 = W*in
   wire signed [14:0] m129_63;
   assign m129_63 =15'b0;

   // m129_64 = W*in
   wire signed [14:0] m129_64;
   assign m129_64 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_65 = W*in
   wire signed [14:0] m129_65;
   assign m129_65 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_66 = W*in
   wire signed [14:0] m129_66;
   assign m129_66 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_67 = W*in
   wire signed [14:0] m129_67;
   assign m129_67 =15'b0;

   // m129_68 = W*in
   wire signed [14:0] m129_68;
   assign m129_68 =15'b0;

   // m129_69 = W*in
   wire signed [14:0] m129_69;
   assign m129_69 ={ {3{in129[14]}} , in129[14:3] };

   // m129_70 = W*in
   wire signed [14:0] m129_70;
   assign m129_70 =15'b0;

   // m129_71 = W*in
   wire signed [14:0] m129_71;
   assign m129_71 =15'b0;

   // m129_72 = W*in
   wire signed [14:0] m129_72;
   assign m129_72 =15'b0;

   // m129_73 = W*in
   wire signed [14:0] m129_73;
   assign m129_73 =15'b0;

   // m129_74 = W*in
   wire signed [14:0] m129_74;
   assign m129_74 =15'b0;

   // m129_75 = W*in
   wire signed [14:0] m129_75;
   assign m129_75 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_76 = W*in
   wire signed [14:0] m129_76;
   assign m129_76 =15'b0;

   // m129_77 = W*in
   wire signed [14:0] m129_77;
   assign m129_77 =15'b0;

   // m129_78 = W*in
   wire signed [14:0] m129_78;
   assign m129_78 =15'b0;

   // m129_79 = W*in
   wire signed [14:0] m129_79;
   assign m129_79 =15'b0;

   // m129_80 = W*in
   wire signed [14:0] m129_80;
   assign m129_80 =15'b0;

   // m129_81 = W*in
   wire signed [14:0] m129_81;
   assign m129_81 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_82 = W*in
   wire signed [14:0] m129_82;
   assign m129_82 =15'b0;

   // m129_83 = W*in
   wire signed [14:0] m129_83;
   assign m129_83 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_84 = W*in
   wire signed [14:0] m129_84;
   assign m129_84 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_85 = W*in
   wire signed [14:0] m129_85;
   assign m129_85 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_86 = W*in
   wire signed [14:0] m129_86;
   assign m129_86 =15'b0;

   // m129_87 = W*in
   wire signed [14:0] m129_87;
   assign m129_87 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_88 = W*in
   wire signed [14:0] m129_88;
   assign m129_88 =15'b0;

   // m129_89 = W*in
   wire signed [14:0] m129_89;
   assign m129_89 =15'b0;

   // m129_90 = W*in
   wire signed [14:0] m129_90;
   assign m129_90 =15'b0;

   // m129_91 = W*in
   wire signed [14:0] m129_91;
   assign m129_91 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_92 = W*in
   wire signed [14:0] m129_92;
   assign m129_92 =15'b0;

   // m129_93 = W*in
   wire signed [14:0] m129_93;
   assign m129_93 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_94 = W*in
   wire signed [14:0] m129_94;
   assign m129_94 =15'b0;

   // m129_95 = W*in
   wire signed [14:0] m129_95;
   assign m129_95 =15'b0;

   // m129_96 = W*in
   wire signed [14:0] m129_96;
   assign m129_96 ={ {4{in129[14]}} , in129[14:4] };

   // m129_97 = W*in
   wire signed [14:0] m129_97;
   assign m129_97 ={ {3{neg129[14]}} , neg129[14:3] };

   // m129_98 = W*in
   wire signed [14:0] m129_98;
   assign m129_98 ={ {3{in129[14]}} , in129[14:3] };

   // m129_99 = W*in
   wire signed [14:0] m129_99;
   assign m129_99 =15'b0;

   // m129_100 = W*in
   wire signed [14:0] m129_100;
   assign m129_100 ={ {3{neg129[14]}} , neg129[14:3] };

   // m130_1 = W*in
   wire signed [14:0] m130_1;
   assign m130_1 =15'b0;

   // m130_2 = W*in
   wire signed [14:0] m130_2;
   assign m130_2 =15'b0;

   // m130_3 = W*in
   wire signed [14:0] m130_3;
   assign m130_3 =15'b0;

   // m130_4 = W*in
   wire signed [14:0] m130_4;
   assign m130_4 =15'b0;

   // m130_5 = W*in
   wire signed [14:0] m130_5;
   assign m130_5 ={ {3{neg130[14]}} , neg130[14:3] };

   // m130_6 = W*in
   wire signed [14:0] m130_6;
   assign m130_6 =15'b0;

   // m130_7 = W*in
   wire signed [14:0] m130_7;
   assign m130_7 =15'b0;

   // m130_8 = W*in
   wire signed [14:0] m130_8;
   assign m130_8 =15'b0;

   // m130_9 = W*in
   wire signed [14:0] m130_9;
   assign m130_9 =15'b0;

   // m130_10 = W*in
   wire signed [14:0] m130_10;
   assign m130_10 =15'b0;

   // m130_11 = W*in
   wire signed [14:0] m130_11;
   assign m130_11 =15'b0;

   // m130_12 = W*in
   wire signed [14:0] m130_12;
   assign m130_12 =15'b0;

   // m130_13 = W*in
   wire signed [14:0] m130_13;
   assign m130_13 =15'b0;

   // m130_14 = W*in
   wire signed [14:0] m130_14;
   assign m130_14 =15'b0;

   // m130_15 = W*in
   wire signed [14:0] m130_15;
   assign m130_15 =15'b0;

   // m130_16 = W*in
   wire signed [14:0] m130_16;
   assign m130_16 =15'b0;

   // m130_17 = W*in
   wire signed [14:0] m130_17;
   assign m130_17 =15'b0;

   // m130_18 = W*in
   wire signed [14:0] m130_18;
   assign m130_18 ={ {4{neg130[14]}} , neg130[14:4] };

   // m130_19 = W*in
   wire signed [14:0] m130_19;
   assign m130_19 =15'b0;

   // m130_20 = W*in
   wire signed [14:0] m130_20;
   assign m130_20 =15'b0;

   // m130_21 = W*in
   wire signed [14:0] m130_21;
   assign m130_21 =15'b0;

   // m130_22 = W*in
   wire signed [14:0] m130_22;
   assign m130_22 =15'b0;

   // m130_23 = W*in
   wire signed [14:0] m130_23;
   assign m130_23 =15'b0;

   // m130_24 = W*in
   wire signed [14:0] m130_24;
   assign m130_24 =15'b0;

   // m130_25 = W*in
   wire signed [14:0] m130_25;
   assign m130_25 =15'b0;

   // m130_26 = W*in
   wire signed [14:0] m130_26;
   assign m130_26 =15'b0;

   // m130_27 = W*in
   wire signed [14:0] m130_27;
   assign m130_27 =15'b0;

   // m130_28 = W*in
   wire signed [14:0] m130_28;
   assign m130_28 =15'b0;

   // m130_29 = W*in
   wire signed [14:0] m130_29;
   assign m130_29 ={ {4{neg130[14]}} , neg130[14:4] };

   // m130_30 = W*in
   wire signed [14:0] m130_30;
   assign m130_30 =15'b0;

   // m130_31 = W*in
   wire signed [14:0] m130_31;
   assign m130_31 ={ {3{neg130[14]}} , neg130[14:3] };

   // m130_32 = W*in
   wire signed [14:0] m130_32;
   assign m130_32 =15'b0;

   // m130_33 = W*in
   wire signed [14:0] m130_33;
   assign m130_33 =15'b0;

   // m130_34 = W*in
   wire signed [14:0] m130_34;
   assign m130_34 =15'b0;

   // m130_35 = W*in
   wire signed [14:0] m130_35;
   assign m130_35 ={ {3{neg130[14]}} , neg130[14:3] };

   // m130_36 = W*in
   wire signed [14:0] m130_36;
   assign m130_36 ={ {3{neg130[14]}} , neg130[14:3] };

   // m130_37 = W*in
   wire signed [14:0] m130_37;
   assign m130_37 =15'b0;

   // m130_38 = W*in
   wire signed [14:0] m130_38;
   assign m130_38 =15'b0;

   // m130_39 = W*in
   wire signed [14:0] m130_39;
   assign m130_39 =15'b0;

   // m130_40 = W*in
   wire signed [14:0] m130_40;
   assign m130_40 =15'b0;

   // m130_41 = W*in
   wire signed [14:0] m130_41;
   assign m130_41 =15'b0;

   // m130_42 = W*in
   wire signed [14:0] m130_42;
   assign m130_42 =15'b0;

   // m130_43 = W*in
   wire signed [14:0] m130_43;
   assign m130_43 =15'b0;

   // m130_44 = W*in
   wire signed [14:0] m130_44;
   assign m130_44 =15'b0;

   // m130_45 = W*in
   wire signed [14:0] m130_45;
   assign m130_45 =15'b0;

   // m130_46 = W*in
   wire signed [14:0] m130_46;
   assign m130_46 =15'b0;

   // m130_47 = W*in
   wire signed [14:0] m130_47;
   assign m130_47 =15'b0;

   // m130_48 = W*in
   wire signed [14:0] m130_48;
   assign m130_48 =15'b0;

   // m130_49 = W*in
   wire signed [14:0] m130_49;
   assign m130_49 =15'b0;

   // m130_50 = W*in
   wire signed [14:0] m130_50;
   assign m130_50 =15'b0;

   // m130_51 = W*in
   wire signed [14:0] m130_51;
   assign m130_51 =15'b0;

   // m130_52 = W*in
   wire signed [14:0] m130_52;
   assign m130_52 =15'b0;

   // m130_53 = W*in
   wire signed [14:0] m130_53;
   assign m130_53 =15'b0;

   // m130_54 = W*in
   wire signed [14:0] m130_54;
   assign m130_54 =15'b0;

   // m130_55 = W*in
   wire signed [14:0] m130_55;
   assign m130_55 =15'b0;

   // m130_56 = W*in
   wire signed [14:0] m130_56;
   assign m130_56 =15'b0;

   // m130_57 = W*in
   wire signed [14:0] m130_57;
   assign m130_57 =15'b0;

   // m130_58 = W*in
   wire signed [14:0] m130_58;
   assign m130_58 =15'b0;

   // m130_59 = W*in
   wire signed [14:0] m130_59;
   assign m130_59 =15'b0;

   // m130_60 = W*in
   wire signed [14:0] m130_60;
   assign m130_60 =15'b0;

   // m130_61 = W*in
   wire signed [14:0] m130_61;
   assign m130_61 =15'b0;

   // m130_62 = W*in
   wire signed [14:0] m130_62;
   assign m130_62 =15'b0;

   // m130_63 = W*in
   wire signed [14:0] m130_63;
   assign m130_63 =15'b0;

   // m130_64 = W*in
   wire signed [14:0] m130_64;
   assign m130_64 =15'b0;

   // m130_65 = W*in
   wire signed [14:0] m130_65;
   assign m130_65 =15'b0;

   // m130_66 = W*in
   wire signed [14:0] m130_66;
   assign m130_66 ={ {4{neg130[14]}} , neg130[14:4] };

   // m130_67 = W*in
   wire signed [14:0] m130_67;
   assign m130_67 =15'b0;

   // m130_68 = W*in
   wire signed [14:0] m130_68;
   assign m130_68 =15'b0;

   // m130_69 = W*in
   wire signed [14:0] m130_69;
   assign m130_69 ={ {3{neg130[14]}} , neg130[14:3] };

   // m130_70 = W*in
   wire signed [14:0] m130_70;
   assign m130_70 ={ {4{in130[14]}} , in130[14:4] };

   // m130_71 = W*in
   wire signed [14:0] m130_71;
   assign m130_71 =15'b0;

   // m130_72 = W*in
   wire signed [14:0] m130_72;
   assign m130_72 =15'b0;

   // m130_73 = W*in
   wire signed [14:0] m130_73;
   assign m130_73 =15'b0;

   // m130_74 = W*in
   wire signed [14:0] m130_74;
   assign m130_74 ={ {4{in130[14]}} , in130[14:4] };

   // m130_75 = W*in
   wire signed [14:0] m130_75;
   assign m130_75 ={ {4{in130[14]}} , in130[14:4] };

   // m130_76 = W*in
   wire signed [14:0] m130_76;
   assign m130_76 =15'b0;

   // m130_77 = W*in
   wire signed [14:0] m130_77;
   assign m130_77 =15'b0;

   // m130_78 = W*in
   wire signed [14:0] m130_78;
   assign m130_78 ={ {4{neg130[14]}} , neg130[14:4] };

   // m130_79 = W*in
   wire signed [14:0] m130_79;
   assign m130_79 =15'b0;

   // m130_80 = W*in
   wire signed [14:0] m130_80;
   assign m130_80 =15'b0;

   // m130_81 = W*in
   wire signed [14:0] m130_81;
   assign m130_81 ={ {3{in130[14]}} , in130[14:3] };

   // m130_82 = W*in
   wire signed [14:0] m130_82;
   assign m130_82 =15'b0;

   // m130_83 = W*in
   wire signed [14:0] m130_83;
   assign m130_83 =15'b0;

   // m130_84 = W*in
   wire signed [14:0] m130_84;
   assign m130_84 =15'b0;

   // m130_85 = W*in
   wire signed [14:0] m130_85;
   assign m130_85 =15'b0;

   // m130_86 = W*in
   wire signed [14:0] m130_86;
   assign m130_86 =15'b0;

   // m130_87 = W*in
   wire signed [14:0] m130_87;
   assign m130_87 =15'b0;

   // m130_88 = W*in
   wire signed [14:0] m130_88;
   assign m130_88 =15'b0;

   // m130_89 = W*in
   wire signed [14:0] m130_89;
   assign m130_89 =15'b0;

   // m130_90 = W*in
   wire signed [14:0] m130_90;
   assign m130_90 =15'b0;

   // m130_91 = W*in
   wire signed [14:0] m130_91;
   assign m130_91 =15'b0;

   // m130_92 = W*in
   wire signed [14:0] m130_92;
   assign m130_92 =15'b0;

   // m130_93 = W*in
   wire signed [14:0] m130_93;
   assign m130_93 =15'b0;

   // m130_94 = W*in
   wire signed [14:0] m130_94;
   assign m130_94 =15'b0;

   // m130_95 = W*in
   wire signed [14:0] m130_95;
   assign m130_95 =15'b0;

   // m130_96 = W*in
   wire signed [14:0] m130_96;
   assign m130_96 =15'b0;

   // m130_97 = W*in
   wire signed [14:0] m130_97;
   assign m130_97 =15'b0;

   // m130_98 = W*in
   wire signed [14:0] m130_98;
   assign m130_98 =15'b0;

   // m130_99 = W*in
   wire signed [14:0] m130_99;
   assign m130_99 ={ {3{in130[14]}} , in130[14:3] };

   // m130_100 = W*in
   wire signed [14:0] m130_100;
   assign m130_100 =15'b0;

   // m131_1 = W*in
   wire signed [14:0] m131_1;
   assign m131_1 =15'b0;

   // m131_2 = W*in
   wire signed [14:0] m131_2;
   assign m131_2 =15'b0;

   // m131_3 = W*in
   wire signed [14:0] m131_3;
   assign m131_3 =15'b0;

   // m131_4 = W*in
   wire signed [14:0] m131_4;
   assign m131_4 =15'b0;

   // m131_5 = W*in
   wire signed [14:0] m131_5;
   assign m131_5 =15'b0;

   // m131_6 = W*in
   wire signed [14:0] m131_6;
   assign m131_6 =15'b0;

   // m131_7 = W*in
   wire signed [14:0] m131_7;
   assign m131_7 =15'b0;

   // m131_8 = W*in
   wire signed [14:0] m131_8;
   assign m131_8 =15'b0;

   // m131_9 = W*in
   wire signed [14:0] m131_9;
   assign m131_9 =15'b0;

   // m131_10 = W*in
   wire signed [14:0] m131_10;
   assign m131_10 ={ {3{neg131[14]}} , neg131[14:3] };

   // m131_11 = W*in
   wire signed [14:0] m131_11;
   assign m131_11 =15'b0;

   // m131_12 = W*in
   wire signed [14:0] m131_12;
   assign m131_12 =15'b0;

   // m131_13 = W*in
   wire signed [14:0] m131_13;
   assign m131_13 =15'b0;

   // m131_14 = W*in
   wire signed [14:0] m131_14;
   assign m131_14 =15'b0;

   // m131_15 = W*in
   wire signed [14:0] m131_15;
   assign m131_15 ={ {4{in131[14]}} , in131[14:4] };

   // m131_16 = W*in
   wire signed [14:0] m131_16;
   assign m131_16 =15'b0;

   // m131_17 = W*in
   wire signed [14:0] m131_17;
   assign m131_17 =15'b0;

   // m131_18 = W*in
   wire signed [14:0] m131_18;
   assign m131_18 =15'b0;

   // m131_19 = W*in
   wire signed [14:0] m131_19;
   assign m131_19 ={ {3{in131[14]}} , in131[14:3] };

   // m131_20 = W*in
   wire signed [14:0] m131_20;
   assign m131_20 =15'b0;

   // m131_21 = W*in
   wire signed [14:0] m131_21;
   assign m131_21 =15'b0;

   // m131_22 = W*in
   wire signed [14:0] m131_22;
   assign m131_22 =15'b0;

   // m131_23 = W*in
   wire signed [14:0] m131_23;
   assign m131_23 =15'b0;

   // m131_24 = W*in
   wire signed [14:0] m131_24;
   assign m131_24 =15'b0;

   // m131_25 = W*in
   wire signed [14:0] m131_25;
   assign m131_25 =15'b0;

   // m131_26 = W*in
   wire signed [14:0] m131_26;
   assign m131_26 =15'b0;

   // m131_27 = W*in
   wire signed [14:0] m131_27;
   assign m131_27 =15'b0;

   // m131_28 = W*in
   wire signed [14:0] m131_28;
   assign m131_28 =15'b0;

   // m131_29 = W*in
   wire signed [14:0] m131_29;
   assign m131_29 =15'b0;

   // m131_30 = W*in
   wire signed [14:0] m131_30;
   assign m131_30 =15'b0;

   // m131_31 = W*in
   wire signed [14:0] m131_31;
   assign m131_31 =15'b0;

   // m131_32 = W*in
   wire signed [14:0] m131_32;
   assign m131_32 =15'b0;

   // m131_33 = W*in
   wire signed [14:0] m131_33;
   assign m131_33 ={ {4{in131[14]}} , in131[14:4] };

   // m131_34 = W*in
   wire signed [14:0] m131_34;
   assign m131_34 =15'b0;

   // m131_35 = W*in
   wire signed [14:0] m131_35;
   assign m131_35 =15'b0;

   // m131_36 = W*in
   wire signed [14:0] m131_36;
   assign m131_36 =15'b0;

   // m131_37 = W*in
   wire signed [14:0] m131_37;
   assign m131_37 =15'b0;

   // m131_38 = W*in
   wire signed [14:0] m131_38;
   assign m131_38 =15'b0;

   // m131_39 = W*in
   wire signed [14:0] m131_39;
   assign m131_39 ={ {3{in131[14]}} , in131[14:3] };

   // m131_40 = W*in
   wire signed [14:0] m131_40;
   assign m131_40 =15'b0;

   // m131_41 = W*in
   wire signed [14:0] m131_41;
   assign m131_41 =15'b0;

   // m131_42 = W*in
   wire signed [14:0] m131_42;
   assign m131_42 =15'b0;

   // m131_43 = W*in
   wire signed [14:0] m131_43;
   assign m131_43 =15'b0;

   // m131_44 = W*in
   wire signed [14:0] m131_44;
   assign m131_44 =15'b0;

   // m131_45 = W*in
   wire signed [14:0] m131_45;
   assign m131_45 =15'b0;

   // m131_46 = W*in
   wire signed [14:0] m131_46;
   assign m131_46 =15'b0;

   // m131_47 = W*in
   wire signed [14:0] m131_47;
   assign m131_47 =15'b0;

   // m131_48 = W*in
   wire signed [14:0] m131_48;
   assign m131_48 =15'b0;

   // m131_49 = W*in
   wire signed [14:0] m131_49;
   assign m131_49 =15'b0;

   // m131_50 = W*in
   wire signed [14:0] m131_50;
   assign m131_50 =15'b0;

   // m131_51 = W*in
   wire signed [14:0] m131_51;
   assign m131_51 =15'b0;

   // m131_52 = W*in
   wire signed [14:0] m131_52;
   assign m131_52 =15'b0;

   // m131_53 = W*in
   wire signed [14:0] m131_53;
   assign m131_53 =15'b0;

   // m131_54 = W*in
   wire signed [14:0] m131_54;
   assign m131_54 =15'b0;

   // m131_55 = W*in
   wire signed [14:0] m131_55;
   assign m131_55 =15'b0;

   // m131_56 = W*in
   wire signed [14:0] m131_56;
   assign m131_56 =15'b0;

   // m131_57 = W*in
   wire signed [14:0] m131_57;
   assign m131_57 =15'b0;

   // m131_58 = W*in
   wire signed [14:0] m131_58;
   assign m131_58 =15'b0;

   // m131_59 = W*in
   wire signed [14:0] m131_59;
   assign m131_59 =15'b0;

   // m131_60 = W*in
   wire signed [14:0] m131_60;
   assign m131_60 =15'b0;

   // m131_61 = W*in
   wire signed [14:0] m131_61;
   assign m131_61 =15'b0;

   // m131_62 = W*in
   wire signed [14:0] m131_62;
   assign m131_62 =15'b0;

   // m131_63 = W*in
   wire signed [14:0] m131_63;
   assign m131_63 ={ {4{in131[14]}} , in131[14:4] };

   // m131_64 = W*in
   wire signed [14:0] m131_64;
   assign m131_64 =15'b0;

   // m131_65 = W*in
   wire signed [14:0] m131_65;
   assign m131_65 =15'b0;

   // m131_66 = W*in
   wire signed [14:0] m131_66;
   assign m131_66 ={ {2{in131[14]}} , in131[14:2] };

   // m131_67 = W*in
   wire signed [14:0] m131_67;
   assign m131_67 =15'b0;

   // m131_68 = W*in
   wire signed [14:0] m131_68;
   assign m131_68 =15'b0;

   // m131_69 = W*in
   wire signed [14:0] m131_69;
   assign m131_69 =15'b0;

   // m131_70 = W*in
   wire signed [14:0] m131_70;
   assign m131_70 =15'b0;

   // m131_71 = W*in
   wire signed [14:0] m131_71;
   assign m131_71 ={ {4{in131[14]}} , in131[14:4] };

   // m131_72 = W*in
   wire signed [14:0] m131_72;
   assign m131_72 =15'b0;

   // m131_73 = W*in
   wire signed [14:0] m131_73;
   assign m131_73 =15'b0;

   // m131_74 = W*in
   wire signed [14:0] m131_74;
   assign m131_74 ={ {3{neg131[14]}} , neg131[14:3] };

   // m131_75 = W*in
   wire signed [14:0] m131_75;
   assign m131_75 =15'b0;

   // m131_76 = W*in
   wire signed [14:0] m131_76;
   assign m131_76 =15'b0;

   // m131_77 = W*in
   wire signed [14:0] m131_77;
   assign m131_77 =15'b0;

   // m131_78 = W*in
   wire signed [14:0] m131_78;
   assign m131_78 =15'b0;

   // m131_79 = W*in
   wire signed [14:0] m131_79;
   assign m131_79 =15'b0;

   // m131_80 = W*in
   wire signed [14:0] m131_80;
   assign m131_80 =15'b0;

   // m131_81 = W*in
   wire signed [14:0] m131_81;
   assign m131_81 =15'b0;

   // m131_82 = W*in
   wire signed [14:0] m131_82;
   assign m131_82 =15'b0;

   // m131_83 = W*in
   wire signed [14:0] m131_83;
   assign m131_83 =15'b0;

   // m131_84 = W*in
   wire signed [14:0] m131_84;
   assign m131_84 =15'b0;

   // m131_85 = W*in
   wire signed [14:0] m131_85;
   assign m131_85 =15'b0;

   // m131_86 = W*in
   wire signed [14:0] m131_86;
   assign m131_86 =15'b0;

   // m131_87 = W*in
   wire signed [14:0] m131_87;
   assign m131_87 =15'b0;

   // m131_88 = W*in
   wire signed [14:0] m131_88;
   assign m131_88 =15'b0;

   // m131_89 = W*in
   wire signed [14:0] m131_89;
   assign m131_89 =15'b0;

   // m131_90 = W*in
   wire signed [14:0] m131_90;
   assign m131_90 =15'b0;

   // m131_91 = W*in
   wire signed [14:0] m131_91;
   assign m131_91 =15'b0;

   // m131_92 = W*in
   wire signed [14:0] m131_92;
   assign m131_92 =15'b0;

   // m131_93 = W*in
   wire signed [14:0] m131_93;
   assign m131_93 =15'b0;

   // m131_94 = W*in
   wire signed [14:0] m131_94;
   assign m131_94 =15'b0;

   // m131_95 = W*in
   wire signed [14:0] m131_95;
   assign m131_95 =15'b0;

   // m131_96 = W*in
   wire signed [14:0] m131_96;
   assign m131_96 =15'b0;

   // m131_97 = W*in
   wire signed [14:0] m131_97;
   assign m131_97 =15'b0;

   // m131_98 = W*in
   wire signed [14:0] m131_98;
   assign m131_98 ={ {3{in131[14]}} , in131[14:3] };

   // m131_99 = W*in
   wire signed [14:0] m131_99;
   assign m131_99 =15'b0;

   // m131_100 = W*in
   wire signed [14:0] m131_100;
   assign m131_100 =15'b0;

   // m132_1 = W*in
   wire signed [14:0] m132_1;
   assign m132_1 =15'b0;

   // m132_2 = W*in
   wire signed [14:0] m132_2;
   assign m132_2 =15'b0;

   // m132_3 = W*in
   wire signed [14:0] m132_3;
   assign m132_3 ={ {4{neg132[14]}} , neg132[14:4] };

   // m132_4 = W*in
   wire signed [14:0] m132_4;
   assign m132_4 =15'b0;

   // m132_5 = W*in
   wire signed [14:0] m132_5;
   assign m132_5 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_6 = W*in
   wire signed [14:0] m132_6;
   assign m132_6 =15'b0;

   // m132_7 = W*in
   wire signed [14:0] m132_7;
   assign m132_7 ={ {3{in132[14]}} , in132[14:3] };

   // m132_8 = W*in
   wire signed [14:0] m132_8;
   assign m132_8 =15'b0;

   // m132_9 = W*in
   wire signed [14:0] m132_9;
   assign m132_9 =15'b0;

   // m132_10 = W*in
   wire signed [14:0] m132_10;
   assign m132_10 =15'b0;

   // m132_11 = W*in
   wire signed [14:0] m132_11;
   assign m132_11 =15'b0;

   // m132_12 = W*in
   wire signed [14:0] m132_12;
   assign m132_12 =15'b0;

   // m132_13 = W*in
   wire signed [14:0] m132_13;
   assign m132_13 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_14 = W*in
   wire signed [14:0] m132_14;
   assign m132_14 =15'b0;

   // m132_15 = W*in
   wire signed [14:0] m132_15;
   assign m132_15 =15'b0;

   // m132_16 = W*in
   wire signed [14:0] m132_16;
   assign m132_16 =15'b0;

   // m132_17 = W*in
   wire signed [14:0] m132_17;
   assign m132_17 =15'b0;

   // m132_18 = W*in
   wire signed [14:0] m132_18;
   assign m132_18 =15'b0;

   // m132_19 = W*in
   wire signed [14:0] m132_19;
   assign m132_19 =15'b0;

   // m132_20 = W*in
   wire signed [14:0] m132_20;
   assign m132_20 =15'b0;

   // m132_21 = W*in
   wire signed [14:0] m132_21;
   assign m132_21 ={ {3{in132[14]}} , in132[14:3] };

   // m132_22 = W*in
   wire signed [14:0] m132_22;
   assign m132_22 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_23 = W*in
   wire signed [14:0] m132_23;
   assign m132_23 =15'b0;

   // m132_24 = W*in
   wire signed [14:0] m132_24;
   assign m132_24 =15'b0;

   // m132_25 = W*in
   wire signed [14:0] m132_25;
   assign m132_25 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_26 = W*in
   wire signed [14:0] m132_26;
   assign m132_26 =15'b0;

   // m132_27 = W*in
   wire signed [14:0] m132_27;
   assign m132_27 =15'b0;

   // m132_28 = W*in
   wire signed [14:0] m132_28;
   assign m132_28 =15'b0;

   // m132_29 = W*in
   wire signed [14:0] m132_29;
   assign m132_29 =15'b0;

   // m132_30 = W*in
   wire signed [14:0] m132_30;
   assign m132_30 ={ {3{in132[14]}} , in132[14:3] };

   // m132_31 = W*in
   wire signed [14:0] m132_31;
   assign m132_31 =15'b0;

   // m132_32 = W*in
   wire signed [14:0] m132_32;
   assign m132_32 =15'b0;

   // m132_33 = W*in
   wire signed [14:0] m132_33;
   assign m132_33 =15'b0;

   // m132_34 = W*in
   wire signed [14:0] m132_34;
   assign m132_34 =15'b0;

   // m132_35 = W*in
   wire signed [14:0] m132_35;
   assign m132_35 =15'b0;

   // m132_36 = W*in
   wire signed [14:0] m132_36;
   assign m132_36 =15'b0;

   // m132_37 = W*in
   wire signed [14:0] m132_37;
   assign m132_37 =15'b0;

   // m132_38 = W*in
   wire signed [14:0] m132_38;
   assign m132_38 =15'b0;

   // m132_39 = W*in
   wire signed [14:0] m132_39;
   assign m132_39 =15'b0;

   // m132_40 = W*in
   wire signed [14:0] m132_40;
   assign m132_40 =15'b0;

   // m132_41 = W*in
   wire signed [14:0] m132_41;
   assign m132_41 =15'b0;

   // m132_42 = W*in
   wire signed [14:0] m132_42;
   assign m132_42 =15'b0;

   // m132_43 = W*in
   wire signed [14:0] m132_43;
   assign m132_43 =15'b0;

   // m132_44 = W*in
   wire signed [14:0] m132_44;
   assign m132_44 ={ {3{in132[14]}} , in132[14:3] };

   // m132_45 = W*in
   wire signed [14:0] m132_45;
   assign m132_45 =15'b0;

   // m132_46 = W*in
   wire signed [14:0] m132_46;
   assign m132_46 =15'b0;

   // m132_47 = W*in
   wire signed [14:0] m132_47;
   assign m132_47 =15'b0;

   // m132_48 = W*in
   wire signed [14:0] m132_48;
   assign m132_48 =15'b0;

   // m132_49 = W*in
   wire signed [14:0] m132_49;
   assign m132_49 =15'b0;

   // m132_50 = W*in
   wire signed [14:0] m132_50;
   assign m132_50 =15'b0;

   // m132_51 = W*in
   wire signed [14:0] m132_51;
   assign m132_51 =15'b0;

   // m132_52 = W*in
   wire signed [14:0] m132_52;
   assign m132_52 =15'b0;

   // m132_53 = W*in
   wire signed [14:0] m132_53;
   assign m132_53 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_54 = W*in
   wire signed [14:0] m132_54;
   assign m132_54 =15'b0;

   // m132_55 = W*in
   wire signed [14:0] m132_55;
   assign m132_55 =15'b0;

   // m132_56 = W*in
   wire signed [14:0] m132_56;
   assign m132_56 =15'b0;

   // m132_57 = W*in
   wire signed [14:0] m132_57;
   assign m132_57 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_58 = W*in
   wire signed [14:0] m132_58;
   assign m132_58 =15'b0;

   // m132_59 = W*in
   wire signed [14:0] m132_59;
   assign m132_59 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_60 = W*in
   wire signed [14:0] m132_60;
   assign m132_60 =15'b0;

   // m132_61 = W*in
   wire signed [14:0] m132_61;
   assign m132_61 ={ {4{neg132[14]}} , neg132[14:4] };

   // m132_62 = W*in
   wire signed [14:0] m132_62;
   assign m132_62 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_63 = W*in
   wire signed [14:0] m132_63;
   assign m132_63 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_64 = W*in
   wire signed [14:0] m132_64;
   assign m132_64 ={ {4{neg132[14]}} , neg132[14:4] };

   // m132_65 = W*in
   wire signed [14:0] m132_65;
   assign m132_65 =15'b0;

   // m132_66 = W*in
   wire signed [14:0] m132_66;
   assign m132_66 =15'b0;

   // m132_67 = W*in
   wire signed [14:0] m132_67;
   assign m132_67 =15'b0;

   // m132_68 = W*in
   wire signed [14:0] m132_68;
   assign m132_68 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_69 = W*in
   wire signed [14:0] m132_69;
   assign m132_69 =15'b0;

   // m132_70 = W*in
   wire signed [14:0] m132_70;
   assign m132_70 =15'b0;

   // m132_71 = W*in
   wire signed [14:0] m132_71;
   assign m132_71 =15'b0;

   // m132_72 = W*in
   wire signed [14:0] m132_72;
   assign m132_72 =15'b0;

   // m132_73 = W*in
   wire signed [14:0] m132_73;
   assign m132_73 =15'b0;

   // m132_74 = W*in
   wire signed [14:0] m132_74;
   assign m132_74 ={ {4{neg132[14]}} , neg132[14:4] };

   // m132_75 = W*in
   wire signed [14:0] m132_75;
   assign m132_75 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_76 = W*in
   wire signed [14:0] m132_76;
   assign m132_76 =15'b0;

   // m132_77 = W*in
   wire signed [14:0] m132_77;
   assign m132_77 =15'b0;

   // m132_78 = W*in
   wire signed [14:0] m132_78;
   assign m132_78 =15'b0;

   // m132_79 = W*in
   wire signed [14:0] m132_79;
   assign m132_79 =15'b0;

   // m132_80 = W*in
   wire signed [14:0] m132_80;
   assign m132_80 =15'b0;

   // m132_81 = W*in
   wire signed [14:0] m132_81;
   assign m132_81 =15'b0;

   // m132_82 = W*in
   wire signed [14:0] m132_82;
   assign m132_82 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_83 = W*in
   wire signed [14:0] m132_83;
   assign m132_83 =15'b0;

   // m132_84 = W*in
   wire signed [14:0] m132_84;
   assign m132_84 =15'b0;

   // m132_85 = W*in
   wire signed [14:0] m132_85;
   assign m132_85 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_86 = W*in
   wire signed [14:0] m132_86;
   assign m132_86 =15'b0;

   // m132_87 = W*in
   wire signed [14:0] m132_87;
   assign m132_87 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_88 = W*in
   wire signed [14:0] m132_88;
   assign m132_88 =15'b0;

   // m132_89 = W*in
   wire signed [14:0] m132_89;
   assign m132_89 =15'b0;

   // m132_90 = W*in
   wire signed [14:0] m132_90;
   assign m132_90 ={ {3{in132[14]}} , in132[14:3] };

   // m132_91 = W*in
   wire signed [14:0] m132_91;
   assign m132_91 =15'b0;

   // m132_92 = W*in
   wire signed [14:0] m132_92;
   assign m132_92 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_93 = W*in
   wire signed [14:0] m132_93;
   assign m132_93 =15'b0;

   // m132_94 = W*in
   wire signed [14:0] m132_94;
   assign m132_94 =15'b0;

   // m132_95 = W*in
   wire signed [14:0] m132_95;
   assign m132_95 =15'b0;

   // m132_96 = W*in
   wire signed [14:0] m132_96;
   assign m132_96 ={ {4{in132[14]}} , in132[14:4] };

   // m132_97 = W*in
   wire signed [14:0] m132_97;
   assign m132_97 =15'b0;

   // m132_98 = W*in
   wire signed [14:0] m132_98;
   assign m132_98 ={ {3{in132[14]}} , in132[14:3] };

   // m132_99 = W*in
   wire signed [14:0] m132_99;
   assign m132_99 ={ {3{neg132[14]}} , neg132[14:3] };

   // m132_100 = W*in
   wire signed [14:0] m132_100;
   assign m132_100 ={ {3{neg132[14]}} , neg132[14:3] };

   // m133_1 = W*in
   wire signed [14:0] m133_1;
   assign m133_1 ={ {3{in133[14]}} , in133[14:3] };

   // m133_2 = W*in
   wire signed [14:0] m133_2;
   assign m133_2 ={ {3{in133[14]}} , in133[14:3] };

   // m133_3 = W*in
   wire signed [14:0] m133_3;
   assign m133_3 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_4 = W*in
   wire signed [14:0] m133_4;
   assign m133_4 =15'b0;

   // m133_5 = W*in
   wire signed [14:0] m133_5;
   assign m133_5 =15'b0;

   // m133_6 = W*in
   wire signed [14:0] m133_6;
   assign m133_6 =15'b0;

   // m133_7 = W*in
   wire signed [14:0] m133_7;
   assign m133_7 =15'b0;

   // m133_8 = W*in
   wire signed [14:0] m133_8;
   assign m133_8 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_9 = W*in
   wire signed [14:0] m133_9;
   assign m133_9 =15'b0;

   // m133_10 = W*in
   wire signed [14:0] m133_10;
   assign m133_10 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_11 = W*in
   wire signed [14:0] m133_11;
   assign m133_11 =15'b0;

   // m133_12 = W*in
   wire signed [14:0] m133_12;
   assign m133_12 =15'b0;

   // m133_13 = W*in
   wire signed [14:0] m133_13;
   assign m133_13 =15'b0;

   // m133_14 = W*in
   wire signed [14:0] m133_14;
   assign m133_14 =15'b0;

   // m133_15 = W*in
   wire signed [14:0] m133_15;
   assign m133_15 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_16 = W*in
   wire signed [14:0] m133_16;
   assign m133_16 =15'b0;

   // m133_17 = W*in
   wire signed [14:0] m133_17;
   assign m133_17 =15'b0;

   // m133_18 = W*in
   wire signed [14:0] m133_18;
   assign m133_18 ={ {4{in133[14]}} , in133[14:4] };

   // m133_19 = W*in
   wire signed [14:0] m133_19;
   assign m133_19 =15'b0;

   // m133_20 = W*in
   wire signed [14:0] m133_20;
   assign m133_20 =15'b0;

   // m133_21 = W*in
   wire signed [14:0] m133_21;
   assign m133_21 =15'b0;

   // m133_22 = W*in
   wire signed [14:0] m133_22;
   assign m133_22 =15'b0;

   // m133_23 = W*in
   wire signed [14:0] m133_23;
   assign m133_23 ={ {3{in133[14]}} , in133[14:3] };

   // m133_24 = W*in
   wire signed [14:0] m133_24;
   assign m133_24 =15'b0;

   // m133_25 = W*in
   wire signed [14:0] m133_25;
   assign m133_25 =15'b0;

   // m133_26 = W*in
   wire signed [14:0] m133_26;
   assign m133_26 =15'b0;

   // m133_27 = W*in
   wire signed [14:0] m133_27;
   assign m133_27 =15'b0;

   // m133_28 = W*in
   wire signed [14:0] m133_28;
   assign m133_28 ={ {4{in133[14]}} , in133[14:4] };

   // m133_29 = W*in
   wire signed [14:0] m133_29;
   assign m133_29 ={ {3{in133[14]}} , in133[14:3] };

   // m133_30 = W*in
   wire signed [14:0] m133_30;
   assign m133_30 =15'b0;

   // m133_31 = W*in
   wire signed [14:0] m133_31;
   assign m133_31 =15'b0;

   // m133_32 = W*in
   wire signed [14:0] m133_32;
   assign m133_32 ={ {3{in133[14]}} , in133[14:3] };

   // m133_33 = W*in
   wire signed [14:0] m133_33;
   assign m133_33 ={ {3{in133[14]}} , in133[14:3] };

   // m133_34 = W*in
   wire signed [14:0] m133_34;
   assign m133_34 =15'b0;

   // m133_35 = W*in
   wire signed [14:0] m133_35;
   assign m133_35 ={ {3{in133[14]}} , in133[14:3] };

   // m133_36 = W*in
   wire signed [14:0] m133_36;
   assign m133_36 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_37 = W*in
   wire signed [14:0] m133_37;
   assign m133_37 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_38 = W*in
   wire signed [14:0] m133_38;
   assign m133_38 ={ {3{in133[14]}} , in133[14:3] };

   // m133_39 = W*in
   wire signed [14:0] m133_39;
   assign m133_39 =15'b0;

   // m133_40 = W*in
   wire signed [14:0] m133_40;
   assign m133_40 =15'b0;

   // m133_41 = W*in
   wire signed [14:0] m133_41;
   assign m133_41 =15'b0;

   // m133_42 = W*in
   wire signed [14:0] m133_42;
   assign m133_42 =15'b0;

   // m133_43 = W*in
   wire signed [14:0] m133_43;
   assign m133_43 =15'b0;

   // m133_44 = W*in
   wire signed [14:0] m133_44;
   assign m133_44 =15'b0;

   // m133_45 = W*in
   wire signed [14:0] m133_45;
   assign m133_45 =15'b0;

   // m133_46 = W*in
   wire signed [14:0] m133_46;
   assign m133_46 ={ {4{neg133[14]}} , neg133[14:4] };

   // m133_47 = W*in
   wire signed [14:0] m133_47;
   assign m133_47 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_48 = W*in
   wire signed [14:0] m133_48;
   assign m133_48 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_49 = W*in
   wire signed [14:0] m133_49;
   assign m133_49 =15'b0;

   // m133_50 = W*in
   wire signed [14:0] m133_50;
   assign m133_50 =15'b0;

   // m133_51 = W*in
   wire signed [14:0] m133_51;
   assign m133_51 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_52 = W*in
   wire signed [14:0] m133_52;
   assign m133_52 =15'b0;

   // m133_53 = W*in
   wire signed [14:0] m133_53;
   assign m133_53 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_54 = W*in
   wire signed [14:0] m133_54;
   assign m133_54 =15'b0;

   // m133_55 = W*in
   wire signed [14:0] m133_55;
   assign m133_55 =15'b0;

   // m133_56 = W*in
   wire signed [14:0] m133_56;
   assign m133_56 =15'b0;

   // m133_57 = W*in
   wire signed [14:0] m133_57;
   assign m133_57 =15'b0;

   // m133_58 = W*in
   wire signed [14:0] m133_58;
   assign m133_58 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_59 = W*in
   wire signed [14:0] m133_59;
   assign m133_59 =15'b0;

   // m133_60 = W*in
   wire signed [14:0] m133_60;
   assign m133_60 =15'b0;

   // m133_61 = W*in
   wire signed [14:0] m133_61;
   assign m133_61 ={ {4{neg133[14]}} , neg133[14:4] };

   // m133_62 = W*in
   wire signed [14:0] m133_62;
   assign m133_62 =15'b0;

   // m133_63 = W*in
   wire signed [14:0] m133_63;
   assign m133_63 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_64 = W*in
   wire signed [14:0] m133_64;
   assign m133_64 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_65 = W*in
   wire signed [14:0] m133_65;
   assign m133_65 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_66 = W*in
   wire signed [14:0] m133_66;
   assign m133_66 ={ {4{neg133[14]}} , neg133[14:4] };

   // m133_67 = W*in
   wire signed [14:0] m133_67;
   assign m133_67 ={ {4{neg133[14]}} , neg133[14:4] };

   // m133_68 = W*in
   wire signed [14:0] m133_68;
   assign m133_68 =15'b0;

   // m133_69 = W*in
   wire signed [14:0] m133_69;
   assign m133_69 =15'b0;

   // m133_70 = W*in
   wire signed [14:0] m133_70;
   assign m133_70 =15'b0;

   // m133_71 = W*in
   wire signed [14:0] m133_71;
   assign m133_71 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_72 = W*in
   wire signed [14:0] m133_72;
   assign m133_72 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_73 = W*in
   wire signed [14:0] m133_73;
   assign m133_73 =15'b0;

   // m133_74 = W*in
   wire signed [14:0] m133_74;
   assign m133_74 ={ {4{in133[14]}} , in133[14:4] };

   // m133_75 = W*in
   wire signed [14:0] m133_75;
   assign m133_75 ={ {3{in133[14]}} , in133[14:3] };

   // m133_76 = W*in
   wire signed [14:0] m133_76;
   assign m133_76 =15'b0;

   // m133_77 = W*in
   wire signed [14:0] m133_77;
   assign m133_77 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_78 = W*in
   wire signed [14:0] m133_78;
   assign m133_78 =15'b0;

   // m133_79 = W*in
   wire signed [14:0] m133_79;
   assign m133_79 =15'b0;

   // m133_80 = W*in
   wire signed [14:0] m133_80;
   assign m133_80 =15'b0;

   // m133_81 = W*in
   wire signed [14:0] m133_81;
   assign m133_81 =15'b0;

   // m133_82 = W*in
   wire signed [14:0] m133_82;
   assign m133_82 =15'b0;

   // m133_83 = W*in
   wire signed [14:0] m133_83;
   assign m133_83 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_84 = W*in
   wire signed [14:0] m133_84;
   assign m133_84 =15'b0;

   // m133_85 = W*in
   wire signed [14:0] m133_85;
   assign m133_85 =15'b0;

   // m133_86 = W*in
   wire signed [14:0] m133_86;
   assign m133_86 =15'b0;

   // m133_87 = W*in
   wire signed [14:0] m133_87;
   assign m133_87 =15'b0;

   // m133_88 = W*in
   wire signed [14:0] m133_88;
   assign m133_88 =15'b0;

   // m133_89 = W*in
   wire signed [14:0] m133_89;
   assign m133_89 ={ {2{neg133[14]}} , neg133[14:2] };

   // m133_90 = W*in
   wire signed [14:0] m133_90;
   assign m133_90 ={ {2{in133[14]}} , in133[14:2] };

   // m133_91 = W*in
   wire signed [14:0] m133_91;
   assign m133_91 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_92 = W*in
   wire signed [14:0] m133_92;
   assign m133_92 =15'b0;

   // m133_93 = W*in
   wire signed [14:0] m133_93;
   assign m133_93 ={ {3{neg133[14]}} , neg133[14:3] };

   // m133_94 = W*in
   wire signed [14:0] m133_94;
   assign m133_94 =15'b0;

   // m133_95 = W*in
   wire signed [14:0] m133_95;
   assign m133_95 =15'b0;

   // m133_96 = W*in
   wire signed [14:0] m133_96;
   assign m133_96 =15'b0;

   // m133_97 = W*in
   wire signed [14:0] m133_97;
   assign m133_97 ={ {3{in133[14]}} , in133[14:3] };

   // m133_98 = W*in
   wire signed [14:0] m133_98;
   assign m133_98 =15'b0;

   // m133_99 = W*in
   wire signed [14:0] m133_99;
   assign m133_99 =15'b0;

   // m133_100 = W*in
   wire signed [14:0] m133_100;
   assign m133_100 =15'b0;

   // m134_1 = W*in
   wire signed [14:0] m134_1;
   assign m134_1 =15'b0;

   // m134_2 = W*in
   wire signed [14:0] m134_2;
   assign m134_2 =15'b0;

   // m134_3 = W*in
   wire signed [14:0] m134_3;
   assign m134_3 =15'b0;

   // m134_4 = W*in
   wire signed [14:0] m134_4;
   assign m134_4 =15'b0;

   // m134_5 = W*in
   wire signed [14:0] m134_5;
   assign m134_5 =15'b0;

   // m134_6 = W*in
   wire signed [14:0] m134_6;
   assign m134_6 =15'b0;

   // m134_7 = W*in
   wire signed [14:0] m134_7;
   assign m134_7 =15'b0;

   // m134_8 = W*in
   wire signed [14:0] m134_8;
   assign m134_8 =15'b0;

   // m134_9 = W*in
   wire signed [14:0] m134_9;
   assign m134_9 =15'b0;

   // m134_10 = W*in
   wire signed [14:0] m134_10;
   assign m134_10 =15'b0;

   // m134_11 = W*in
   wire signed [14:0] m134_11;
   assign m134_11 =15'b0;

   // m134_12 = W*in
   wire signed [14:0] m134_12;
   assign m134_12 =15'b0;

   // m134_13 = W*in
   wire signed [14:0] m134_13;
   assign m134_13 =15'b0;

   // m134_14 = W*in
   wire signed [14:0] m134_14;
   assign m134_14 ={ {3{neg134[14]}} , neg134[14:3] };

   // m134_15 = W*in
   wire signed [14:0] m134_15;
   assign m134_15 ={ {4{in134[14]}} , in134[14:4] };

   // m134_16 = W*in
   wire signed [14:0] m134_16;
   assign m134_16 =15'b0;

   // m134_17 = W*in
   wire signed [14:0] m134_17;
   assign m134_17 =15'b0;

   // m134_18 = W*in
   wire signed [14:0] m134_18;
   assign m134_18 =15'b0;

   // m134_19 = W*in
   wire signed [14:0] m134_19;
   assign m134_19 =15'b0;

   // m134_20 = W*in
   wire signed [14:0] m134_20;
   assign m134_20 =15'b0;

   // m134_21 = W*in
   wire signed [14:0] m134_21;
   assign m134_21 =15'b0;

   // m134_22 = W*in
   wire signed [14:0] m134_22;
   assign m134_22 =15'b0;

   // m134_23 = W*in
   wire signed [14:0] m134_23;
   assign m134_23 =15'b0;

   // m134_24 = W*in
   wire signed [14:0] m134_24;
   assign m134_24 =15'b0;

   // m134_25 = W*in
   wire signed [14:0] m134_25;
   assign m134_25 =15'b0;

   // m134_26 = W*in
   wire signed [14:0] m134_26;
   assign m134_26 =15'b0;

   // m134_27 = W*in
   wire signed [14:0] m134_27;
   assign m134_27 ={ {3{in134[14]}} , in134[14:3] };

   // m134_28 = W*in
   wire signed [14:0] m134_28;
   assign m134_28 =15'b0;

   // m134_29 = W*in
   wire signed [14:0] m134_29;
   assign m134_29 =15'b0;

   // m134_30 = W*in
   wire signed [14:0] m134_30;
   assign m134_30 =15'b0;

   // m134_31 = W*in
   wire signed [14:0] m134_31;
   assign m134_31 =15'b0;

   // m134_32 = W*in
   wire signed [14:0] m134_32;
   assign m134_32 ={ {4{neg134[14]}} , neg134[14:4] };

   // m134_33 = W*in
   wire signed [14:0] m134_33;
   assign m134_33 ={ {4{neg134[14]}} , neg134[14:4] };

   // m134_34 = W*in
   wire signed [14:0] m134_34;
   assign m134_34 =15'b0;

   // m134_35 = W*in
   wire signed [14:0] m134_35;
   assign m134_35 =15'b0;

   // m134_36 = W*in
   wire signed [14:0] m134_36;
   assign m134_36 =15'b0;

   // m134_37 = W*in
   wire signed [14:0] m134_37;
   assign m134_37 ={ {3{neg134[14]}} , neg134[14:3] };

   // m134_38 = W*in
   wire signed [14:0] m134_38;
   assign m134_38 =15'b0;

   // m134_39 = W*in
   wire signed [14:0] m134_39;
   assign m134_39 =15'b0;

   // m134_40 = W*in
   wire signed [14:0] m134_40;
   assign m134_40 ={ {4{in134[14]}} , in134[14:4] };

   // m134_41 = W*in
   wire signed [14:0] m134_41;
   assign m134_41 =15'b0;

   // m134_42 = W*in
   wire signed [14:0] m134_42;
   assign m134_42 =15'b0;

   // m134_43 = W*in
   wire signed [14:0] m134_43;
   assign m134_43 =15'b0;

   // m134_44 = W*in
   wire signed [14:0] m134_44;
   assign m134_44 =15'b0;

   // m134_45 = W*in
   wire signed [14:0] m134_45;
   assign m134_45 =15'b0;

   // m134_46 = W*in
   wire signed [14:0] m134_46;
   assign m134_46 =15'b0;

   // m134_47 = W*in
   wire signed [14:0] m134_47;
   assign m134_47 ={ {4{neg134[14]}} , neg134[14:4] };

   // m134_48 = W*in
   wire signed [14:0] m134_48;
   assign m134_48 ={ {2{in134[14]}} , in134[14:2] };

   // m134_49 = W*in
   wire signed [14:0] m134_49;
   assign m134_49 =15'b0;

   // m134_50 = W*in
   wire signed [14:0] m134_50;
   assign m134_50 =15'b0;

   // m134_51 = W*in
   wire signed [14:0] m134_51;
   assign m134_51 =15'b0;

   // m134_52 = W*in
   wire signed [14:0] m134_52;
   assign m134_52 =15'b0;

   // m134_53 = W*in
   wire signed [14:0] m134_53;
   assign m134_53 =15'b0;

   // m134_54 = W*in
   wire signed [14:0] m134_54;
   assign m134_54 =15'b0;

   // m134_55 = W*in
   wire signed [14:0] m134_55;
   assign m134_55 =15'b0;

   // m134_56 = W*in
   wire signed [14:0] m134_56;
   assign m134_56 =15'b0;

   // m134_57 = W*in
   wire signed [14:0] m134_57;
   assign m134_57 =15'b0;

   // m134_58 = W*in
   wire signed [14:0] m134_58;
   assign m134_58 =15'b0;

   // m134_59 = W*in
   wire signed [14:0] m134_59;
   assign m134_59 =15'b0;

   // m134_60 = W*in
   wire signed [14:0] m134_60;
   assign m134_60 ={ {4{in134[14]}} , in134[14:4] };

   // m134_61 = W*in
   wire signed [14:0] m134_61;
   assign m134_61 =15'b0;

   // m134_62 = W*in
   wire signed [14:0] m134_62;
   assign m134_62 =15'b0;

   // m134_63 = W*in
   wire signed [14:0] m134_63;
   assign m134_63 =15'b0;

   // m134_64 = W*in
   wire signed [14:0] m134_64;
   assign m134_64 =15'b0;

   // m134_65 = W*in
   wire signed [14:0] m134_65;
   assign m134_65 ={ {3{in134[14]}} , in134[14:3] };

   // m134_66 = W*in
   wire signed [14:0] m134_66;
   assign m134_66 ={ {4{neg134[14]}} , neg134[14:4] };

   // m134_67 = W*in
   wire signed [14:0] m134_67;
   assign m134_67 =15'b0;

   // m134_68 = W*in
   wire signed [14:0] m134_68;
   assign m134_68 =15'b0;

   // m134_69 = W*in
   wire signed [14:0] m134_69;
   assign m134_69 =15'b0;

   // m134_70 = W*in
   wire signed [14:0] m134_70;
   assign m134_70 =15'b0;

   // m134_71 = W*in
   wire signed [14:0] m134_71;
   assign m134_71 =15'b0;

   // m134_72 = W*in
   wire signed [14:0] m134_72;
   assign m134_72 =15'b0;

   // m134_73 = W*in
   wire signed [14:0] m134_73;
   assign m134_73 ={ {4{neg134[14]}} , neg134[14:4] };

   // m134_74 = W*in
   wire signed [14:0] m134_74;
   assign m134_74 ={ {3{neg134[14]}} , neg134[14:3] };

   // m134_75 = W*in
   wire signed [14:0] m134_75;
   assign m134_75 =15'b0;

   // m134_76 = W*in
   wire signed [14:0] m134_76;
   assign m134_76 ={ {3{neg134[14]}} , neg134[14:3] };

   // m134_77 = W*in
   wire signed [14:0] m134_77;
   assign m134_77 =15'b0;

   // m134_78 = W*in
   wire signed [14:0] m134_78;
   assign m134_78 =15'b0;

   // m134_79 = W*in
   wire signed [14:0] m134_79;
   assign m134_79 =15'b0;

   // m134_80 = W*in
   wire signed [14:0] m134_80;
   assign m134_80 =15'b0;

   // m134_81 = W*in
   wire signed [14:0] m134_81;
   assign m134_81 =15'b0;

   // m134_82 = W*in
   wire signed [14:0] m134_82;
   assign m134_82 =15'b0;

   // m134_83 = W*in
   wire signed [14:0] m134_83;
   assign m134_83 =15'b0;

   // m134_84 = W*in
   wire signed [14:0] m134_84;
   assign m134_84 =15'b0;

   // m134_85 = W*in
   wire signed [14:0] m134_85;
   assign m134_85 =15'b0;

   // m134_86 = W*in
   wire signed [14:0] m134_86;
   assign m134_86 =15'b0;

   // m134_87 = W*in
   wire signed [14:0] m134_87;
   assign m134_87 =15'b0;

   // m134_88 = W*in
   wire signed [14:0] m134_88;
   assign m134_88 =15'b0;

   // m134_89 = W*in
   wire signed [14:0] m134_89;
   assign m134_89 ={ {3{neg134[14]}} , neg134[14:3] };

   // m134_90 = W*in
   wire signed [14:0] m134_90;
   assign m134_90 =15'b0;

   // m134_91 = W*in
   wire signed [14:0] m134_91;
   assign m134_91 =15'b0;

   // m134_92 = W*in
   wire signed [14:0] m134_92;
   assign m134_92 =15'b0;

   // m134_93 = W*in
   wire signed [14:0] m134_93;
   assign m134_93 =15'b0;

   // m134_94 = W*in
   wire signed [14:0] m134_94;
   assign m134_94 =15'b0;

   // m134_95 = W*in
   wire signed [14:0] m134_95;
   assign m134_95 =15'b0;

   // m134_96 = W*in
   wire signed [14:0] m134_96;
   assign m134_96 =15'b0;

   // m134_97 = W*in
   wire signed [14:0] m134_97;
   assign m134_97 =15'b0;

   // m134_98 = W*in
   wire signed [14:0] m134_98;
   assign m134_98 =15'b0;

   // m134_99 = W*in
   wire signed [14:0] m134_99;
   assign m134_99 =15'b0;

   // m134_100 = W*in
   wire signed [14:0] m134_100;
   assign m134_100 =15'b0;

   // m135_1 = W*in
   wire signed [14:0] m135_1;
   assign m135_1 =15'b0;

   // m135_2 = W*in
   wire signed [14:0] m135_2;
   assign m135_2 =15'b0;

   // m135_3 = W*in
   wire signed [14:0] m135_3;
   assign m135_3 =15'b0;

   // m135_4 = W*in
   wire signed [14:0] m135_4;
   assign m135_4 =15'b0;

   // m135_5 = W*in
   wire signed [14:0] m135_5;
   assign m135_5 =15'b0;

   // m135_6 = W*in
   wire signed [14:0] m135_6;
   assign m135_6 =15'b0;

   // m135_7 = W*in
   wire signed [14:0] m135_7;
   assign m135_7 =15'b0;

   // m135_8 = W*in
   wire signed [14:0] m135_8;
   assign m135_8 =15'b0;

   // m135_9 = W*in
   wire signed [14:0] m135_9;
   assign m135_9 =15'b0;

   // m135_10 = W*in
   wire signed [14:0] m135_10;
   assign m135_10 =15'b0;

   // m135_11 = W*in
   wire signed [14:0] m135_11;
   assign m135_11 =15'b0;

   // m135_12 = W*in
   wire signed [14:0] m135_12;
   assign m135_12 ={ {3{in135[14]}} , in135[14:3] };

   // m135_13 = W*in
   wire signed [14:0] m135_13;
   assign m135_13 =15'b0;

   // m135_14 = W*in
   wire signed [14:0] m135_14;
   assign m135_14 =15'b0;

   // m135_15 = W*in
   wire signed [14:0] m135_15;
   assign m135_15 =15'b0;

   // m135_16 = W*in
   wire signed [14:0] m135_16;
   assign m135_16 =15'b0;

   // m135_17 = W*in
   wire signed [14:0] m135_17;
   assign m135_17 ={ {4{neg135[14]}} , neg135[14:4] };

   // m135_18 = W*in
   wire signed [14:0] m135_18;
   assign m135_18 ={ {4{in135[14]}} , in135[14:4] };

   // m135_19 = W*in
   wire signed [14:0] m135_19;
   assign m135_19 ={ {3{neg135[14]}} , neg135[14:3] };

   // m135_20 = W*in
   wire signed [14:0] m135_20;
   assign m135_20 =15'b0;

   // m135_21 = W*in
   wire signed [14:0] m135_21;
   assign m135_21 =15'b0;

   // m135_22 = W*in
   wire signed [14:0] m135_22;
   assign m135_22 =15'b0;

   // m135_23 = W*in
   wire signed [14:0] m135_23;
   assign m135_23 =15'b0;

   // m135_24 = W*in
   wire signed [14:0] m135_24;
   assign m135_24 =15'b0;

   // m135_25 = W*in
   wire signed [14:0] m135_25;
   assign m135_25 ={ {3{neg135[14]}} , neg135[14:3] };

   // m135_26 = W*in
   wire signed [14:0] m135_26;
   assign m135_26 =15'b0;

   // m135_27 = W*in
   wire signed [14:0] m135_27;
   assign m135_27 =15'b0;

   // m135_28 = W*in
   wire signed [14:0] m135_28;
   assign m135_28 =15'b0;

   // m135_29 = W*in
   wire signed [14:0] m135_29;
   assign m135_29 ={ {3{in135[14]}} , in135[14:3] };

   // m135_30 = W*in
   wire signed [14:0] m135_30;
   assign m135_30 =15'b0;

   // m135_31 = W*in
   wire signed [14:0] m135_31;
   assign m135_31 ={ {3{in135[14]}} , in135[14:3] };

   // m135_32 = W*in
   wire signed [14:0] m135_32;
   assign m135_32 =15'b0;

   // m135_33 = W*in
   wire signed [14:0] m135_33;
   assign m135_33 =15'b0;

   // m135_34 = W*in
   wire signed [14:0] m135_34;
   assign m135_34 =15'b0;

   // m135_35 = W*in
   wire signed [14:0] m135_35;
   assign m135_35 =15'b0;

   // m135_36 = W*in
   wire signed [14:0] m135_36;
   assign m135_36 =15'b0;

   // m135_37 = W*in
   wire signed [14:0] m135_37;
   assign m135_37 =15'b0;

   // m135_38 = W*in
   wire signed [14:0] m135_38;
   assign m135_38 =15'b0;

   // m135_39 = W*in
   wire signed [14:0] m135_39;
   assign m135_39 =15'b0;

   // m135_40 = W*in
   wire signed [14:0] m135_40;
   assign m135_40 =15'b0;

   // m135_41 = W*in
   wire signed [14:0] m135_41;
   assign m135_41 =15'b0;

   // m135_42 = W*in
   wire signed [14:0] m135_42;
   assign m135_42 =15'b0;

   // m135_43 = W*in
   wire signed [14:0] m135_43;
   assign m135_43 =15'b0;

   // m135_44 = W*in
   wire signed [14:0] m135_44;
   assign m135_44 =15'b0;

   // m135_45 = W*in
   wire signed [14:0] m135_45;
   assign m135_45 =15'b0;

   // m135_46 = W*in
   wire signed [14:0] m135_46;
   assign m135_46 =15'b0;

   // m135_47 = W*in
   wire signed [14:0] m135_47;
   assign m135_47 =15'b0;

   // m135_48 = W*in
   wire signed [14:0] m135_48;
   assign m135_48 =15'b0;

   // m135_49 = W*in
   wire signed [14:0] m135_49;
   assign m135_49 =15'b0;

   // m135_50 = W*in
   wire signed [14:0] m135_50;
   assign m135_50 =15'b0;

   // m135_51 = W*in
   wire signed [14:0] m135_51;
   assign m135_51 =15'b0;

   // m135_52 = W*in
   wire signed [14:0] m135_52;
   assign m135_52 ={ {3{in135[14]}} , in135[14:3] };

   // m135_53 = W*in
   wire signed [14:0] m135_53;
   assign m135_53 =15'b0;

   // m135_54 = W*in
   wire signed [14:0] m135_54;
   assign m135_54 =15'b0;

   // m135_55 = W*in
   wire signed [14:0] m135_55;
   assign m135_55 =15'b0;

   // m135_56 = W*in
   wire signed [14:0] m135_56;
   assign m135_56 =15'b0;

   // m135_57 = W*in
   wire signed [14:0] m135_57;
   assign m135_57 =15'b0;

   // m135_58 = W*in
   wire signed [14:0] m135_58;
   assign m135_58 =15'b0;

   // m135_59 = W*in
   wire signed [14:0] m135_59;
   assign m135_59 =15'b0;

   // m135_60 = W*in
   wire signed [14:0] m135_60;
   assign m135_60 ={ {4{in135[14]}} , in135[14:4] };

   // m135_61 = W*in
   wire signed [14:0] m135_61;
   assign m135_61 =15'b0;

   // m135_62 = W*in
   wire signed [14:0] m135_62;
   assign m135_62 =15'b0;

   // m135_63 = W*in
   wire signed [14:0] m135_63;
   assign m135_63 =15'b0;

   // m135_64 = W*in
   wire signed [14:0] m135_64;
   assign m135_64 =15'b0;

   // m135_65 = W*in
   wire signed [14:0] m135_65;
   assign m135_65 =15'b0;

   // m135_66 = W*in
   wire signed [14:0] m135_66;
   assign m135_66 =15'b0;

   // m135_67 = W*in
   wire signed [14:0] m135_67;
   assign m135_67 =15'b0;

   // m135_68 = W*in
   wire signed [14:0] m135_68;
   assign m135_68 =15'b0;

   // m135_69 = W*in
   wire signed [14:0] m135_69;
   assign m135_69 =15'b0;

   // m135_70 = W*in
   wire signed [14:0] m135_70;
   assign m135_70 =15'b0;

   // m135_71 = W*in
   wire signed [14:0] m135_71;
   assign m135_71 =15'b0;

   // m135_72 = W*in
   wire signed [14:0] m135_72;
   assign m135_72 ={ {3{neg135[14]}} , neg135[14:3] };

   // m135_73 = W*in
   wire signed [14:0] m135_73;
   assign m135_73 ={ {4{in135[14]}} , in135[14:4] };

   // m135_74 = W*in
   wire signed [14:0] m135_74;
   assign m135_74 =15'b0;

   // m135_75 = W*in
   wire signed [14:0] m135_75;
   assign m135_75 =15'b0;

   // m135_76 = W*in
   wire signed [14:0] m135_76;
   assign m135_76 =15'b0;

   // m135_77 = W*in
   wire signed [14:0] m135_77;
   assign m135_77 =15'b0;

   // m135_78 = W*in
   wire signed [14:0] m135_78;
   assign m135_78 =15'b0;

   // m135_79 = W*in
   wire signed [14:0] m135_79;
   assign m135_79 =15'b0;

   // m135_80 = W*in
   wire signed [14:0] m135_80;
   assign m135_80 =15'b0;

   // m135_81 = W*in
   wire signed [14:0] m135_81;
   assign m135_81 ={ {4{in135[14]}} , in135[14:4] };

   // m135_82 = W*in
   wire signed [14:0] m135_82;
   assign m135_82 =15'b0;

   // m135_83 = W*in
   wire signed [14:0] m135_83;
   assign m135_83 =15'b0;

   // m135_84 = W*in
   wire signed [14:0] m135_84;
   assign m135_84 =15'b0;

   // m135_85 = W*in
   wire signed [14:0] m135_85;
   assign m135_85 =15'b0;

   // m135_86 = W*in
   wire signed [14:0] m135_86;
   assign m135_86 =15'b0;

   // m135_87 = W*in
   wire signed [14:0] m135_87;
   assign m135_87 =15'b0;

   // m135_88 = W*in
   wire signed [14:0] m135_88;
   assign m135_88 =15'b0;

   // m135_89 = W*in
   wire signed [14:0] m135_89;
   assign m135_89 =15'b0;

   // m135_90 = W*in
   wire signed [14:0] m135_90;
   assign m135_90 ={ {4{neg135[14]}} , neg135[14:4] };

   // m135_91 = W*in
   wire signed [14:0] m135_91;
   assign m135_91 =15'b0;

   // m135_92 = W*in
   wire signed [14:0] m135_92;
   assign m135_92 =15'b0;

   // m135_93 = W*in
   wire signed [14:0] m135_93;
   assign m135_93 =15'b0;

   // m135_94 = W*in
   wire signed [14:0] m135_94;
   assign m135_94 =15'b0;

   // m135_95 = W*in
   wire signed [14:0] m135_95;
   assign m135_95 =15'b0;

   // m135_96 = W*in
   wire signed [14:0] m135_96;
   assign m135_96 =15'b0;

   // m135_97 = W*in
   wire signed [14:0] m135_97;
   assign m135_97 =15'b0;

   // m135_98 = W*in
   wire signed [14:0] m135_98;
   assign m135_98 =15'b0;

   // m135_99 = W*in
   wire signed [14:0] m135_99;
   assign m135_99 =15'b0;

   // m135_100 = W*in
   wire signed [14:0] m135_100;
   assign m135_100 =15'b0;

   // m136_1 = W*in
   wire signed [14:0] m136_1;
   assign m136_1 =15'b0;

   // m136_2 = W*in
   wire signed [14:0] m136_2;
   assign m136_2 =15'b0;

   // m136_3 = W*in
   wire signed [14:0] m136_3;
   assign m136_3 =15'b0;

   // m136_4 = W*in
   wire signed [14:0] m136_4;
   assign m136_4 =15'b0;

   // m136_5 = W*in
   wire signed [14:0] m136_5;
   assign m136_5 ={ {3{neg136[14]}} , neg136[14:3] };

   // m136_6 = W*in
   wire signed [14:0] m136_6;
   assign m136_6 =15'b0;

   // m136_7 = W*in
   wire signed [14:0] m136_7;
   assign m136_7 =15'b0;

   // m136_8 = W*in
   wire signed [14:0] m136_8;
   assign m136_8 =15'b0;

   // m136_9 = W*in
   wire signed [14:0] m136_9;
   assign m136_9 =15'b0;

   // m136_10 = W*in
   wire signed [14:0] m136_10;
   assign m136_10 =15'b0;

   // m136_11 = W*in
   wire signed [14:0] m136_11;
   assign m136_11 =15'b0;

   // m136_12 = W*in
   wire signed [14:0] m136_12;
   assign m136_12 ={ {3{neg136[14]}} , neg136[14:3] };

   // m136_13 = W*in
   wire signed [14:0] m136_13;
   assign m136_13 =15'b0;

   // m136_14 = W*in
   wire signed [14:0] m136_14;
   assign m136_14 =15'b0;

   // m136_15 = W*in
   wire signed [14:0] m136_15;
   assign m136_15 =15'b0;

   // m136_16 = W*in
   wire signed [14:0] m136_16;
   assign m136_16 =15'b0;

   // m136_17 = W*in
   wire signed [14:0] m136_17;
   assign m136_17 =15'b0;

   // m136_18 = W*in
   wire signed [14:0] m136_18;
   assign m136_18 =15'b0;

   // m136_19 = W*in
   wire signed [14:0] m136_19;
   assign m136_19 =15'b0;

   // m136_20 = W*in
   wire signed [14:0] m136_20;
   assign m136_20 ={ {3{neg136[14]}} , neg136[14:3] };

   // m136_21 = W*in
   wire signed [14:0] m136_21;
   assign m136_21 =15'b0;

   // m136_22 = W*in
   wire signed [14:0] m136_22;
   assign m136_22 ={ {3{neg136[14]}} , neg136[14:3] };

   // m136_23 = W*in
   wire signed [14:0] m136_23;
   assign m136_23 =15'b0;

   // m136_24 = W*in
   wire signed [14:0] m136_24;
   assign m136_24 =15'b0;

   // m136_25 = W*in
   wire signed [14:0] m136_25;
   assign m136_25 ={ {4{in136[14]}} , in136[14:4] };

   // m136_26 = W*in
   wire signed [14:0] m136_26;
   assign m136_26 =15'b0;

   // m136_27 = W*in
   wire signed [14:0] m136_27;
   assign m136_27 =15'b0;

   // m136_28 = W*in
   wire signed [14:0] m136_28;
   assign m136_28 ={ {4{in136[14]}} , in136[14:4] };

   // m136_29 = W*in
   wire signed [14:0] m136_29;
   assign m136_29 =15'b0;

   // m136_30 = W*in
   wire signed [14:0] m136_30;
   assign m136_30 =15'b0;

   // m136_31 = W*in
   wire signed [14:0] m136_31;
   assign m136_31 =15'b0;

   // m136_32 = W*in
   wire signed [14:0] m136_32;
   assign m136_32 =15'b0;

   // m136_33 = W*in
   wire signed [14:0] m136_33;
   assign m136_33 =15'b0;

   // m136_34 = W*in
   wire signed [14:0] m136_34;
   assign m136_34 =15'b0;

   // m136_35 = W*in
   wire signed [14:0] m136_35;
   assign m136_35 =15'b0;

   // m136_36 = W*in
   wire signed [14:0] m136_36;
   assign m136_36 =15'b0;

   // m136_37 = W*in
   wire signed [14:0] m136_37;
   assign m136_37 =15'b0;

   // m136_38 = W*in
   wire signed [14:0] m136_38;
   assign m136_38 =15'b0;

   // m136_39 = W*in
   wire signed [14:0] m136_39;
   assign m136_39 =15'b0;

   // m136_40 = W*in
   wire signed [14:0] m136_40;
   assign m136_40 =15'b0;

   // m136_41 = W*in
   wire signed [14:0] m136_41;
   assign m136_41 =15'b0;

   // m136_42 = W*in
   wire signed [14:0] m136_42;
   assign m136_42 =15'b0;

   // m136_43 = W*in
   wire signed [14:0] m136_43;
   assign m136_43 =15'b0;

   // m136_44 = W*in
   wire signed [14:0] m136_44;
   assign m136_44 =15'b0;

   // m136_45 = W*in
   wire signed [14:0] m136_45;
   assign m136_45 =15'b0;

   // m136_46 = W*in
   wire signed [14:0] m136_46;
   assign m136_46 =15'b0;

   // m136_47 = W*in
   wire signed [14:0] m136_47;
   assign m136_47 =15'b0;

   // m136_48 = W*in
   wire signed [14:0] m136_48;
   assign m136_48 =15'b0;

   // m136_49 = W*in
   wire signed [14:0] m136_49;
   assign m136_49 =15'b0;

   // m136_50 = W*in
   wire signed [14:0] m136_50;
   assign m136_50 ={ {3{in136[14]}} , in136[14:3] };

   // m136_51 = W*in
   wire signed [14:0] m136_51;
   assign m136_51 =15'b0;

   // m136_52 = W*in
   wire signed [14:0] m136_52;
   assign m136_52 =15'b0;

   // m136_53 = W*in
   wire signed [14:0] m136_53;
   assign m136_53 =15'b0;

   // m136_54 = W*in
   wire signed [14:0] m136_54;
   assign m136_54 ={ {3{in136[14]}} , in136[14:3] };

   // m136_55 = W*in
   wire signed [14:0] m136_55;
   assign m136_55 ={ {3{in136[14]}} , in136[14:3] };

   // m136_56 = W*in
   wire signed [14:0] m136_56;
   assign m136_56 ={ {4{in136[14]}} , in136[14:4] };

   // m136_57 = W*in
   wire signed [14:0] m136_57;
   assign m136_57 =15'b0;

   // m136_58 = W*in
   wire signed [14:0] m136_58;
   assign m136_58 ={ {4{neg136[14]}} , neg136[14:4] };

   // m136_59 = W*in
   wire signed [14:0] m136_59;
   assign m136_59 =15'b0;

   // m136_60 = W*in
   wire signed [14:0] m136_60;
   assign m136_60 =15'b0;

   // m136_61 = W*in
   wire signed [14:0] m136_61;
   assign m136_61 ={ {4{neg136[14]}} , neg136[14:4] };

   // m136_62 = W*in
   wire signed [14:0] m136_62;
   assign m136_62 =15'b0;

   // m136_63 = W*in
   wire signed [14:0] m136_63;
   assign m136_63 =15'b0;

   // m136_64 = W*in
   wire signed [14:0] m136_64;
   assign m136_64 =15'b0;

   // m136_65 = W*in
   wire signed [14:0] m136_65;
   assign m136_65 =15'b0;

   // m136_66 = W*in
   wire signed [14:0] m136_66;
   assign m136_66 =15'b0;

   // m136_67 = W*in
   wire signed [14:0] m136_67;
   assign m136_67 ={ {4{in136[14]}} , in136[14:4] };

   // m136_68 = W*in
   wire signed [14:0] m136_68;
   assign m136_68 =15'b0;

   // m136_69 = W*in
   wire signed [14:0] m136_69;
   assign m136_69 ={ {4{in136[14]}} , in136[14:4] };

   // m136_70 = W*in
   wire signed [14:0] m136_70;
   assign m136_70 ={ {3{in136[14]}} , in136[14:3] };

   // m136_71 = W*in
   wire signed [14:0] m136_71;
   assign m136_71 =15'b0;

   // m136_72 = W*in
   wire signed [14:0] m136_72;
   assign m136_72 =15'b0;

   // m136_73 = W*in
   wire signed [14:0] m136_73;
   assign m136_73 =15'b0;

   // m136_74 = W*in
   wire signed [14:0] m136_74;
   assign m136_74 ={ {4{neg136[14]}} , neg136[14:4] };

   // m136_75 = W*in
   wire signed [14:0] m136_75;
   assign m136_75 =15'b0;

   // m136_76 = W*in
   wire signed [14:0] m136_76;
   assign m136_76 =15'b0;

   // m136_77 = W*in
   wire signed [14:0] m136_77;
   assign m136_77 =15'b0;

   // m136_78 = W*in
   wire signed [14:0] m136_78;
   assign m136_78 =15'b0;

   // m136_79 = W*in
   wire signed [14:0] m136_79;
   assign m136_79 =15'b0;

   // m136_80 = W*in
   wire signed [14:0] m136_80;
   assign m136_80 =15'b0;

   // m136_81 = W*in
   wire signed [14:0] m136_81;
   assign m136_81 =15'b0;

   // m136_82 = W*in
   wire signed [14:0] m136_82;
   assign m136_82 =15'b0;

   // m136_83 = W*in
   wire signed [14:0] m136_83;
   assign m136_83 =15'b0;

   // m136_84 = W*in
   wire signed [14:0] m136_84;
   assign m136_84 =15'b0;

   // m136_85 = W*in
   wire signed [14:0] m136_85;
   assign m136_85 =15'b0;

   // m136_86 = W*in
   wire signed [14:0] m136_86;
   assign m136_86 =15'b0;

   // m136_87 = W*in
   wire signed [14:0] m136_87;
   assign m136_87 =15'b0;

   // m136_88 = W*in
   wire signed [14:0] m136_88;
   assign m136_88 =15'b0;

   // m136_89 = W*in
   wire signed [14:0] m136_89;
   assign m136_89 =15'b0;

   // m136_90 = W*in
   wire signed [14:0] m136_90;
   assign m136_90 =15'b0;

   // m136_91 = W*in
   wire signed [14:0] m136_91;
   assign m136_91 =15'b0;

   // m136_92 = W*in
   wire signed [14:0] m136_92;
   assign m136_92 =15'b0;

   // m136_93 = W*in
   wire signed [14:0] m136_93;
   assign m136_93 =15'b0;

   // m136_94 = W*in
   wire signed [14:0] m136_94;
   assign m136_94 =15'b0;

   // m136_95 = W*in
   wire signed [14:0] m136_95;
   assign m136_95 ={ {4{in136[14]}} , in136[14:4] };

   // m136_96 = W*in
   wire signed [14:0] m136_96;
   assign m136_96 =15'b0;

   // m136_97 = W*in
   wire signed [14:0] m136_97;
   assign m136_97 ={ {4{neg136[14]}} , neg136[14:4] };

   // m136_98 = W*in
   wire signed [14:0] m136_98;
   assign m136_98 =15'b0;

   // m136_99 = W*in
   wire signed [14:0] m136_99;
   assign m136_99 =15'b0;

   // m136_100 = W*in
   wire signed [14:0] m136_100;
   assign m136_100 =15'b0;

   // m137_1 = W*in
   wire signed [14:0] m137_1;
   assign m137_1 =15'b0;

   // m137_2 = W*in
   wire signed [14:0] m137_2;
   assign m137_2 =15'b0;

   // m137_3 = W*in
   wire signed [14:0] m137_3;
   assign m137_3 =15'b0;

   // m137_4 = W*in
   wire signed [14:0] m137_4;
   assign m137_4 ={ {3{in137[14]}} , in137[14:3] };

   // m137_5 = W*in
   wire signed [14:0] m137_5;
   assign m137_5 =15'b0;

   // m137_6 = W*in
   wire signed [14:0] m137_6;
   assign m137_6 =15'b0;

   // m137_7 = W*in
   wire signed [14:0] m137_7;
   assign m137_7 =15'b0;

   // m137_8 = W*in
   wire signed [14:0] m137_8;
   assign m137_8 =15'b0;

   // m137_9 = W*in
   wire signed [14:0] m137_9;
   assign m137_9 =15'b0;

   // m137_10 = W*in
   wire signed [14:0] m137_10;
   assign m137_10 =15'b0;

   // m137_11 = W*in
   wire signed [14:0] m137_11;
   assign m137_11 =15'b0;

   // m137_12 = W*in
   wire signed [14:0] m137_12;
   assign m137_12 =15'b0;

   // m137_13 = W*in
   wire signed [14:0] m137_13;
   assign m137_13 =15'b0;

   // m137_14 = W*in
   wire signed [14:0] m137_14;
   assign m137_14 =15'b0;

   // m137_15 = W*in
   wire signed [14:0] m137_15;
   assign m137_15 =15'b0;

   // m137_16 = W*in
   wire signed [14:0] m137_16;
   assign m137_16 =15'b0;

   // m137_17 = W*in
   wire signed [14:0] m137_17;
   assign m137_17 =15'b0;

   // m137_18 = W*in
   wire signed [14:0] m137_18;
   assign m137_18 =15'b0;

   // m137_19 = W*in
   wire signed [14:0] m137_19;
   assign m137_19 =15'b0;

   // m137_20 = W*in
   wire signed [14:0] m137_20;
   assign m137_20 ={ {4{neg137[14]}} , neg137[14:4] };

   // m137_21 = W*in
   wire signed [14:0] m137_21;
   assign m137_21 ={ {4{neg137[14]}} , neg137[14:4] };

   // m137_22 = W*in
   wire signed [14:0] m137_22;
   assign m137_22 =15'b0;

   // m137_23 = W*in
   wire signed [14:0] m137_23;
   assign m137_23 =15'b0;

   // m137_24 = W*in
   wire signed [14:0] m137_24;
   assign m137_24 =15'b0;

   // m137_25 = W*in
   wire signed [14:0] m137_25;
   assign m137_25 ={ {4{in137[14]}} , in137[14:4] };

   // m137_26 = W*in
   wire signed [14:0] m137_26;
   assign m137_26 ={ {4{neg137[14]}} , neg137[14:4] };

   // m137_27 = W*in
   wire signed [14:0] m137_27;
   assign m137_27 =15'b0;

   // m137_28 = W*in
   wire signed [14:0] m137_28;
   assign m137_28 =15'b0;

   // m137_29 = W*in
   wire signed [14:0] m137_29;
   assign m137_29 =15'b0;

   // m137_30 = W*in
   wire signed [14:0] m137_30;
   assign m137_30 =15'b0;

   // m137_31 = W*in
   wire signed [14:0] m137_31;
   assign m137_31 =15'b0;

   // m137_32 = W*in
   wire signed [14:0] m137_32;
   assign m137_32 =15'b0;

   // m137_33 = W*in
   wire signed [14:0] m137_33;
   assign m137_33 =15'b0;

   // m137_34 = W*in
   wire signed [14:0] m137_34;
   assign m137_34 =15'b0;

   // m137_35 = W*in
   wire signed [14:0] m137_35;
   assign m137_35 =15'b0;

   // m137_36 = W*in
   wire signed [14:0] m137_36;
   assign m137_36 =15'b0;

   // m137_37 = W*in
   wire signed [14:0] m137_37;
   assign m137_37 =15'b0;

   // m137_38 = W*in
   wire signed [14:0] m137_38;
   assign m137_38 =15'b0;

   // m137_39 = W*in
   wire signed [14:0] m137_39;
   assign m137_39 ={ {3{in137[14]}} , in137[14:3] };

   // m137_40 = W*in
   wire signed [14:0] m137_40;
   assign m137_40 =15'b0;

   // m137_41 = W*in
   wire signed [14:0] m137_41;
   assign m137_41 =15'b0;

   // m137_42 = W*in
   wire signed [14:0] m137_42;
   assign m137_42 =15'b0;

   // m137_43 = W*in
   wire signed [14:0] m137_43;
   assign m137_43 =15'b0;

   // m137_44 = W*in
   wire signed [14:0] m137_44;
   assign m137_44 =15'b0;

   // m137_45 = W*in
   wire signed [14:0] m137_45;
   assign m137_45 =15'b0;

   // m137_46 = W*in
   wire signed [14:0] m137_46;
   assign m137_46 =15'b0;

   // m137_47 = W*in
   wire signed [14:0] m137_47;
   assign m137_47 =15'b0;

   // m137_48 = W*in
   wire signed [14:0] m137_48;
   assign m137_48 =15'b0;

   // m137_49 = W*in
   wire signed [14:0] m137_49;
   assign m137_49 =15'b0;

   // m137_50 = W*in
   wire signed [14:0] m137_50;
   assign m137_50 =15'b0;

   // m137_51 = W*in
   wire signed [14:0] m137_51;
   assign m137_51 =15'b0;

   // m137_52 = W*in
   wire signed [14:0] m137_52;
   assign m137_52 =15'b0;

   // m137_53 = W*in
   wire signed [14:0] m137_53;
   assign m137_53 =15'b0;

   // m137_54 = W*in
   wire signed [14:0] m137_54;
   assign m137_54 ={ {3{in137[14]}} , in137[14:3] };

   // m137_55 = W*in
   wire signed [14:0] m137_55;
   assign m137_55 =15'b0;

   // m137_56 = W*in
   wire signed [14:0] m137_56;
   assign m137_56 =15'b0;

   // m137_57 = W*in
   wire signed [14:0] m137_57;
   assign m137_57 =15'b0;

   // m137_58 = W*in
   wire signed [14:0] m137_58;
   assign m137_58 =15'b0;

   // m137_59 = W*in
   wire signed [14:0] m137_59;
   assign m137_59 =15'b0;

   // m137_60 = W*in
   wire signed [14:0] m137_60;
   assign m137_60 =15'b0;

   // m137_61 = W*in
   wire signed [14:0] m137_61;
   assign m137_61 ={ {4{neg137[14]}} , neg137[14:4] };

   // m137_62 = W*in
   wire signed [14:0] m137_62;
   assign m137_62 =15'b0;

   // m137_63 = W*in
   wire signed [14:0] m137_63;
   assign m137_63 =15'b0;

   // m137_64 = W*in
   wire signed [14:0] m137_64;
   assign m137_64 =15'b0;

   // m137_65 = W*in
   wire signed [14:0] m137_65;
   assign m137_65 =15'b0;

   // m137_66 = W*in
   wire signed [14:0] m137_66;
   assign m137_66 ={ {4{in137[14]}} , in137[14:4] };

   // m137_67 = W*in
   wire signed [14:0] m137_67;
   assign m137_67 =15'b0;

   // m137_68 = W*in
   wire signed [14:0] m137_68;
   assign m137_68 =15'b0;

   // m137_69 = W*in
   wire signed [14:0] m137_69;
   assign m137_69 =15'b0;

   // m137_70 = W*in
   wire signed [14:0] m137_70;
   assign m137_70 =15'b0;

   // m137_71 = W*in
   wire signed [14:0] m137_71;
   assign m137_71 =15'b0;

   // m137_72 = W*in
   wire signed [14:0] m137_72;
   assign m137_72 ={ {3{in137[14]}} , in137[14:3] };

   // m137_73 = W*in
   wire signed [14:0] m137_73;
   assign m137_73 =15'b0;

   // m137_74 = W*in
   wire signed [14:0] m137_74;
   assign m137_74 =15'b0;

   // m137_75 = W*in
   wire signed [14:0] m137_75;
   assign m137_75 =15'b0;

   // m137_76 = W*in
   wire signed [14:0] m137_76;
   assign m137_76 =15'b0;

   // m137_77 = W*in
   wire signed [14:0] m137_77;
   assign m137_77 =15'b0;

   // m137_78 = W*in
   wire signed [14:0] m137_78;
   assign m137_78 =15'b0;

   // m137_79 = W*in
   wire signed [14:0] m137_79;
   assign m137_79 =15'b0;

   // m137_80 = W*in
   wire signed [14:0] m137_80;
   assign m137_80 =15'b0;

   // m137_81 = W*in
   wire signed [14:0] m137_81;
   assign m137_81 =15'b0;

   // m137_82 = W*in
   wire signed [14:0] m137_82;
   assign m137_82 =15'b0;

   // m137_83 = W*in
   wire signed [14:0] m137_83;
   assign m137_83 =15'b0;

   // m137_84 = W*in
   wire signed [14:0] m137_84;
   assign m137_84 =15'b0;

   // m137_85 = W*in
   wire signed [14:0] m137_85;
   assign m137_85 =15'b0;

   // m137_86 = W*in
   wire signed [14:0] m137_86;
   assign m137_86 =15'b0;

   // m137_87 = W*in
   wire signed [14:0] m137_87;
   assign m137_87 =15'b0;

   // m137_88 = W*in
   wire signed [14:0] m137_88;
   assign m137_88 =15'b0;

   // m137_89 = W*in
   wire signed [14:0] m137_89;
   assign m137_89 =15'b0;

   // m137_90 = W*in
   wire signed [14:0] m137_90;
   assign m137_90 =15'b0;

   // m137_91 = W*in
   wire signed [14:0] m137_91;
   assign m137_91 =15'b0;

   // m137_92 = W*in
   wire signed [14:0] m137_92;
   assign m137_92 =15'b0;

   // m137_93 = W*in
   wire signed [14:0] m137_93;
   assign m137_93 =15'b0;

   // m137_94 = W*in
   wire signed [14:0] m137_94;
   assign m137_94 =15'b0;

   // m137_95 = W*in
   wire signed [14:0] m137_95;
   assign m137_95 =15'b0;

   // m137_96 = W*in
   wire signed [14:0] m137_96;
   assign m137_96 =15'b0;

   // m137_97 = W*in
   wire signed [14:0] m137_97;
   assign m137_97 =15'b0;

   // m137_98 = W*in
   wire signed [14:0] m137_98;
   assign m137_98 =15'b0;

   // m137_99 = W*in
   wire signed [14:0] m137_99;
   assign m137_99 =15'b0;

   // m137_100 = W*in
   wire signed [14:0] m137_100;
   assign m137_100 =15'b0;

   // m138_1 = W*in
   wire signed [14:0] m138_1;
   assign m138_1 ={ {3{in138[14]}} , in138[14:3] };

   // m138_2 = W*in
   wire signed [14:0] m138_2;
   assign m138_2 =15'b0;

   // m138_3 = W*in
   wire signed [14:0] m138_3;
   assign m138_3 =15'b0;

   // m138_4 = W*in
   wire signed [14:0] m138_4;
   assign m138_4 =15'b0;

   // m138_5 = W*in
   wire signed [14:0] m138_5;
   assign m138_5 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_6 = W*in
   wire signed [14:0] m138_6;
   assign m138_6 =15'b0;

   // m138_7 = W*in
   wire signed [14:0] m138_7;
   assign m138_7 ={ {4{in138[14]}} , in138[14:4] };

   // m138_8 = W*in
   wire signed [14:0] m138_8;
   assign m138_8 ={ {4{in138[14]}} , in138[14:4] };

   // m138_9 = W*in
   wire signed [14:0] m138_9;
   assign m138_9 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_10 = W*in
   wire signed [14:0] m138_10;
   assign m138_10 =15'b0;

   // m138_11 = W*in
   wire signed [14:0] m138_11;
   assign m138_11 =15'b0;

   // m138_12 = W*in
   wire signed [14:0] m138_12;
   assign m138_12 =15'b0;

   // m138_13 = W*in
   wire signed [14:0] m138_13;
   assign m138_13 =15'b0;

   // m138_14 = W*in
   wire signed [14:0] m138_14;
   assign m138_14 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_15 = W*in
   wire signed [14:0] m138_15;
   assign m138_15 =15'b0;

   // m138_16 = W*in
   wire signed [14:0] m138_16;
   assign m138_16 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_17 = W*in
   wire signed [14:0] m138_17;
   assign m138_17 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_18 = W*in
   wire signed [14:0] m138_18;
   assign m138_18 =15'b0;

   // m138_19 = W*in
   wire signed [14:0] m138_19;
   assign m138_19 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_20 = W*in
   wire signed [14:0] m138_20;
   assign m138_20 =15'b0;

   // m138_21 = W*in
   wire signed [14:0] m138_21;
   assign m138_21 =15'b0;

   // m138_22 = W*in
   wire signed [14:0] m138_22;
   assign m138_22 ={ {4{in138[14]}} , in138[14:4] };

   // m138_23 = W*in
   wire signed [14:0] m138_23;
   assign m138_23 =15'b0;

   // m138_24 = W*in
   wire signed [14:0] m138_24;
   assign m138_24 =15'b0;

   // m138_25 = W*in
   wire signed [14:0] m138_25;
   assign m138_25 =15'b0;

   // m138_26 = W*in
   wire signed [14:0] m138_26;
   assign m138_26 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_27 = W*in
   wire signed [14:0] m138_27;
   assign m138_27 =15'b0;

   // m138_28 = W*in
   wire signed [14:0] m138_28;
   assign m138_28 =15'b0;

   // m138_29 = W*in
   wire signed [14:0] m138_29;
   assign m138_29 =15'b0;

   // m138_30 = W*in
   wire signed [14:0] m138_30;
   assign m138_30 =15'b0;

   // m138_31 = W*in
   wire signed [14:0] m138_31;
   assign m138_31 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_32 = W*in
   wire signed [14:0] m138_32;
   assign m138_32 =15'b0;

   // m138_33 = W*in
   wire signed [14:0] m138_33;
   assign m138_33 =15'b0;

   // m138_34 = W*in
   wire signed [14:0] m138_34;
   assign m138_34 =15'b0;

   // m138_35 = W*in
   wire signed [14:0] m138_35;
   assign m138_35 =15'b0;

   // m138_36 = W*in
   wire signed [14:0] m138_36;
   assign m138_36 =15'b0;

   // m138_37 = W*in
   wire signed [14:0] m138_37;
   assign m138_37 =15'b0;

   // m138_38 = W*in
   wire signed [14:0] m138_38;
   assign m138_38 =15'b0;

   // m138_39 = W*in
   wire signed [14:0] m138_39;
   assign m138_39 =15'b0;

   // m138_40 = W*in
   wire signed [14:0] m138_40;
   assign m138_40 =15'b0;

   // m138_41 = W*in
   wire signed [14:0] m138_41;
   assign m138_41 =15'b0;

   // m138_42 = W*in
   wire signed [14:0] m138_42;
   assign m138_42 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_43 = W*in
   wire signed [14:0] m138_43;
   assign m138_43 =15'b0;

   // m138_44 = W*in
   wire signed [14:0] m138_44;
   assign m138_44 =15'b0;

   // m138_45 = W*in
   wire signed [14:0] m138_45;
   assign m138_45 =15'b0;

   // m138_46 = W*in
   wire signed [14:0] m138_46;
   assign m138_46 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_47 = W*in
   wire signed [14:0] m138_47;
   assign m138_47 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_48 = W*in
   wire signed [14:0] m138_48;
   assign m138_48 =15'b0;

   // m138_49 = W*in
   wire signed [14:0] m138_49;
   assign m138_49 =15'b0;

   // m138_50 = W*in
   wire signed [14:0] m138_50;
   assign m138_50 =15'b0;

   // m138_51 = W*in
   wire signed [14:0] m138_51;
   assign m138_51 =15'b0;

   // m138_52 = W*in
   wire signed [14:0] m138_52;
   assign m138_52 =15'b0;

   // m138_53 = W*in
   wire signed [14:0] m138_53;
   assign m138_53 =15'b0;

   // m138_54 = W*in
   wire signed [14:0] m138_54;
   assign m138_54 =15'b0;

   // m138_55 = W*in
   wire signed [14:0] m138_55;
   assign m138_55 =15'b0;

   // m138_56 = W*in
   wire signed [14:0] m138_56;
   assign m138_56 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_57 = W*in
   wire signed [14:0] m138_57;
   assign m138_57 =15'b0;

   // m138_58 = W*in
   wire signed [14:0] m138_58;
   assign m138_58 =15'b0;

   // m138_59 = W*in
   wire signed [14:0] m138_59;
   assign m138_59 =15'b0;

   // m138_60 = W*in
   wire signed [14:0] m138_60;
   assign m138_60 =15'b0;

   // m138_61 = W*in
   wire signed [14:0] m138_61;
   assign m138_61 =15'b0;

   // m138_62 = W*in
   wire signed [14:0] m138_62;
   assign m138_62 =15'b0;

   // m138_63 = W*in
   wire signed [14:0] m138_63;
   assign m138_63 =15'b0;

   // m138_64 = W*in
   wire signed [14:0] m138_64;
   assign m138_64 =15'b0;

   // m138_65 = W*in
   wire signed [14:0] m138_65;
   assign m138_65 ={ {3{in138[14]}} , in138[14:3] };

   // m138_66 = W*in
   wire signed [14:0] m138_66;
   assign m138_66 =15'b0;

   // m138_67 = W*in
   wire signed [14:0] m138_67;
   assign m138_67 =15'b0;

   // m138_68 = W*in
   wire signed [14:0] m138_68;
   assign m138_68 =15'b0;

   // m138_69 = W*in
   wire signed [14:0] m138_69;
   assign m138_69 =15'b0;

   // m138_70 = W*in
   wire signed [14:0] m138_70;
   assign m138_70 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_71 = W*in
   wire signed [14:0] m138_71;
   assign m138_71 =15'b0;

   // m138_72 = W*in
   wire signed [14:0] m138_72;
   assign m138_72 =15'b0;

   // m138_73 = W*in
   wire signed [14:0] m138_73;
   assign m138_73 =15'b0;

   // m138_74 = W*in
   wire signed [14:0] m138_74;
   assign m138_74 ={ {4{neg138[14]}} , neg138[14:4] };

   // m138_75 = W*in
   wire signed [14:0] m138_75;
   assign m138_75 =15'b0;

   // m138_76 = W*in
   wire signed [14:0] m138_76;
   assign m138_76 =15'b0;

   // m138_77 = W*in
   wire signed [14:0] m138_77;
   assign m138_77 =15'b0;

   // m138_78 = W*in
   wire signed [14:0] m138_78;
   assign m138_78 =15'b0;

   // m138_79 = W*in
   wire signed [14:0] m138_79;
   assign m138_79 =15'b0;

   // m138_80 = W*in
   wire signed [14:0] m138_80;
   assign m138_80 ={ {4{in138[14]}} , in138[14:4] };

   // m138_81 = W*in
   wire signed [14:0] m138_81;
   assign m138_81 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_82 = W*in
   wire signed [14:0] m138_82;
   assign m138_82 =15'b0;

   // m138_83 = W*in
   wire signed [14:0] m138_83;
   assign m138_83 =15'b0;

   // m138_84 = W*in
   wire signed [14:0] m138_84;
   assign m138_84 =15'b0;

   // m138_85 = W*in
   wire signed [14:0] m138_85;
   assign m138_85 =15'b0;

   // m138_86 = W*in
   wire signed [14:0] m138_86;
   assign m138_86 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_87 = W*in
   wire signed [14:0] m138_87;
   assign m138_87 =15'b0;

   // m138_88 = W*in
   wire signed [14:0] m138_88;
   assign m138_88 =15'b0;

   // m138_89 = W*in
   wire signed [14:0] m138_89;
   assign m138_89 =15'b0;

   // m138_90 = W*in
   wire signed [14:0] m138_90;
   assign m138_90 =15'b0;

   // m138_91 = W*in
   wire signed [14:0] m138_91;
   assign m138_91 =15'b0;

   // m138_92 = W*in
   wire signed [14:0] m138_92;
   assign m138_92 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_93 = W*in
   wire signed [14:0] m138_93;
   assign m138_93 =15'b0;

   // m138_94 = W*in
   wire signed [14:0] m138_94;
   assign m138_94 ={ {3{neg138[14]}} , neg138[14:3] };

   // m138_95 = W*in
   wire signed [14:0] m138_95;
   assign m138_95 =15'b0;

   // m138_96 = W*in
   wire signed [14:0] m138_96;
   assign m138_96 =15'b0;

   // m138_97 = W*in
   wire signed [14:0] m138_97;
   assign m138_97 =15'b0;

   // m138_98 = W*in
   wire signed [14:0] m138_98;
   assign m138_98 =15'b0;

   // m138_99 = W*in
   wire signed [14:0] m138_99;
   assign m138_99 =15'b0;

   // m138_100 = W*in
   wire signed [14:0] m138_100;
   assign m138_100 =15'b0;

   // m139_1 = W*in
   wire signed [14:0] m139_1;
   assign m139_1 =15'b0;

   // m139_2 = W*in
   wire signed [14:0] m139_2;
   assign m139_2 =15'b0;

   // m139_3 = W*in
   wire signed [14:0] m139_3;
   assign m139_3 =15'b0;

   // m139_4 = W*in
   wire signed [14:0] m139_4;
   assign m139_4 =15'b0;

   // m139_5 = W*in
   wire signed [14:0] m139_5;
   assign m139_5 =15'b0;

   // m139_6 = W*in
   wire signed [14:0] m139_6;
   assign m139_6 =15'b0;

   // m139_7 = W*in
   wire signed [14:0] m139_7;
   assign m139_7 ={ {4{neg139[14]}} , neg139[14:4] };

   // m139_8 = W*in
   wire signed [14:0] m139_8;
   assign m139_8 =15'b0;

   // m139_9 = W*in
   wire signed [14:0] m139_9;
   assign m139_9 =15'b0;

   // m139_10 = W*in
   wire signed [14:0] m139_10;
   assign m139_10 ={ {3{neg139[14]}} , neg139[14:3] };

   // m139_11 = W*in
   wire signed [14:0] m139_11;
   assign m139_11 =15'b0;

   // m139_12 = W*in
   wire signed [14:0] m139_12;
   assign m139_12 =15'b0;

   // m139_13 = W*in
   wire signed [14:0] m139_13;
   assign m139_13 =15'b0;

   // m139_14 = W*in
   wire signed [14:0] m139_14;
   assign m139_14 =15'b0;

   // m139_15 = W*in
   wire signed [14:0] m139_15;
   assign m139_15 =15'b0;

   // m139_16 = W*in
   wire signed [14:0] m139_16;
   assign m139_16 =15'b0;

   // m139_17 = W*in
   wire signed [14:0] m139_17;
   assign m139_17 =15'b0;

   // m139_18 = W*in
   wire signed [14:0] m139_18;
   assign m139_18 =15'b0;

   // m139_19 = W*in
   wire signed [14:0] m139_19;
   assign m139_19 =15'b0;

   // m139_20 = W*in
   wire signed [14:0] m139_20;
   assign m139_20 =15'b0;

   // m139_21 = W*in
   wire signed [14:0] m139_21;
   assign m139_21 =15'b0;

   // m139_22 = W*in
   wire signed [14:0] m139_22;
   assign m139_22 =15'b0;

   // m139_23 = W*in
   wire signed [14:0] m139_23;
   assign m139_23 =15'b0;

   // m139_24 = W*in
   wire signed [14:0] m139_24;
   assign m139_24 =15'b0;

   // m139_25 = W*in
   wire signed [14:0] m139_25;
   assign m139_25 =15'b0;

   // m139_26 = W*in
   wire signed [14:0] m139_26;
   assign m139_26 =15'b0;

   // m139_27 = W*in
   wire signed [14:0] m139_27;
   assign m139_27 =15'b0;

   // m139_28 = W*in
   wire signed [14:0] m139_28;
   assign m139_28 =15'b0;

   // m139_29 = W*in
   wire signed [14:0] m139_29;
   assign m139_29 =15'b0;

   // m139_30 = W*in
   wire signed [14:0] m139_30;
   assign m139_30 =15'b0;

   // m139_31 = W*in
   wire signed [14:0] m139_31;
   assign m139_31 =15'b0;

   // m139_32 = W*in
   wire signed [14:0] m139_32;
   assign m139_32 =15'b0;

   // m139_33 = W*in
   wire signed [14:0] m139_33;
   assign m139_33 ={ {4{neg139[14]}} , neg139[14:4] };

   // m139_34 = W*in
   wire signed [14:0] m139_34;
   assign m139_34 =15'b0;

   // m139_35 = W*in
   wire signed [14:0] m139_35;
   assign m139_35 =15'b0;

   // m139_36 = W*in
   wire signed [14:0] m139_36;
   assign m139_36 =15'b0;

   // m139_37 = W*in
   wire signed [14:0] m139_37;
   assign m139_37 =15'b0;

   // m139_38 = W*in
   wire signed [14:0] m139_38;
   assign m139_38 =15'b0;

   // m139_39 = W*in
   wire signed [14:0] m139_39;
   assign m139_39 =15'b0;

   // m139_40 = W*in
   wire signed [14:0] m139_40;
   assign m139_40 =15'b0;

   // m139_41 = W*in
   wire signed [14:0] m139_41;
   assign m139_41 =15'b0;

   // m139_42 = W*in
   wire signed [14:0] m139_42;
   assign m139_42 =15'b0;

   // m139_43 = W*in
   wire signed [14:0] m139_43;
   assign m139_43 =15'b0;

   // m139_44 = W*in
   wire signed [14:0] m139_44;
   assign m139_44 ={ {3{in139[14]}} , in139[14:3] };

   // m139_45 = W*in
   wire signed [14:0] m139_45;
   assign m139_45 =15'b0;

   // m139_46 = W*in
   wire signed [14:0] m139_46;
   assign m139_46 =15'b0;

   // m139_47 = W*in
   wire signed [14:0] m139_47;
   assign m139_47 =15'b0;

   // m139_48 = W*in
   wire signed [14:0] m139_48;
   assign m139_48 =15'b0;

   // m139_49 = W*in
   wire signed [14:0] m139_49;
   assign m139_49 =15'b0;

   // m139_50 = W*in
   wire signed [14:0] m139_50;
   assign m139_50 =15'b0;

   // m139_51 = W*in
   wire signed [14:0] m139_51;
   assign m139_51 =15'b0;

   // m139_52 = W*in
   wire signed [14:0] m139_52;
   assign m139_52 =15'b0;

   // m139_53 = W*in
   wire signed [14:0] m139_53;
   assign m139_53 =15'b0;

   // m139_54 = W*in
   wire signed [14:0] m139_54;
   assign m139_54 =15'b0;

   // m139_55 = W*in
   wire signed [14:0] m139_55;
   assign m139_55 =15'b0;

   // m139_56 = W*in
   wire signed [14:0] m139_56;
   assign m139_56 =15'b0;

   // m139_57 = W*in
   wire signed [14:0] m139_57;
   assign m139_57 =15'b0;

   // m139_58 = W*in
   wire signed [14:0] m139_58;
   assign m139_58 =15'b0;

   // m139_59 = W*in
   wire signed [14:0] m139_59;
   assign m139_59 =15'b0;

   // m139_60 = W*in
   wire signed [14:0] m139_60;
   assign m139_60 =15'b0;

   // m139_61 = W*in
   wire signed [14:0] m139_61;
   assign m139_61 =15'b0;

   // m139_62 = W*in
   wire signed [14:0] m139_62;
   assign m139_62 =15'b0;

   // m139_63 = W*in
   wire signed [14:0] m139_63;
   assign m139_63 ={ {3{neg139[14]}} , neg139[14:3] };

   // m139_64 = W*in
   wire signed [14:0] m139_64;
   assign m139_64 =15'b0;

   // m139_65 = W*in
   wire signed [14:0] m139_65;
   assign m139_65 =15'b0;

   // m139_66 = W*in
   wire signed [14:0] m139_66;
   assign m139_66 =15'b0;

   // m139_67 = W*in
   wire signed [14:0] m139_67;
   assign m139_67 =15'b0;

   // m139_68 = W*in
   wire signed [14:0] m139_68;
   assign m139_68 =15'b0;

   // m139_69 = W*in
   wire signed [14:0] m139_69;
   assign m139_69 =15'b0;

   // m139_70 = W*in
   wire signed [14:0] m139_70;
   assign m139_70 =15'b0;

   // m139_71 = W*in
   wire signed [14:0] m139_71;
   assign m139_71 =15'b0;

   // m139_72 = W*in
   wire signed [14:0] m139_72;
   assign m139_72 =15'b0;

   // m139_73 = W*in
   wire signed [14:0] m139_73;
   assign m139_73 =15'b0;

   // m139_74 = W*in
   wire signed [14:0] m139_74;
   assign m139_74 ={ {3{neg139[14]}} , neg139[14:3] };

   // m139_75 = W*in
   wire signed [14:0] m139_75;
   assign m139_75 =15'b0;

   // m139_76 = W*in
   wire signed [14:0] m139_76;
   assign m139_76 =15'b0;

   // m139_77 = W*in
   wire signed [14:0] m139_77;
   assign m139_77 =15'b0;

   // m139_78 = W*in
   wire signed [14:0] m139_78;
   assign m139_78 =15'b0;

   // m139_79 = W*in
   wire signed [14:0] m139_79;
   assign m139_79 =15'b0;

   // m139_80 = W*in
   wire signed [14:0] m139_80;
   assign m139_80 =15'b0;

   // m139_81 = W*in
   wire signed [14:0] m139_81;
   assign m139_81 =15'b0;

   // m139_82 = W*in
   wire signed [14:0] m139_82;
   assign m139_82 =15'b0;

   // m139_83 = W*in
   wire signed [14:0] m139_83;
   assign m139_83 =15'b0;

   // m139_84 = W*in
   wire signed [14:0] m139_84;
   assign m139_84 =15'b0;

   // m139_85 = W*in
   wire signed [14:0] m139_85;
   assign m139_85 =15'b0;

   // m139_86 = W*in
   wire signed [14:0] m139_86;
   assign m139_86 =15'b0;

   // m139_87 = W*in
   wire signed [14:0] m139_87;
   assign m139_87 =15'b0;

   // m139_88 = W*in
   wire signed [14:0] m139_88;
   assign m139_88 ={ {4{neg139[14]}} , neg139[14:4] };

   // m139_89 = W*in
   wire signed [14:0] m139_89;
   assign m139_89 =15'b0;

   // m139_90 = W*in
   wire signed [14:0] m139_90;
   assign m139_90 =15'b0;

   // m139_91 = W*in
   wire signed [14:0] m139_91;
   assign m139_91 =15'b0;

   // m139_92 = W*in
   wire signed [14:0] m139_92;
   assign m139_92 =15'b0;

   // m139_93 = W*in
   wire signed [14:0] m139_93;
   assign m139_93 =15'b0;

   // m139_94 = W*in
   wire signed [14:0] m139_94;
   assign m139_94 =15'b0;

   // m139_95 = W*in
   wire signed [14:0] m139_95;
   assign m139_95 =15'b0;

   // m139_96 = W*in
   wire signed [14:0] m139_96;
   assign m139_96 =15'b0;

   // m139_97 = W*in
   wire signed [14:0] m139_97;
   assign m139_97 =15'b0;

   // m139_98 = W*in
   wire signed [14:0] m139_98;
   assign m139_98 =15'b0;

   // m139_99 = W*in
   wire signed [14:0] m139_99;
   assign m139_99 =15'b0;

   // m139_100 = W*in
   wire signed [14:0] m139_100;
   assign m139_100 =15'b0;

   // m140_1 = W*in
   wire signed [14:0] m140_1;
   assign m140_1 =15'b0;

   // m140_2 = W*in
   wire signed [14:0] m140_2;
   assign m140_2 =15'b0;

   // m140_3 = W*in
   wire signed [14:0] m140_3;
   assign m140_3 =15'b0;

   // m140_4 = W*in
   wire signed [14:0] m140_4;
   assign m140_4 =15'b0;

   // m140_5 = W*in
   wire signed [14:0] m140_5;
   assign m140_5 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_6 = W*in
   wire signed [14:0] m140_6;
   assign m140_6 =15'b0;

   // m140_7 = W*in
   wire signed [14:0] m140_7;
   assign m140_7 =15'b0;

   // m140_8 = W*in
   wire signed [14:0] m140_8;
   assign m140_8 ={ {3{in140[14]}} , in140[14:3] };

   // m140_9 = W*in
   wire signed [14:0] m140_9;
   assign m140_9 =15'b0;

   // m140_10 = W*in
   wire signed [14:0] m140_10;
   assign m140_10 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_11 = W*in
   wire signed [14:0] m140_11;
   assign m140_11 =15'b0;

   // m140_12 = W*in
   wire signed [14:0] m140_12;
   assign m140_12 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_13 = W*in
   wire signed [14:0] m140_13;
   assign m140_13 ={ {3{in140[14]}} , in140[14:3] };

   // m140_14 = W*in
   wire signed [14:0] m140_14;
   assign m140_14 =15'b0;

   // m140_15 = W*in
   wire signed [14:0] m140_15;
   assign m140_15 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_16 = W*in
   wire signed [14:0] m140_16;
   assign m140_16 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_17 = W*in
   wire signed [14:0] m140_17;
   assign m140_17 ={ {3{in140[14]}} , in140[14:3] };

   // m140_18 = W*in
   wire signed [14:0] m140_18;
   assign m140_18 =15'b0;

   // m140_19 = W*in
   wire signed [14:0] m140_19;
   assign m140_19 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_20 = W*in
   wire signed [14:0] m140_20;
   assign m140_20 =15'b0;

   // m140_21 = W*in
   wire signed [14:0] m140_21;
   assign m140_21 ={ {4{in140[14]}} , in140[14:4] };

   // m140_22 = W*in
   wire signed [14:0] m140_22;
   assign m140_22 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_23 = W*in
   wire signed [14:0] m140_23;
   assign m140_23 ={ {3{in140[14]}} , in140[14:3] };

   // m140_24 = W*in
   wire signed [14:0] m140_24;
   assign m140_24 =15'b0;

   // m140_25 = W*in
   wire signed [14:0] m140_25;
   assign m140_25 ={ {4{in140[14]}} , in140[14:4] };

   // m140_26 = W*in
   wire signed [14:0] m140_26;
   assign m140_26 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_27 = W*in
   wire signed [14:0] m140_27;
   assign m140_27 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_28 = W*in
   wire signed [14:0] m140_28;
   assign m140_28 ={ {4{in140[14]}} , in140[14:4] };

   // m140_29 = W*in
   wire signed [14:0] m140_29;
   assign m140_29 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_30 = W*in
   wire signed [14:0] m140_30;
   assign m140_30 =15'b0;

   // m140_31 = W*in
   wire signed [14:0] m140_31;
   assign m140_31 =15'b0;

   // m140_32 = W*in
   wire signed [14:0] m140_32;
   assign m140_32 ={ {4{neg140[14]}} , neg140[14:4] };

   // m140_33 = W*in
   wire signed [14:0] m140_33;
   assign m140_33 =15'b0;

   // m140_34 = W*in
   wire signed [14:0] m140_34;
   assign m140_34 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_35 = W*in
   wire signed [14:0] m140_35;
   assign m140_35 =15'b0;

   // m140_36 = W*in
   wire signed [14:0] m140_36;
   assign m140_36 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_37 = W*in
   wire signed [14:0] m140_37;
   assign m140_37 ={ {3{in140[14]}} , in140[14:3] };

   // m140_38 = W*in
   wire signed [14:0] m140_38;
   assign m140_38 =15'b0;

   // m140_39 = W*in
   wire signed [14:0] m140_39;
   assign m140_39 =15'b0;

   // m140_40 = W*in
   wire signed [14:0] m140_40;
   assign m140_40 =15'b0;

   // m140_41 = W*in
   wire signed [14:0] m140_41;
   assign m140_41 ={ {3{in140[14]}} , in140[14:3] };

   // m140_42 = W*in
   wire signed [14:0] m140_42;
   assign m140_42 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_43 = W*in
   wire signed [14:0] m140_43;
   assign m140_43 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_44 = W*in
   wire signed [14:0] m140_44;
   assign m140_44 =15'b0;

   // m140_45 = W*in
   wire signed [14:0] m140_45;
   assign m140_45 ={ {3{in140[14]}} , in140[14:3] };

   // m140_46 = W*in
   wire signed [14:0] m140_46;
   assign m140_46 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_47 = W*in
   wire signed [14:0] m140_47;
   assign m140_47 =15'b0;

   // m140_48 = W*in
   wire signed [14:0] m140_48;
   assign m140_48 =15'b0;

   // m140_49 = W*in
   wire signed [14:0] m140_49;
   assign m140_49 =15'b0;

   // m140_50 = W*in
   wire signed [14:0] m140_50;
   assign m140_50 =15'b0;

   // m140_51 = W*in
   wire signed [14:0] m140_51;
   assign m140_51 =15'b0;

   // m140_52 = W*in
   wire signed [14:0] m140_52;
   assign m140_52 =15'b0;

   // m140_53 = W*in
   wire signed [14:0] m140_53;
   assign m140_53 =15'b0;

   // m140_54 = W*in
   wire signed [14:0] m140_54;
   assign m140_54 =15'b0;

   // m140_55 = W*in
   wire signed [14:0] m140_55;
   assign m140_55 =15'b0;

   // m140_56 = W*in
   wire signed [14:0] m140_56;
   assign m140_56 ={ {3{in140[14]}} , in140[14:3] };

   // m140_57 = W*in
   wire signed [14:0] m140_57;
   assign m140_57 =15'b0;

   // m140_58 = W*in
   wire signed [14:0] m140_58;
   assign m140_58 =15'b0;

   // m140_59 = W*in
   wire signed [14:0] m140_59;
   assign m140_59 =15'b0;

   // m140_60 = W*in
   wire signed [14:0] m140_60;
   assign m140_60 =15'b0;

   // m140_61 = W*in
   wire signed [14:0] m140_61;
   assign m140_61 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_62 = W*in
   wire signed [14:0] m140_62;
   assign m140_62 =15'b0;

   // m140_63 = W*in
   wire signed [14:0] m140_63;
   assign m140_63 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_64 = W*in
   wire signed [14:0] m140_64;
   assign m140_64 =15'b0;

   // m140_65 = W*in
   wire signed [14:0] m140_65;
   assign m140_65 ={ {2{neg140[14]}} , neg140[14:2] };

   // m140_66 = W*in
   wire signed [14:0] m140_66;
   assign m140_66 ={ {4{neg140[14]}} , neg140[14:4] };

   // m140_67 = W*in
   wire signed [14:0] m140_67;
   assign m140_67 =15'b0;

   // m140_68 = W*in
   wire signed [14:0] m140_68;
   assign m140_68 ={ {4{in140[14]}} , in140[14:4] };

   // m140_69 = W*in
   wire signed [14:0] m140_69;
   assign m140_69 ={ {4{neg140[14]}} , neg140[14:4] };

   // m140_70 = W*in
   wire signed [14:0] m140_70;
   assign m140_70 ={ {2{in140[14]}} , in140[14:2] };

   // m140_71 = W*in
   wire signed [14:0] m140_71;
   assign m140_71 =15'b0;

   // m140_72 = W*in
   wire signed [14:0] m140_72;
   assign m140_72 =15'b0;

   // m140_73 = W*in
   wire signed [14:0] m140_73;
   assign m140_73 =15'b0;

   // m140_74 = W*in
   wire signed [14:0] m140_74;
   assign m140_74 ={ {4{in140[14]}} , in140[14:4] };

   // m140_75 = W*in
   wire signed [14:0] m140_75;
   assign m140_75 =15'b0;

   // m140_76 = W*in
   wire signed [14:0] m140_76;
   assign m140_76 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_77 = W*in
   wire signed [14:0] m140_77;
   assign m140_77 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_78 = W*in
   wire signed [14:0] m140_78;
   assign m140_78 =15'b0;

   // m140_79 = W*in
   wire signed [14:0] m140_79;
   assign m140_79 =15'b0;

   // m140_80 = W*in
   wire signed [14:0] m140_80;
   assign m140_80 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_81 = W*in
   wire signed [14:0] m140_81;
   assign m140_81 =15'b0;

   // m140_82 = W*in
   wire signed [14:0] m140_82;
   assign m140_82 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_83 = W*in
   wire signed [14:0] m140_83;
   assign m140_83 =15'b0;

   // m140_84 = W*in
   wire signed [14:0] m140_84;
   assign m140_84 =15'b0;

   // m140_85 = W*in
   wire signed [14:0] m140_85;
   assign m140_85 =15'b0;

   // m140_86 = W*in
   wire signed [14:0] m140_86;
   assign m140_86 =15'b0;

   // m140_87 = W*in
   wire signed [14:0] m140_87;
   assign m140_87 =15'b0;

   // m140_88 = W*in
   wire signed [14:0] m140_88;
   assign m140_88 =15'b0;

   // m140_89 = W*in
   wire signed [14:0] m140_89;
   assign m140_89 =15'b0;

   // m140_90 = W*in
   wire signed [14:0] m140_90;
   assign m140_90 =15'b0;

   // m140_91 = W*in
   wire signed [14:0] m140_91;
   assign m140_91 =15'b0;

   // m140_92 = W*in
   wire signed [14:0] m140_92;
   assign m140_92 =15'b0;

   // m140_93 = W*in
   wire signed [14:0] m140_93;
   assign m140_93 =15'b0;

   // m140_94 = W*in
   wire signed [14:0] m140_94;
   assign m140_94 =15'b0;

   // m140_95 = W*in
   wire signed [14:0] m140_95;
   assign m140_95 =15'b0;

   // m140_96 = W*in
   wire signed [14:0] m140_96;
   assign m140_96 =15'b0;

   // m140_97 = W*in
   wire signed [14:0] m140_97;
   assign m140_97 ={ {3{neg140[14]}} , neg140[14:3] };

   // m140_98 = W*in
   wire signed [14:0] m140_98;
   assign m140_98 =15'b0;

   // m140_99 = W*in
   wire signed [14:0] m140_99;
   assign m140_99 =15'b0;

   // m140_100 = W*in
   wire signed [14:0] m140_100;
   assign m140_100 =15'b0;

   // m141_1 = W*in
   wire signed [14:0] m141_1;
   assign m141_1 =15'b0;

   // m141_2 = W*in
   wire signed [14:0] m141_2;
   assign m141_2 =15'b0;

   // m141_3 = W*in
   wire signed [14:0] m141_3;
   assign m141_3 =15'b0;

   // m141_4 = W*in
   wire signed [14:0] m141_4;
   assign m141_4 =15'b0;

   // m141_5 = W*in
   wire signed [14:0] m141_5;
   assign m141_5 =15'b0;

   // m141_6 = W*in
   wire signed [14:0] m141_6;
   assign m141_6 =15'b0;

   // m141_7 = W*in
   wire signed [14:0] m141_7;
   assign m141_7 =15'b0;

   // m141_8 = W*in
   wire signed [14:0] m141_8;
   assign m141_8 =15'b0;

   // m141_9 = W*in
   wire signed [14:0] m141_9;
   assign m141_9 =15'b0;

   // m141_10 = W*in
   wire signed [14:0] m141_10;
   assign m141_10 =15'b0;

   // m141_11 = W*in
   wire signed [14:0] m141_11;
   assign m141_11 ={ {3{neg141[14]}} , neg141[14:3] };

   // m141_12 = W*in
   wire signed [14:0] m141_12;
   assign m141_12 =15'b0;

   // m141_13 = W*in
   wire signed [14:0] m141_13;
   assign m141_13 =15'b0;

   // m141_14 = W*in
   wire signed [14:0] m141_14;
   assign m141_14 =15'b0;

   // m141_15 = W*in
   wire signed [14:0] m141_15;
   assign m141_15 ={ {3{neg141[14]}} , neg141[14:3] };

   // m141_16 = W*in
   wire signed [14:0] m141_16;
   assign m141_16 =15'b0;

   // m141_17 = W*in
   wire signed [14:0] m141_17;
   assign m141_17 =15'b0;

   // m141_18 = W*in
   wire signed [14:0] m141_18;
   assign m141_18 =15'b0;

   // m141_19 = W*in
   wire signed [14:0] m141_19;
   assign m141_19 =15'b0;

   // m141_20 = W*in
   wire signed [14:0] m141_20;
   assign m141_20 =15'b0;

   // m141_21 = W*in
   wire signed [14:0] m141_21;
   assign m141_21 =15'b0;

   // m141_22 = W*in
   wire signed [14:0] m141_22;
   assign m141_22 =15'b0;

   // m141_23 = W*in
   wire signed [14:0] m141_23;
   assign m141_23 =15'b0;

   // m141_24 = W*in
   wire signed [14:0] m141_24;
   assign m141_24 =15'b0;

   // m141_25 = W*in
   wire signed [14:0] m141_25;
   assign m141_25 =15'b0;

   // m141_26 = W*in
   wire signed [14:0] m141_26;
   assign m141_26 =15'b0;

   // m141_27 = W*in
   wire signed [14:0] m141_27;
   assign m141_27 ={ {4{in141[14]}} , in141[14:4] };

   // m141_28 = W*in
   wire signed [14:0] m141_28;
   assign m141_28 =15'b0;

   // m141_29 = W*in
   wire signed [14:0] m141_29;
   assign m141_29 =15'b0;

   // m141_30 = W*in
   wire signed [14:0] m141_30;
   assign m141_30 ={ {3{neg141[14]}} , neg141[14:3] };

   // m141_31 = W*in
   wire signed [14:0] m141_31;
   assign m141_31 ={ {3{in141[14]}} , in141[14:3] };

   // m141_32 = W*in
   wire signed [14:0] m141_32;
   assign m141_32 =15'b0;

   // m141_33 = W*in
   wire signed [14:0] m141_33;
   assign m141_33 =15'b0;

   // m141_34 = W*in
   wire signed [14:0] m141_34;
   assign m141_34 =15'b0;

   // m141_35 = W*in
   wire signed [14:0] m141_35;
   assign m141_35 =15'b0;

   // m141_36 = W*in
   wire signed [14:0] m141_36;
   assign m141_36 =15'b0;

   // m141_37 = W*in
   wire signed [14:0] m141_37;
   assign m141_37 =15'b0;

   // m141_38 = W*in
   wire signed [14:0] m141_38;
   assign m141_38 =15'b0;

   // m141_39 = W*in
   wire signed [14:0] m141_39;
   assign m141_39 =15'b0;

   // m141_40 = W*in
   wire signed [14:0] m141_40;
   assign m141_40 =15'b0;

   // m141_41 = W*in
   wire signed [14:0] m141_41;
   assign m141_41 =15'b0;

   // m141_42 = W*in
   wire signed [14:0] m141_42;
   assign m141_42 =15'b0;

   // m141_43 = W*in
   wire signed [14:0] m141_43;
   assign m141_43 =15'b0;

   // m141_44 = W*in
   wire signed [14:0] m141_44;
   assign m141_44 =15'b0;

   // m141_45 = W*in
   wire signed [14:0] m141_45;
   assign m141_45 ={ {3{in141[14]}} , in141[14:3] };

   // m141_46 = W*in
   wire signed [14:0] m141_46;
   assign m141_46 =15'b0;

   // m141_47 = W*in
   wire signed [14:0] m141_47;
   assign m141_47 =15'b0;

   // m141_48 = W*in
   wire signed [14:0] m141_48;
   assign m141_48 =15'b0;

   // m141_49 = W*in
   wire signed [14:0] m141_49;
   assign m141_49 =15'b0;

   // m141_50 = W*in
   wire signed [14:0] m141_50;
   assign m141_50 =15'b0;

   // m141_51 = W*in
   wire signed [14:0] m141_51;
   assign m141_51 =15'b0;

   // m141_52 = W*in
   wire signed [14:0] m141_52;
   assign m141_52 =15'b0;

   // m141_53 = W*in
   wire signed [14:0] m141_53;
   assign m141_53 =15'b0;

   // m141_54 = W*in
   wire signed [14:0] m141_54;
   assign m141_54 =15'b0;

   // m141_55 = W*in
   wire signed [14:0] m141_55;
   assign m141_55 =15'b0;

   // m141_56 = W*in
   wire signed [14:0] m141_56;
   assign m141_56 =15'b0;

   // m141_57 = W*in
   wire signed [14:0] m141_57;
   assign m141_57 ={ {3{neg141[14]}} , neg141[14:3] };

   // m141_58 = W*in
   wire signed [14:0] m141_58;
   assign m141_58 =15'b0;

   // m141_59 = W*in
   wire signed [14:0] m141_59;
   assign m141_59 =15'b0;

   // m141_60 = W*in
   wire signed [14:0] m141_60;
   assign m141_60 =15'b0;

   // m141_61 = W*in
   wire signed [14:0] m141_61;
   assign m141_61 =15'b0;

   // m141_62 = W*in
   wire signed [14:0] m141_62;
   assign m141_62 =15'b0;

   // m141_63 = W*in
   wire signed [14:0] m141_63;
   assign m141_63 ={ {3{neg141[14]}} , neg141[14:3] };

   // m141_64 = W*in
   wire signed [14:0] m141_64;
   assign m141_64 =15'b0;

   // m141_65 = W*in
   wire signed [14:0] m141_65;
   assign m141_65 =15'b0;

   // m141_66 = W*in
   wire signed [14:0] m141_66;
   assign m141_66 =15'b0;

   // m141_67 = W*in
   wire signed [14:0] m141_67;
   assign m141_67 ={ {3{neg141[14]}} , neg141[14:3] };

   // m141_68 = W*in
   wire signed [14:0] m141_68;
   assign m141_68 =15'b0;

   // m141_69 = W*in
   wire signed [14:0] m141_69;
   assign m141_69 =15'b0;

   // m141_70 = W*in
   wire signed [14:0] m141_70;
   assign m141_70 ={ {4{neg141[14]}} , neg141[14:4] };

   // m141_71 = W*in
   wire signed [14:0] m141_71;
   assign m141_71 =15'b0;

   // m141_72 = W*in
   wire signed [14:0] m141_72;
   assign m141_72 =15'b0;

   // m141_73 = W*in
   wire signed [14:0] m141_73;
   assign m141_73 =15'b0;

   // m141_74 = W*in
   wire signed [14:0] m141_74;
   assign m141_74 =15'b0;

   // m141_75 = W*in
   wire signed [14:0] m141_75;
   assign m141_75 =15'b0;

   // m141_76 = W*in
   wire signed [14:0] m141_76;
   assign m141_76 =15'b0;

   // m141_77 = W*in
   wire signed [14:0] m141_77;
   assign m141_77 =15'b0;

   // m141_78 = W*in
   wire signed [14:0] m141_78;
   assign m141_78 =15'b0;

   // m141_79 = W*in
   wire signed [14:0] m141_79;
   assign m141_79 =15'b0;

   // m141_80 = W*in
   wire signed [14:0] m141_80;
   assign m141_80 ={ {4{neg141[14]}} , neg141[14:4] };

   // m141_81 = W*in
   wire signed [14:0] m141_81;
   assign m141_81 =15'b0;

   // m141_82 = W*in
   wire signed [14:0] m141_82;
   assign m141_82 =15'b0;

   // m141_83 = W*in
   wire signed [14:0] m141_83;
   assign m141_83 ={ {3{in141[14]}} , in141[14:3] };

   // m141_84 = W*in
   wire signed [14:0] m141_84;
   assign m141_84 =15'b0;

   // m141_85 = W*in
   wire signed [14:0] m141_85;
   assign m141_85 =15'b0;

   // m141_86 = W*in
   wire signed [14:0] m141_86;
   assign m141_86 =15'b0;

   // m141_87 = W*in
   wire signed [14:0] m141_87;
   assign m141_87 =15'b0;

   // m141_88 = W*in
   wire signed [14:0] m141_88;
   assign m141_88 =15'b0;

   // m141_89 = W*in
   wire signed [14:0] m141_89;
   assign m141_89 =15'b0;

   // m141_90 = W*in
   wire signed [14:0] m141_90;
   assign m141_90 =15'b0;

   // m141_91 = W*in
   wire signed [14:0] m141_91;
   assign m141_91 =15'b0;

   // m141_92 = W*in
   wire signed [14:0] m141_92;
   assign m141_92 =15'b0;

   // m141_93 = W*in
   wire signed [14:0] m141_93;
   assign m141_93 =15'b0;

   // m141_94 = W*in
   wire signed [14:0] m141_94;
   assign m141_94 =15'b0;

   // m141_95 = W*in
   wire signed [14:0] m141_95;
   assign m141_95 =15'b0;

   // m141_96 = W*in
   wire signed [14:0] m141_96;
   assign m141_96 =15'b0;

   // m141_97 = W*in
   wire signed [14:0] m141_97;
   assign m141_97 =15'b0;

   // m141_98 = W*in
   wire signed [14:0] m141_98;
   assign m141_98 =15'b0;

   // m141_99 = W*in
   wire signed [14:0] m141_99;
   assign m141_99 =15'b0;

   // m141_100 = W*in
   wire signed [14:0] m141_100;
   assign m141_100 =15'b0;

   // m142_1 = W*in
   wire signed [14:0] m142_1;
   assign m142_1 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_2 = W*in
   wire signed [14:0] m142_2;
   assign m142_2 =15'b0;

   // m142_3 = W*in
   wire signed [14:0] m142_3;
   assign m142_3 =15'b0;

   // m142_4 = W*in
   wire signed [14:0] m142_4;
   assign m142_4 =15'b0;

   // m142_5 = W*in
   wire signed [14:0] m142_5;
   assign m142_5 =15'b0;

   // m142_6 = W*in
   wire signed [14:0] m142_6;
   assign m142_6 =15'b0;

   // m142_7 = W*in
   wire signed [14:0] m142_7;
   assign m142_7 =15'b0;

   // m142_8 = W*in
   wire signed [14:0] m142_8;
   assign m142_8 =15'b0;

   // m142_9 = W*in
   wire signed [14:0] m142_9;
   assign m142_9 =15'b0;

   // m142_10 = W*in
   wire signed [14:0] m142_10;
   assign m142_10 =15'b0;

   // m142_11 = W*in
   wire signed [14:0] m142_11;
   assign m142_11 =15'b0;

   // m142_12 = W*in
   wire signed [14:0] m142_12;
   assign m142_12 =15'b0;

   // m142_13 = W*in
   wire signed [14:0] m142_13;
   assign m142_13 =15'b0;

   // m142_14 = W*in
   wire signed [14:0] m142_14;
   assign m142_14 =15'b0;

   // m142_15 = W*in
   wire signed [14:0] m142_15;
   assign m142_15 =15'b0;

   // m142_16 = W*in
   wire signed [14:0] m142_16;
   assign m142_16 =15'b0;

   // m142_17 = W*in
   wire signed [14:0] m142_17;
   assign m142_17 ={ {3{in142[14]}} , in142[14:3] };

   // m142_18 = W*in
   wire signed [14:0] m142_18;
   assign m142_18 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_19 = W*in
   wire signed [14:0] m142_19;
   assign m142_19 =15'b0;

   // m142_20 = W*in
   wire signed [14:0] m142_20;
   assign m142_20 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_21 = W*in
   wire signed [14:0] m142_21;
   assign m142_21 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_22 = W*in
   wire signed [14:0] m142_22;
   assign m142_22 =15'b0;

   // m142_23 = W*in
   wire signed [14:0] m142_23;
   assign m142_23 =15'b0;

   // m142_24 = W*in
   wire signed [14:0] m142_24;
   assign m142_24 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_25 = W*in
   wire signed [14:0] m142_25;
   assign m142_25 ={ {4{in142[14]}} , in142[14:4] };

   // m142_26 = W*in
   wire signed [14:0] m142_26;
   assign m142_26 =15'b0;

   // m142_27 = W*in
   wire signed [14:0] m142_27;
   assign m142_27 =15'b0;

   // m142_28 = W*in
   wire signed [14:0] m142_28;
   assign m142_28 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_29 = W*in
   wire signed [14:0] m142_29;
   assign m142_29 =15'b0;

   // m142_30 = W*in
   wire signed [14:0] m142_30;
   assign m142_30 =15'b0;

   // m142_31 = W*in
   wire signed [14:0] m142_31;
   assign m142_31 =15'b0;

   // m142_32 = W*in
   wire signed [14:0] m142_32;
   assign m142_32 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_33 = W*in
   wire signed [14:0] m142_33;
   assign m142_33 ={ {4{in142[14]}} , in142[14:4] };

   // m142_34 = W*in
   wire signed [14:0] m142_34;
   assign m142_34 =15'b0;

   // m142_35 = W*in
   wire signed [14:0] m142_35;
   assign m142_35 =15'b0;

   // m142_36 = W*in
   wire signed [14:0] m142_36;
   assign m142_36 =15'b0;

   // m142_37 = W*in
   wire signed [14:0] m142_37;
   assign m142_37 =15'b0;

   // m142_38 = W*in
   wire signed [14:0] m142_38;
   assign m142_38 =15'b0;

   // m142_39 = W*in
   wire signed [14:0] m142_39;
   assign m142_39 ={ {2{in142[14]}} , in142[14:2] };

   // m142_40 = W*in
   wire signed [14:0] m142_40;
   assign m142_40 =15'b0;

   // m142_41 = W*in
   wire signed [14:0] m142_41;
   assign m142_41 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_42 = W*in
   wire signed [14:0] m142_42;
   assign m142_42 =15'b0;

   // m142_43 = W*in
   wire signed [14:0] m142_43;
   assign m142_43 =15'b0;

   // m142_44 = W*in
   wire signed [14:0] m142_44;
   assign m142_44 ={ {3{in142[14]}} , in142[14:3] };

   // m142_45 = W*in
   wire signed [14:0] m142_45;
   assign m142_45 =15'b0;

   // m142_46 = W*in
   wire signed [14:0] m142_46;
   assign m142_46 =15'b0;

   // m142_47 = W*in
   wire signed [14:0] m142_47;
   assign m142_47 =15'b0;

   // m142_48 = W*in
   wire signed [14:0] m142_48;
   assign m142_48 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_49 = W*in
   wire signed [14:0] m142_49;
   assign m142_49 =15'b0;

   // m142_50 = W*in
   wire signed [14:0] m142_50;
   assign m142_50 =15'b0;

   // m142_51 = W*in
   wire signed [14:0] m142_51;
   assign m142_51 =15'b0;

   // m142_52 = W*in
   wire signed [14:0] m142_52;
   assign m142_52 =15'b0;

   // m142_53 = W*in
   wire signed [14:0] m142_53;
   assign m142_53 =15'b0;

   // m142_54 = W*in
   wire signed [14:0] m142_54;
   assign m142_54 ={ {3{in142[14]}} , in142[14:3] };

   // m142_55 = W*in
   wire signed [14:0] m142_55;
   assign m142_55 =15'b0;

   // m142_56 = W*in
   wire signed [14:0] m142_56;
   assign m142_56 ={ {3{in142[14]}} , in142[14:3] };

   // m142_57 = W*in
   wire signed [14:0] m142_57;
   assign m142_57 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_58 = W*in
   wire signed [14:0] m142_58;
   assign m142_58 =15'b0;

   // m142_59 = W*in
   wire signed [14:0] m142_59;
   assign m142_59 =15'b0;

   // m142_60 = W*in
   wire signed [14:0] m142_60;
   assign m142_60 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_61 = W*in
   wire signed [14:0] m142_61;
   assign m142_61 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_62 = W*in
   wire signed [14:0] m142_62;
   assign m142_62 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_63 = W*in
   wire signed [14:0] m142_63;
   assign m142_63 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_64 = W*in
   wire signed [14:0] m142_64;
   assign m142_64 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_65 = W*in
   wire signed [14:0] m142_65;
   assign m142_65 =15'b0;

   // m142_66 = W*in
   wire signed [14:0] m142_66;
   assign m142_66 ={ {3{in142[14]}} , in142[14:3] };

   // m142_67 = W*in
   wire signed [14:0] m142_67;
   assign m142_67 =15'b0;

   // m142_68 = W*in
   wire signed [14:0] m142_68;
   assign m142_68 ={ {4{neg142[14]}} , neg142[14:4] };

   // m142_69 = W*in
   wire signed [14:0] m142_69;
   assign m142_69 =15'b0;

   // m142_70 = W*in
   wire signed [14:0] m142_70;
   assign m142_70 =15'b0;

   // m142_71 = W*in
   wire signed [14:0] m142_71;
   assign m142_71 =15'b0;

   // m142_72 = W*in
   wire signed [14:0] m142_72;
   assign m142_72 =15'b0;

   // m142_73 = W*in
   wire signed [14:0] m142_73;
   assign m142_73 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_74 = W*in
   wire signed [14:0] m142_74;
   assign m142_74 =15'b0;

   // m142_75 = W*in
   wire signed [14:0] m142_75;
   assign m142_75 =15'b0;

   // m142_76 = W*in
   wire signed [14:0] m142_76;
   assign m142_76 =15'b0;

   // m142_77 = W*in
   wire signed [14:0] m142_77;
   assign m142_77 =15'b0;

   // m142_78 = W*in
   wire signed [14:0] m142_78;
   assign m142_78 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_79 = W*in
   wire signed [14:0] m142_79;
   assign m142_79 =15'b0;

   // m142_80 = W*in
   wire signed [14:0] m142_80;
   assign m142_80 =15'b0;

   // m142_81 = W*in
   wire signed [14:0] m142_81;
   assign m142_81 =15'b0;

   // m142_82 = W*in
   wire signed [14:0] m142_82;
   assign m142_82 =15'b0;

   // m142_83 = W*in
   wire signed [14:0] m142_83;
   assign m142_83 =15'b0;

   // m142_84 = W*in
   wire signed [14:0] m142_84;
   assign m142_84 =15'b0;

   // m142_85 = W*in
   wire signed [14:0] m142_85;
   assign m142_85 =15'b0;

   // m142_86 = W*in
   wire signed [14:0] m142_86;
   assign m142_86 =15'b0;

   // m142_87 = W*in
   wire signed [14:0] m142_87;
   assign m142_87 =15'b0;

   // m142_88 = W*in
   wire signed [14:0] m142_88;
   assign m142_88 ={ {3{neg142[14]}} , neg142[14:3] };

   // m142_89 = W*in
   wire signed [14:0] m142_89;
   assign m142_89 =15'b0;

   // m142_90 = W*in
   wire signed [14:0] m142_90;
   assign m142_90 =15'b0;

   // m142_91 = W*in
   wire signed [14:0] m142_91;
   assign m142_91 =15'b0;

   // m142_92 = W*in
   wire signed [14:0] m142_92;
   assign m142_92 =15'b0;

   // m142_93 = W*in
   wire signed [14:0] m142_93;
   assign m142_93 =15'b0;

   // m142_94 = W*in
   wire signed [14:0] m142_94;
   assign m142_94 =15'b0;

   // m142_95 = W*in
   wire signed [14:0] m142_95;
   assign m142_95 =15'b0;

   // m142_96 = W*in
   wire signed [14:0] m142_96;
   assign m142_96 =15'b0;

   // m142_97 = W*in
   wire signed [14:0] m142_97;
   assign m142_97 =15'b0;

   // m142_98 = W*in
   wire signed [14:0] m142_98;
   assign m142_98 =15'b0;

   // m142_99 = W*in
   wire signed [14:0] m142_99;
   assign m142_99 =15'b0;

   // m142_100 = W*in
   wire signed [14:0] m142_100;
   assign m142_100 =15'b0;

   // m143_1 = W*in
   wire signed [14:0] m143_1;
   assign m143_1 =15'b0;

   // m143_2 = W*in
   wire signed [14:0] m143_2;
   assign m143_2 =15'b0;

   // m143_3 = W*in
   wire signed [14:0] m143_3;
   assign m143_3 =15'b0;

   // m143_4 = W*in
   wire signed [14:0] m143_4;
   assign m143_4 =15'b0;

   // m143_5 = W*in
   wire signed [14:0] m143_5;
   assign m143_5 =15'b0;

   // m143_6 = W*in
   wire signed [14:0] m143_6;
   assign m143_6 =15'b0;

   // m143_7 = W*in
   wire signed [14:0] m143_7;
   assign m143_7 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_8 = W*in
   wire signed [14:0] m143_8;
   assign m143_8 =15'b0;

   // m143_9 = W*in
   wire signed [14:0] m143_9;
   assign m143_9 =15'b0;

   // m143_10 = W*in
   wire signed [14:0] m143_10;
   assign m143_10 =15'b0;

   // m143_11 = W*in
   wire signed [14:0] m143_11;
   assign m143_11 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_12 = W*in
   wire signed [14:0] m143_12;
   assign m143_12 =15'b0;

   // m143_13 = W*in
   wire signed [14:0] m143_13;
   assign m143_13 =15'b0;

   // m143_14 = W*in
   wire signed [14:0] m143_14;
   assign m143_14 ={ {3{in143[14]}} , in143[14:3] };

   // m143_15 = W*in
   wire signed [14:0] m143_15;
   assign m143_15 =15'b0;

   // m143_16 = W*in
   wire signed [14:0] m143_16;
   assign m143_16 =15'b0;

   // m143_17 = W*in
   wire signed [14:0] m143_17;
   assign m143_17 =15'b0;

   // m143_18 = W*in
   wire signed [14:0] m143_18;
   assign m143_18 =15'b0;

   // m143_19 = W*in
   wire signed [14:0] m143_19;
   assign m143_19 =15'b0;

   // m143_20 = W*in
   wire signed [14:0] m143_20;
   assign m143_20 =15'b0;

   // m143_21 = W*in
   wire signed [14:0] m143_21;
   assign m143_21 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_22 = W*in
   wire signed [14:0] m143_22;
   assign m143_22 =15'b0;

   // m143_23 = W*in
   wire signed [14:0] m143_23;
   assign m143_23 =15'b0;

   // m143_24 = W*in
   wire signed [14:0] m143_24;
   assign m143_24 =15'b0;

   // m143_25 = W*in
   wire signed [14:0] m143_25;
   assign m143_25 ={ {4{neg143[14]}} , neg143[14:4] };

   // m143_26 = W*in
   wire signed [14:0] m143_26;
   assign m143_26 =15'b0;

   // m143_27 = W*in
   wire signed [14:0] m143_27;
   assign m143_27 =15'b0;

   // m143_28 = W*in
   wire signed [14:0] m143_28;
   assign m143_28 =15'b0;

   // m143_29 = W*in
   wire signed [14:0] m143_29;
   assign m143_29 =15'b0;

   // m143_30 = W*in
   wire signed [14:0] m143_30;
   assign m143_30 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_31 = W*in
   wire signed [14:0] m143_31;
   assign m143_31 =15'b0;

   // m143_32 = W*in
   wire signed [14:0] m143_32;
   assign m143_32 =15'b0;

   // m143_33 = W*in
   wire signed [14:0] m143_33;
   assign m143_33 =15'b0;

   // m143_34 = W*in
   wire signed [14:0] m143_34;
   assign m143_34 =15'b0;

   // m143_35 = W*in
   wire signed [14:0] m143_35;
   assign m143_35 =15'b0;

   // m143_36 = W*in
   wire signed [14:0] m143_36;
   assign m143_36 =15'b0;

   // m143_37 = W*in
   wire signed [14:0] m143_37;
   assign m143_37 ={ {3{in143[14]}} , in143[14:3] };

   // m143_38 = W*in
   wire signed [14:0] m143_38;
   assign m143_38 ={ {3{in143[14]}} , in143[14:3] };

   // m143_39 = W*in
   wire signed [14:0] m143_39;
   assign m143_39 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_40 = W*in
   wire signed [14:0] m143_40;
   assign m143_40 =15'b0;

   // m143_41 = W*in
   wire signed [14:0] m143_41;
   assign m143_41 =15'b0;

   // m143_42 = W*in
   wire signed [14:0] m143_42;
   assign m143_42 =15'b0;

   // m143_43 = W*in
   wire signed [14:0] m143_43;
   assign m143_43 =15'b0;

   // m143_44 = W*in
   wire signed [14:0] m143_44;
   assign m143_44 =15'b0;

   // m143_45 = W*in
   wire signed [14:0] m143_45;
   assign m143_45 =15'b0;

   // m143_46 = W*in
   wire signed [14:0] m143_46;
   assign m143_46 ={ {3{in143[14]}} , in143[14:3] };

   // m143_47 = W*in
   wire signed [14:0] m143_47;
   assign m143_47 =15'b0;

   // m143_48 = W*in
   wire signed [14:0] m143_48;
   assign m143_48 =15'b0;

   // m143_49 = W*in
   wire signed [14:0] m143_49;
   assign m143_49 =15'b0;

   // m143_50 = W*in
   wire signed [14:0] m143_50;
   assign m143_50 =15'b0;

   // m143_51 = W*in
   wire signed [14:0] m143_51;
   assign m143_51 =15'b0;

   // m143_52 = W*in
   wire signed [14:0] m143_52;
   assign m143_52 =15'b0;

   // m143_53 = W*in
   wire signed [14:0] m143_53;
   assign m143_53 =15'b0;

   // m143_54 = W*in
   wire signed [14:0] m143_54;
   assign m143_54 =15'b0;

   // m143_55 = W*in
   wire signed [14:0] m143_55;
   assign m143_55 =15'b0;

   // m143_56 = W*in
   wire signed [14:0] m143_56;
   assign m143_56 =15'b0;

   // m143_57 = W*in
   wire signed [14:0] m143_57;
   assign m143_57 =15'b0;

   // m143_58 = W*in
   wire signed [14:0] m143_58;
   assign m143_58 =15'b0;

   // m143_59 = W*in
   wire signed [14:0] m143_59;
   assign m143_59 =15'b0;

   // m143_60 = W*in
   wire signed [14:0] m143_60;
   assign m143_60 =15'b0;

   // m143_61 = W*in
   wire signed [14:0] m143_61;
   assign m143_61 =15'b0;

   // m143_62 = W*in
   wire signed [14:0] m143_62;
   assign m143_62 =15'b0;

   // m143_63 = W*in
   wire signed [14:0] m143_63;
   assign m143_63 =15'b0;

   // m143_64 = W*in
   wire signed [14:0] m143_64;
   assign m143_64 =15'b0;

   // m143_65 = W*in
   wire signed [14:0] m143_65;
   assign m143_65 =15'b0;

   // m143_66 = W*in
   wire signed [14:0] m143_66;
   assign m143_66 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_67 = W*in
   wire signed [14:0] m143_67;
   assign m143_67 =15'b0;

   // m143_68 = W*in
   wire signed [14:0] m143_68;
   assign m143_68 =15'b0;

   // m143_69 = W*in
   wire signed [14:0] m143_69;
   assign m143_69 =15'b0;

   // m143_70 = W*in
   wire signed [14:0] m143_70;
   assign m143_70 =15'b0;

   // m143_71 = W*in
   wire signed [14:0] m143_71;
   assign m143_71 =15'b0;

   // m143_72 = W*in
   wire signed [14:0] m143_72;
   assign m143_72 =15'b0;

   // m143_73 = W*in
   wire signed [14:0] m143_73;
   assign m143_73 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_74 = W*in
   wire signed [14:0] m143_74;
   assign m143_74 =15'b0;

   // m143_75 = W*in
   wire signed [14:0] m143_75;
   assign m143_75 ={ {3{in143[14]}} , in143[14:3] };

   // m143_76 = W*in
   wire signed [14:0] m143_76;
   assign m143_76 =15'b0;

   // m143_77 = W*in
   wire signed [14:0] m143_77;
   assign m143_77 =15'b0;

   // m143_78 = W*in
   wire signed [14:0] m143_78;
   assign m143_78 =15'b0;

   // m143_79 = W*in
   wire signed [14:0] m143_79;
   assign m143_79 =15'b0;

   // m143_80 = W*in
   wire signed [14:0] m143_80;
   assign m143_80 =15'b0;

   // m143_81 = W*in
   wire signed [14:0] m143_81;
   assign m143_81 ={ {3{in143[14]}} , in143[14:3] };

   // m143_82 = W*in
   wire signed [14:0] m143_82;
   assign m143_82 =15'b0;

   // m143_83 = W*in
   wire signed [14:0] m143_83;
   assign m143_83 =15'b0;

   // m143_84 = W*in
   wire signed [14:0] m143_84;
   assign m143_84 =15'b0;

   // m143_85 = W*in
   wire signed [14:0] m143_85;
   assign m143_85 ={ {3{in143[14]}} , in143[14:3] };

   // m143_86 = W*in
   wire signed [14:0] m143_86;
   assign m143_86 =15'b0;

   // m143_87 = W*in
   wire signed [14:0] m143_87;
   assign m143_87 =15'b0;

   // m143_88 = W*in
   wire signed [14:0] m143_88;
   assign m143_88 =15'b0;

   // m143_89 = W*in
   wire signed [14:0] m143_89;
   assign m143_89 =15'b0;

   // m143_90 = W*in
   wire signed [14:0] m143_90;
   assign m143_90 =15'b0;

   // m143_91 = W*in
   wire signed [14:0] m143_91;
   assign m143_91 =15'b0;

   // m143_92 = W*in
   wire signed [14:0] m143_92;
   assign m143_92 =15'b0;

   // m143_93 = W*in
   wire signed [14:0] m143_93;
   assign m143_93 ={ {3{in143[14]}} , in143[14:3] };

   // m143_94 = W*in
   wire signed [14:0] m143_94;
   assign m143_94 =15'b0;

   // m143_95 = W*in
   wire signed [14:0] m143_95;
   assign m143_95 =15'b0;

   // m143_96 = W*in
   wire signed [14:0] m143_96;
   assign m143_96 =15'b0;

   // m143_97 = W*in
   wire signed [14:0] m143_97;
   assign m143_97 =15'b0;

   // m143_98 = W*in
   wire signed [14:0] m143_98;
   assign m143_98 ={ {3{neg143[14]}} , neg143[14:3] };

   // m143_99 = W*in
   wire signed [14:0] m143_99;
   assign m143_99 ={ {3{in143[14]}} , in143[14:3] };

   // m143_100 = W*in
   wire signed [14:0] m143_100;
   assign m143_100 ={ {3{in143[14]}} , in143[14:3] };

   // m144_1 = W*in
   wire signed [14:0] m144_1;
   assign m144_1 =15'b0;

   // m144_2 = W*in
   wire signed [14:0] m144_2;
   assign m144_2 ={ {3{in144[14]}} , in144[14:3] };

   // m144_3 = W*in
   wire signed [14:0] m144_3;
   assign m144_3 =15'b0;

   // m144_4 = W*in
   wire signed [14:0] m144_4;
   assign m144_4 =15'b0;

   // m144_5 = W*in
   wire signed [14:0] m144_5;
   assign m144_5 =15'b0;

   // m144_6 = W*in
   wire signed [14:0] m144_6;
   assign m144_6 =15'b0;

   // m144_7 = W*in
   wire signed [14:0] m144_7;
   assign m144_7 =15'b0;

   // m144_8 = W*in
   wire signed [14:0] m144_8;
   assign m144_8 =15'b0;

   // m144_9 = W*in
   wire signed [14:0] m144_9;
   assign m144_9 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_10 = W*in
   wire signed [14:0] m144_10;
   assign m144_10 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_11 = W*in
   wire signed [14:0] m144_11;
   assign m144_11 =15'b0;

   // m144_12 = W*in
   wire signed [14:0] m144_12;
   assign m144_12 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_13 = W*in
   wire signed [14:0] m144_13;
   assign m144_13 ={ {3{in144[14]}} , in144[14:3] };

   // m144_14 = W*in
   wire signed [14:0] m144_14;
   assign m144_14 =15'b0;

   // m144_15 = W*in
   wire signed [14:0] m144_15;
   assign m144_15 =15'b0;

   // m144_16 = W*in
   wire signed [14:0] m144_16;
   assign m144_16 =15'b0;

   // m144_17 = W*in
   wire signed [14:0] m144_17;
   assign m144_17 =15'b0;

   // m144_18 = W*in
   wire signed [14:0] m144_18;
   assign m144_18 ={ {2{in144[14]}} , in144[14:2] };

   // m144_19 = W*in
   wire signed [14:0] m144_19;
   assign m144_19 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_20 = W*in
   wire signed [14:0] m144_20;
   assign m144_20 =15'b0;

   // m144_21 = W*in
   wire signed [14:0] m144_21;
   assign m144_21 =15'b0;

   // m144_22 = W*in
   wire signed [14:0] m144_22;
   assign m144_22 =15'b0;

   // m144_23 = W*in
   wire signed [14:0] m144_23;
   assign m144_23 =15'b0;

   // m144_24 = W*in
   wire signed [14:0] m144_24;
   assign m144_24 =15'b0;

   // m144_25 = W*in
   wire signed [14:0] m144_25;
   assign m144_25 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_26 = W*in
   wire signed [14:0] m144_26;
   assign m144_26 =15'b0;

   // m144_27 = W*in
   wire signed [14:0] m144_27;
   assign m144_27 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_28 = W*in
   wire signed [14:0] m144_28;
   assign m144_28 ={ {2{in144[14]}} , in144[14:2] };

   // m144_29 = W*in
   wire signed [14:0] m144_29;
   assign m144_29 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_30 = W*in
   wire signed [14:0] m144_30;
   assign m144_30 =15'b0;

   // m144_31 = W*in
   wire signed [14:0] m144_31;
   assign m144_31 =15'b0;

   // m144_32 = W*in
   wire signed [14:0] m144_32;
   assign m144_32 =15'b0;

   // m144_33 = W*in
   wire signed [14:0] m144_33;
   assign m144_33 ={ {4{in144[14]}} , in144[14:4] };

   // m144_34 = W*in
   wire signed [14:0] m144_34;
   assign m144_34 =15'b0;

   // m144_35 = W*in
   wire signed [14:0] m144_35;
   assign m144_35 =15'b0;

   // m144_36 = W*in
   wire signed [14:0] m144_36;
   assign m144_36 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_37 = W*in
   wire signed [14:0] m144_37;
   assign m144_37 =15'b0;

   // m144_38 = W*in
   wire signed [14:0] m144_38;
   assign m144_38 =15'b0;

   // m144_39 = W*in
   wire signed [14:0] m144_39;
   assign m144_39 =15'b0;

   // m144_40 = W*in
   wire signed [14:0] m144_40;
   assign m144_40 ={ {3{in144[14]}} , in144[14:3] };

   // m144_41 = W*in
   wire signed [14:0] m144_41;
   assign m144_41 =15'b0;

   // m144_42 = W*in
   wire signed [14:0] m144_42;
   assign m144_42 =15'b0;

   // m144_43 = W*in
   wire signed [14:0] m144_43;
   assign m144_43 =15'b0;

   // m144_44 = W*in
   wire signed [14:0] m144_44;
   assign m144_44 =15'b0;

   // m144_45 = W*in
   wire signed [14:0] m144_45;
   assign m144_45 ={ {4{in144[14]}} , in144[14:4] };

   // m144_46 = W*in
   wire signed [14:0] m144_46;
   assign m144_46 ={ {4{neg144[14]}} , neg144[14:4] };

   // m144_47 = W*in
   wire signed [14:0] m144_47;
   assign m144_47 =15'b0;

   // m144_48 = W*in
   wire signed [14:0] m144_48;
   assign m144_48 ={ {3{in144[14]}} , in144[14:3] };

   // m144_49 = W*in
   wire signed [14:0] m144_49;
   assign m144_49 =15'b0;

   // m144_50 = W*in
   wire signed [14:0] m144_50;
   assign m144_50 =15'b0;

   // m144_51 = W*in
   wire signed [14:0] m144_51;
   assign m144_51 =15'b0;

   // m144_52 = W*in
   wire signed [14:0] m144_52;
   assign m144_52 =15'b0;

   // m144_53 = W*in
   wire signed [14:0] m144_53;
   assign m144_53 =15'b0;

   // m144_54 = W*in
   wire signed [14:0] m144_54;
   assign m144_54 =15'b0;

   // m144_55 = W*in
   wire signed [14:0] m144_55;
   assign m144_55 ={ {3{in144[14]}} , in144[14:3] };

   // m144_56 = W*in
   wire signed [14:0] m144_56;
   assign m144_56 ={ {3{in144[14]}} , in144[14:3] };

   // m144_57 = W*in
   wire signed [14:0] m144_57;
   assign m144_57 =15'b0;

   // m144_58 = W*in
   wire signed [14:0] m144_58;
   assign m144_58 =15'b0;

   // m144_59 = W*in
   wire signed [14:0] m144_59;
   assign m144_59 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_60 = W*in
   wire signed [14:0] m144_60;
   assign m144_60 =15'b0;

   // m144_61 = W*in
   wire signed [14:0] m144_61;
   assign m144_61 =15'b0;

   // m144_62 = W*in
   wire signed [14:0] m144_62;
   assign m144_62 =15'b0;

   // m144_63 = W*in
   wire signed [14:0] m144_63;
   assign m144_63 =15'b0;

   // m144_64 = W*in
   wire signed [14:0] m144_64;
   assign m144_64 =15'b0;

   // m144_65 = W*in
   wire signed [14:0] m144_65;
   assign m144_65 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_66 = W*in
   wire signed [14:0] m144_66;
   assign m144_66 =15'b0;

   // m144_67 = W*in
   wire signed [14:0] m144_67;
   assign m144_67 =15'b0;

   // m144_68 = W*in
   wire signed [14:0] m144_68;
   assign m144_68 =15'b0;

   // m144_69 = W*in
   wire signed [14:0] m144_69;
   assign m144_69 ={ {4{neg144[14]}} , neg144[14:4] };

   // m144_70 = W*in
   wire signed [14:0] m144_70;
   assign m144_70 =15'b0;

   // m144_71 = W*in
   wire signed [14:0] m144_71;
   assign m144_71 =15'b0;

   // m144_72 = W*in
   wire signed [14:0] m144_72;
   assign m144_72 =15'b0;

   // m144_73 = W*in
   wire signed [14:0] m144_73;
   assign m144_73 =15'b0;

   // m144_74 = W*in
   wire signed [14:0] m144_74;
   assign m144_74 =15'b0;

   // m144_75 = W*in
   wire signed [14:0] m144_75;
   assign m144_75 =15'b0;

   // m144_76 = W*in
   wire signed [14:0] m144_76;
   assign m144_76 =15'b0;

   // m144_77 = W*in
   wire signed [14:0] m144_77;
   assign m144_77 =15'b0;

   // m144_78 = W*in
   wire signed [14:0] m144_78;
   assign m144_78 =15'b0;

   // m144_79 = W*in
   wire signed [14:0] m144_79;
   assign m144_79 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_80 = W*in
   wire signed [14:0] m144_80;
   assign m144_80 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_81 = W*in
   wire signed [14:0] m144_81;
   assign m144_81 =15'b0;

   // m144_82 = W*in
   wire signed [14:0] m144_82;
   assign m144_82 =15'b0;

   // m144_83 = W*in
   wire signed [14:0] m144_83;
   assign m144_83 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_84 = W*in
   wire signed [14:0] m144_84;
   assign m144_84 =15'b0;

   // m144_85 = W*in
   wire signed [14:0] m144_85;
   assign m144_85 =15'b0;

   // m144_86 = W*in
   wire signed [14:0] m144_86;
   assign m144_86 =15'b0;

   // m144_87 = W*in
   wire signed [14:0] m144_87;
   assign m144_87 =15'b0;

   // m144_88 = W*in
   wire signed [14:0] m144_88;
   assign m144_88 =15'b0;

   // m144_89 = W*in
   wire signed [14:0] m144_89;
   assign m144_89 =15'b0;

   // m144_90 = W*in
   wire signed [14:0] m144_90;
   assign m144_90 ={ {3{in144[14]}} , in144[14:3] };

   // m144_91 = W*in
   wire signed [14:0] m144_91;
   assign m144_91 =15'b0;

   // m144_92 = W*in
   wire signed [14:0] m144_92;
   assign m144_92 ={ {3{neg144[14]}} , neg144[14:3] };

   // m144_93 = W*in
   wire signed [14:0] m144_93;
   assign m144_93 =15'b0;

   // m144_94 = W*in
   wire signed [14:0] m144_94;
   assign m144_94 ={ {3{in144[14]}} , in144[14:3] };

   // m144_95 = W*in
   wire signed [14:0] m144_95;
   assign m144_95 =15'b0;

   // m144_96 = W*in
   wire signed [14:0] m144_96;
   assign m144_96 =15'b0;

   // m144_97 = W*in
   wire signed [14:0] m144_97;
   assign m144_97 =15'b0;

   // m144_98 = W*in
   wire signed [14:0] m144_98;
   assign m144_98 =15'b0;

   // m144_99 = W*in
   wire signed [14:0] m144_99;
   assign m144_99 =15'b0;

   // m144_100 = W*in
   wire signed [14:0] m144_100;
   assign m144_100 =15'b0;

   // m145_1 = W*in
   wire signed [14:0] m145_1;
   assign m145_1 =15'b0;

   // m145_2 = W*in
   wire signed [14:0] m145_2;
   assign m145_2 =15'b0;

   // m145_3 = W*in
   wire signed [14:0] m145_3;
   assign m145_3 ={ {3{in145[14]}} , in145[14:3] };

   // m145_4 = W*in
   wire signed [14:0] m145_4;
   assign m145_4 =15'b0;

   // m145_5 = W*in
   wire signed [14:0] m145_5;
   assign m145_5 ={ {3{neg145[14]}} , neg145[14:3] };

   // m145_6 = W*in
   wire signed [14:0] m145_6;
   assign m145_6 =15'b0;

   // m145_7 = W*in
   wire signed [14:0] m145_7;
   assign m145_7 =15'b0;

   // m145_8 = W*in
   wire signed [14:0] m145_8;
   assign m145_8 ={ {3{in145[14]}} , in145[14:3] };

   // m145_9 = W*in
   wire signed [14:0] m145_9;
   assign m145_9 =15'b0;

   // m145_10 = W*in
   wire signed [14:0] m145_10;
   assign m145_10 =15'b0;

   // m145_11 = W*in
   wire signed [14:0] m145_11;
   assign m145_11 =15'b0;

   // m145_12 = W*in
   wire signed [14:0] m145_12;
   assign m145_12 =15'b0;

   // m145_13 = W*in
   wire signed [14:0] m145_13;
   assign m145_13 =15'b0;

   // m145_14 = W*in
   wire signed [14:0] m145_14;
   assign m145_14 =15'b0;

   // m145_15 = W*in
   wire signed [14:0] m145_15;
   assign m145_15 =15'b0;

   // m145_16 = W*in
   wire signed [14:0] m145_16;
   assign m145_16 =15'b0;

   // m145_17 = W*in
   wire signed [14:0] m145_17;
   assign m145_17 =15'b0;

   // m145_18 = W*in
   wire signed [14:0] m145_18;
   assign m145_18 =15'b0;

   // m145_19 = W*in
   wire signed [14:0] m145_19;
   assign m145_19 =15'b0;

   // m145_20 = W*in
   wire signed [14:0] m145_20;
   assign m145_20 =15'b0;

   // m145_21 = W*in
   wire signed [14:0] m145_21;
   assign m145_21 =15'b0;

   // m145_22 = W*in
   wire signed [14:0] m145_22;
   assign m145_22 =15'b0;

   // m145_23 = W*in
   wire signed [14:0] m145_23;
   assign m145_23 =15'b0;

   // m145_24 = W*in
   wire signed [14:0] m145_24;
   assign m145_24 =15'b0;

   // m145_25 = W*in
   wire signed [14:0] m145_25;
   assign m145_25 =15'b0;

   // m145_26 = W*in
   wire signed [14:0] m145_26;
   assign m145_26 =15'b0;

   // m145_27 = W*in
   wire signed [14:0] m145_27;
   assign m145_27 =15'b0;

   // m145_28 = W*in
   wire signed [14:0] m145_28;
   assign m145_28 =15'b0;

   // m145_29 = W*in
   wire signed [14:0] m145_29;
   assign m145_29 ={ {4{in145[14]}} , in145[14:4] };

   // m145_30 = W*in
   wire signed [14:0] m145_30;
   assign m145_30 =15'b0;

   // m145_31 = W*in
   wire signed [14:0] m145_31;
   assign m145_31 ={ {3{in145[14]}} , in145[14:3] };

   // m145_32 = W*in
   wire signed [14:0] m145_32;
   assign m145_32 =15'b0;

   // m145_33 = W*in
   wire signed [14:0] m145_33;
   assign m145_33 =15'b0;

   // m145_34 = W*in
   wire signed [14:0] m145_34;
   assign m145_34 =15'b0;

   // m145_35 = W*in
   wire signed [14:0] m145_35;
   assign m145_35 =15'b0;

   // m145_36 = W*in
   wire signed [14:0] m145_36;
   assign m145_36 =15'b0;

   // m145_37 = W*in
   wire signed [14:0] m145_37;
   assign m145_37 =15'b0;

   // m145_38 = W*in
   wire signed [14:0] m145_38;
   assign m145_38 =15'b0;

   // m145_39 = W*in
   wire signed [14:0] m145_39;
   assign m145_39 =15'b0;

   // m145_40 = W*in
   wire signed [14:0] m145_40;
   assign m145_40 =15'b0;

   // m145_41 = W*in
   wire signed [14:0] m145_41;
   assign m145_41 =15'b0;

   // m145_42 = W*in
   wire signed [14:0] m145_42;
   assign m145_42 =15'b0;

   // m145_43 = W*in
   wire signed [14:0] m145_43;
   assign m145_43 =15'b0;

   // m145_44 = W*in
   wire signed [14:0] m145_44;
   assign m145_44 =15'b0;

   // m145_45 = W*in
   wire signed [14:0] m145_45;
   assign m145_45 =15'b0;

   // m145_46 = W*in
   wire signed [14:0] m145_46;
   assign m145_46 =15'b0;

   // m145_47 = W*in
   wire signed [14:0] m145_47;
   assign m145_47 =15'b0;

   // m145_48 = W*in
   wire signed [14:0] m145_48;
   assign m145_48 =15'b0;

   // m145_49 = W*in
   wire signed [14:0] m145_49;
   assign m145_49 ={ {3{neg145[14]}} , neg145[14:3] };

   // m145_50 = W*in
   wire signed [14:0] m145_50;
   assign m145_50 =15'b0;

   // m145_51 = W*in
   wire signed [14:0] m145_51;
   assign m145_51 =15'b0;

   // m145_52 = W*in
   wire signed [14:0] m145_52;
   assign m145_52 ={ {3{in145[14]}} , in145[14:3] };

   // m145_53 = W*in
   wire signed [14:0] m145_53;
   assign m145_53 =15'b0;

   // m145_54 = W*in
   wire signed [14:0] m145_54;
   assign m145_54 =15'b0;

   // m145_55 = W*in
   wire signed [14:0] m145_55;
   assign m145_55 ={ {3{neg145[14]}} , neg145[14:3] };

   // m145_56 = W*in
   wire signed [14:0] m145_56;
   assign m145_56 =15'b0;

   // m145_57 = W*in
   wire signed [14:0] m145_57;
   assign m145_57 =15'b0;

   // m145_58 = W*in
   wire signed [14:0] m145_58;
   assign m145_58 =15'b0;

   // m145_59 = W*in
   wire signed [14:0] m145_59;
   assign m145_59 =15'b0;

   // m145_60 = W*in
   wire signed [14:0] m145_60;
   assign m145_60 ={ {3{in145[14]}} , in145[14:3] };

   // m145_61 = W*in
   wire signed [14:0] m145_61;
   assign m145_61 =15'b0;

   // m145_62 = W*in
   wire signed [14:0] m145_62;
   assign m145_62 =15'b0;

   // m145_63 = W*in
   wire signed [14:0] m145_63;
   assign m145_63 =15'b0;

   // m145_64 = W*in
   wire signed [14:0] m145_64;
   assign m145_64 =15'b0;

   // m145_65 = W*in
   wire signed [14:0] m145_65;
   assign m145_65 =15'b0;

   // m145_66 = W*in
   wire signed [14:0] m145_66;
   assign m145_66 =15'b0;

   // m145_67 = W*in
   wire signed [14:0] m145_67;
   assign m145_67 =15'b0;

   // m145_68 = W*in
   wire signed [14:0] m145_68;
   assign m145_68 =15'b0;

   // m145_69 = W*in
   wire signed [14:0] m145_69;
   assign m145_69 ={ {4{in145[14]}} , in145[14:4] };

   // m145_70 = W*in
   wire signed [14:0] m145_70;
   assign m145_70 =15'b0;

   // m145_71 = W*in
   wire signed [14:0] m145_71;
   assign m145_71 =15'b0;

   // m145_72 = W*in
   wire signed [14:0] m145_72;
   assign m145_72 =15'b0;

   // m145_73 = W*in
   wire signed [14:0] m145_73;
   assign m145_73 =15'b0;

   // m145_74 = W*in
   wire signed [14:0] m145_74;
   assign m145_74 =15'b0;

   // m145_75 = W*in
   wire signed [14:0] m145_75;
   assign m145_75 =15'b0;

   // m145_76 = W*in
   wire signed [14:0] m145_76;
   assign m145_76 =15'b0;

   // m145_77 = W*in
   wire signed [14:0] m145_77;
   assign m145_77 ={ {3{in145[14]}} , in145[14:3] };

   // m145_78 = W*in
   wire signed [14:0] m145_78;
   assign m145_78 =15'b0;

   // m145_79 = W*in
   wire signed [14:0] m145_79;
   assign m145_79 =15'b0;

   // m145_80 = W*in
   wire signed [14:0] m145_80;
   assign m145_80 =15'b0;

   // m145_81 = W*in
   wire signed [14:0] m145_81;
   assign m145_81 =15'b0;

   // m145_82 = W*in
   wire signed [14:0] m145_82;
   assign m145_82 =15'b0;

   // m145_83 = W*in
   wire signed [14:0] m145_83;
   assign m145_83 =15'b0;

   // m145_84 = W*in
   wire signed [14:0] m145_84;
   assign m145_84 =15'b0;

   // m145_85 = W*in
   wire signed [14:0] m145_85;
   assign m145_85 =15'b0;

   // m145_86 = W*in
   wire signed [14:0] m145_86;
   assign m145_86 ={ {3{neg145[14]}} , neg145[14:3] };

   // m145_87 = W*in
   wire signed [14:0] m145_87;
   assign m145_87 ={ {3{neg145[14]}} , neg145[14:3] };

   // m145_88 = W*in
   wire signed [14:0] m145_88;
   assign m145_88 =15'b0;

   // m145_89 = W*in
   wire signed [14:0] m145_89;
   assign m145_89 =15'b0;

   // m145_90 = W*in
   wire signed [14:0] m145_90;
   assign m145_90 =15'b0;

   // m145_91 = W*in
   wire signed [14:0] m145_91;
   assign m145_91 =15'b0;

   // m145_92 = W*in
   wire signed [14:0] m145_92;
   assign m145_92 =15'b0;

   // m145_93 = W*in
   wire signed [14:0] m145_93;
   assign m145_93 =15'b0;

   // m145_94 = W*in
   wire signed [14:0] m145_94;
   assign m145_94 =15'b0;

   // m145_95 = W*in
   wire signed [14:0] m145_95;
   assign m145_95 =15'b0;

   // m145_96 = W*in
   wire signed [14:0] m145_96;
   assign m145_96 =15'b0;

   // m145_97 = W*in
   wire signed [14:0] m145_97;
   assign m145_97 =15'b0;

   // m145_98 = W*in
   wire signed [14:0] m145_98;
   assign m145_98 =15'b0;

   // m145_99 = W*in
   wire signed [14:0] m145_99;
   assign m145_99 =15'b0;

   // m145_100 = W*in
   wire signed [14:0] m145_100;
   assign m145_100 =15'b0;

   // m146_1 = W*in
   wire signed [14:0] m146_1;
   assign m146_1 =15'b0;

   // m146_2 = W*in
   wire signed [14:0] m146_2;
   assign m146_2 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_3 = W*in
   wire signed [14:0] m146_3;
   assign m146_3 =15'b0;

   // m146_4 = W*in
   wire signed [14:0] m146_4;
   assign m146_4 =15'b0;

   // m146_5 = W*in
   wire signed [14:0] m146_5;
   assign m146_5 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_6 = W*in
   wire signed [14:0] m146_6;
   assign m146_6 =15'b0;

   // m146_7 = W*in
   wire signed [14:0] m146_7;
   assign m146_7 =15'b0;

   // m146_8 = W*in
   wire signed [14:0] m146_8;
   assign m146_8 ={ {3{in146[14]}} , in146[14:3] };

   // m146_9 = W*in
   wire signed [14:0] m146_9;
   assign m146_9 =15'b0;

   // m146_10 = W*in
   wire signed [14:0] m146_10;
   assign m146_10 =15'b0;

   // m146_11 = W*in
   wire signed [14:0] m146_11;
   assign m146_11 =15'b0;

   // m146_12 = W*in
   wire signed [14:0] m146_12;
   assign m146_12 =15'b0;

   // m146_13 = W*in
   wire signed [14:0] m146_13;
   assign m146_13 =15'b0;

   // m146_14 = W*in
   wire signed [14:0] m146_14;
   assign m146_14 =15'b0;

   // m146_15 = W*in
   wire signed [14:0] m146_15;
   assign m146_15 =15'b0;

   // m146_16 = W*in
   wire signed [14:0] m146_16;
   assign m146_16 =15'b0;

   // m146_17 = W*in
   wire signed [14:0] m146_17;
   assign m146_17 =15'b0;

   // m146_18 = W*in
   wire signed [14:0] m146_18;
   assign m146_18 =15'b0;

   // m146_19 = W*in
   wire signed [14:0] m146_19;
   assign m146_19 =15'b0;

   // m146_20 = W*in
   wire signed [14:0] m146_20;
   assign m146_20 =15'b0;

   // m146_21 = W*in
   wire signed [14:0] m146_21;
   assign m146_21 ={ {4{in146[14]}} , in146[14:4] };

   // m146_22 = W*in
   wire signed [14:0] m146_22;
   assign m146_22 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_23 = W*in
   wire signed [14:0] m146_23;
   assign m146_23 =15'b0;

   // m146_24 = W*in
   wire signed [14:0] m146_24;
   assign m146_24 =15'b0;

   // m146_25 = W*in
   wire signed [14:0] m146_25;
   assign m146_25 ={ {2{in146[14]}} , in146[14:2] };

   // m146_26 = W*in
   wire signed [14:0] m146_26;
   assign m146_26 ={ {4{in146[14]}} , in146[14:4] };

   // m146_27 = W*in
   wire signed [14:0] m146_27;
   assign m146_27 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_28 = W*in
   wire signed [14:0] m146_28;
   assign m146_28 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_29 = W*in
   wire signed [14:0] m146_29;
   assign m146_29 ={ {4{in146[14]}} , in146[14:4] };

   // m146_30 = W*in
   wire signed [14:0] m146_30;
   assign m146_30 =15'b0;

   // m146_31 = W*in
   wire signed [14:0] m146_31;
   assign m146_31 ={ {4{in146[14]}} , in146[14:4] };

   // m146_32 = W*in
   wire signed [14:0] m146_32;
   assign m146_32 ={ {4{in146[14]}} , in146[14:4] };

   // m146_33 = W*in
   wire signed [14:0] m146_33;
   assign m146_33 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_34 = W*in
   wire signed [14:0] m146_34;
   assign m146_34 =15'b0;

   // m146_35 = W*in
   wire signed [14:0] m146_35;
   assign m146_35 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_36 = W*in
   wire signed [14:0] m146_36;
   assign m146_36 =15'b0;

   // m146_37 = W*in
   wire signed [14:0] m146_37;
   assign m146_37 =15'b0;

   // m146_38 = W*in
   wire signed [14:0] m146_38;
   assign m146_38 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_39 = W*in
   wire signed [14:0] m146_39;
   assign m146_39 =15'b0;

   // m146_40 = W*in
   wire signed [14:0] m146_40;
   assign m146_40 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_41 = W*in
   wire signed [14:0] m146_41;
   assign m146_41 =15'b0;

   // m146_42 = W*in
   wire signed [14:0] m146_42;
   assign m146_42 =15'b0;

   // m146_43 = W*in
   wire signed [14:0] m146_43;
   assign m146_43 =15'b0;

   // m146_44 = W*in
   wire signed [14:0] m146_44;
   assign m146_44 =15'b0;

   // m146_45 = W*in
   wire signed [14:0] m146_45;
   assign m146_45 =15'b0;

   // m146_46 = W*in
   wire signed [14:0] m146_46;
   assign m146_46 =15'b0;

   // m146_47 = W*in
   wire signed [14:0] m146_47;
   assign m146_47 =15'b0;

   // m146_48 = W*in
   wire signed [14:0] m146_48;
   assign m146_48 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_49 = W*in
   wire signed [14:0] m146_49;
   assign m146_49 =15'b0;

   // m146_50 = W*in
   wire signed [14:0] m146_50;
   assign m146_50 =15'b0;

   // m146_51 = W*in
   wire signed [14:0] m146_51;
   assign m146_51 =15'b0;

   // m146_52 = W*in
   wire signed [14:0] m146_52;
   assign m146_52 =15'b0;

   // m146_53 = W*in
   wire signed [14:0] m146_53;
   assign m146_53 =15'b0;

   // m146_54 = W*in
   wire signed [14:0] m146_54;
   assign m146_54 =15'b0;

   // m146_55 = W*in
   wire signed [14:0] m146_55;
   assign m146_55 =15'b0;

   // m146_56 = W*in
   wire signed [14:0] m146_56;
   assign m146_56 =15'b0;

   // m146_57 = W*in
   wire signed [14:0] m146_57;
   assign m146_57 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_58 = W*in
   wire signed [14:0] m146_58;
   assign m146_58 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_59 = W*in
   wire signed [14:0] m146_59;
   assign m146_59 ={ {4{in146[14]}} , in146[14:4] };

   // m146_60 = W*in
   wire signed [14:0] m146_60;
   assign m146_60 =15'b0;

   // m146_61 = W*in
   wire signed [14:0] m146_61;
   assign m146_61 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_62 = W*in
   wire signed [14:0] m146_62;
   assign m146_62 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_63 = W*in
   wire signed [14:0] m146_63;
   assign m146_63 =15'b0;

   // m146_64 = W*in
   wire signed [14:0] m146_64;
   assign m146_64 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_65 = W*in
   wire signed [14:0] m146_65;
   assign m146_65 ={ {4{in146[14]}} , in146[14:4] };

   // m146_66 = W*in
   wire signed [14:0] m146_66;
   assign m146_66 =15'b0;

   // m146_67 = W*in
   wire signed [14:0] m146_67;
   assign m146_67 ={ {4{in146[14]}} , in146[14:4] };

   // m146_68 = W*in
   wire signed [14:0] m146_68;
   assign m146_68 ={ {3{in146[14]}} , in146[14:3] };

   // m146_69 = W*in
   wire signed [14:0] m146_69;
   assign m146_69 ={ {3{in146[14]}} , in146[14:3] };

   // m146_70 = W*in
   wire signed [14:0] m146_70;
   assign m146_70 ={ {4{neg146[14]}} , neg146[14:4] };

   // m146_71 = W*in
   wire signed [14:0] m146_71;
   assign m146_71 =15'b0;

   // m146_72 = W*in
   wire signed [14:0] m146_72;
   assign m146_72 =15'b0;

   // m146_73 = W*in
   wire signed [14:0] m146_73;
   assign m146_73 ={ {3{in146[14]}} , in146[14:3] };

   // m146_74 = W*in
   wire signed [14:0] m146_74;
   assign m146_74 =15'b0;

   // m146_75 = W*in
   wire signed [14:0] m146_75;
   assign m146_75 =15'b0;

   // m146_76 = W*in
   wire signed [14:0] m146_76;
   assign m146_76 =15'b0;

   // m146_77 = W*in
   wire signed [14:0] m146_77;
   assign m146_77 ={ {3{in146[14]}} , in146[14:3] };

   // m146_78 = W*in
   wire signed [14:0] m146_78;
   assign m146_78 =15'b0;

   // m146_79 = W*in
   wire signed [14:0] m146_79;
   assign m146_79 =15'b0;

   // m146_80 = W*in
   wire signed [14:0] m146_80;
   assign m146_80 ={ {3{in146[14]}} , in146[14:3] };

   // m146_81 = W*in
   wire signed [14:0] m146_81;
   assign m146_81 =15'b0;

   // m146_82 = W*in
   wire signed [14:0] m146_82;
   assign m146_82 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_83 = W*in
   wire signed [14:0] m146_83;
   assign m146_83 =15'b0;

   // m146_84 = W*in
   wire signed [14:0] m146_84;
   assign m146_84 =15'b0;

   // m146_85 = W*in
   wire signed [14:0] m146_85;
   assign m146_85 =15'b0;

   // m146_86 = W*in
   wire signed [14:0] m146_86;
   assign m146_86 =15'b0;

   // m146_87 = W*in
   wire signed [14:0] m146_87;
   assign m146_87 =15'b0;

   // m146_88 = W*in
   wire signed [14:0] m146_88;
   assign m146_88 =15'b0;

   // m146_89 = W*in
   wire signed [14:0] m146_89;
   assign m146_89 =15'b0;

   // m146_90 = W*in
   wire signed [14:0] m146_90;
   assign m146_90 =15'b0;

   // m146_91 = W*in
   wire signed [14:0] m146_91;
   assign m146_91 =15'b0;

   // m146_92 = W*in
   wire signed [14:0] m146_92;
   assign m146_92 =15'b0;

   // m146_93 = W*in
   wire signed [14:0] m146_93;
   assign m146_93 =15'b0;

   // m146_94 = W*in
   wire signed [14:0] m146_94;
   assign m146_94 =15'b0;

   // m146_95 = W*in
   wire signed [14:0] m146_95;
   assign m146_95 =15'b0;

   // m146_96 = W*in
   wire signed [14:0] m146_96;
   assign m146_96 ={ {4{in146[14]}} , in146[14:4] };

   // m146_97 = W*in
   wire signed [14:0] m146_97;
   assign m146_97 ={ {3{neg146[14]}} , neg146[14:3] };

   // m146_98 = W*in
   wire signed [14:0] m146_98;
   assign m146_98 =15'b0;

   // m146_99 = W*in
   wire signed [14:0] m146_99;
   assign m146_99 =15'b0;

   // m146_100 = W*in
   wire signed [14:0] m146_100;
   assign m146_100 =15'b0;

   // m147_1 = W*in
   wire signed [14:0] m147_1;
   assign m147_1 ={ {3{in147[14]}} , in147[14:3] };

   // m147_2 = W*in
   wire signed [14:0] m147_2;
   assign m147_2 =15'b0;

   // m147_3 = W*in
   wire signed [14:0] m147_3;
   assign m147_3 =15'b0;

   // m147_4 = W*in
   wire signed [14:0] m147_4;
   assign m147_4 ={ {3{in147[14]}} , in147[14:3] };

   // m147_5 = W*in
   wire signed [14:0] m147_5;
   assign m147_5 =15'b0;

   // m147_6 = W*in
   wire signed [14:0] m147_6;
   assign m147_6 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_7 = W*in
   wire signed [14:0] m147_7;
   assign m147_7 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_8 = W*in
   wire signed [14:0] m147_8;
   assign m147_8 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_9 = W*in
   wire signed [14:0] m147_9;
   assign m147_9 =15'b0;

   // m147_10 = W*in
   wire signed [14:0] m147_10;
   assign m147_10 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_11 = W*in
   wire signed [14:0] m147_11;
   assign m147_11 =15'b0;

   // m147_12 = W*in
   wire signed [14:0] m147_12;
   assign m147_12 =15'b0;

   // m147_13 = W*in
   wire signed [14:0] m147_13;
   assign m147_13 =15'b0;

   // m147_14 = W*in
   wire signed [14:0] m147_14;
   assign m147_14 =15'b0;

   // m147_15 = W*in
   wire signed [14:0] m147_15;
   assign m147_15 =15'b0;

   // m147_16 = W*in
   wire signed [14:0] m147_16;
   assign m147_16 =15'b0;

   // m147_17 = W*in
   wire signed [14:0] m147_17;
   assign m147_17 =15'b0;

   // m147_18 = W*in
   wire signed [14:0] m147_18;
   assign m147_18 =15'b0;

   // m147_19 = W*in
   wire signed [14:0] m147_19;
   assign m147_19 =15'b0;

   // m147_20 = W*in
   wire signed [14:0] m147_20;
   assign m147_20 =15'b0;

   // m147_21 = W*in
   wire signed [14:0] m147_21;
   assign m147_21 =15'b0;

   // m147_22 = W*in
   wire signed [14:0] m147_22;
   assign m147_22 =15'b0;

   // m147_23 = W*in
   wire signed [14:0] m147_23;
   assign m147_23 ={ {3{in147[14]}} , in147[14:3] };

   // m147_24 = W*in
   wire signed [14:0] m147_24;
   assign m147_24 =15'b0;

   // m147_25 = W*in
   wire signed [14:0] m147_25;
   assign m147_25 =15'b0;

   // m147_26 = W*in
   wire signed [14:0] m147_26;
   assign m147_26 =15'b0;

   // m147_27 = W*in
   wire signed [14:0] m147_27;
   assign m147_27 =15'b0;

   // m147_28 = W*in
   wire signed [14:0] m147_28;
   assign m147_28 =15'b0;

   // m147_29 = W*in
   wire signed [14:0] m147_29;
   assign m147_29 =15'b0;

   // m147_30 = W*in
   wire signed [14:0] m147_30;
   assign m147_30 ={ {3{in147[14]}} , in147[14:3] };

   // m147_31 = W*in
   wire signed [14:0] m147_31;
   assign m147_31 =15'b0;

   // m147_32 = W*in
   wire signed [14:0] m147_32;
   assign m147_32 =15'b0;

   // m147_33 = W*in
   wire signed [14:0] m147_33;
   assign m147_33 ={ {4{neg147[14]}} , neg147[14:4] };

   // m147_34 = W*in
   wire signed [14:0] m147_34;
   assign m147_34 =15'b0;

   // m147_35 = W*in
   wire signed [14:0] m147_35;
   assign m147_35 =15'b0;

   // m147_36 = W*in
   wire signed [14:0] m147_36;
   assign m147_36 =15'b0;

   // m147_37 = W*in
   wire signed [14:0] m147_37;
   assign m147_37 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_38 = W*in
   wire signed [14:0] m147_38;
   assign m147_38 ={ {3{in147[14]}} , in147[14:3] };

   // m147_39 = W*in
   wire signed [14:0] m147_39;
   assign m147_39 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_40 = W*in
   wire signed [14:0] m147_40;
   assign m147_40 =15'b0;

   // m147_41 = W*in
   wire signed [14:0] m147_41;
   assign m147_41 ={ {3{in147[14]}} , in147[14:3] };

   // m147_42 = W*in
   wire signed [14:0] m147_42;
   assign m147_42 =15'b0;

   // m147_43 = W*in
   wire signed [14:0] m147_43;
   assign m147_43 ={ {3{in147[14]}} , in147[14:3] };

   // m147_44 = W*in
   wire signed [14:0] m147_44;
   assign m147_44 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_45 = W*in
   wire signed [14:0] m147_45;
   assign m147_45 ={ {3{in147[14]}} , in147[14:3] };

   // m147_46 = W*in
   wire signed [14:0] m147_46;
   assign m147_46 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_47 = W*in
   wire signed [14:0] m147_47;
   assign m147_47 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_48 = W*in
   wire signed [14:0] m147_48;
   assign m147_48 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_49 = W*in
   wire signed [14:0] m147_49;
   assign m147_49 =15'b0;

   // m147_50 = W*in
   wire signed [14:0] m147_50;
   assign m147_50 ={ {3{in147[14]}} , in147[14:3] };

   // m147_51 = W*in
   wire signed [14:0] m147_51;
   assign m147_51 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_52 = W*in
   wire signed [14:0] m147_52;
   assign m147_52 =15'b0;

   // m147_53 = W*in
   wire signed [14:0] m147_53;
   assign m147_53 =15'b0;

   // m147_54 = W*in
   wire signed [14:0] m147_54;
   assign m147_54 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_55 = W*in
   wire signed [14:0] m147_55;
   assign m147_55 ={ {3{in147[14]}} , in147[14:3] };

   // m147_56 = W*in
   wire signed [14:0] m147_56;
   assign m147_56 =15'b0;

   // m147_57 = W*in
   wire signed [14:0] m147_57;
   assign m147_57 =15'b0;

   // m147_58 = W*in
   wire signed [14:0] m147_58;
   assign m147_58 =15'b0;

   // m147_59 = W*in
   wire signed [14:0] m147_59;
   assign m147_59 =15'b0;

   // m147_60 = W*in
   wire signed [14:0] m147_60;
   assign m147_60 ={ {4{neg147[14]}} , neg147[14:4] };

   // m147_61 = W*in
   wire signed [14:0] m147_61;
   assign m147_61 =15'b0;

   // m147_62 = W*in
   wire signed [14:0] m147_62;
   assign m147_62 ={ {3{in147[14]}} , in147[14:3] };

   // m147_63 = W*in
   wire signed [14:0] m147_63;
   assign m147_63 =15'b0;

   // m147_64 = W*in
   wire signed [14:0] m147_64;
   assign m147_64 =15'b0;

   // m147_65 = W*in
   wire signed [14:0] m147_65;
   assign m147_65 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_66 = W*in
   wire signed [14:0] m147_66;
   assign m147_66 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_67 = W*in
   wire signed [14:0] m147_67;
   assign m147_67 ={ {4{in147[14]}} , in147[14:4] };

   // m147_68 = W*in
   wire signed [14:0] m147_68;
   assign m147_68 =15'b0;

   // m147_69 = W*in
   wire signed [14:0] m147_69;
   assign m147_69 =15'b0;

   // m147_70 = W*in
   wire signed [14:0] m147_70;
   assign m147_70 ={ {4{in147[14]}} , in147[14:4] };

   // m147_71 = W*in
   wire signed [14:0] m147_71;
   assign m147_71 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_72 = W*in
   wire signed [14:0] m147_72;
   assign m147_72 =15'b0;

   // m147_73 = W*in
   wire signed [14:0] m147_73;
   assign m147_73 =15'b0;

   // m147_74 = W*in
   wire signed [14:0] m147_74;
   assign m147_74 =15'b0;

   // m147_75 = W*in
   wire signed [14:0] m147_75;
   assign m147_75 ={ {3{in147[14]}} , in147[14:3] };

   // m147_76 = W*in
   wire signed [14:0] m147_76;
   assign m147_76 =15'b0;

   // m147_77 = W*in
   wire signed [14:0] m147_77;
   assign m147_77 =15'b0;

   // m147_78 = W*in
   wire signed [14:0] m147_78;
   assign m147_78 ={ {3{in147[14]}} , in147[14:3] };

   // m147_79 = W*in
   wire signed [14:0] m147_79;
   assign m147_79 =15'b0;

   // m147_80 = W*in
   wire signed [14:0] m147_80;
   assign m147_80 =15'b0;

   // m147_81 = W*in
   wire signed [14:0] m147_81;
   assign m147_81 =15'b0;

   // m147_82 = W*in
   wire signed [14:0] m147_82;
   assign m147_82 =15'b0;

   // m147_83 = W*in
   wire signed [14:0] m147_83;
   assign m147_83 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_84 = W*in
   wire signed [14:0] m147_84;
   assign m147_84 =15'b0;

   // m147_85 = W*in
   wire signed [14:0] m147_85;
   assign m147_85 =15'b0;

   // m147_86 = W*in
   wire signed [14:0] m147_86;
   assign m147_86 =15'b0;

   // m147_87 = W*in
   wire signed [14:0] m147_87;
   assign m147_87 =15'b0;

   // m147_88 = W*in
   wire signed [14:0] m147_88;
   assign m147_88 =15'b0;

   // m147_89 = W*in
   wire signed [14:0] m147_89;
   assign m147_89 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_90 = W*in
   wire signed [14:0] m147_90;
   assign m147_90 =15'b0;

   // m147_91 = W*in
   wire signed [14:0] m147_91;
   assign m147_91 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_92 = W*in
   wire signed [14:0] m147_92;
   assign m147_92 =15'b0;

   // m147_93 = W*in
   wire signed [14:0] m147_93;
   assign m147_93 ={ {3{neg147[14]}} , neg147[14:3] };

   // m147_94 = W*in
   wire signed [14:0] m147_94;
   assign m147_94 =15'b0;

   // m147_95 = W*in
   wire signed [14:0] m147_95;
   assign m147_95 =15'b0;

   // m147_96 = W*in
   wire signed [14:0] m147_96;
   assign m147_96 =15'b0;

   // m147_97 = W*in
   wire signed [14:0] m147_97;
   assign m147_97 ={ {3{in147[14]}} , in147[14:3] };

   // m147_98 = W*in
   wire signed [14:0] m147_98;
   assign m147_98 =15'b0;

   // m147_99 = W*in
   wire signed [14:0] m147_99;
   assign m147_99 =15'b0;

   // m147_100 = W*in
   wire signed [14:0] m147_100;
   assign m147_100 ={ {3{neg147[14]}} , neg147[14:3] };

   // m148_1 = W*in
   wire signed [14:0] m148_1;
   assign m148_1 =15'b0;

   // m148_2 = W*in
   wire signed [14:0] m148_2;
   assign m148_2 =15'b0;

   // m148_3 = W*in
   wire signed [14:0] m148_3;
   assign m148_3 =15'b0;

   // m148_4 = W*in
   wire signed [14:0] m148_4;
   assign m148_4 =15'b0;

   // m148_5 = W*in
   wire signed [14:0] m148_5;
   assign m148_5 ={ {4{neg148[14]}} , neg148[14:4] };

   // m148_6 = W*in
   wire signed [14:0] m148_6;
   assign m148_6 =15'b0;

   // m148_7 = W*in
   wire signed [14:0] m148_7;
   assign m148_7 =15'b0;

   // m148_8 = W*in
   wire signed [14:0] m148_8;
   assign m148_8 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_9 = W*in
   wire signed [14:0] m148_9;
   assign m148_9 =15'b0;

   // m148_10 = W*in
   wire signed [14:0] m148_10;
   assign m148_10 =15'b0;

   // m148_11 = W*in
   wire signed [14:0] m148_11;
   assign m148_11 ={ {3{in148[14]}} , in148[14:3] };

   // m148_12 = W*in
   wire signed [14:0] m148_12;
   assign m148_12 ={ {3{in148[14]}} , in148[14:3] };

   // m148_13 = W*in
   wire signed [14:0] m148_13;
   assign m148_13 =15'b0;

   // m148_14 = W*in
   wire signed [14:0] m148_14;
   assign m148_14 =15'b0;

   // m148_15 = W*in
   wire signed [14:0] m148_15;
   assign m148_15 =15'b0;

   // m148_16 = W*in
   wire signed [14:0] m148_16;
   assign m148_16 =15'b0;

   // m148_17 = W*in
   wire signed [14:0] m148_17;
   assign m148_17 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_18 = W*in
   wire signed [14:0] m148_18;
   assign m148_18 =15'b0;

   // m148_19 = W*in
   wire signed [14:0] m148_19;
   assign m148_19 =15'b0;

   // m148_20 = W*in
   wire signed [14:0] m148_20;
   assign m148_20 =15'b0;

   // m148_21 = W*in
   wire signed [14:0] m148_21;
   assign m148_21 =15'b0;

   // m148_22 = W*in
   wire signed [14:0] m148_22;
   assign m148_22 =15'b0;

   // m148_23 = W*in
   wire signed [14:0] m148_23;
   assign m148_23 ={ {4{in148[14]}} , in148[14:4] };

   // m148_24 = W*in
   wire signed [14:0] m148_24;
   assign m148_24 =15'b0;

   // m148_25 = W*in
   wire signed [14:0] m148_25;
   assign m148_25 =15'b0;

   // m148_26 = W*in
   wire signed [14:0] m148_26;
   assign m148_26 =15'b0;

   // m148_27 = W*in
   wire signed [14:0] m148_27;
   assign m148_27 =15'b0;

   // m148_28 = W*in
   wire signed [14:0] m148_28;
   assign m148_28 =15'b0;

   // m148_29 = W*in
   wire signed [14:0] m148_29;
   assign m148_29 =15'b0;

   // m148_30 = W*in
   wire signed [14:0] m148_30;
   assign m148_30 ={ {3{in148[14]}} , in148[14:3] };

   // m148_31 = W*in
   wire signed [14:0] m148_31;
   assign m148_31 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_32 = W*in
   wire signed [14:0] m148_32;
   assign m148_32 =15'b0;

   // m148_33 = W*in
   wire signed [14:0] m148_33;
   assign m148_33 =15'b0;

   // m148_34 = W*in
   wire signed [14:0] m148_34;
   assign m148_34 ={ {2{in148[14]}} , in148[14:2] };

   // m148_35 = W*in
   wire signed [14:0] m148_35;
   assign m148_35 =15'b0;

   // m148_36 = W*in
   wire signed [14:0] m148_36;
   assign m148_36 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_37 = W*in
   wire signed [14:0] m148_37;
   assign m148_37 =15'b0;

   // m148_38 = W*in
   wire signed [14:0] m148_38;
   assign m148_38 =15'b0;

   // m148_39 = W*in
   wire signed [14:0] m148_39;
   assign m148_39 =15'b0;

   // m148_40 = W*in
   wire signed [14:0] m148_40;
   assign m148_40 =15'b0;

   // m148_41 = W*in
   wire signed [14:0] m148_41;
   assign m148_41 =15'b0;

   // m148_42 = W*in
   wire signed [14:0] m148_42;
   assign m148_42 =15'b0;

   // m148_43 = W*in
   wire signed [14:0] m148_43;
   assign m148_43 =15'b0;

   // m148_44 = W*in
   wire signed [14:0] m148_44;
   assign m148_44 ={ {4{neg148[14]}} , neg148[14:4] };

   // m148_45 = W*in
   wire signed [14:0] m148_45;
   assign m148_45 ={ {4{in148[14]}} , in148[14:4] };

   // m148_46 = W*in
   wire signed [14:0] m148_46;
   assign m148_46 =15'b0;

   // m148_47 = W*in
   wire signed [14:0] m148_47;
   assign m148_47 =15'b0;

   // m148_48 = W*in
   wire signed [14:0] m148_48;
   assign m148_48 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_49 = W*in
   wire signed [14:0] m148_49;
   assign m148_49 =15'b0;

   // m148_50 = W*in
   wire signed [14:0] m148_50;
   assign m148_50 =15'b0;

   // m148_51 = W*in
   wire signed [14:0] m148_51;
   assign m148_51 =15'b0;

   // m148_52 = W*in
   wire signed [14:0] m148_52;
   assign m148_52 =15'b0;

   // m148_53 = W*in
   wire signed [14:0] m148_53;
   assign m148_53 =15'b0;

   // m148_54 = W*in
   wire signed [14:0] m148_54;
   assign m148_54 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_55 = W*in
   wire signed [14:0] m148_55;
   assign m148_55 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_56 = W*in
   wire signed [14:0] m148_56;
   assign m148_56 =15'b0;

   // m148_57 = W*in
   wire signed [14:0] m148_57;
   assign m148_57 ={ {4{in148[14]}} , in148[14:4] };

   // m148_58 = W*in
   wire signed [14:0] m148_58;
   assign m148_58 =15'b0;

   // m148_59 = W*in
   wire signed [14:0] m148_59;
   assign m148_59 =15'b0;

   // m148_60 = W*in
   wire signed [14:0] m148_60;
   assign m148_60 =15'b0;

   // m148_61 = W*in
   wire signed [14:0] m148_61;
   assign m148_61 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_62 = W*in
   wire signed [14:0] m148_62;
   assign m148_62 =15'b0;

   // m148_63 = W*in
   wire signed [14:0] m148_63;
   assign m148_63 =15'b0;

   // m148_64 = W*in
   wire signed [14:0] m148_64;
   assign m148_64 =15'b0;

   // m148_65 = W*in
   wire signed [14:0] m148_65;
   assign m148_65 =15'b0;

   // m148_66 = W*in
   wire signed [14:0] m148_66;
   assign m148_66 =15'b0;

   // m148_67 = W*in
   wire signed [14:0] m148_67;
   assign m148_67 =15'b0;

   // m148_68 = W*in
   wire signed [14:0] m148_68;
   assign m148_68 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_69 = W*in
   wire signed [14:0] m148_69;
   assign m148_69 =15'b0;

   // m148_70 = W*in
   wire signed [14:0] m148_70;
   assign m148_70 =15'b0;

   // m148_71 = W*in
   wire signed [14:0] m148_71;
   assign m148_71 =15'b0;

   // m148_72 = W*in
   wire signed [14:0] m148_72;
   assign m148_72 =15'b0;

   // m148_73 = W*in
   wire signed [14:0] m148_73;
   assign m148_73 =15'b0;

   // m148_74 = W*in
   wire signed [14:0] m148_74;
   assign m148_74 =15'b0;

   // m148_75 = W*in
   wire signed [14:0] m148_75;
   assign m148_75 =15'b0;

   // m148_76 = W*in
   wire signed [14:0] m148_76;
   assign m148_76 =15'b0;

   // m148_77 = W*in
   wire signed [14:0] m148_77;
   assign m148_77 =15'b0;

   // m148_78 = W*in
   wire signed [14:0] m148_78;
   assign m148_78 =15'b0;

   // m148_79 = W*in
   wire signed [14:0] m148_79;
   assign m148_79 =15'b0;

   // m148_80 = W*in
   wire signed [14:0] m148_80;
   assign m148_80 =15'b0;

   // m148_81 = W*in
   wire signed [14:0] m148_81;
   assign m148_81 =15'b0;

   // m148_82 = W*in
   wire signed [14:0] m148_82;
   assign m148_82 =15'b0;

   // m148_83 = W*in
   wire signed [14:0] m148_83;
   assign m148_83 =15'b0;

   // m148_84 = W*in
   wire signed [14:0] m148_84;
   assign m148_84 =15'b0;

   // m148_85 = W*in
   wire signed [14:0] m148_85;
   assign m148_85 =15'b0;

   // m148_86 = W*in
   wire signed [14:0] m148_86;
   assign m148_86 =15'b0;

   // m148_87 = W*in
   wire signed [14:0] m148_87;
   assign m148_87 =15'b0;

   // m148_88 = W*in
   wire signed [14:0] m148_88;
   assign m148_88 ={ {3{in148[14]}} , in148[14:3] };

   // m148_89 = W*in
   wire signed [14:0] m148_89;
   assign m148_89 ={ {3{neg148[14]}} , neg148[14:3] };

   // m148_90 = W*in
   wire signed [14:0] m148_90;
   assign m148_90 =15'b0;

   // m148_91 = W*in
   wire signed [14:0] m148_91;
   assign m148_91 =15'b0;

   // m148_92 = W*in
   wire signed [14:0] m148_92;
   assign m148_92 =15'b0;

   // m148_93 = W*in
   wire signed [14:0] m148_93;
   assign m148_93 =15'b0;

   // m148_94 = W*in
   wire signed [14:0] m148_94;
   assign m148_94 =15'b0;

   // m148_95 = W*in
   wire signed [14:0] m148_95;
   assign m148_95 =15'b0;

   // m148_96 = W*in
   wire signed [14:0] m148_96;
   assign m148_96 ={ {4{in148[14]}} , in148[14:4] };

   // m148_97 = W*in
   wire signed [14:0] m148_97;
   assign m148_97 =15'b0;

   // m148_98 = W*in
   wire signed [14:0] m148_98;
   assign m148_98 =15'b0;

   // m148_99 = W*in
   wire signed [14:0] m148_99;
   assign m148_99 =15'b0;

   // m148_100 = W*in
   wire signed [14:0] m148_100;
   assign m148_100 =15'b0;

   // m149_1 = W*in
   wire signed [14:0] m149_1;
   assign m149_1 =15'b0;

   // m149_2 = W*in
   wire signed [14:0] m149_2;
   assign m149_2 ={ {4{neg149[14]}} , neg149[14:4] };

   // m149_3 = W*in
   wire signed [14:0] m149_3;
   assign m149_3 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_4 = W*in
   wire signed [14:0] m149_4;
   assign m149_4 =15'b0;

   // m149_5 = W*in
   wire signed [14:0] m149_5;
   assign m149_5 =15'b0;

   // m149_6 = W*in
   wire signed [14:0] m149_6;
   assign m149_6 =15'b0;

   // m149_7 = W*in
   wire signed [14:0] m149_7;
   assign m149_7 =15'b0;

   // m149_8 = W*in
   wire signed [14:0] m149_8;
   assign m149_8 =15'b0;

   // m149_9 = W*in
   wire signed [14:0] m149_9;
   assign m149_9 =15'b0;

   // m149_10 = W*in
   wire signed [14:0] m149_10;
   assign m149_10 ={ {3{in149[14]}} , in149[14:3] };

   // m149_11 = W*in
   wire signed [14:0] m149_11;
   assign m149_11 =15'b0;

   // m149_12 = W*in
   wire signed [14:0] m149_12;
   assign m149_12 =15'b0;

   // m149_13 = W*in
   wire signed [14:0] m149_13;
   assign m149_13 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_14 = W*in
   wire signed [14:0] m149_14;
   assign m149_14 =15'b0;

   // m149_15 = W*in
   wire signed [14:0] m149_15;
   assign m149_15 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_16 = W*in
   wire signed [14:0] m149_16;
   assign m149_16 ={ {3{in149[14]}} , in149[14:3] };

   // m149_17 = W*in
   wire signed [14:0] m149_17;
   assign m149_17 =15'b0;

   // m149_18 = W*in
   wire signed [14:0] m149_18;
   assign m149_18 ={ {4{neg149[14]}} , neg149[14:4] };

   // m149_19 = W*in
   wire signed [14:0] m149_19;
   assign m149_19 ={ {3{in149[14]}} , in149[14:3] };

   // m149_20 = W*in
   wire signed [14:0] m149_20;
   assign m149_20 ={ {4{neg149[14]}} , neg149[14:4] };

   // m149_21 = W*in
   wire signed [14:0] m149_21;
   assign m149_21 =15'b0;

   // m149_22 = W*in
   wire signed [14:0] m149_22;
   assign m149_22 =15'b0;

   // m149_23 = W*in
   wire signed [14:0] m149_23;
   assign m149_23 =15'b0;

   // m149_24 = W*in
   wire signed [14:0] m149_24;
   assign m149_24 =15'b0;

   // m149_25 = W*in
   wire signed [14:0] m149_25;
   assign m149_25 =15'b0;

   // m149_26 = W*in
   wire signed [14:0] m149_26;
   assign m149_26 ={ {3{in149[14]}} , in149[14:3] };

   // m149_27 = W*in
   wire signed [14:0] m149_27;
   assign m149_27 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_28 = W*in
   wire signed [14:0] m149_28;
   assign m149_28 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_29 = W*in
   wire signed [14:0] m149_29;
   assign m149_29 =15'b0;

   // m149_30 = W*in
   wire signed [14:0] m149_30;
   assign m149_30 =15'b0;

   // m149_31 = W*in
   wire signed [14:0] m149_31;
   assign m149_31 ={ {3{in149[14]}} , in149[14:3] };

   // m149_32 = W*in
   wire signed [14:0] m149_32;
   assign m149_32 ={ {4{in149[14]}} , in149[14:4] };

   // m149_33 = W*in
   wire signed [14:0] m149_33;
   assign m149_33 =15'b0;

   // m149_34 = W*in
   wire signed [14:0] m149_34;
   assign m149_34 =15'b0;

   // m149_35 = W*in
   wire signed [14:0] m149_35;
   assign m149_35 =15'b0;

   // m149_36 = W*in
   wire signed [14:0] m149_36;
   assign m149_36 =15'b0;

   // m149_37 = W*in
   wire signed [14:0] m149_37;
   assign m149_37 =15'b0;

   // m149_38 = W*in
   wire signed [14:0] m149_38;
   assign m149_38 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_39 = W*in
   wire signed [14:0] m149_39;
   assign m149_39 ={ {3{in149[14]}} , in149[14:3] };

   // m149_40 = W*in
   wire signed [14:0] m149_40;
   assign m149_40 =15'b0;

   // m149_41 = W*in
   wire signed [14:0] m149_41;
   assign m149_41 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_42 = W*in
   wire signed [14:0] m149_42;
   assign m149_42 =15'b0;

   // m149_43 = W*in
   wire signed [14:0] m149_43;
   assign m149_43 =15'b0;

   // m149_44 = W*in
   wire signed [14:0] m149_44;
   assign m149_44 =15'b0;

   // m149_45 = W*in
   wire signed [14:0] m149_45;
   assign m149_45 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_46 = W*in
   wire signed [14:0] m149_46;
   assign m149_46 ={ {3{in149[14]}} , in149[14:3] };

   // m149_47 = W*in
   wire signed [14:0] m149_47;
   assign m149_47 ={ {2{in149[14]}} , in149[14:2] };

   // m149_48 = W*in
   wire signed [14:0] m149_48;
   assign m149_48 =15'b0;

   // m149_49 = W*in
   wire signed [14:0] m149_49;
   assign m149_49 =15'b0;

   // m149_50 = W*in
   wire signed [14:0] m149_50;
   assign m149_50 =15'b0;

   // m149_51 = W*in
   wire signed [14:0] m149_51;
   assign m149_51 =15'b0;

   // m149_52 = W*in
   wire signed [14:0] m149_52;
   assign m149_52 =15'b0;

   // m149_53 = W*in
   wire signed [14:0] m149_53;
   assign m149_53 =15'b0;

   // m149_54 = W*in
   wire signed [14:0] m149_54;
   assign m149_54 =15'b0;

   // m149_55 = W*in
   wire signed [14:0] m149_55;
   assign m149_55 =15'b0;

   // m149_56 = W*in
   wire signed [14:0] m149_56;
   assign m149_56 =15'b0;

   // m149_57 = W*in
   wire signed [14:0] m149_57;
   assign m149_57 =15'b0;

   // m149_58 = W*in
   wire signed [14:0] m149_58;
   assign m149_58 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_59 = W*in
   wire signed [14:0] m149_59;
   assign m149_59 =15'b0;

   // m149_60 = W*in
   wire signed [14:0] m149_60;
   assign m149_60 ={ {4{neg149[14]}} , neg149[14:4] };

   // m149_61 = W*in
   wire signed [14:0] m149_61;
   assign m149_61 =15'b0;

   // m149_62 = W*in
   wire signed [14:0] m149_62;
   assign m149_62 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_63 = W*in
   wire signed [14:0] m149_63;
   assign m149_63 =15'b0;

   // m149_64 = W*in
   wire signed [14:0] m149_64;
   assign m149_64 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_65 = W*in
   wire signed [14:0] m149_65;
   assign m149_65 ={ {3{in149[14]}} , in149[14:3] };

   // m149_66 = W*in
   wire signed [14:0] m149_66;
   assign m149_66 =15'b0;

   // m149_67 = W*in
   wire signed [14:0] m149_67;
   assign m149_67 =15'b0;

   // m149_68 = W*in
   wire signed [14:0] m149_68;
   assign m149_68 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_69 = W*in
   wire signed [14:0] m149_69;
   assign m149_69 =15'b0;

   // m149_70 = W*in
   wire signed [14:0] m149_70;
   assign m149_70 =15'b0;

   // m149_71 = W*in
   wire signed [14:0] m149_71;
   assign m149_71 =15'b0;

   // m149_72 = W*in
   wire signed [14:0] m149_72;
   assign m149_72 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_73 = W*in
   wire signed [14:0] m149_73;
   assign m149_73 =15'b0;

   // m149_74 = W*in
   wire signed [14:0] m149_74;
   assign m149_74 ={ {4{neg149[14]}} , neg149[14:4] };

   // m149_75 = W*in
   wire signed [14:0] m149_75;
   assign m149_75 =15'b0;

   // m149_76 = W*in
   wire signed [14:0] m149_76;
   assign m149_76 =15'b0;

   // m149_77 = W*in
   wire signed [14:0] m149_77;
   assign m149_77 =15'b0;

   // m149_78 = W*in
   wire signed [14:0] m149_78;
   assign m149_78 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_79 = W*in
   wire signed [14:0] m149_79;
   assign m149_79 ={ {3{in149[14]}} , in149[14:3] };

   // m149_80 = W*in
   wire signed [14:0] m149_80;
   assign m149_80 =15'b0;

   // m149_81 = W*in
   wire signed [14:0] m149_81;
   assign m149_81 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_82 = W*in
   wire signed [14:0] m149_82;
   assign m149_82 =15'b0;

   // m149_83 = W*in
   wire signed [14:0] m149_83;
   assign m149_83 =15'b0;

   // m149_84 = W*in
   wire signed [14:0] m149_84;
   assign m149_84 =15'b0;

   // m149_85 = W*in
   wire signed [14:0] m149_85;
   assign m149_85 =15'b0;

   // m149_86 = W*in
   wire signed [14:0] m149_86;
   assign m149_86 =15'b0;

   // m149_87 = W*in
   wire signed [14:0] m149_87;
   assign m149_87 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_88 = W*in
   wire signed [14:0] m149_88;
   assign m149_88 =15'b0;

   // m149_89 = W*in
   wire signed [14:0] m149_89;
   assign m149_89 =15'b0;

   // m149_90 = W*in
   wire signed [14:0] m149_90;
   assign m149_90 =15'b0;

   // m149_91 = W*in
   wire signed [14:0] m149_91;
   assign m149_91 =15'b0;

   // m149_92 = W*in
   wire signed [14:0] m149_92;
   assign m149_92 =15'b0;

   // m149_93 = W*in
   wire signed [14:0] m149_93;
   assign m149_93 =15'b0;

   // m149_94 = W*in
   wire signed [14:0] m149_94;
   assign m149_94 =15'b0;

   // m149_95 = W*in
   wire signed [14:0] m149_95;
   assign m149_95 =15'b0;

   // m149_96 = W*in
   wire signed [14:0] m149_96;
   assign m149_96 ={ {3{neg149[14]}} , neg149[14:3] };

   // m149_97 = W*in
   wire signed [14:0] m149_97;
   assign m149_97 =15'b0;

   // m149_98 = W*in
   wire signed [14:0] m149_98;
   assign m149_98 =15'b0;

   // m149_99 = W*in
   wire signed [14:0] m149_99;
   assign m149_99 =15'b0;

   // m149_100 = W*in
   wire signed [14:0] m149_100;
   assign m149_100 =15'b0;

   // m150_1 = W*in
   wire signed [14:0] m150_1;
   assign m150_1 =15'b0;

   // m150_2 = W*in
   wire signed [14:0] m150_2;
   assign m150_2 =15'b0;

   // m150_3 = W*in
   wire signed [14:0] m150_3;
   assign m150_3 =15'b0;

   // m150_4 = W*in
   wire signed [14:0] m150_4;
   assign m150_4 =15'b0;

   // m150_5 = W*in
   wire signed [14:0] m150_5;
   assign m150_5 =15'b0;

   // m150_6 = W*in
   wire signed [14:0] m150_6;
   assign m150_6 ={ {4{in150[14]}} , in150[14:4] };

   // m150_7 = W*in
   wire signed [14:0] m150_7;
   assign m150_7 =15'b0;

   // m150_8 = W*in
   wire signed [14:0] m150_8;
   assign m150_8 =15'b0;

   // m150_9 = W*in
   wire signed [14:0] m150_9;
   assign m150_9 =15'b0;

   // m150_10 = W*in
   wire signed [14:0] m150_10;
   assign m150_10 =15'b0;

   // m150_11 = W*in
   wire signed [14:0] m150_11;
   assign m150_11 =15'b0;

   // m150_12 = W*in
   wire signed [14:0] m150_12;
   assign m150_12 =15'b0;

   // m150_13 = W*in
   wire signed [14:0] m150_13;
   assign m150_13 =15'b0;

   // m150_14 = W*in
   wire signed [14:0] m150_14;
   assign m150_14 ={ {4{neg150[14]}} , neg150[14:4] };

   // m150_15 = W*in
   wire signed [14:0] m150_15;
   assign m150_15 =15'b0;

   // m150_16 = W*in
   wire signed [14:0] m150_16;
   assign m150_16 ={ {3{neg150[14]}} , neg150[14:3] };

   // m150_17 = W*in
   wire signed [14:0] m150_17;
   assign m150_17 =15'b0;

   // m150_18 = W*in
   wire signed [14:0] m150_18;
   assign m150_18 =15'b0;

   // m150_19 = W*in
   wire signed [14:0] m150_19;
   assign m150_19 =15'b0;

   // m150_20 = W*in
   wire signed [14:0] m150_20;
   assign m150_20 =15'b0;

   // m150_21 = W*in
   wire signed [14:0] m150_21;
   assign m150_21 =15'b0;

   // m150_22 = W*in
   wire signed [14:0] m150_22;
   assign m150_22 =15'b0;

   // m150_23 = W*in
   wire signed [14:0] m150_23;
   assign m150_23 =15'b0;

   // m150_24 = W*in
   wire signed [14:0] m150_24;
   assign m150_24 =15'b0;

   // m150_25 = W*in
   wire signed [14:0] m150_25;
   assign m150_25 =15'b0;

   // m150_26 = W*in
   wire signed [14:0] m150_26;
   assign m150_26 ={ {4{in150[14]}} , in150[14:4] };

   // m150_27 = W*in
   wire signed [14:0] m150_27;
   assign m150_27 =15'b0;

   // m150_28 = W*in
   wire signed [14:0] m150_28;
   assign m150_28 =15'b0;

   // m150_29 = W*in
   wire signed [14:0] m150_29;
   assign m150_29 =15'b0;

   // m150_30 = W*in
   wire signed [14:0] m150_30;
   assign m150_30 =15'b0;

   // m150_31 = W*in
   wire signed [14:0] m150_31;
   assign m150_31 =15'b0;

   // m150_32 = W*in
   wire signed [14:0] m150_32;
   assign m150_32 ={ {3{neg150[14]}} , neg150[14:3] };

   // m150_33 = W*in
   wire signed [14:0] m150_33;
   assign m150_33 =15'b0;

   // m150_34 = W*in
   wire signed [14:0] m150_34;
   assign m150_34 =15'b0;

   // m150_35 = W*in
   wire signed [14:0] m150_35;
   assign m150_35 =15'b0;

   // m150_36 = W*in
   wire signed [14:0] m150_36;
   assign m150_36 =15'b0;

   // m150_37 = W*in
   wire signed [14:0] m150_37;
   assign m150_37 ={ {4{neg150[14]}} , neg150[14:4] };

   // m150_38 = W*in
   wire signed [14:0] m150_38;
   assign m150_38 =15'b0;

   // m150_39 = W*in
   wire signed [14:0] m150_39;
   assign m150_39 =15'b0;

   // m150_40 = W*in
   wire signed [14:0] m150_40;
   assign m150_40 ={ {4{neg150[14]}} , neg150[14:4] };

   // m150_41 = W*in
   wire signed [14:0] m150_41;
   assign m150_41 =15'b0;

   // m150_42 = W*in
   wire signed [14:0] m150_42;
   assign m150_42 ={ {3{neg150[14]}} , neg150[14:3] };

   // m150_43 = W*in
   wire signed [14:0] m150_43;
   assign m150_43 =15'b0;

   // m150_44 = W*in
   wire signed [14:0] m150_44;
   assign m150_44 =15'b0;

   // m150_45 = W*in
   wire signed [14:0] m150_45;
   assign m150_45 =15'b0;

   // m150_46 = W*in
   wire signed [14:0] m150_46;
   assign m150_46 ={ {2{in150[14]}} , in150[14:2] };

   // m150_47 = W*in
   wire signed [14:0] m150_47;
   assign m150_47 =15'b0;

   // m150_48 = W*in
   wire signed [14:0] m150_48;
   assign m150_48 =15'b0;

   // m150_49 = W*in
   wire signed [14:0] m150_49;
   assign m150_49 =15'b0;

   // m150_50 = W*in
   wire signed [14:0] m150_50;
   assign m150_50 =15'b0;

   // m150_51 = W*in
   wire signed [14:0] m150_51;
   assign m150_51 =15'b0;

   // m150_52 = W*in
   wire signed [14:0] m150_52;
   assign m150_52 =15'b0;

   // m150_53 = W*in
   wire signed [14:0] m150_53;
   assign m150_53 =15'b0;

   // m150_54 = W*in
   wire signed [14:0] m150_54;
   assign m150_54 ={ {4{neg150[14]}} , neg150[14:4] };

   // m150_55 = W*in
   wire signed [14:0] m150_55;
   assign m150_55 =15'b0;

   // m150_56 = W*in
   wire signed [14:0] m150_56;
   assign m150_56 =15'b0;

   // m150_57 = W*in
   wire signed [14:0] m150_57;
   assign m150_57 =15'b0;

   // m150_58 = W*in
   wire signed [14:0] m150_58;
   assign m150_58 =15'b0;

   // m150_59 = W*in
   wire signed [14:0] m150_59;
   assign m150_59 ={ {3{in150[14]}} , in150[14:3] };

   // m150_60 = W*in
   wire signed [14:0] m150_60;
   assign m150_60 =15'b0;

   // m150_61 = W*in
   wire signed [14:0] m150_61;
   assign m150_61 ={ {4{in150[14]}} , in150[14:4] };

   // m150_62 = W*in
   wire signed [14:0] m150_62;
   assign m150_62 =15'b0;

   // m150_63 = W*in
   wire signed [14:0] m150_63;
   assign m150_63 =15'b0;

   // m150_64 = W*in
   wire signed [14:0] m150_64;
   assign m150_64 =15'b0;

   // m150_65 = W*in
   wire signed [14:0] m150_65;
   assign m150_65 =15'b0;

   // m150_66 = W*in
   wire signed [14:0] m150_66;
   assign m150_66 =15'b0;

   // m150_67 = W*in
   wire signed [14:0] m150_67;
   assign m150_67 =15'b0;

   // m150_68 = W*in
   wire signed [14:0] m150_68;
   assign m150_68 =15'b0;

   // m150_69 = W*in
   wire signed [14:0] m150_69;
   assign m150_69 ={ {3{neg150[14]}} , neg150[14:3] };

   // m150_70 = W*in
   wire signed [14:0] m150_70;
   assign m150_70 =15'b0;

   // m150_71 = W*in
   wire signed [14:0] m150_71;
   assign m150_71 =15'b0;

   // m150_72 = W*in
   wire signed [14:0] m150_72;
   assign m150_72 =15'b0;

   // m150_73 = W*in
   wire signed [14:0] m150_73;
   assign m150_73 =15'b0;

   // m150_74 = W*in
   wire signed [14:0] m150_74;
   assign m150_74 =15'b0;

   // m150_75 = W*in
   wire signed [14:0] m150_75;
   assign m150_75 =15'b0;

   // m150_76 = W*in
   wire signed [14:0] m150_76;
   assign m150_76 =15'b0;

   // m150_77 = W*in
   wire signed [14:0] m150_77;
   assign m150_77 =15'b0;

   // m150_78 = W*in
   wire signed [14:0] m150_78;
   assign m150_78 =15'b0;

   // m150_79 = W*in
   wire signed [14:0] m150_79;
   assign m150_79 =15'b0;

   // m150_80 = W*in
   wire signed [14:0] m150_80;
   assign m150_80 =15'b0;

   // m150_81 = W*in
   wire signed [14:0] m150_81;
   assign m150_81 ={ {4{in150[14]}} , in150[14:4] };

   // m150_82 = W*in
   wire signed [14:0] m150_82;
   assign m150_82 =15'b0;

   // m150_83 = W*in
   wire signed [14:0] m150_83;
   assign m150_83 =15'b0;

   // m150_84 = W*in
   wire signed [14:0] m150_84;
   assign m150_84 =15'b0;

   // m150_85 = W*in
   wire signed [14:0] m150_85;
   assign m150_85 =15'b0;

   // m150_86 = W*in
   wire signed [14:0] m150_86;
   assign m150_86 =15'b0;

   // m150_87 = W*in
   wire signed [14:0] m150_87;
   assign m150_87 =15'b0;

   // m150_88 = W*in
   wire signed [14:0] m150_88;
   assign m150_88 =15'b0;

   // m150_89 = W*in
   wire signed [14:0] m150_89;
   assign m150_89 =15'b0;

   // m150_90 = W*in
   wire signed [14:0] m150_90;
   assign m150_90 =15'b0;

   // m150_91 = W*in
   wire signed [14:0] m150_91;
   assign m150_91 ={ {4{in150[14]}} , in150[14:4] };

   // m150_92 = W*in
   wire signed [14:0] m150_92;
   assign m150_92 ={ {4{neg150[14]}} , neg150[14:4] };

   // m150_93 = W*in
   wire signed [14:0] m150_93;
   assign m150_93 =15'b0;

   // m150_94 = W*in
   wire signed [14:0] m150_94;
   assign m150_94 =15'b0;

   // m150_95 = W*in
   wire signed [14:0] m150_95;
   assign m150_95 =15'b0;

   // m150_96 = W*in
   wire signed [14:0] m150_96;
   assign m150_96 =15'b0;

   // m150_97 = W*in
   wire signed [14:0] m150_97;
   assign m150_97 =15'b0;

   // m150_98 = W*in
   wire signed [14:0] m150_98;
   assign m150_98 =15'b0;

   // m150_99 = W*in
   wire signed [14:0] m150_99;
   assign m150_99 =15'b0;

   // m150_100 = W*in
   wire signed [14:0] m150_100;
   assign m150_100 =15'b0;

   // m151_1 = W*in
   wire signed [14:0] m151_1;
   assign m151_1 =15'b0;

   // m151_2 = W*in
   wire signed [14:0] m151_2;
   assign m151_2 =15'b0;

   // m151_3 = W*in
   wire signed [14:0] m151_3;
   assign m151_3 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_4 = W*in
   wire signed [14:0] m151_4;
   assign m151_4 ={ {3{in151[14]}} , in151[14:3] };

   // m151_5 = W*in
   wire signed [14:0] m151_5;
   assign m151_5 =15'b0;

   // m151_6 = W*in
   wire signed [14:0] m151_6;
   assign m151_6 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_7 = W*in
   wire signed [14:0] m151_7;
   assign m151_7 =15'b0;

   // m151_8 = W*in
   wire signed [14:0] m151_8;
   assign m151_8 =15'b0;

   // m151_9 = W*in
   wire signed [14:0] m151_9;
   assign m151_9 =15'b0;

   // m151_10 = W*in
   wire signed [14:0] m151_10;
   assign m151_10 =15'b0;

   // m151_11 = W*in
   wire signed [14:0] m151_11;
   assign m151_11 =15'b0;

   // m151_12 = W*in
   wire signed [14:0] m151_12;
   assign m151_12 =15'b0;

   // m151_13 = W*in
   wire signed [14:0] m151_13;
   assign m151_13 =15'b0;

   // m151_14 = W*in
   wire signed [14:0] m151_14;
   assign m151_14 ={ {3{in151[14]}} , in151[14:3] };

   // m151_15 = W*in
   wire signed [14:0] m151_15;
   assign m151_15 =15'b0;

   // m151_16 = W*in
   wire signed [14:0] m151_16;
   assign m151_16 =15'b0;

   // m151_17 = W*in
   wire signed [14:0] m151_17;
   assign m151_17 =15'b0;

   // m151_18 = W*in
   wire signed [14:0] m151_18;
   assign m151_18 =15'b0;

   // m151_19 = W*in
   wire signed [14:0] m151_19;
   assign m151_19 =15'b0;

   // m151_20 = W*in
   wire signed [14:0] m151_20;
   assign m151_20 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_21 = W*in
   wire signed [14:0] m151_21;
   assign m151_21 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_22 = W*in
   wire signed [14:0] m151_22;
   assign m151_22 =15'b0;

   // m151_23 = W*in
   wire signed [14:0] m151_23;
   assign m151_23 =15'b0;

   // m151_24 = W*in
   wire signed [14:0] m151_24;
   assign m151_24 =15'b0;

   // m151_25 = W*in
   wire signed [14:0] m151_25;
   assign m151_25 ={ {4{neg151[14]}} , neg151[14:4] };

   // m151_26 = W*in
   wire signed [14:0] m151_26;
   assign m151_26 =15'b0;

   // m151_27 = W*in
   wire signed [14:0] m151_27;
   assign m151_27 =15'b0;

   // m151_28 = W*in
   wire signed [14:0] m151_28;
   assign m151_28 =15'b0;

   // m151_29 = W*in
   wire signed [14:0] m151_29;
   assign m151_29 =15'b0;

   // m151_30 = W*in
   wire signed [14:0] m151_30;
   assign m151_30 =15'b0;

   // m151_31 = W*in
   wire signed [14:0] m151_31;
   assign m151_31 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_32 = W*in
   wire signed [14:0] m151_32;
   assign m151_32 ={ {3{in151[14]}} , in151[14:3] };

   // m151_33 = W*in
   wire signed [14:0] m151_33;
   assign m151_33 ={ {3{in151[14]}} , in151[14:3] };

   // m151_34 = W*in
   wire signed [14:0] m151_34;
   assign m151_34 =15'b0;

   // m151_35 = W*in
   wire signed [14:0] m151_35;
   assign m151_35 =15'b0;

   // m151_36 = W*in
   wire signed [14:0] m151_36;
   assign m151_36 =15'b0;

   // m151_37 = W*in
   wire signed [14:0] m151_37;
   assign m151_37 =15'b0;

   // m151_38 = W*in
   wire signed [14:0] m151_38;
   assign m151_38 =15'b0;

   // m151_39 = W*in
   wire signed [14:0] m151_39;
   assign m151_39 =15'b0;

   // m151_40 = W*in
   wire signed [14:0] m151_40;
   assign m151_40 ={ {3{in151[14]}} , in151[14:3] };

   // m151_41 = W*in
   wire signed [14:0] m151_41;
   assign m151_41 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_42 = W*in
   wire signed [14:0] m151_42;
   assign m151_42 ={ {2{in151[14]}} , in151[14:2] };

   // m151_43 = W*in
   wire signed [14:0] m151_43;
   assign m151_43 =15'b0;

   // m151_44 = W*in
   wire signed [14:0] m151_44;
   assign m151_44 =15'b0;

   // m151_45 = W*in
   wire signed [14:0] m151_45;
   assign m151_45 =15'b0;

   // m151_46 = W*in
   wire signed [14:0] m151_46;
   assign m151_46 =15'b0;

   // m151_47 = W*in
   wire signed [14:0] m151_47;
   assign m151_47 =15'b0;

   // m151_48 = W*in
   wire signed [14:0] m151_48;
   assign m151_48 ={ {3{in151[14]}} , in151[14:3] };

   // m151_49 = W*in
   wire signed [14:0] m151_49;
   assign m151_49 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_50 = W*in
   wire signed [14:0] m151_50;
   assign m151_50 =15'b0;

   // m151_51 = W*in
   wire signed [14:0] m151_51;
   assign m151_51 =15'b0;

   // m151_52 = W*in
   wire signed [14:0] m151_52;
   assign m151_52 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_53 = W*in
   wire signed [14:0] m151_53;
   assign m151_53 =15'b0;

   // m151_54 = W*in
   wire signed [14:0] m151_54;
   assign m151_54 =15'b0;

   // m151_55 = W*in
   wire signed [14:0] m151_55;
   assign m151_55 =15'b0;

   // m151_56 = W*in
   wire signed [14:0] m151_56;
   assign m151_56 =15'b0;

   // m151_57 = W*in
   wire signed [14:0] m151_57;
   assign m151_57 ={ {3{in151[14]}} , in151[14:3] };

   // m151_58 = W*in
   wire signed [14:0] m151_58;
   assign m151_58 =15'b0;

   // m151_59 = W*in
   wire signed [14:0] m151_59;
   assign m151_59 =15'b0;

   // m151_60 = W*in
   wire signed [14:0] m151_60;
   assign m151_60 =15'b0;

   // m151_61 = W*in
   wire signed [14:0] m151_61;
   assign m151_61 =15'b0;

   // m151_62 = W*in
   wire signed [14:0] m151_62;
   assign m151_62 =15'b0;

   // m151_63 = W*in
   wire signed [14:0] m151_63;
   assign m151_63 ={ {3{in151[14]}} , in151[14:3] };

   // m151_64 = W*in
   wire signed [14:0] m151_64;
   assign m151_64 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_65 = W*in
   wire signed [14:0] m151_65;
   assign m151_65 =15'b0;

   // m151_66 = W*in
   wire signed [14:0] m151_66;
   assign m151_66 ={ {3{in151[14]}} , in151[14:3] };

   // m151_67 = W*in
   wire signed [14:0] m151_67;
   assign m151_67 =15'b0;

   // m151_68 = W*in
   wire signed [14:0] m151_68;
   assign m151_68 =15'b0;

   // m151_69 = W*in
   wire signed [14:0] m151_69;
   assign m151_69 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_70 = W*in
   wire signed [14:0] m151_70;
   assign m151_70 =15'b0;

   // m151_71 = W*in
   wire signed [14:0] m151_71;
   assign m151_71 =15'b0;

   // m151_72 = W*in
   wire signed [14:0] m151_72;
   assign m151_72 =15'b0;

   // m151_73 = W*in
   wire signed [14:0] m151_73;
   assign m151_73 =15'b0;

   // m151_74 = W*in
   wire signed [14:0] m151_74;
   assign m151_74 ={ {4{neg151[14]}} , neg151[14:4] };

   // m151_75 = W*in
   wire signed [14:0] m151_75;
   assign m151_75 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_76 = W*in
   wire signed [14:0] m151_76;
   assign m151_76 =15'b0;

   // m151_77 = W*in
   wire signed [14:0] m151_77;
   assign m151_77 ={ {4{neg151[14]}} , neg151[14:4] };

   // m151_78 = W*in
   wire signed [14:0] m151_78;
   assign m151_78 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_79 = W*in
   wire signed [14:0] m151_79;
   assign m151_79 ={ {4{neg151[14]}} , neg151[14:4] };

   // m151_80 = W*in
   wire signed [14:0] m151_80;
   assign m151_80 =15'b0;

   // m151_81 = W*in
   wire signed [14:0] m151_81;
   assign m151_81 =15'b0;

   // m151_82 = W*in
   wire signed [14:0] m151_82;
   assign m151_82 ={ {3{in151[14]}} , in151[14:3] };

   // m151_83 = W*in
   wire signed [14:0] m151_83;
   assign m151_83 =15'b0;

   // m151_84 = W*in
   wire signed [14:0] m151_84;
   assign m151_84 =15'b0;

   // m151_85 = W*in
   wire signed [14:0] m151_85;
   assign m151_85 =15'b0;

   // m151_86 = W*in
   wire signed [14:0] m151_86;
   assign m151_86 =15'b0;

   // m151_87 = W*in
   wire signed [14:0] m151_87;
   assign m151_87 =15'b0;

   // m151_88 = W*in
   wire signed [14:0] m151_88;
   assign m151_88 =15'b0;

   // m151_89 = W*in
   wire signed [14:0] m151_89;
   assign m151_89 =15'b0;

   // m151_90 = W*in
   wire signed [14:0] m151_90;
   assign m151_90 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_91 = W*in
   wire signed [14:0] m151_91;
   assign m151_91 =15'b0;

   // m151_92 = W*in
   wire signed [14:0] m151_92;
   assign m151_92 =15'b0;

   // m151_93 = W*in
   wire signed [14:0] m151_93;
   assign m151_93 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_94 = W*in
   wire signed [14:0] m151_94;
   assign m151_94 ={ {4{neg151[14]}} , neg151[14:4] };

   // m151_95 = W*in
   wire signed [14:0] m151_95;
   assign m151_95 =15'b0;

   // m151_96 = W*in
   wire signed [14:0] m151_96;
   assign m151_96 ={ {3{neg151[14]}} , neg151[14:3] };

   // m151_97 = W*in
   wire signed [14:0] m151_97;
   assign m151_97 =15'b0;

   // m151_98 = W*in
   wire signed [14:0] m151_98;
   assign m151_98 =15'b0;

   // m151_99 = W*in
   wire signed [14:0] m151_99;
   assign m151_99 =15'b0;

   // m151_100 = W*in
   wire signed [14:0] m151_100;
   assign m151_100 =15'b0;

   // m152_1 = W*in
   wire signed [14:0] m152_1;
   assign m152_1 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_2 = W*in
   wire signed [14:0] m152_2;
   assign m152_2 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_3 = W*in
   wire signed [14:0] m152_3;
   assign m152_3 =15'b0;

   // m152_4 = W*in
   wire signed [14:0] m152_4;
   assign m152_4 =15'b0;

   // m152_5 = W*in
   wire signed [14:0] m152_5;
   assign m152_5 =15'b0;

   // m152_6 = W*in
   wire signed [14:0] m152_6;
   assign m152_6 =15'b0;

   // m152_7 = W*in
   wire signed [14:0] m152_7;
   assign m152_7 =15'b0;

   // m152_8 = W*in
   wire signed [14:0] m152_8;
   assign m152_8 ={ {3{in152[14]}} , in152[14:3] };

   // m152_9 = W*in
   wire signed [14:0] m152_9;
   assign m152_9 =15'b0;

   // m152_10 = W*in
   wire signed [14:0] m152_10;
   assign m152_10 =15'b0;

   // m152_11 = W*in
   wire signed [14:0] m152_11;
   assign m152_11 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_12 = W*in
   wire signed [14:0] m152_12;
   assign m152_12 =15'b0;

   // m152_13 = W*in
   wire signed [14:0] m152_13;
   assign m152_13 =15'b0;

   // m152_14 = W*in
   wire signed [14:0] m152_14;
   assign m152_14 =15'b0;

   // m152_15 = W*in
   wire signed [14:0] m152_15;
   assign m152_15 =15'b0;

   // m152_16 = W*in
   wire signed [14:0] m152_16;
   assign m152_16 =15'b0;

   // m152_17 = W*in
   wire signed [14:0] m152_17;
   assign m152_17 =15'b0;

   // m152_18 = W*in
   wire signed [14:0] m152_18;
   assign m152_18 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_19 = W*in
   wire signed [14:0] m152_19;
   assign m152_19 =15'b0;

   // m152_20 = W*in
   wire signed [14:0] m152_20;
   assign m152_20 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_21 = W*in
   wire signed [14:0] m152_21;
   assign m152_21 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_22 = W*in
   wire signed [14:0] m152_22;
   assign m152_22 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_23 = W*in
   wire signed [14:0] m152_23;
   assign m152_23 =15'b0;

   // m152_24 = W*in
   wire signed [14:0] m152_24;
   assign m152_24 =15'b0;

   // m152_25 = W*in
   wire signed [14:0] m152_25;
   assign m152_25 =15'b0;

   // m152_26 = W*in
   wire signed [14:0] m152_26;
   assign m152_26 =15'b0;

   // m152_27 = W*in
   wire signed [14:0] m152_27;
   assign m152_27 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_28 = W*in
   wire signed [14:0] m152_28;
   assign m152_28 =15'b0;

   // m152_29 = W*in
   wire signed [14:0] m152_29;
   assign m152_29 =15'b0;

   // m152_30 = W*in
   wire signed [14:0] m152_30;
   assign m152_30 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_31 = W*in
   wire signed [14:0] m152_31;
   assign m152_31 ={ {3{in152[14]}} , in152[14:3] };

   // m152_32 = W*in
   wire signed [14:0] m152_32;
   assign m152_32 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_33 = W*in
   wire signed [14:0] m152_33;
   assign m152_33 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_34 = W*in
   wire signed [14:0] m152_34;
   assign m152_34 =15'b0;

   // m152_35 = W*in
   wire signed [14:0] m152_35;
   assign m152_35 =15'b0;

   // m152_36 = W*in
   wire signed [14:0] m152_36;
   assign m152_36 =15'b0;

   // m152_37 = W*in
   wire signed [14:0] m152_37;
   assign m152_37 ={ {3{in152[14]}} , in152[14:3] };

   // m152_38 = W*in
   wire signed [14:0] m152_38;
   assign m152_38 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_39 = W*in
   wire signed [14:0] m152_39;
   assign m152_39 =15'b0;

   // m152_40 = W*in
   wire signed [14:0] m152_40;
   assign m152_40 =15'b0;

   // m152_41 = W*in
   wire signed [14:0] m152_41;
   assign m152_41 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_42 = W*in
   wire signed [14:0] m152_42;
   assign m152_42 =15'b0;

   // m152_43 = W*in
   wire signed [14:0] m152_43;
   assign m152_43 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_44 = W*in
   wire signed [14:0] m152_44;
   assign m152_44 =15'b0;

   // m152_45 = W*in
   wire signed [14:0] m152_45;
   assign m152_45 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_46 = W*in
   wire signed [14:0] m152_46;
   assign m152_46 =15'b0;

   // m152_47 = W*in
   wire signed [14:0] m152_47;
   assign m152_47 =15'b0;

   // m152_48 = W*in
   wire signed [14:0] m152_48;
   assign m152_48 ={ {4{in152[14]}} , in152[14:4] };

   // m152_49 = W*in
   wire signed [14:0] m152_49;
   assign m152_49 =15'b0;

   // m152_50 = W*in
   wire signed [14:0] m152_50;
   assign m152_50 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_51 = W*in
   wire signed [14:0] m152_51;
   assign m152_51 ={ {3{in152[14]}} , in152[14:3] };

   // m152_52 = W*in
   wire signed [14:0] m152_52;
   assign m152_52 =15'b0;

   // m152_53 = W*in
   wire signed [14:0] m152_53;
   assign m152_53 =15'b0;

   // m152_54 = W*in
   wire signed [14:0] m152_54;
   assign m152_54 ={ {3{in152[14]}} , in152[14:3] };

   // m152_55 = W*in
   wire signed [14:0] m152_55;
   assign m152_55 =15'b0;

   // m152_56 = W*in
   wire signed [14:0] m152_56;
   assign m152_56 =15'b0;

   // m152_57 = W*in
   wire signed [14:0] m152_57;
   assign m152_57 =15'b0;

   // m152_58 = W*in
   wire signed [14:0] m152_58;
   assign m152_58 =15'b0;

   // m152_59 = W*in
   wire signed [14:0] m152_59;
   assign m152_59 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_60 = W*in
   wire signed [14:0] m152_60;
   assign m152_60 =15'b0;

   // m152_61 = W*in
   wire signed [14:0] m152_61;
   assign m152_61 =15'b0;

   // m152_62 = W*in
   wire signed [14:0] m152_62;
   assign m152_62 =15'b0;

   // m152_63 = W*in
   wire signed [14:0] m152_63;
   assign m152_63 ={ {3{in152[14]}} , in152[14:3] };

   // m152_64 = W*in
   wire signed [14:0] m152_64;
   assign m152_64 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_65 = W*in
   wire signed [14:0] m152_65;
   assign m152_65 =15'b0;

   // m152_66 = W*in
   wire signed [14:0] m152_66;
   assign m152_66 ={ {4{in152[14]}} , in152[14:4] };

   // m152_67 = W*in
   wire signed [14:0] m152_67;
   assign m152_67 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_68 = W*in
   wire signed [14:0] m152_68;
   assign m152_68 =15'b0;

   // m152_69 = W*in
   wire signed [14:0] m152_69;
   assign m152_69 =15'b0;

   // m152_70 = W*in
   wire signed [14:0] m152_70;
   assign m152_70 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_71 = W*in
   wire signed [14:0] m152_71;
   assign m152_71 ={ {3{in152[14]}} , in152[14:3] };

   // m152_72 = W*in
   wire signed [14:0] m152_72;
   assign m152_72 =15'b0;

   // m152_73 = W*in
   wire signed [14:0] m152_73;
   assign m152_73 =15'b0;

   // m152_74 = W*in
   wire signed [14:0] m152_74;
   assign m152_74 =15'b0;

   // m152_75 = W*in
   wire signed [14:0] m152_75;
   assign m152_75 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_76 = W*in
   wire signed [14:0] m152_76;
   assign m152_76 =15'b0;

   // m152_77 = W*in
   wire signed [14:0] m152_77;
   assign m152_77 =15'b0;

   // m152_78 = W*in
   wire signed [14:0] m152_78;
   assign m152_78 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_79 = W*in
   wire signed [14:0] m152_79;
   assign m152_79 =15'b0;

   // m152_80 = W*in
   wire signed [14:0] m152_80;
   assign m152_80 ={ {3{in152[14]}} , in152[14:3] };

   // m152_81 = W*in
   wire signed [14:0] m152_81;
   assign m152_81 =15'b0;

   // m152_82 = W*in
   wire signed [14:0] m152_82;
   assign m152_82 =15'b0;

   // m152_83 = W*in
   wire signed [14:0] m152_83;
   assign m152_83 ={ {3{in152[14]}} , in152[14:3] };

   // m152_84 = W*in
   wire signed [14:0] m152_84;
   assign m152_84 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_85 = W*in
   wire signed [14:0] m152_85;
   assign m152_85 =15'b0;

   // m152_86 = W*in
   wire signed [14:0] m152_86;
   assign m152_86 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_87 = W*in
   wire signed [14:0] m152_87;
   assign m152_87 =15'b0;

   // m152_88 = W*in
   wire signed [14:0] m152_88;
   assign m152_88 =15'b0;

   // m152_89 = W*in
   wire signed [14:0] m152_89;
   assign m152_89 ={ {3{in152[14]}} , in152[14:3] };

   // m152_90 = W*in
   wire signed [14:0] m152_90;
   assign m152_90 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_91 = W*in
   wire signed [14:0] m152_91;
   assign m152_91 ={ {3{in152[14]}} , in152[14:3] };

   // m152_92 = W*in
   wire signed [14:0] m152_92;
   assign m152_92 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_93 = W*in
   wire signed [14:0] m152_93;
   assign m152_93 =15'b0;

   // m152_94 = W*in
   wire signed [14:0] m152_94;
   assign m152_94 ={ {4{neg152[14]}} , neg152[14:4] };

   // m152_95 = W*in
   wire signed [14:0] m152_95;
   assign m152_95 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_96 = W*in
   wire signed [14:0] m152_96;
   assign m152_96 =15'b0;

   // m152_97 = W*in
   wire signed [14:0] m152_97;
   assign m152_97 =15'b0;

   // m152_98 = W*in
   wire signed [14:0] m152_98;
   assign m152_98 ={ {3{neg152[14]}} , neg152[14:3] };

   // m152_99 = W*in
   wire signed [14:0] m152_99;
   assign m152_99 =15'b0;

   // m152_100 = W*in
   wire signed [14:0] m152_100;
   assign m152_100 ={ {3{in152[14]}} , in152[14:3] };

   // m153_1 = W*in
   wire signed [14:0] m153_1;
   assign m153_1 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_2 = W*in
   wire signed [14:0] m153_2;
   assign m153_2 =15'b0;

   // m153_3 = W*in
   wire signed [14:0] m153_3;
   assign m153_3 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_4 = W*in
   wire signed [14:0] m153_4;
   assign m153_4 =15'b0;

   // m153_5 = W*in
   wire signed [14:0] m153_5;
   assign m153_5 =15'b0;

   // m153_6 = W*in
   wire signed [14:0] m153_6;
   assign m153_6 =15'b0;

   // m153_7 = W*in
   wire signed [14:0] m153_7;
   assign m153_7 =15'b0;

   // m153_8 = W*in
   wire signed [14:0] m153_8;
   assign m153_8 =15'b0;

   // m153_9 = W*in
   wire signed [14:0] m153_9;
   assign m153_9 =15'b0;

   // m153_10 = W*in
   wire signed [14:0] m153_10;
   assign m153_10 =15'b0;

   // m153_11 = W*in
   wire signed [14:0] m153_11;
   assign m153_11 =15'b0;

   // m153_12 = W*in
   wire signed [14:0] m153_12;
   assign m153_12 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_13 = W*in
   wire signed [14:0] m153_13;
   assign m153_13 =15'b0;

   // m153_14 = W*in
   wire signed [14:0] m153_14;
   assign m153_14 =15'b0;

   // m153_15 = W*in
   wire signed [14:0] m153_15;
   assign m153_15 =15'b0;

   // m153_16 = W*in
   wire signed [14:0] m153_16;
   assign m153_16 =15'b0;

   // m153_17 = W*in
   wire signed [14:0] m153_17;
   assign m153_17 =15'b0;

   // m153_18 = W*in
   wire signed [14:0] m153_18;
   assign m153_18 =15'b0;

   // m153_19 = W*in
   wire signed [14:0] m153_19;
   assign m153_19 =15'b0;

   // m153_20 = W*in
   wire signed [14:0] m153_20;
   assign m153_20 =15'b0;

   // m153_21 = W*in
   wire signed [14:0] m153_21;
   assign m153_21 ={ {4{neg153[14]}} , neg153[14:4] };

   // m153_22 = W*in
   wire signed [14:0] m153_22;
   assign m153_22 =15'b0;

   // m153_23 = W*in
   wire signed [14:0] m153_23;
   assign m153_23 =15'b0;

   // m153_24 = W*in
   wire signed [14:0] m153_24;
   assign m153_24 =15'b0;

   // m153_25 = W*in
   wire signed [14:0] m153_25;
   assign m153_25 =15'b0;

   // m153_26 = W*in
   wire signed [14:0] m153_26;
   assign m153_26 =15'b0;

   // m153_27 = W*in
   wire signed [14:0] m153_27;
   assign m153_27 =15'b0;

   // m153_28 = W*in
   wire signed [14:0] m153_28;
   assign m153_28 =15'b0;

   // m153_29 = W*in
   wire signed [14:0] m153_29;
   assign m153_29 ={ {4{neg153[14]}} , neg153[14:4] };

   // m153_30 = W*in
   wire signed [14:0] m153_30;
   assign m153_30 =15'b0;

   // m153_31 = W*in
   wire signed [14:0] m153_31;
   assign m153_31 =15'b0;

   // m153_32 = W*in
   wire signed [14:0] m153_32;
   assign m153_32 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_33 = W*in
   wire signed [14:0] m153_33;
   assign m153_33 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_34 = W*in
   wire signed [14:0] m153_34;
   assign m153_34 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_35 = W*in
   wire signed [14:0] m153_35;
   assign m153_35 =15'b0;

   // m153_36 = W*in
   wire signed [14:0] m153_36;
   assign m153_36 =15'b0;

   // m153_37 = W*in
   wire signed [14:0] m153_37;
   assign m153_37 ={ {3{in153[14]}} , in153[14:3] };

   // m153_38 = W*in
   wire signed [14:0] m153_38;
   assign m153_38 =15'b0;

   // m153_39 = W*in
   wire signed [14:0] m153_39;
   assign m153_39 =15'b0;

   // m153_40 = W*in
   wire signed [14:0] m153_40;
   assign m153_40 =15'b0;

   // m153_41 = W*in
   wire signed [14:0] m153_41;
   assign m153_41 =15'b0;

   // m153_42 = W*in
   wire signed [14:0] m153_42;
   assign m153_42 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_43 = W*in
   wire signed [14:0] m153_43;
   assign m153_43 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_44 = W*in
   wire signed [14:0] m153_44;
   assign m153_44 ={ {4{neg153[14]}} , neg153[14:4] };

   // m153_45 = W*in
   wire signed [14:0] m153_45;
   assign m153_45 =15'b0;

   // m153_46 = W*in
   wire signed [14:0] m153_46;
   assign m153_46 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_47 = W*in
   wire signed [14:0] m153_47;
   assign m153_47 =15'b0;

   // m153_48 = W*in
   wire signed [14:0] m153_48;
   assign m153_48 =15'b0;

   // m153_49 = W*in
   wire signed [14:0] m153_49;
   assign m153_49 =15'b0;

   // m153_50 = W*in
   wire signed [14:0] m153_50;
   assign m153_50 =15'b0;

   // m153_51 = W*in
   wire signed [14:0] m153_51;
   assign m153_51 =15'b0;

   // m153_52 = W*in
   wire signed [14:0] m153_52;
   assign m153_52 ={ {3{in153[14]}} , in153[14:3] };

   // m153_53 = W*in
   wire signed [14:0] m153_53;
   assign m153_53 ={ {3{in153[14]}} , in153[14:3] };

   // m153_54 = W*in
   wire signed [14:0] m153_54;
   assign m153_54 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_55 = W*in
   wire signed [14:0] m153_55;
   assign m153_55 =15'b0;

   // m153_56 = W*in
   wire signed [14:0] m153_56;
   assign m153_56 =15'b0;

   // m153_57 = W*in
   wire signed [14:0] m153_57;
   assign m153_57 =15'b0;

   // m153_58 = W*in
   wire signed [14:0] m153_58;
   assign m153_58 ={ {3{in153[14]}} , in153[14:3] };

   // m153_59 = W*in
   wire signed [14:0] m153_59;
   assign m153_59 =15'b0;

   // m153_60 = W*in
   wire signed [14:0] m153_60;
   assign m153_60 ={ {3{in153[14]}} , in153[14:3] };

   // m153_61 = W*in
   wire signed [14:0] m153_61;
   assign m153_61 ={ {3{in153[14]}} , in153[14:3] };

   // m153_62 = W*in
   wire signed [14:0] m153_62;
   assign m153_62 =15'b0;

   // m153_63 = W*in
   wire signed [14:0] m153_63;
   assign m153_63 =15'b0;

   // m153_64 = W*in
   wire signed [14:0] m153_64;
   assign m153_64 =15'b0;

   // m153_65 = W*in
   wire signed [14:0] m153_65;
   assign m153_65 =15'b0;

   // m153_66 = W*in
   wire signed [14:0] m153_66;
   assign m153_66 =15'b0;

   // m153_67 = W*in
   wire signed [14:0] m153_67;
   assign m153_67 =15'b0;

   // m153_68 = W*in
   wire signed [14:0] m153_68;
   assign m153_68 ={ {3{in153[14]}} , in153[14:3] };

   // m153_69 = W*in
   wire signed [14:0] m153_69;
   assign m153_69 =15'b0;

   // m153_70 = W*in
   wire signed [14:0] m153_70;
   assign m153_70 ={ {4{neg153[14]}} , neg153[14:4] };

   // m153_71 = W*in
   wire signed [14:0] m153_71;
   assign m153_71 =15'b0;

   // m153_72 = W*in
   wire signed [14:0] m153_72;
   assign m153_72 =15'b0;

   // m153_73 = W*in
   wire signed [14:0] m153_73;
   assign m153_73 =15'b0;

   // m153_74 = W*in
   wire signed [14:0] m153_74;
   assign m153_74 =15'b0;

   // m153_75 = W*in
   wire signed [14:0] m153_75;
   assign m153_75 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_76 = W*in
   wire signed [14:0] m153_76;
   assign m153_76 =15'b0;

   // m153_77 = W*in
   wire signed [14:0] m153_77;
   assign m153_77 =15'b0;

   // m153_78 = W*in
   wire signed [14:0] m153_78;
   assign m153_78 =15'b0;

   // m153_79 = W*in
   wire signed [14:0] m153_79;
   assign m153_79 =15'b0;

   // m153_80 = W*in
   wire signed [14:0] m153_80;
   assign m153_80 =15'b0;

   // m153_81 = W*in
   wire signed [14:0] m153_81;
   assign m153_81 =15'b0;

   // m153_82 = W*in
   wire signed [14:0] m153_82;
   assign m153_82 =15'b0;

   // m153_83 = W*in
   wire signed [14:0] m153_83;
   assign m153_83 =15'b0;

   // m153_84 = W*in
   wire signed [14:0] m153_84;
   assign m153_84 =15'b0;

   // m153_85 = W*in
   wire signed [14:0] m153_85;
   assign m153_85 =15'b0;

   // m153_86 = W*in
   wire signed [14:0] m153_86;
   assign m153_86 =15'b0;

   // m153_87 = W*in
   wire signed [14:0] m153_87;
   assign m153_87 =15'b0;

   // m153_88 = W*in
   wire signed [14:0] m153_88;
   assign m153_88 =15'b0;

   // m153_89 = W*in
   wire signed [14:0] m153_89;
   assign m153_89 =15'b0;

   // m153_90 = W*in
   wire signed [14:0] m153_90;
   assign m153_90 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_91 = W*in
   wire signed [14:0] m153_91;
   assign m153_91 =15'b0;

   // m153_92 = W*in
   wire signed [14:0] m153_92;
   assign m153_92 =15'b0;

   // m153_93 = W*in
   wire signed [14:0] m153_93;
   assign m153_93 =15'b0;

   // m153_94 = W*in
   wire signed [14:0] m153_94;
   assign m153_94 =15'b0;

   // m153_95 = W*in
   wire signed [14:0] m153_95;
   assign m153_95 ={ {3{neg153[14]}} , neg153[14:3] };

   // m153_96 = W*in
   wire signed [14:0] m153_96;
   assign m153_96 ={ {4{in153[14]}} , in153[14:4] };

   // m153_97 = W*in
   wire signed [14:0] m153_97;
   assign m153_97 =15'b0;

   // m153_98 = W*in
   wire signed [14:0] m153_98;
   assign m153_98 =15'b0;

   // m153_99 = W*in
   wire signed [14:0] m153_99;
   assign m153_99 =15'b0;

   // m153_100 = W*in
   wire signed [14:0] m153_100;
   assign m153_100 =15'b0;

   // m154_1 = W*in
   wire signed [14:0] m154_1;
   assign m154_1 =15'b0;

   // m154_2 = W*in
   wire signed [14:0] m154_2;
   assign m154_2 =15'b0;

   // m154_3 = W*in
   wire signed [14:0] m154_3;
   assign m154_3 =15'b0;

   // m154_4 = W*in
   wire signed [14:0] m154_4;
   assign m154_4 =15'b0;

   // m154_5 = W*in
   wire signed [14:0] m154_5;
   assign m154_5 =15'b0;

   // m154_6 = W*in
   wire signed [14:0] m154_6;
   assign m154_6 =15'b0;

   // m154_7 = W*in
   wire signed [14:0] m154_7;
   assign m154_7 =15'b0;

   // m154_8 = W*in
   wire signed [14:0] m154_8;
   assign m154_8 =15'b0;

   // m154_9 = W*in
   wire signed [14:0] m154_9;
   assign m154_9 =15'b0;

   // m154_10 = W*in
   wire signed [14:0] m154_10;
   assign m154_10 =15'b0;

   // m154_11 = W*in
   wire signed [14:0] m154_11;
   assign m154_11 ={ {3{neg154[14]}} , neg154[14:3] };

   // m154_12 = W*in
   wire signed [14:0] m154_12;
   assign m154_12 =15'b0;

   // m154_13 = W*in
   wire signed [14:0] m154_13;
   assign m154_13 =15'b0;

   // m154_14 = W*in
   wire signed [14:0] m154_14;
   assign m154_14 ={ {3{in154[14]}} , in154[14:3] };

   // m154_15 = W*in
   wire signed [14:0] m154_15;
   assign m154_15 =15'b0;

   // m154_16 = W*in
   wire signed [14:0] m154_16;
   assign m154_16 =15'b0;

   // m154_17 = W*in
   wire signed [14:0] m154_17;
   assign m154_17 =15'b0;

   // m154_18 = W*in
   wire signed [14:0] m154_18;
   assign m154_18 ={ {4{in154[14]}} , in154[14:4] };

   // m154_19 = W*in
   wire signed [14:0] m154_19;
   assign m154_19 =15'b0;

   // m154_20 = W*in
   wire signed [14:0] m154_20;
   assign m154_20 =15'b0;

   // m154_21 = W*in
   wire signed [14:0] m154_21;
   assign m154_21 =15'b0;

   // m154_22 = W*in
   wire signed [14:0] m154_22;
   assign m154_22 =15'b0;

   // m154_23 = W*in
   wire signed [14:0] m154_23;
   assign m154_23 =15'b0;

   // m154_24 = W*in
   wire signed [14:0] m154_24;
   assign m154_24 =15'b0;

   // m154_25 = W*in
   wire signed [14:0] m154_25;
   assign m154_25 =15'b0;

   // m154_26 = W*in
   wire signed [14:0] m154_26;
   assign m154_26 =15'b0;

   // m154_27 = W*in
   wire signed [14:0] m154_27;
   assign m154_27 =15'b0;

   // m154_28 = W*in
   wire signed [14:0] m154_28;
   assign m154_28 =15'b0;

   // m154_29 = W*in
   wire signed [14:0] m154_29;
   assign m154_29 =15'b0;

   // m154_30 = W*in
   wire signed [14:0] m154_30;
   assign m154_30 =15'b0;

   // m154_31 = W*in
   wire signed [14:0] m154_31;
   assign m154_31 ={ {3{neg154[14]}} , neg154[14:3] };

   // m154_32 = W*in
   wire signed [14:0] m154_32;
   assign m154_32 =15'b0;

   // m154_33 = W*in
   wire signed [14:0] m154_33;
   assign m154_33 =15'b0;

   // m154_34 = W*in
   wire signed [14:0] m154_34;
   assign m154_34 ={ {4{neg154[14]}} , neg154[14:4] };

   // m154_35 = W*in
   wire signed [14:0] m154_35;
   assign m154_35 =15'b0;

   // m154_36 = W*in
   wire signed [14:0] m154_36;
   assign m154_36 =15'b0;

   // m154_37 = W*in
   wire signed [14:0] m154_37;
   assign m154_37 =15'b0;

   // m154_38 = W*in
   wire signed [14:0] m154_38;
   assign m154_38 =15'b0;

   // m154_39 = W*in
   wire signed [14:0] m154_39;
   assign m154_39 =15'b0;

   // m154_40 = W*in
   wire signed [14:0] m154_40;
   assign m154_40 =15'b0;

   // m154_41 = W*in
   wire signed [14:0] m154_41;
   assign m154_41 =15'b0;

   // m154_42 = W*in
   wire signed [14:0] m154_42;
   assign m154_42 ={ {3{neg154[14]}} , neg154[14:3] };

   // m154_43 = W*in
   wire signed [14:0] m154_43;
   assign m154_43 =15'b0;

   // m154_44 = W*in
   wire signed [14:0] m154_44;
   assign m154_44 =15'b0;

   // m154_45 = W*in
   wire signed [14:0] m154_45;
   assign m154_45 =15'b0;

   // m154_46 = W*in
   wire signed [14:0] m154_46;
   assign m154_46 =15'b0;

   // m154_47 = W*in
   wire signed [14:0] m154_47;
   assign m154_47 =15'b0;

   // m154_48 = W*in
   wire signed [14:0] m154_48;
   assign m154_48 =15'b0;

   // m154_49 = W*in
   wire signed [14:0] m154_49;
   assign m154_49 =15'b0;

   // m154_50 = W*in
   wire signed [14:0] m154_50;
   assign m154_50 =15'b0;

   // m154_51 = W*in
   wire signed [14:0] m154_51;
   assign m154_51 =15'b0;

   // m154_52 = W*in
   wire signed [14:0] m154_52;
   assign m154_52 =15'b0;

   // m154_53 = W*in
   wire signed [14:0] m154_53;
   assign m154_53 =15'b0;

   // m154_54 = W*in
   wire signed [14:0] m154_54;
   assign m154_54 =15'b0;

   // m154_55 = W*in
   wire signed [14:0] m154_55;
   assign m154_55 =15'b0;

   // m154_56 = W*in
   wire signed [14:0] m154_56;
   assign m154_56 ={ {4{in154[14]}} , in154[14:4] };

   // m154_57 = W*in
   wire signed [14:0] m154_57;
   assign m154_57 =15'b0;

   // m154_58 = W*in
   wire signed [14:0] m154_58;
   assign m154_58 =15'b0;

   // m154_59 = W*in
   wire signed [14:0] m154_59;
   assign m154_59 ={ {2{in154[14]}} , in154[14:2] };

   // m154_60 = W*in
   wire signed [14:0] m154_60;
   assign m154_60 =15'b0;

   // m154_61 = W*in
   wire signed [14:0] m154_61;
   assign m154_61 =15'b0;

   // m154_62 = W*in
   wire signed [14:0] m154_62;
   assign m154_62 =15'b0;

   // m154_63 = W*in
   wire signed [14:0] m154_63;
   assign m154_63 =15'b0;

   // m154_64 = W*in
   wire signed [14:0] m154_64;
   assign m154_64 =15'b0;

   // m154_65 = W*in
   wire signed [14:0] m154_65;
   assign m154_65 =15'b0;

   // m154_66 = W*in
   wire signed [14:0] m154_66;
   assign m154_66 =15'b0;

   // m154_67 = W*in
   wire signed [14:0] m154_67;
   assign m154_67 =15'b0;

   // m154_68 = W*in
   wire signed [14:0] m154_68;
   assign m154_68 =15'b0;

   // m154_69 = W*in
   wire signed [14:0] m154_69;
   assign m154_69 =15'b0;

   // m154_70 = W*in
   wire signed [14:0] m154_70;
   assign m154_70 =15'b0;

   // m154_71 = W*in
   wire signed [14:0] m154_71;
   assign m154_71 =15'b0;

   // m154_72 = W*in
   wire signed [14:0] m154_72;
   assign m154_72 =15'b0;

   // m154_73 = W*in
   wire signed [14:0] m154_73;
   assign m154_73 =15'b0;

   // m154_74 = W*in
   wire signed [14:0] m154_74;
   assign m154_74 =15'b0;

   // m154_75 = W*in
   wire signed [14:0] m154_75;
   assign m154_75 =15'b0;

   // m154_76 = W*in
   wire signed [14:0] m154_76;
   assign m154_76 =15'b0;

   // m154_77 = W*in
   wire signed [14:0] m154_77;
   assign m154_77 =15'b0;

   // m154_78 = W*in
   wire signed [14:0] m154_78;
   assign m154_78 =15'b0;

   // m154_79 = W*in
   wire signed [14:0] m154_79;
   assign m154_79 =15'b0;

   // m154_80 = W*in
   wire signed [14:0] m154_80;
   assign m154_80 =15'b0;

   // m154_81 = W*in
   wire signed [14:0] m154_81;
   assign m154_81 =15'b0;

   // m154_82 = W*in
   wire signed [14:0] m154_82;
   assign m154_82 =15'b0;

   // m154_83 = W*in
   wire signed [14:0] m154_83;
   assign m154_83 =15'b0;

   // m154_84 = W*in
   wire signed [14:0] m154_84;
   assign m154_84 =15'b0;

   // m154_85 = W*in
   wire signed [14:0] m154_85;
   assign m154_85 =15'b0;

   // m154_86 = W*in
   wire signed [14:0] m154_86;
   assign m154_86 =15'b0;

   // m154_87 = W*in
   wire signed [14:0] m154_87;
   assign m154_87 =15'b0;

   // m154_88 = W*in
   wire signed [14:0] m154_88;
   assign m154_88 =15'b0;

   // m154_89 = W*in
   wire signed [14:0] m154_89;
   assign m154_89 =15'b0;

   // m154_90 = W*in
   wire signed [14:0] m154_90;
   assign m154_90 =15'b0;

   // m154_91 = W*in
   wire signed [14:0] m154_91;
   assign m154_91 =15'b0;

   // m154_92 = W*in
   wire signed [14:0] m154_92;
   assign m154_92 =15'b0;

   // m154_93 = W*in
   wire signed [14:0] m154_93;
   assign m154_93 =15'b0;

   // m154_94 = W*in
   wire signed [14:0] m154_94;
   assign m154_94 =15'b0;

   // m154_95 = W*in
   wire signed [14:0] m154_95;
   assign m154_95 =15'b0;

   // m154_96 = W*in
   wire signed [14:0] m154_96;
   assign m154_96 =15'b0;

   // m154_97 = W*in
   wire signed [14:0] m154_97;
   assign m154_97 =15'b0;

   // m154_98 = W*in
   wire signed [14:0] m154_98;
   assign m154_98 =15'b0;

   // m154_99 = W*in
   wire signed [14:0] m154_99;
   assign m154_99 ={ {4{in154[14]}} , in154[14:4] };

   // m154_100 = W*in
   wire signed [14:0] m154_100;
   assign m154_100 ={ {3{in154[14]}} , in154[14:3] };

   // m155_1 = W*in
   wire signed [14:0] m155_1;
   assign m155_1 =15'b0;

   // m155_2 = W*in
   wire signed [14:0] m155_2;
   assign m155_2 ={ {3{in155[14]}} , in155[14:3] };

   // m155_3 = W*in
   wire signed [14:0] m155_3;
   assign m155_3 ={ {3{in155[14]}} , in155[14:3] };

   // m155_4 = W*in
   wire signed [14:0] m155_4;
   assign m155_4 ={ {3{in155[14]}} , in155[14:3] };

   // m155_5 = W*in
   wire signed [14:0] m155_5;
   assign m155_5 =15'b0;

   // m155_6 = W*in
   wire signed [14:0] m155_6;
   assign m155_6 ={ {3{in155[14]}} , in155[14:3] };

   // m155_7 = W*in
   wire signed [14:0] m155_7;
   assign m155_7 =15'b0;

   // m155_8 = W*in
   wire signed [14:0] m155_8;
   assign m155_8 =15'b0;

   // m155_9 = W*in
   wire signed [14:0] m155_9;
   assign m155_9 =15'b0;

   // m155_10 = W*in
   wire signed [14:0] m155_10;
   assign m155_10 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_11 = W*in
   wire signed [14:0] m155_11;
   assign m155_11 =15'b0;

   // m155_12 = W*in
   wire signed [14:0] m155_12;
   assign m155_12 =15'b0;

   // m155_13 = W*in
   wire signed [14:0] m155_13;
   assign m155_13 ={ {3{in155[14]}} , in155[14:3] };

   // m155_14 = W*in
   wire signed [14:0] m155_14;
   assign m155_14 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_15 = W*in
   wire signed [14:0] m155_15;
   assign m155_15 =15'b0;

   // m155_16 = W*in
   wire signed [14:0] m155_16;
   assign m155_16 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_17 = W*in
   wire signed [14:0] m155_17;
   assign m155_17 =15'b0;

   // m155_18 = W*in
   wire signed [14:0] m155_18;
   assign m155_18 ={ {3{in155[14]}} , in155[14:3] };

   // m155_19 = W*in
   wire signed [14:0] m155_19;
   assign m155_19 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_20 = W*in
   wire signed [14:0] m155_20;
   assign m155_20 =15'b0;

   // m155_21 = W*in
   wire signed [14:0] m155_21;
   assign m155_21 =15'b0;

   // m155_22 = W*in
   wire signed [14:0] m155_22;
   assign m155_22 ={ {4{in155[14]}} , in155[14:4] };

   // m155_23 = W*in
   wire signed [14:0] m155_23;
   assign m155_23 =15'b0;

   // m155_24 = W*in
   wire signed [14:0] m155_24;
   assign m155_24 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_25 = W*in
   wire signed [14:0] m155_25;
   assign m155_25 ={ {3{in155[14]}} , in155[14:3] };

   // m155_26 = W*in
   wire signed [14:0] m155_26;
   assign m155_26 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_27 = W*in
   wire signed [14:0] m155_27;
   assign m155_27 =15'b0;

   // m155_28 = W*in
   wire signed [14:0] m155_28;
   assign m155_28 ={ {3{in155[14]}} , in155[14:3] };

   // m155_29 = W*in
   wire signed [14:0] m155_29;
   assign m155_29 =15'b0;

   // m155_30 = W*in
   wire signed [14:0] m155_30;
   assign m155_30 =15'b0;

   // m155_31 = W*in
   wire signed [14:0] m155_31;
   assign m155_31 =15'b0;

   // m155_32 = W*in
   wire signed [14:0] m155_32;
   assign m155_32 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_33 = W*in
   wire signed [14:0] m155_33;
   assign m155_33 =15'b0;

   // m155_34 = W*in
   wire signed [14:0] m155_34;
   assign m155_34 ={ {3{in155[14]}} , in155[14:3] };

   // m155_35 = W*in
   wire signed [14:0] m155_35;
   assign m155_35 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_36 = W*in
   wire signed [14:0] m155_36;
   assign m155_36 =15'b0;

   // m155_37 = W*in
   wire signed [14:0] m155_37;
   assign m155_37 =15'b0;

   // m155_38 = W*in
   wire signed [14:0] m155_38;
   assign m155_38 ={ {3{in155[14]}} , in155[14:3] };

   // m155_39 = W*in
   wire signed [14:0] m155_39;
   assign m155_39 =15'b0;

   // m155_40 = W*in
   wire signed [14:0] m155_40;
   assign m155_40 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_41 = W*in
   wire signed [14:0] m155_41;
   assign m155_41 ={ {3{in155[14]}} , in155[14:3] };

   // m155_42 = W*in
   wire signed [14:0] m155_42;
   assign m155_42 =15'b0;

   // m155_43 = W*in
   wire signed [14:0] m155_43;
   assign m155_43 =15'b0;

   // m155_44 = W*in
   wire signed [14:0] m155_44;
   assign m155_44 =15'b0;

   // m155_45 = W*in
   wire signed [14:0] m155_45;
   assign m155_45 ={ {3{in155[14]}} , in155[14:3] };

   // m155_46 = W*in
   wire signed [14:0] m155_46;
   assign m155_46 ={ {4{neg155[14]}} , neg155[14:4] };

   // m155_47 = W*in
   wire signed [14:0] m155_47;
   assign m155_47 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_48 = W*in
   wire signed [14:0] m155_48;
   assign m155_48 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_49 = W*in
   wire signed [14:0] m155_49;
   assign m155_49 =15'b0;

   // m155_50 = W*in
   wire signed [14:0] m155_50;
   assign m155_50 =15'b0;

   // m155_51 = W*in
   wire signed [14:0] m155_51;
   assign m155_51 =15'b0;

   // m155_52 = W*in
   wire signed [14:0] m155_52;
   assign m155_52 =15'b0;

   // m155_53 = W*in
   wire signed [14:0] m155_53;
   assign m155_53 =15'b0;

   // m155_54 = W*in
   wire signed [14:0] m155_54;
   assign m155_54 =15'b0;

   // m155_55 = W*in
   wire signed [14:0] m155_55;
   assign m155_55 =15'b0;

   // m155_56 = W*in
   wire signed [14:0] m155_56;
   assign m155_56 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_57 = W*in
   wire signed [14:0] m155_57;
   assign m155_57 =15'b0;

   // m155_58 = W*in
   wire signed [14:0] m155_58;
   assign m155_58 ={ {4{neg155[14]}} , neg155[14:4] };

   // m155_59 = W*in
   wire signed [14:0] m155_59;
   assign m155_59 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_60 = W*in
   wire signed [14:0] m155_60;
   assign m155_60 ={ {3{in155[14]}} , in155[14:3] };

   // m155_61 = W*in
   wire signed [14:0] m155_61;
   assign m155_61 =15'b0;

   // m155_62 = W*in
   wire signed [14:0] m155_62;
   assign m155_62 =15'b0;

   // m155_63 = W*in
   wire signed [14:0] m155_63;
   assign m155_63 =15'b0;

   // m155_64 = W*in
   wire signed [14:0] m155_64;
   assign m155_64 =15'b0;

   // m155_65 = W*in
   wire signed [14:0] m155_65;
   assign m155_65 =15'b0;

   // m155_66 = W*in
   wire signed [14:0] m155_66;
   assign m155_66 =15'b0;

   // m155_67 = W*in
   wire signed [14:0] m155_67;
   assign m155_67 =15'b0;

   // m155_68 = W*in
   wire signed [14:0] m155_68;
   assign m155_68 ={ {4{in155[14]}} , in155[14:4] };

   // m155_69 = W*in
   wire signed [14:0] m155_69;
   assign m155_69 ={ {3{in155[14]}} , in155[14:3] };

   // m155_70 = W*in
   wire signed [14:0] m155_70;
   assign m155_70 ={ {2{neg155[14]}} , neg155[14:2] };

   // m155_71 = W*in
   wire signed [14:0] m155_71;
   assign m155_71 =15'b0;

   // m155_72 = W*in
   wire signed [14:0] m155_72;
   assign m155_72 ={ {3{in155[14]}} , in155[14:3] };

   // m155_73 = W*in
   wire signed [14:0] m155_73;
   assign m155_73 =15'b0;

   // m155_74 = W*in
   wire signed [14:0] m155_74;
   assign m155_74 =15'b0;

   // m155_75 = W*in
   wire signed [14:0] m155_75;
   assign m155_75 =15'b0;

   // m155_76 = W*in
   wire signed [14:0] m155_76;
   assign m155_76 =15'b0;

   // m155_77 = W*in
   wire signed [14:0] m155_77;
   assign m155_77 =15'b0;

   // m155_78 = W*in
   wire signed [14:0] m155_78;
   assign m155_78 =15'b0;

   // m155_79 = W*in
   wire signed [14:0] m155_79;
   assign m155_79 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_80 = W*in
   wire signed [14:0] m155_80;
   assign m155_80 =15'b0;

   // m155_81 = W*in
   wire signed [14:0] m155_81;
   assign m155_81 =15'b0;

   // m155_82 = W*in
   wire signed [14:0] m155_82;
   assign m155_82 =15'b0;

   // m155_83 = W*in
   wire signed [14:0] m155_83;
   assign m155_83 =15'b0;

   // m155_84 = W*in
   wire signed [14:0] m155_84;
   assign m155_84 =15'b0;

   // m155_85 = W*in
   wire signed [14:0] m155_85;
   assign m155_85 =15'b0;

   // m155_86 = W*in
   wire signed [14:0] m155_86;
   assign m155_86 =15'b0;

   // m155_87 = W*in
   wire signed [14:0] m155_87;
   assign m155_87 =15'b0;

   // m155_88 = W*in
   wire signed [14:0] m155_88;
   assign m155_88 =15'b0;

   // m155_89 = W*in
   wire signed [14:0] m155_89;
   assign m155_89 =15'b0;

   // m155_90 = W*in
   wire signed [14:0] m155_90;
   assign m155_90 =15'b0;

   // m155_91 = W*in
   wire signed [14:0] m155_91;
   assign m155_91 =15'b0;

   // m155_92 = W*in
   wire signed [14:0] m155_92;
   assign m155_92 =15'b0;

   // m155_93 = W*in
   wire signed [14:0] m155_93;
   assign m155_93 =15'b0;

   // m155_94 = W*in
   wire signed [14:0] m155_94;
   assign m155_94 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_95 = W*in
   wire signed [14:0] m155_95;
   assign m155_95 =15'b0;

   // m155_96 = W*in
   wire signed [14:0] m155_96;
   assign m155_96 ={ {3{in155[14]}} , in155[14:3] };

   // m155_97 = W*in
   wire signed [14:0] m155_97;
   assign m155_97 ={ {3{in155[14]}} , in155[14:3] };

   // m155_98 = W*in
   wire signed [14:0] m155_98;
   assign m155_98 ={ {3{neg155[14]}} , neg155[14:3] };

   // m155_99 = W*in
   wire signed [14:0] m155_99;
   assign m155_99 =15'b0;

   // m155_100 = W*in
   wire signed [14:0] m155_100;
   assign m155_100 =15'b0;

   // m156_1 = W*in
   wire signed [14:0] m156_1;
   assign m156_1 =15'b0;

   // m156_2 = W*in
   wire signed [14:0] m156_2;
   assign m156_2 =15'b0;

   // m156_3 = W*in
   wire signed [14:0] m156_3;
   assign m156_3 ={ {4{in156[14]}} , in156[14:4] };

   // m156_4 = W*in
   wire signed [14:0] m156_4;
   assign m156_4 ={ {3{in156[14]}} , in156[14:3] };

   // m156_5 = W*in
   wire signed [14:0] m156_5;
   assign m156_5 =15'b0;

   // m156_6 = W*in
   wire signed [14:0] m156_6;
   assign m156_6 =15'b0;

   // m156_7 = W*in
   wire signed [14:0] m156_7;
   assign m156_7 =15'b0;

   // m156_8 = W*in
   wire signed [14:0] m156_8;
   assign m156_8 =15'b0;

   // m156_9 = W*in
   wire signed [14:0] m156_9;
   assign m156_9 =15'b0;

   // m156_10 = W*in
   wire signed [14:0] m156_10;
   assign m156_10 =15'b0;

   // m156_11 = W*in
   wire signed [14:0] m156_11;
   assign m156_11 =15'b0;

   // m156_12 = W*in
   wire signed [14:0] m156_12;
   assign m156_12 =15'b0;

   // m156_13 = W*in
   wire signed [14:0] m156_13;
   assign m156_13 ={ {3{in156[14]}} , in156[14:3] };

   // m156_14 = W*in
   wire signed [14:0] m156_14;
   assign m156_14 =15'b0;

   // m156_15 = W*in
   wire signed [14:0] m156_15;
   assign m156_15 =15'b0;

   // m156_16 = W*in
   wire signed [14:0] m156_16;
   assign m156_16 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_17 = W*in
   wire signed [14:0] m156_17;
   assign m156_17 =15'b0;

   // m156_18 = W*in
   wire signed [14:0] m156_18;
   assign m156_18 =15'b0;

   // m156_19 = W*in
   wire signed [14:0] m156_19;
   assign m156_19 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_20 = W*in
   wire signed [14:0] m156_20;
   assign m156_20 =15'b0;

   // m156_21 = W*in
   wire signed [14:0] m156_21;
   assign m156_21 =15'b0;

   // m156_22 = W*in
   wire signed [14:0] m156_22;
   assign m156_22 =15'b0;

   // m156_23 = W*in
   wire signed [14:0] m156_23;
   assign m156_23 =15'b0;

   // m156_24 = W*in
   wire signed [14:0] m156_24;
   assign m156_24 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_25 = W*in
   wire signed [14:0] m156_25;
   assign m156_25 ={ {2{in156[14]}} , in156[14:2] };

   // m156_26 = W*in
   wire signed [14:0] m156_26;
   assign m156_26 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_27 = W*in
   wire signed [14:0] m156_27;
   assign m156_27 =15'b0;

   // m156_28 = W*in
   wire signed [14:0] m156_28;
   assign m156_28 =15'b0;

   // m156_29 = W*in
   wire signed [14:0] m156_29;
   assign m156_29 =15'b0;

   // m156_30 = W*in
   wire signed [14:0] m156_30;
   assign m156_30 =15'b0;

   // m156_31 = W*in
   wire signed [14:0] m156_31;
   assign m156_31 =15'b0;

   // m156_32 = W*in
   wire signed [14:0] m156_32;
   assign m156_32 =15'b0;

   // m156_33 = W*in
   wire signed [14:0] m156_33;
   assign m156_33 =15'b0;

   // m156_34 = W*in
   wire signed [14:0] m156_34;
   assign m156_34 ={ {3{in156[14]}} , in156[14:3] };

   // m156_35 = W*in
   wire signed [14:0] m156_35;
   assign m156_35 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_36 = W*in
   wire signed [14:0] m156_36;
   assign m156_36 =15'b0;

   // m156_37 = W*in
   wire signed [14:0] m156_37;
   assign m156_37 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_38 = W*in
   wire signed [14:0] m156_38;
   assign m156_38 =15'b0;

   // m156_39 = W*in
   wire signed [14:0] m156_39;
   assign m156_39 =15'b0;

   // m156_40 = W*in
   wire signed [14:0] m156_40;
   assign m156_40 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_41 = W*in
   wire signed [14:0] m156_41;
   assign m156_41 =15'b0;

   // m156_42 = W*in
   wire signed [14:0] m156_42;
   assign m156_42 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_43 = W*in
   wire signed [14:0] m156_43;
   assign m156_43 =15'b0;

   // m156_44 = W*in
   wire signed [14:0] m156_44;
   assign m156_44 =15'b0;

   // m156_45 = W*in
   wire signed [14:0] m156_45;
   assign m156_45 =15'b0;

   // m156_46 = W*in
   wire signed [14:0] m156_46;
   assign m156_46 =15'b0;

   // m156_47 = W*in
   wire signed [14:0] m156_47;
   assign m156_47 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_48 = W*in
   wire signed [14:0] m156_48;
   assign m156_48 ={ {4{neg156[14]}} , neg156[14:4] };

   // m156_49 = W*in
   wire signed [14:0] m156_49;
   assign m156_49 =15'b0;

   // m156_50 = W*in
   wire signed [14:0] m156_50;
   assign m156_50 =15'b0;

   // m156_51 = W*in
   wire signed [14:0] m156_51;
   assign m156_51 =15'b0;

   // m156_52 = W*in
   wire signed [14:0] m156_52;
   assign m156_52 =15'b0;

   // m156_53 = W*in
   wire signed [14:0] m156_53;
   assign m156_53 =15'b0;

   // m156_54 = W*in
   wire signed [14:0] m156_54;
   assign m156_54 =15'b0;

   // m156_55 = W*in
   wire signed [14:0] m156_55;
   assign m156_55 =15'b0;

   // m156_56 = W*in
   wire signed [14:0] m156_56;
   assign m156_56 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_57 = W*in
   wire signed [14:0] m156_57;
   assign m156_57 =15'b0;

   // m156_58 = W*in
   wire signed [14:0] m156_58;
   assign m156_58 ={ {4{in156[14]}} , in156[14:4] };

   // m156_59 = W*in
   wire signed [14:0] m156_59;
   assign m156_59 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_60 = W*in
   wire signed [14:0] m156_60;
   assign m156_60 =15'b0;

   // m156_61 = W*in
   wire signed [14:0] m156_61;
   assign m156_61 =15'b0;

   // m156_62 = W*in
   wire signed [14:0] m156_62;
   assign m156_62 =15'b0;

   // m156_63 = W*in
   wire signed [14:0] m156_63;
   assign m156_63 =15'b0;

   // m156_64 = W*in
   wire signed [14:0] m156_64;
   assign m156_64 ={ {4{in156[14]}} , in156[14:4] };

   // m156_65 = W*in
   wire signed [14:0] m156_65;
   assign m156_65 =15'b0;

   // m156_66 = W*in
   wire signed [14:0] m156_66;
   assign m156_66 =15'b0;

   // m156_67 = W*in
   wire signed [14:0] m156_67;
   assign m156_67 =15'b0;

   // m156_68 = W*in
   wire signed [14:0] m156_68;
   assign m156_68 ={ {3{in156[14]}} , in156[14:3] };

   // m156_69 = W*in
   wire signed [14:0] m156_69;
   assign m156_69 ={ {3{in156[14]}} , in156[14:3] };

   // m156_70 = W*in
   wire signed [14:0] m156_70;
   assign m156_70 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_71 = W*in
   wire signed [14:0] m156_71;
   assign m156_71 =15'b0;

   // m156_72 = W*in
   wire signed [14:0] m156_72;
   assign m156_72 ={ {3{in156[14]}} , in156[14:3] };

   // m156_73 = W*in
   wire signed [14:0] m156_73;
   assign m156_73 =15'b0;

   // m156_74 = W*in
   wire signed [14:0] m156_74;
   assign m156_74 ={ {4{neg156[14]}} , neg156[14:4] };

   // m156_75 = W*in
   wire signed [14:0] m156_75;
   assign m156_75 =15'b0;

   // m156_76 = W*in
   wire signed [14:0] m156_76;
   assign m156_76 =15'b0;

   // m156_77 = W*in
   wire signed [14:0] m156_77;
   assign m156_77 =15'b0;

   // m156_78 = W*in
   wire signed [14:0] m156_78;
   assign m156_78 =15'b0;

   // m156_79 = W*in
   wire signed [14:0] m156_79;
   assign m156_79 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_80 = W*in
   wire signed [14:0] m156_80;
   assign m156_80 ={ {3{in156[14]}} , in156[14:3] };

   // m156_81 = W*in
   wire signed [14:0] m156_81;
   assign m156_81 =15'b0;

   // m156_82 = W*in
   wire signed [14:0] m156_82;
   assign m156_82 =15'b0;

   // m156_83 = W*in
   wire signed [14:0] m156_83;
   assign m156_83 =15'b0;

   // m156_84 = W*in
   wire signed [14:0] m156_84;
   assign m156_84 =15'b0;

   // m156_85 = W*in
   wire signed [14:0] m156_85;
   assign m156_85 =15'b0;

   // m156_86 = W*in
   wire signed [14:0] m156_86;
   assign m156_86 =15'b0;

   // m156_87 = W*in
   wire signed [14:0] m156_87;
   assign m156_87 =15'b0;

   // m156_88 = W*in
   wire signed [14:0] m156_88;
   assign m156_88 =15'b0;

   // m156_89 = W*in
   wire signed [14:0] m156_89;
   assign m156_89 =15'b0;

   // m156_90 = W*in
   wire signed [14:0] m156_90;
   assign m156_90 =15'b0;

   // m156_91 = W*in
   wire signed [14:0] m156_91;
   assign m156_91 =15'b0;

   // m156_92 = W*in
   wire signed [14:0] m156_92;
   assign m156_92 =15'b0;

   // m156_93 = W*in
   wire signed [14:0] m156_93;
   assign m156_93 =15'b0;

   // m156_94 = W*in
   wire signed [14:0] m156_94;
   assign m156_94 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_95 = W*in
   wire signed [14:0] m156_95;
   assign m156_95 =15'b0;

   // m156_96 = W*in
   wire signed [14:0] m156_96;
   assign m156_96 =15'b0;

   // m156_97 = W*in
   wire signed [14:0] m156_97;
   assign m156_97 =15'b0;

   // m156_98 = W*in
   wire signed [14:0] m156_98;
   assign m156_98 ={ {3{neg156[14]}} , neg156[14:3] };

   // m156_99 = W*in
   wire signed [14:0] m156_99;
   assign m156_99 =15'b0;

   // m156_100 = W*in
   wire signed [14:0] m156_100;
   assign m156_100 ={ {4{in156[14]}} , in156[14:4] };

   // m157_1 = W*in
   wire signed [14:0] m157_1;
   assign m157_1 ={ {3{in157[14]}} , in157[14:3] };

   // m157_2 = W*in
   wire signed [14:0] m157_2;
   assign m157_2 ={ {3{in157[14]}} , in157[14:3] };

   // m157_3 = W*in
   wire signed [14:0] m157_3;
   assign m157_3 =15'b0;

   // m157_4 = W*in
   wire signed [14:0] m157_4;
   assign m157_4 =15'b0;

   // m157_5 = W*in
   wire signed [14:0] m157_5;
   assign m157_5 =15'b0;

   // m157_6 = W*in
   wire signed [14:0] m157_6;
   assign m157_6 =15'b0;

   // m157_7 = W*in
   wire signed [14:0] m157_7;
   assign m157_7 =15'b0;

   // m157_8 = W*in
   wire signed [14:0] m157_8;
   assign m157_8 =15'b0;

   // m157_9 = W*in
   wire signed [14:0] m157_9;
   assign m157_9 ={ {3{in157[14]}} , in157[14:3] };

   // m157_10 = W*in
   wire signed [14:0] m157_10;
   assign m157_10 =15'b0;

   // m157_11 = W*in
   wire signed [14:0] m157_11;
   assign m157_11 =15'b0;

   // m157_12 = W*in
   wire signed [14:0] m157_12;
   assign m157_12 =15'b0;

   // m157_13 = W*in
   wire signed [14:0] m157_13;
   assign m157_13 =15'b0;

   // m157_14 = W*in
   wire signed [14:0] m157_14;
   assign m157_14 =15'b0;

   // m157_15 = W*in
   wire signed [14:0] m157_15;
   assign m157_15 =15'b0;

   // m157_16 = W*in
   wire signed [14:0] m157_16;
   assign m157_16 =15'b0;

   // m157_17 = W*in
   wire signed [14:0] m157_17;
   assign m157_17 =15'b0;

   // m157_18 = W*in
   wire signed [14:0] m157_18;
   assign m157_18 =15'b0;

   // m157_19 = W*in
   wire signed [14:0] m157_19;
   assign m157_19 =15'b0;

   // m157_20 = W*in
   wire signed [14:0] m157_20;
   assign m157_20 =15'b0;

   // m157_21 = W*in
   wire signed [14:0] m157_21;
   assign m157_21 =15'b0;

   // m157_22 = W*in
   wire signed [14:0] m157_22;
   assign m157_22 ={ {4{in157[14]}} , in157[14:4] };

   // m157_23 = W*in
   wire signed [14:0] m157_23;
   assign m157_23 =15'b0;

   // m157_24 = W*in
   wire signed [14:0] m157_24;
   assign m157_24 =15'b0;

   // m157_25 = W*in
   wire signed [14:0] m157_25;
   assign m157_25 =15'b0;

   // m157_26 = W*in
   wire signed [14:0] m157_26;
   assign m157_26 =15'b0;

   // m157_27 = W*in
   wire signed [14:0] m157_27;
   assign m157_27 =15'b0;

   // m157_28 = W*in
   wire signed [14:0] m157_28;
   assign m157_28 =15'b0;

   // m157_29 = W*in
   wire signed [14:0] m157_29;
   assign m157_29 =15'b0;

   // m157_30 = W*in
   wire signed [14:0] m157_30;
   assign m157_30 =15'b0;

   // m157_31 = W*in
   wire signed [14:0] m157_31;
   assign m157_31 ={ {3{neg157[14]}} , neg157[14:3] };

   // m157_32 = W*in
   wire signed [14:0] m157_32;
   assign m157_32 ={ {3{in157[14]}} , in157[14:3] };

   // m157_33 = W*in
   wire signed [14:0] m157_33;
   assign m157_33 =15'b0;

   // m157_34 = W*in
   wire signed [14:0] m157_34;
   assign m157_34 =15'b0;

   // m157_35 = W*in
   wire signed [14:0] m157_35;
   assign m157_35 ={ {3{in157[14]}} , in157[14:3] };

   // m157_36 = W*in
   wire signed [14:0] m157_36;
   assign m157_36 =15'b0;

   // m157_37 = W*in
   wire signed [14:0] m157_37;
   assign m157_37 ={ {3{neg157[14]}} , neg157[14:3] };

   // m157_38 = W*in
   wire signed [14:0] m157_38;
   assign m157_38 =15'b0;

   // m157_39 = W*in
   wire signed [14:0] m157_39;
   assign m157_39 =15'b0;

   // m157_40 = W*in
   wire signed [14:0] m157_40;
   assign m157_40 =15'b0;

   // m157_41 = W*in
   wire signed [14:0] m157_41;
   assign m157_41 =15'b0;

   // m157_42 = W*in
   wire signed [14:0] m157_42;
   assign m157_42 ={ {3{in157[14]}} , in157[14:3] };

   // m157_43 = W*in
   wire signed [14:0] m157_43;
   assign m157_43 =15'b0;

   // m157_44 = W*in
   wire signed [14:0] m157_44;
   assign m157_44 =15'b0;

   // m157_45 = W*in
   wire signed [14:0] m157_45;
   assign m157_45 =15'b0;

   // m157_46 = W*in
   wire signed [14:0] m157_46;
   assign m157_46 =15'b0;

   // m157_47 = W*in
   wire signed [14:0] m157_47;
   assign m157_47 =15'b0;

   // m157_48 = W*in
   wire signed [14:0] m157_48;
   assign m157_48 =15'b0;

   // m157_49 = W*in
   wire signed [14:0] m157_49;
   assign m157_49 =15'b0;

   // m157_50 = W*in
   wire signed [14:0] m157_50;
   assign m157_50 =15'b0;

   // m157_51 = W*in
   wire signed [14:0] m157_51;
   assign m157_51 ={ {3{neg157[14]}} , neg157[14:3] };

   // m157_52 = W*in
   wire signed [14:0] m157_52;
   assign m157_52 =15'b0;

   // m157_53 = W*in
   wire signed [14:0] m157_53;
   assign m157_53 =15'b0;

   // m157_54 = W*in
   wire signed [14:0] m157_54;
   assign m157_54 =15'b0;

   // m157_55 = W*in
   wire signed [14:0] m157_55;
   assign m157_55 =15'b0;

   // m157_56 = W*in
   wire signed [14:0] m157_56;
   assign m157_56 =15'b0;

   // m157_57 = W*in
   wire signed [14:0] m157_57;
   assign m157_57 =15'b0;

   // m157_58 = W*in
   wire signed [14:0] m157_58;
   assign m157_58 =15'b0;

   // m157_59 = W*in
   wire signed [14:0] m157_59;
   assign m157_59 =15'b0;

   // m157_60 = W*in
   wire signed [14:0] m157_60;
   assign m157_60 =15'b0;

   // m157_61 = W*in
   wire signed [14:0] m157_61;
   assign m157_61 =15'b0;

   // m157_62 = W*in
   wire signed [14:0] m157_62;
   assign m157_62 =15'b0;

   // m157_63 = W*in
   wire signed [14:0] m157_63;
   assign m157_63 =15'b0;

   // m157_64 = W*in
   wire signed [14:0] m157_64;
   assign m157_64 =15'b0;

   // m157_65 = W*in
   wire signed [14:0] m157_65;
   assign m157_65 =15'b0;

   // m157_66 = W*in
   wire signed [14:0] m157_66;
   assign m157_66 =15'b0;

   // m157_67 = W*in
   wire signed [14:0] m157_67;
   assign m157_67 =15'b0;

   // m157_68 = W*in
   wire signed [14:0] m157_68;
   assign m157_68 =15'b0;

   // m157_69 = W*in
   wire signed [14:0] m157_69;
   assign m157_69 =15'b0;

   // m157_70 = W*in
   wire signed [14:0] m157_70;
   assign m157_70 ={ {4{neg157[14]}} , neg157[14:4] };

   // m157_71 = W*in
   wire signed [14:0] m157_71;
   assign m157_71 =15'b0;

   // m157_72 = W*in
   wire signed [14:0] m157_72;
   assign m157_72 =15'b0;

   // m157_73 = W*in
   wire signed [14:0] m157_73;
   assign m157_73 =15'b0;

   // m157_74 = W*in
   wire signed [14:0] m157_74;
   assign m157_74 ={ {4{neg157[14]}} , neg157[14:4] };

   // m157_75 = W*in
   wire signed [14:0] m157_75;
   assign m157_75 =15'b0;

   // m157_76 = W*in
   wire signed [14:0] m157_76;
   assign m157_76 =15'b0;

   // m157_77 = W*in
   wire signed [14:0] m157_77;
   assign m157_77 =15'b0;

   // m157_78 = W*in
   wire signed [14:0] m157_78;
   assign m157_78 =15'b0;

   // m157_79 = W*in
   wire signed [14:0] m157_79;
   assign m157_79 =15'b0;

   // m157_80 = W*in
   wire signed [14:0] m157_80;
   assign m157_80 =15'b0;

   // m157_81 = W*in
   wire signed [14:0] m157_81;
   assign m157_81 =15'b0;

   // m157_82 = W*in
   wire signed [14:0] m157_82;
   assign m157_82 ={ {3{in157[14]}} , in157[14:3] };

   // m157_83 = W*in
   wire signed [14:0] m157_83;
   assign m157_83 =15'b0;

   // m157_84 = W*in
   wire signed [14:0] m157_84;
   assign m157_84 =15'b0;

   // m157_85 = W*in
   wire signed [14:0] m157_85;
   assign m157_85 =15'b0;

   // m157_86 = W*in
   wire signed [14:0] m157_86;
   assign m157_86 =15'b0;

   // m157_87 = W*in
   wire signed [14:0] m157_87;
   assign m157_87 =15'b0;

   // m157_88 = W*in
   wire signed [14:0] m157_88;
   assign m157_88 =15'b0;

   // m157_89 = W*in
   wire signed [14:0] m157_89;
   assign m157_89 =15'b0;

   // m157_90 = W*in
   wire signed [14:0] m157_90;
   assign m157_90 =15'b0;

   // m157_91 = W*in
   wire signed [14:0] m157_91;
   assign m157_91 =15'b0;

   // m157_92 = W*in
   wire signed [14:0] m157_92;
   assign m157_92 =15'b0;

   // m157_93 = W*in
   wire signed [14:0] m157_93;
   assign m157_93 =15'b0;

   // m157_94 = W*in
   wire signed [14:0] m157_94;
   assign m157_94 =15'b0;

   // m157_95 = W*in
   wire signed [14:0] m157_95;
   assign m157_95 =15'b0;

   // m157_96 = W*in
   wire signed [14:0] m157_96;
   assign m157_96 =15'b0;

   // m157_97 = W*in
   wire signed [14:0] m157_97;
   assign m157_97 =15'b0;

   // m157_98 = W*in
   wire signed [14:0] m157_98;
   assign m157_98 =15'b0;

   // m157_99 = W*in
   wire signed [14:0] m157_99;
   assign m157_99 =15'b0;

   // m157_100 = W*in
   wire signed [14:0] m157_100;
   assign m157_100 =15'b0;

   // m158_1 = W*in
   wire signed [14:0] m158_1;
   assign m158_1 =15'b0;

   // m158_2 = W*in
   wire signed [14:0] m158_2;
   assign m158_2 ={ {3{in158[14]}} , in158[14:3] };

   // m158_3 = W*in
   wire signed [14:0] m158_3;
   assign m158_3 =15'b0;

   // m158_4 = W*in
   wire signed [14:0] m158_4;
   assign m158_4 =15'b0;

   // m158_5 = W*in
   wire signed [14:0] m158_5;
   assign m158_5 =15'b0;

   // m158_6 = W*in
   wire signed [14:0] m158_6;
   assign m158_6 =15'b0;

   // m158_7 = W*in
   wire signed [14:0] m158_7;
   assign m158_7 ={ {3{in158[14]}} , in158[14:3] };

   // m158_8 = W*in
   wire signed [14:0] m158_8;
   assign m158_8 =15'b0;

   // m158_9 = W*in
   wire signed [14:0] m158_9;
   assign m158_9 =15'b0;

   // m158_10 = W*in
   wire signed [14:0] m158_10;
   assign m158_10 =15'b0;

   // m158_11 = W*in
   wire signed [14:0] m158_11;
   assign m158_11 ={ {3{in158[14]}} , in158[14:3] };

   // m158_12 = W*in
   wire signed [14:0] m158_12;
   assign m158_12 =15'b0;

   // m158_13 = W*in
   wire signed [14:0] m158_13;
   assign m158_13 =15'b0;

   // m158_14 = W*in
   wire signed [14:0] m158_14;
   assign m158_14 =15'b0;

   // m158_15 = W*in
   wire signed [14:0] m158_15;
   assign m158_15 =15'b0;

   // m158_16 = W*in
   wire signed [14:0] m158_16;
   assign m158_16 ={ {3{in158[14]}} , in158[14:3] };

   // m158_17 = W*in
   wire signed [14:0] m158_17;
   assign m158_17 =15'b0;

   // m158_18 = W*in
   wire signed [14:0] m158_18;
   assign m158_18 ={ {3{in158[14]}} , in158[14:3] };

   // m158_19 = W*in
   wire signed [14:0] m158_19;
   assign m158_19 =15'b0;

   // m158_20 = W*in
   wire signed [14:0] m158_20;
   assign m158_20 =15'b0;

   // m158_21 = W*in
   wire signed [14:0] m158_21;
   assign m158_21 ={ {3{in158[14]}} , in158[14:3] };

   // m158_22 = W*in
   wire signed [14:0] m158_22;
   assign m158_22 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_23 = W*in
   wire signed [14:0] m158_23;
   assign m158_23 =15'b0;

   // m158_24 = W*in
   wire signed [14:0] m158_24;
   assign m158_24 =15'b0;

   // m158_25 = W*in
   wire signed [14:0] m158_25;
   assign m158_25 =15'b0;

   // m158_26 = W*in
   wire signed [14:0] m158_26;
   assign m158_26 =15'b0;

   // m158_27 = W*in
   wire signed [14:0] m158_27;
   assign m158_27 =15'b0;

   // m158_28 = W*in
   wire signed [14:0] m158_28;
   assign m158_28 =15'b0;

   // m158_29 = W*in
   wire signed [14:0] m158_29;
   assign m158_29 ={ {4{in158[14]}} , in158[14:4] };

   // m158_30 = W*in
   wire signed [14:0] m158_30;
   assign m158_30 ={ {3{in158[14]}} , in158[14:3] };

   // m158_31 = W*in
   wire signed [14:0] m158_31;
   assign m158_31 ={ {4{neg158[14]}} , neg158[14:4] };

   // m158_32 = W*in
   wire signed [14:0] m158_32;
   assign m158_32 =15'b0;

   // m158_33 = W*in
   wire signed [14:0] m158_33;
   assign m158_33 =15'b0;

   // m158_34 = W*in
   wire signed [14:0] m158_34;
   assign m158_34 =15'b0;

   // m158_35 = W*in
   wire signed [14:0] m158_35;
   assign m158_35 =15'b0;

   // m158_36 = W*in
   wire signed [14:0] m158_36;
   assign m158_36 =15'b0;

   // m158_37 = W*in
   wire signed [14:0] m158_37;
   assign m158_37 =15'b0;

   // m158_38 = W*in
   wire signed [14:0] m158_38;
   assign m158_38 =15'b0;

   // m158_39 = W*in
   wire signed [14:0] m158_39;
   assign m158_39 =15'b0;

   // m158_40 = W*in
   wire signed [14:0] m158_40;
   assign m158_40 =15'b0;

   // m158_41 = W*in
   wire signed [14:0] m158_41;
   assign m158_41 =15'b0;

   // m158_42 = W*in
   wire signed [14:0] m158_42;
   assign m158_42 =15'b0;

   // m158_43 = W*in
   wire signed [14:0] m158_43;
   assign m158_43 =15'b0;

   // m158_44 = W*in
   wire signed [14:0] m158_44;
   assign m158_44 ={ {3{in158[14]}} , in158[14:3] };

   // m158_45 = W*in
   wire signed [14:0] m158_45;
   assign m158_45 =15'b0;

   // m158_46 = W*in
   wire signed [14:0] m158_46;
   assign m158_46 =15'b0;

   // m158_47 = W*in
   wire signed [14:0] m158_47;
   assign m158_47 =15'b0;

   // m158_48 = W*in
   wire signed [14:0] m158_48;
   assign m158_48 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_49 = W*in
   wire signed [14:0] m158_49;
   assign m158_49 =15'b0;

   // m158_50 = W*in
   wire signed [14:0] m158_50;
   assign m158_50 =15'b0;

   // m158_51 = W*in
   wire signed [14:0] m158_51;
   assign m158_51 =15'b0;

   // m158_52 = W*in
   wire signed [14:0] m158_52;
   assign m158_52 =15'b0;

   // m158_53 = W*in
   wire signed [14:0] m158_53;
   assign m158_53 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_54 = W*in
   wire signed [14:0] m158_54;
   assign m158_54 =15'b0;

   // m158_55 = W*in
   wire signed [14:0] m158_55;
   assign m158_55 =15'b0;

   // m158_56 = W*in
   wire signed [14:0] m158_56;
   assign m158_56 =15'b0;

   // m158_57 = W*in
   wire signed [14:0] m158_57;
   assign m158_57 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_58 = W*in
   wire signed [14:0] m158_58;
   assign m158_58 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_59 = W*in
   wire signed [14:0] m158_59;
   assign m158_59 ={ {4{neg158[14]}} , neg158[14:4] };

   // m158_60 = W*in
   wire signed [14:0] m158_60;
   assign m158_60 =15'b0;

   // m158_61 = W*in
   wire signed [14:0] m158_61;
   assign m158_61 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_62 = W*in
   wire signed [14:0] m158_62;
   assign m158_62 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_63 = W*in
   wire signed [14:0] m158_63;
   assign m158_63 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_64 = W*in
   wire signed [14:0] m158_64;
   assign m158_64 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_65 = W*in
   wire signed [14:0] m158_65;
   assign m158_65 ={ {3{in158[14]}} , in158[14:3] };

   // m158_66 = W*in
   wire signed [14:0] m158_66;
   assign m158_66 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_67 = W*in
   wire signed [14:0] m158_67;
   assign m158_67 =15'b0;

   // m158_68 = W*in
   wire signed [14:0] m158_68;
   assign m158_68 ={ {4{neg158[14]}} , neg158[14:4] };

   // m158_69 = W*in
   wire signed [14:0] m158_69;
   assign m158_69 =15'b0;

   // m158_70 = W*in
   wire signed [14:0] m158_70;
   assign m158_70 =15'b0;

   // m158_71 = W*in
   wire signed [14:0] m158_71;
   assign m158_71 =15'b0;

   // m158_72 = W*in
   wire signed [14:0] m158_72;
   assign m158_72 =15'b0;

   // m158_73 = W*in
   wire signed [14:0] m158_73;
   assign m158_73 =15'b0;

   // m158_74 = W*in
   wire signed [14:0] m158_74;
   assign m158_74 =15'b0;

   // m158_75 = W*in
   wire signed [14:0] m158_75;
   assign m158_75 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_76 = W*in
   wire signed [14:0] m158_76;
   assign m158_76 =15'b0;

   // m158_77 = W*in
   wire signed [14:0] m158_77;
   assign m158_77 ={ {3{in158[14]}} , in158[14:3] };

   // m158_78 = W*in
   wire signed [14:0] m158_78;
   assign m158_78 ={ {3{in158[14]}} , in158[14:3] };

   // m158_79 = W*in
   wire signed [14:0] m158_79;
   assign m158_79 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_80 = W*in
   wire signed [14:0] m158_80;
   assign m158_80 =15'b0;

   // m158_81 = W*in
   wire signed [14:0] m158_81;
   assign m158_81 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_82 = W*in
   wire signed [14:0] m158_82;
   assign m158_82 =15'b0;

   // m158_83 = W*in
   wire signed [14:0] m158_83;
   assign m158_83 =15'b0;

   // m158_84 = W*in
   wire signed [14:0] m158_84;
   assign m158_84 ={ {3{in158[14]}} , in158[14:3] };

   // m158_85 = W*in
   wire signed [14:0] m158_85;
   assign m158_85 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_86 = W*in
   wire signed [14:0] m158_86;
   assign m158_86 =15'b0;

   // m158_87 = W*in
   wire signed [14:0] m158_87;
   assign m158_87 =15'b0;

   // m158_88 = W*in
   wire signed [14:0] m158_88;
   assign m158_88 =15'b0;

   // m158_89 = W*in
   wire signed [14:0] m158_89;
   assign m158_89 =15'b0;

   // m158_90 = W*in
   wire signed [14:0] m158_90;
   assign m158_90 ={ {3{in158[14]}} , in158[14:3] };

   // m158_91 = W*in
   wire signed [14:0] m158_91;
   assign m158_91 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_92 = W*in
   wire signed [14:0] m158_92;
   assign m158_92 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_93 = W*in
   wire signed [14:0] m158_93;
   assign m158_93 =15'b0;

   // m158_94 = W*in
   wire signed [14:0] m158_94;
   assign m158_94 =15'b0;

   // m158_95 = W*in
   wire signed [14:0] m158_95;
   assign m158_95 ={ {3{in158[14]}} , in158[14:3] };

   // m158_96 = W*in
   wire signed [14:0] m158_96;
   assign m158_96 ={ {4{in158[14]}} , in158[14:4] };

   // m158_97 = W*in
   wire signed [14:0] m158_97;
   assign m158_97 =15'b0;

   // m158_98 = W*in
   wire signed [14:0] m158_98;
   assign m158_98 ={ {3{in158[14]}} , in158[14:3] };

   // m158_99 = W*in
   wire signed [14:0] m158_99;
   assign m158_99 ={ {3{neg158[14]}} , neg158[14:3] };

   // m158_100 = W*in
   wire signed [14:0] m158_100;
   assign m158_100 ={ {3{neg158[14]}} , neg158[14:3] };

   // m159_1 = W*in
   wire signed [14:0] m159_1;
   assign m159_1 ={ {3{in159[14]}} , in159[14:3] };

   // m159_2 = W*in
   wire signed [14:0] m159_2;
   assign m159_2 ={ {3{in159[14]}} , in159[14:3] };

   // m159_3 = W*in
   wire signed [14:0] m159_3;
   assign m159_3 =15'b0;

   // m159_4 = W*in
   wire signed [14:0] m159_4;
   assign m159_4 =15'b0;

   // m159_5 = W*in
   wire signed [14:0] m159_5;
   assign m159_5 =15'b0;

   // m159_6 = W*in
   wire signed [14:0] m159_6;
   assign m159_6 =15'b0;

   // m159_7 = W*in
   wire signed [14:0] m159_7;
   assign m159_7 =15'b0;

   // m159_8 = W*in
   wire signed [14:0] m159_8;
   assign m159_8 =15'b0;

   // m159_9 = W*in
   wire signed [14:0] m159_9;
   assign m159_9 ={ {3{in159[14]}} , in159[14:3] };

   // m159_10 = W*in
   wire signed [14:0] m159_10;
   assign m159_10 =15'b0;

   // m159_11 = W*in
   wire signed [14:0] m159_11;
   assign m159_11 =15'b0;

   // m159_12 = W*in
   wire signed [14:0] m159_12;
   assign m159_12 =15'b0;

   // m159_13 = W*in
   wire signed [14:0] m159_13;
   assign m159_13 ={ {3{in159[14]}} , in159[14:3] };

   // m159_14 = W*in
   wire signed [14:0] m159_14;
   assign m159_14 =15'b0;

   // m159_15 = W*in
   wire signed [14:0] m159_15;
   assign m159_15 =15'b0;

   // m159_16 = W*in
   wire signed [14:0] m159_16;
   assign m159_16 =15'b0;

   // m159_17 = W*in
   wire signed [14:0] m159_17;
   assign m159_17 =15'b0;

   // m159_18 = W*in
   wire signed [14:0] m159_18;
   assign m159_18 =15'b0;

   // m159_19 = W*in
   wire signed [14:0] m159_19;
   assign m159_19 ={ {3{in159[14]}} , in159[14:3] };

   // m159_20 = W*in
   wire signed [14:0] m159_20;
   assign m159_20 =15'b0;

   // m159_21 = W*in
   wire signed [14:0] m159_21;
   assign m159_21 ={ {4{in159[14]}} , in159[14:4] };

   // m159_22 = W*in
   wire signed [14:0] m159_22;
   assign m159_22 =15'b0;

   // m159_23 = W*in
   wire signed [14:0] m159_23;
   assign m159_23 =15'b0;

   // m159_24 = W*in
   wire signed [14:0] m159_24;
   assign m159_24 =15'b0;

   // m159_25 = W*in
   wire signed [14:0] m159_25;
   assign m159_25 =15'b0;

   // m159_26 = W*in
   wire signed [14:0] m159_26;
   assign m159_26 =15'b0;

   // m159_27 = W*in
   wire signed [14:0] m159_27;
   assign m159_27 ={ {3{in159[14]}} , in159[14:3] };

   // m159_28 = W*in
   wire signed [14:0] m159_28;
   assign m159_28 =15'b0;

   // m159_29 = W*in
   wire signed [14:0] m159_29;
   assign m159_29 ={ {4{in159[14]}} , in159[14:4] };

   // m159_30 = W*in
   wire signed [14:0] m159_30;
   assign m159_30 =15'b0;

   // m159_31 = W*in
   wire signed [14:0] m159_31;
   assign m159_31 =15'b0;

   // m159_32 = W*in
   wire signed [14:0] m159_32;
   assign m159_32 ={ {3{in159[14]}} , in159[14:3] };

   // m159_33 = W*in
   wire signed [14:0] m159_33;
   assign m159_33 ={ {3{in159[14]}} , in159[14:3] };

   // m159_34 = W*in
   wire signed [14:0] m159_34;
   assign m159_34 ={ {3{in159[14]}} , in159[14:3] };

   // m159_35 = W*in
   wire signed [14:0] m159_35;
   assign m159_35 =15'b0;

   // m159_36 = W*in
   wire signed [14:0] m159_36;
   assign m159_36 =15'b0;

   // m159_37 = W*in
   wire signed [14:0] m159_37;
   assign m159_37 ={ {2{neg159[14]}} , neg159[14:2] };

   // m159_38 = W*in
   wire signed [14:0] m159_38;
   assign m159_38 =15'b0;

   // m159_39 = W*in
   wire signed [14:0] m159_39;
   assign m159_39 =15'b0;

   // m159_40 = W*in
   wire signed [14:0] m159_40;
   assign m159_40 =15'b0;

   // m159_41 = W*in
   wire signed [14:0] m159_41;
   assign m159_41 =15'b0;

   // m159_42 = W*in
   wire signed [14:0] m159_42;
   assign m159_42 =15'b0;

   // m159_43 = W*in
   wire signed [14:0] m159_43;
   assign m159_43 =15'b0;

   // m159_44 = W*in
   wire signed [14:0] m159_44;
   assign m159_44 =15'b0;

   // m159_45 = W*in
   wire signed [14:0] m159_45;
   assign m159_45 =15'b0;

   // m159_46 = W*in
   wire signed [14:0] m159_46;
   assign m159_46 ={ {4{neg159[14]}} , neg159[14:4] };

   // m159_47 = W*in
   wire signed [14:0] m159_47;
   assign m159_47 =15'b0;

   // m159_48 = W*in
   wire signed [14:0] m159_48;
   assign m159_48 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_49 = W*in
   wire signed [14:0] m159_49;
   assign m159_49 =15'b0;

   // m159_50 = W*in
   wire signed [14:0] m159_50;
   assign m159_50 =15'b0;

   // m159_51 = W*in
   wire signed [14:0] m159_51;
   assign m159_51 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_52 = W*in
   wire signed [14:0] m159_52;
   assign m159_52 =15'b0;

   // m159_53 = W*in
   wire signed [14:0] m159_53;
   assign m159_53 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_54 = W*in
   wire signed [14:0] m159_54;
   assign m159_54 =15'b0;

   // m159_55 = W*in
   wire signed [14:0] m159_55;
   assign m159_55 =15'b0;

   // m159_56 = W*in
   wire signed [14:0] m159_56;
   assign m159_56 =15'b0;

   // m159_57 = W*in
   wire signed [14:0] m159_57;
   assign m159_57 =15'b0;

   // m159_58 = W*in
   wire signed [14:0] m159_58;
   assign m159_58 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_59 = W*in
   wire signed [14:0] m159_59;
   assign m159_59 =15'b0;

   // m159_60 = W*in
   wire signed [14:0] m159_60;
   assign m159_60 =15'b0;

   // m159_61 = W*in
   wire signed [14:0] m159_61;
   assign m159_61 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_62 = W*in
   wire signed [14:0] m159_62;
   assign m159_62 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_63 = W*in
   wire signed [14:0] m159_63;
   assign m159_63 =15'b0;

   // m159_64 = W*in
   wire signed [14:0] m159_64;
   assign m159_64 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_65 = W*in
   wire signed [14:0] m159_65;
   assign m159_65 =15'b0;

   // m159_66 = W*in
   wire signed [14:0] m159_66;
   assign m159_66 ={ {4{neg159[14]}} , neg159[14:4] };

   // m159_67 = W*in
   wire signed [14:0] m159_67;
   assign m159_67 =15'b0;

   // m159_68 = W*in
   wire signed [14:0] m159_68;
   assign m159_68 =15'b0;

   // m159_69 = W*in
   wire signed [14:0] m159_69;
   assign m159_69 =15'b0;

   // m159_70 = W*in
   wire signed [14:0] m159_70;
   assign m159_70 ={ {4{in159[14]}} , in159[14:4] };

   // m159_71 = W*in
   wire signed [14:0] m159_71;
   assign m159_71 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_72 = W*in
   wire signed [14:0] m159_72;
   assign m159_72 =15'b0;

   // m159_73 = W*in
   wire signed [14:0] m159_73;
   assign m159_73 =15'b0;

   // m159_74 = W*in
   wire signed [14:0] m159_74;
   assign m159_74 =15'b0;

   // m159_75 = W*in
   wire signed [14:0] m159_75;
   assign m159_75 =15'b0;

   // m159_76 = W*in
   wire signed [14:0] m159_76;
   assign m159_76 =15'b0;

   // m159_77 = W*in
   wire signed [14:0] m159_77;
   assign m159_77 =15'b0;

   // m159_78 = W*in
   wire signed [14:0] m159_78;
   assign m159_78 =15'b0;

   // m159_79 = W*in
   wire signed [14:0] m159_79;
   assign m159_79 =15'b0;

   // m159_80 = W*in
   wire signed [14:0] m159_80;
   assign m159_80 =15'b0;

   // m159_81 = W*in
   wire signed [14:0] m159_81;
   assign m159_81 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_82 = W*in
   wire signed [14:0] m159_82;
   assign m159_82 =15'b0;

   // m159_83 = W*in
   wire signed [14:0] m159_83;
   assign m159_83 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_84 = W*in
   wire signed [14:0] m159_84;
   assign m159_84 =15'b0;

   // m159_85 = W*in
   wire signed [14:0] m159_85;
   assign m159_85 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_86 = W*in
   wire signed [14:0] m159_86;
   assign m159_86 =15'b0;

   // m159_87 = W*in
   wire signed [14:0] m159_87;
   assign m159_87 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_88 = W*in
   wire signed [14:0] m159_88;
   assign m159_88 =15'b0;

   // m159_89 = W*in
   wire signed [14:0] m159_89;
   assign m159_89 ={ {2{neg159[14]}} , neg159[14:2] };

   // m159_90 = W*in
   wire signed [14:0] m159_90;
   assign m159_90 ={ {2{in159[14]}} , in159[14:2] };

   // m159_91 = W*in
   wire signed [14:0] m159_91;
   assign m159_91 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_92 = W*in
   wire signed [14:0] m159_92;
   assign m159_92 =15'b0;

   // m159_93 = W*in
   wire signed [14:0] m159_93;
   assign m159_93 ={ {3{neg159[14]}} , neg159[14:3] };

   // m159_94 = W*in
   wire signed [14:0] m159_94;
   assign m159_94 =15'b0;

   // m159_95 = W*in
   wire signed [14:0] m159_95;
   assign m159_95 =15'b0;

   // m159_96 = W*in
   wire signed [14:0] m159_96;
   assign m159_96 =15'b0;

   // m159_97 = W*in
   wire signed [14:0] m159_97;
   assign m159_97 =15'b0;

   // m159_98 = W*in
   wire signed [14:0] m159_98;
   assign m159_98 =15'b0;

   // m159_99 = W*in
   wire signed [14:0] m159_99;
   assign m159_99 =15'b0;

   // m159_100 = W*in
   wire signed [14:0] m159_100;
   assign m159_100 =15'b0;

   // m160_1 = W*in
   wire signed [14:0] m160_1;
   assign m160_1 =15'b0;

   // m160_2 = W*in
   wire signed [14:0] m160_2;
   assign m160_2 =15'b0;

   // m160_3 = W*in
   wire signed [14:0] m160_3;
   assign m160_3 ={ {3{in160[14]}} , in160[14:3] };

   // m160_4 = W*in
   wire signed [14:0] m160_4;
   assign m160_4 =15'b0;

   // m160_5 = W*in
   wire signed [14:0] m160_5;
   assign m160_5 =15'b0;

   // m160_6 = W*in
   wire signed [14:0] m160_6;
   assign m160_6 =15'b0;

   // m160_7 = W*in
   wire signed [14:0] m160_7;
   assign m160_7 =15'b0;

   // m160_8 = W*in
   wire signed [14:0] m160_8;
   assign m160_8 =15'b0;

   // m160_9 = W*in
   wire signed [14:0] m160_9;
   assign m160_9 ={ {3{neg160[14]}} , neg160[14:3] };

   // m160_10 = W*in
   wire signed [14:0] m160_10;
   assign m160_10 =15'b0;

   // m160_11 = W*in
   wire signed [14:0] m160_11;
   assign m160_11 =15'b0;

   // m160_12 = W*in
   wire signed [14:0] m160_12;
   assign m160_12 =15'b0;

   // m160_13 = W*in
   wire signed [14:0] m160_13;
   assign m160_13 =15'b0;

   // m160_14 = W*in
   wire signed [14:0] m160_14;
   assign m160_14 ={ {3{neg160[14]}} , neg160[14:3] };

   // m160_15 = W*in
   wire signed [14:0] m160_15;
   assign m160_15 =15'b0;

   // m160_16 = W*in
   wire signed [14:0] m160_16;
   assign m160_16 =15'b0;

   // m160_17 = W*in
   wire signed [14:0] m160_17;
   assign m160_17 =15'b0;

   // m160_18 = W*in
   wire signed [14:0] m160_18;
   assign m160_18 =15'b0;

   // m160_19 = W*in
   wire signed [14:0] m160_19;
   assign m160_19 =15'b0;

   // m160_20 = W*in
   wire signed [14:0] m160_20;
   assign m160_20 =15'b0;

   // m160_21 = W*in
   wire signed [14:0] m160_21;
   assign m160_21 =15'b0;

   // m160_22 = W*in
   wire signed [14:0] m160_22;
   assign m160_22 ={ {3{in160[14]}} , in160[14:3] };

   // m160_23 = W*in
   wire signed [14:0] m160_23;
   assign m160_23 =15'b0;

   // m160_24 = W*in
   wire signed [14:0] m160_24;
   assign m160_24 =15'b0;

   // m160_25 = W*in
   wire signed [14:0] m160_25;
   assign m160_25 =15'b0;

   // m160_26 = W*in
   wire signed [14:0] m160_26;
   assign m160_26 =15'b0;

   // m160_27 = W*in
   wire signed [14:0] m160_27;
   assign m160_27 =15'b0;

   // m160_28 = W*in
   wire signed [14:0] m160_28;
   assign m160_28 =15'b0;

   // m160_29 = W*in
   wire signed [14:0] m160_29;
   assign m160_29 =15'b0;

   // m160_30 = W*in
   wire signed [14:0] m160_30;
   assign m160_30 =15'b0;

   // m160_31 = W*in
   wire signed [14:0] m160_31;
   assign m160_31 =15'b0;

   // m160_32 = W*in
   wire signed [14:0] m160_32;
   assign m160_32 =15'b0;

   // m160_33 = W*in
   wire signed [14:0] m160_33;
   assign m160_33 =15'b0;

   // m160_34 = W*in
   wire signed [14:0] m160_34;
   assign m160_34 =15'b0;

   // m160_35 = W*in
   wire signed [14:0] m160_35;
   assign m160_35 =15'b0;

   // m160_36 = W*in
   wire signed [14:0] m160_36;
   assign m160_36 =15'b0;

   // m160_37 = W*in
   wire signed [14:0] m160_37;
   assign m160_37 =15'b0;

   // m160_38 = W*in
   wire signed [14:0] m160_38;
   assign m160_38 =15'b0;

   // m160_39 = W*in
   wire signed [14:0] m160_39;
   assign m160_39 =15'b0;

   // m160_40 = W*in
   wire signed [14:0] m160_40;
   assign m160_40 =15'b0;

   // m160_41 = W*in
   wire signed [14:0] m160_41;
   assign m160_41 =15'b0;

   // m160_42 = W*in
   wire signed [14:0] m160_42;
   assign m160_42 =15'b0;

   // m160_43 = W*in
   wire signed [14:0] m160_43;
   assign m160_43 =15'b0;

   // m160_44 = W*in
   wire signed [14:0] m160_44;
   assign m160_44 =15'b0;

   // m160_45 = W*in
   wire signed [14:0] m160_45;
   assign m160_45 =15'b0;

   // m160_46 = W*in
   wire signed [14:0] m160_46;
   assign m160_46 =15'b0;

   // m160_47 = W*in
   wire signed [14:0] m160_47;
   assign m160_47 =15'b0;

   // m160_48 = W*in
   wire signed [14:0] m160_48;
   assign m160_48 =15'b0;

   // m160_49 = W*in
   wire signed [14:0] m160_49;
   assign m160_49 =15'b0;

   // m160_50 = W*in
   wire signed [14:0] m160_50;
   assign m160_50 =15'b0;

   // m160_51 = W*in
   wire signed [14:0] m160_51;
   assign m160_51 ={ {3{in160[14]}} , in160[14:3] };

   // m160_52 = W*in
   wire signed [14:0] m160_52;
   assign m160_52 =15'b0;

   // m160_53 = W*in
   wire signed [14:0] m160_53;
   assign m160_53 =15'b0;

   // m160_54 = W*in
   wire signed [14:0] m160_54;
   assign m160_54 =15'b0;

   // m160_55 = W*in
   wire signed [14:0] m160_55;
   assign m160_55 =15'b0;

   // m160_56 = W*in
   wire signed [14:0] m160_56;
   assign m160_56 =15'b0;

   // m160_57 = W*in
   wire signed [14:0] m160_57;
   assign m160_57 =15'b0;

   // m160_58 = W*in
   wire signed [14:0] m160_58;
   assign m160_58 ={ {4{in160[14]}} , in160[14:4] };

   // m160_59 = W*in
   wire signed [14:0] m160_59;
   assign m160_59 =15'b0;

   // m160_60 = W*in
   wire signed [14:0] m160_60;
   assign m160_60 =15'b0;

   // m160_61 = W*in
   wire signed [14:0] m160_61;
   assign m160_61 =15'b0;

   // m160_62 = W*in
   wire signed [14:0] m160_62;
   assign m160_62 =15'b0;

   // m160_63 = W*in
   wire signed [14:0] m160_63;
   assign m160_63 =15'b0;

   // m160_64 = W*in
   wire signed [14:0] m160_64;
   assign m160_64 ={ {3{in160[14]}} , in160[14:3] };

   // m160_65 = W*in
   wire signed [14:0] m160_65;
   assign m160_65 =15'b0;

   // m160_66 = W*in
   wire signed [14:0] m160_66;
   assign m160_66 =15'b0;

   // m160_67 = W*in
   wire signed [14:0] m160_67;
   assign m160_67 ={ {3{neg160[14]}} , neg160[14:3] };

   // m160_68 = W*in
   wire signed [14:0] m160_68;
   assign m160_68 =15'b0;

   // m160_69 = W*in
   wire signed [14:0] m160_69;
   assign m160_69 =15'b0;

   // m160_70 = W*in
   wire signed [14:0] m160_70;
   assign m160_70 =15'b0;

   // m160_71 = W*in
   wire signed [14:0] m160_71;
   assign m160_71 =15'b0;

   // m160_72 = W*in
   wire signed [14:0] m160_72;
   assign m160_72 =15'b0;

   // m160_73 = W*in
   wire signed [14:0] m160_73;
   assign m160_73 =15'b0;

   // m160_74 = W*in
   wire signed [14:0] m160_74;
   assign m160_74 =15'b0;

   // m160_75 = W*in
   wire signed [14:0] m160_75;
   assign m160_75 =15'b0;

   // m160_76 = W*in
   wire signed [14:0] m160_76;
   assign m160_76 =15'b0;

   // m160_77 = W*in
   wire signed [14:0] m160_77;
   assign m160_77 =15'b0;

   // m160_78 = W*in
   wire signed [14:0] m160_78;
   assign m160_78 =15'b0;

   // m160_79 = W*in
   wire signed [14:0] m160_79;
   assign m160_79 =15'b0;

   // m160_80 = W*in
   wire signed [14:0] m160_80;
   assign m160_80 =15'b0;

   // m160_81 = W*in
   wire signed [14:0] m160_81;
   assign m160_81 =15'b0;

   // m160_82 = W*in
   wire signed [14:0] m160_82;
   assign m160_82 =15'b0;

   // m160_83 = W*in
   wire signed [14:0] m160_83;
   assign m160_83 =15'b0;

   // m160_84 = W*in
   wire signed [14:0] m160_84;
   assign m160_84 =15'b0;

   // m160_85 = W*in
   wire signed [14:0] m160_85;
   assign m160_85 =15'b0;

   // m160_86 = W*in
   wire signed [14:0] m160_86;
   assign m160_86 =15'b0;

   // m160_87 = W*in
   wire signed [14:0] m160_87;
   assign m160_87 =15'b0;

   // m160_88 = W*in
   wire signed [14:0] m160_88;
   assign m160_88 =15'b0;

   // m160_89 = W*in
   wire signed [14:0] m160_89;
   assign m160_89 ={ {3{in160[14]}} , in160[14:3] };

   // m160_90 = W*in
   wire signed [14:0] m160_90;
   assign m160_90 =15'b0;

   // m160_91 = W*in
   wire signed [14:0] m160_91;
   assign m160_91 =15'b0;

   // m160_92 = W*in
   wire signed [14:0] m160_92;
   assign m160_92 =15'b0;

   // m160_93 = W*in
   wire signed [14:0] m160_93;
   assign m160_93 =15'b0;

   // m160_94 = W*in
   wire signed [14:0] m160_94;
   assign m160_94 ={ {3{neg160[14]}} , neg160[14:3] };

   // m160_95 = W*in
   wire signed [14:0] m160_95;
   assign m160_95 =15'b0;

   // m160_96 = W*in
   wire signed [14:0] m160_96;
   assign m160_96 =15'b0;

   // m160_97 = W*in
   wire signed [14:0] m160_97;
   assign m160_97 =15'b0;

   // m160_98 = W*in
   wire signed [14:0] m160_98;
   assign m160_98 ={ {4{neg160[14]}} , neg160[14:4] };

   // m160_99 = W*in
   wire signed [14:0] m160_99;
   assign m160_99 =15'b0;

   // m160_100 = W*in
   wire signed [14:0] m160_100;
   assign m160_100 =15'b0;

   // m161_1 = W*in
   wire signed [14:0] m161_1;
   assign m161_1 =15'b0;

   // m161_2 = W*in
   wire signed [14:0] m161_2;
   assign m161_2 =15'b0;

   // m161_3 = W*in
   wire signed [14:0] m161_3;
   assign m161_3 =15'b0;

   // m161_4 = W*in
   wire signed [14:0] m161_4;
   assign m161_4 =15'b0;

   // m161_5 = W*in
   wire signed [14:0] m161_5;
   assign m161_5 =15'b0;

   // m161_6 = W*in
   wire signed [14:0] m161_6;
   assign m161_6 ={ {4{neg161[14]}} , neg161[14:4] };

   // m161_7 = W*in
   wire signed [14:0] m161_7;
   assign m161_7 =15'b0;

   // m161_8 = W*in
   wire signed [14:0] m161_8;
   assign m161_8 =15'b0;

   // m161_9 = W*in
   wire signed [14:0] m161_9;
   assign m161_9 =15'b0;

   // m161_10 = W*in
   wire signed [14:0] m161_10;
   assign m161_10 =15'b0;

   // m161_11 = W*in
   wire signed [14:0] m161_11;
   assign m161_11 ={ {3{in161[14]}} , in161[14:3] };

   // m161_12 = W*in
   wire signed [14:0] m161_12;
   assign m161_12 ={ {3{in161[14]}} , in161[14:3] };

   // m161_13 = W*in
   wire signed [14:0] m161_13;
   assign m161_13 =15'b0;

   // m161_14 = W*in
   wire signed [14:0] m161_14;
   assign m161_14 =15'b0;

   // m161_15 = W*in
   wire signed [14:0] m161_15;
   assign m161_15 =15'b0;

   // m161_16 = W*in
   wire signed [14:0] m161_16;
   assign m161_16 =15'b0;

   // m161_17 = W*in
   wire signed [14:0] m161_17;
   assign m161_17 =15'b0;

   // m161_18 = W*in
   wire signed [14:0] m161_18;
   assign m161_18 =15'b0;

   // m161_19 = W*in
   wire signed [14:0] m161_19;
   assign m161_19 ={ {4{neg161[14]}} , neg161[14:4] };

   // m161_20 = W*in
   wire signed [14:0] m161_20;
   assign m161_20 =15'b0;

   // m161_21 = W*in
   wire signed [14:0] m161_21;
   assign m161_21 =15'b0;

   // m161_22 = W*in
   wire signed [14:0] m161_22;
   assign m161_22 =15'b0;

   // m161_23 = W*in
   wire signed [14:0] m161_23;
   assign m161_23 =15'b0;

   // m161_24 = W*in
   wire signed [14:0] m161_24;
   assign m161_24 =15'b0;

   // m161_25 = W*in
   wire signed [14:0] m161_25;
   assign m161_25 =15'b0;

   // m161_26 = W*in
   wire signed [14:0] m161_26;
   assign m161_26 ={ {4{neg161[14]}} , neg161[14:4] };

   // m161_27 = W*in
   wire signed [14:0] m161_27;
   assign m161_27 =15'b0;

   // m161_28 = W*in
   wire signed [14:0] m161_28;
   assign m161_28 =15'b0;

   // m161_29 = W*in
   wire signed [14:0] m161_29;
   assign m161_29 =15'b0;

   // m161_30 = W*in
   wire signed [14:0] m161_30;
   assign m161_30 =15'b0;

   // m161_31 = W*in
   wire signed [14:0] m161_31;
   assign m161_31 =15'b0;

   // m161_32 = W*in
   wire signed [14:0] m161_32;
   assign m161_32 =15'b0;

   // m161_33 = W*in
   wire signed [14:0] m161_33;
   assign m161_33 =15'b0;

   // m161_34 = W*in
   wire signed [14:0] m161_34;
   assign m161_34 =15'b0;

   // m161_35 = W*in
   wire signed [14:0] m161_35;
   assign m161_35 =15'b0;

   // m161_36 = W*in
   wire signed [14:0] m161_36;
   assign m161_36 =15'b0;

   // m161_37 = W*in
   wire signed [14:0] m161_37;
   assign m161_37 =15'b0;

   // m161_38 = W*in
   wire signed [14:0] m161_38;
   assign m161_38 =15'b0;

   // m161_39 = W*in
   wire signed [14:0] m161_39;
   assign m161_39 =15'b0;

   // m161_40 = W*in
   wire signed [14:0] m161_40;
   assign m161_40 =15'b0;

   // m161_41 = W*in
   wire signed [14:0] m161_41;
   assign m161_41 =15'b0;

   // m161_42 = W*in
   wire signed [14:0] m161_42;
   assign m161_42 =15'b0;

   // m161_43 = W*in
   wire signed [14:0] m161_43;
   assign m161_43 =15'b0;

   // m161_44 = W*in
   wire signed [14:0] m161_44;
   assign m161_44 =15'b0;

   // m161_45 = W*in
   wire signed [14:0] m161_45;
   assign m161_45 =15'b0;

   // m161_46 = W*in
   wire signed [14:0] m161_46;
   assign m161_46 =15'b0;

   // m161_47 = W*in
   wire signed [14:0] m161_47;
   assign m161_47 =15'b0;

   // m161_48 = W*in
   wire signed [14:0] m161_48;
   assign m161_48 ={ {3{neg161[14]}} , neg161[14:3] };

   // m161_49 = W*in
   wire signed [14:0] m161_49;
   assign m161_49 =15'b0;

   // m161_50 = W*in
   wire signed [14:0] m161_50;
   assign m161_50 =15'b0;

   // m161_51 = W*in
   wire signed [14:0] m161_51;
   assign m161_51 ={ {3{neg161[14]}} , neg161[14:3] };

   // m161_52 = W*in
   wire signed [14:0] m161_52;
   assign m161_52 =15'b0;

   // m161_53 = W*in
   wire signed [14:0] m161_53;
   assign m161_53 =15'b0;

   // m161_54 = W*in
   wire signed [14:0] m161_54;
   assign m161_54 =15'b0;

   // m161_55 = W*in
   wire signed [14:0] m161_55;
   assign m161_55 =15'b0;

   // m161_56 = W*in
   wire signed [14:0] m161_56;
   assign m161_56 =15'b0;

   // m161_57 = W*in
   wire signed [14:0] m161_57;
   assign m161_57 =15'b0;

   // m161_58 = W*in
   wire signed [14:0] m161_58;
   assign m161_58 ={ {3{neg161[14]}} , neg161[14:3] };

   // m161_59 = W*in
   wire signed [14:0] m161_59;
   assign m161_59 =15'b0;

   // m161_60 = W*in
   wire signed [14:0] m161_60;
   assign m161_60 ={ {3{in161[14]}} , in161[14:3] };

   // m161_61 = W*in
   wire signed [14:0] m161_61;
   assign m161_61 =15'b0;

   // m161_62 = W*in
   wire signed [14:0] m161_62;
   assign m161_62 =15'b0;

   // m161_63 = W*in
   wire signed [14:0] m161_63;
   assign m161_63 =15'b0;

   // m161_64 = W*in
   wire signed [14:0] m161_64;
   assign m161_64 ={ {4{in161[14]}} , in161[14:4] };

   // m161_65 = W*in
   wire signed [14:0] m161_65;
   assign m161_65 =15'b0;

   // m161_66 = W*in
   wire signed [14:0] m161_66;
   assign m161_66 =15'b0;

   // m161_67 = W*in
   wire signed [14:0] m161_67;
   assign m161_67 =15'b0;

   // m161_68 = W*in
   wire signed [14:0] m161_68;
   assign m161_68 =15'b0;

   // m161_69 = W*in
   wire signed [14:0] m161_69;
   assign m161_69 =15'b0;

   // m161_70 = W*in
   wire signed [14:0] m161_70;
   assign m161_70 =15'b0;

   // m161_71 = W*in
   wire signed [14:0] m161_71;
   assign m161_71 =15'b0;

   // m161_72 = W*in
   wire signed [14:0] m161_72;
   assign m161_72 =15'b0;

   // m161_73 = W*in
   wire signed [14:0] m161_73;
   assign m161_73 ={ {3{neg161[14]}} , neg161[14:3] };

   // m161_74 = W*in
   wire signed [14:0] m161_74;
   assign m161_74 =15'b0;

   // m161_75 = W*in
   wire signed [14:0] m161_75;
   assign m161_75 =15'b0;

   // m161_76 = W*in
   wire signed [14:0] m161_76;
   assign m161_76 =15'b0;

   // m161_77 = W*in
   wire signed [14:0] m161_77;
   assign m161_77 =15'b0;

   // m161_78 = W*in
   wire signed [14:0] m161_78;
   assign m161_78 =15'b0;

   // m161_79 = W*in
   wire signed [14:0] m161_79;
   assign m161_79 ={ {4{neg161[14]}} , neg161[14:4] };

   // m161_80 = W*in
   wire signed [14:0] m161_80;
   assign m161_80 =15'b0;

   // m161_81 = W*in
   wire signed [14:0] m161_81;
   assign m161_81 =15'b0;

   // m161_82 = W*in
   wire signed [14:0] m161_82;
   assign m161_82 =15'b0;

   // m161_83 = W*in
   wire signed [14:0] m161_83;
   assign m161_83 =15'b0;

   // m161_84 = W*in
   wire signed [14:0] m161_84;
   assign m161_84 =15'b0;

   // m161_85 = W*in
   wire signed [14:0] m161_85;
   assign m161_85 =15'b0;

   // m161_86 = W*in
   wire signed [14:0] m161_86;
   assign m161_86 =15'b0;

   // m161_87 = W*in
   wire signed [14:0] m161_87;
   assign m161_87 =15'b0;

   // m161_88 = W*in
   wire signed [14:0] m161_88;
   assign m161_88 =15'b0;

   // m161_89 = W*in
   wire signed [14:0] m161_89;
   assign m161_89 =15'b0;

   // m161_90 = W*in
   wire signed [14:0] m161_90;
   assign m161_90 =15'b0;

   // m161_91 = W*in
   wire signed [14:0] m161_91;
   assign m161_91 =15'b0;

   // m161_92 = W*in
   wire signed [14:0] m161_92;
   assign m161_92 =15'b0;

   // m161_93 = W*in
   wire signed [14:0] m161_93;
   assign m161_93 =15'b0;

   // m161_94 = W*in
   wire signed [14:0] m161_94;
   assign m161_94 ={ {3{neg161[14]}} , neg161[14:3] };

   // m161_95 = W*in
   wire signed [14:0] m161_95;
   assign m161_95 =15'b0;

   // m161_96 = W*in
   wire signed [14:0] m161_96;
   assign m161_96 =15'b0;

   // m161_97 = W*in
   wire signed [14:0] m161_97;
   assign m161_97 =15'b0;

   // m161_98 = W*in
   wire signed [14:0] m161_98;
   assign m161_98 =15'b0;

   // m161_99 = W*in
   wire signed [14:0] m161_99;
   assign m161_99 =15'b0;

   // m161_100 = W*in
   wire signed [14:0] m161_100;
   assign m161_100 =15'b0;

   // m162_1 = W*in
   wire signed [14:0] m162_1;
   assign m162_1 =15'b0;

   // m162_2 = W*in
   wire signed [14:0] m162_2;
   assign m162_2 ={ {3{in162[14]}} , in162[14:3] };

   // m162_3 = W*in
   wire signed [14:0] m162_3;
   assign m162_3 ={ {3{in162[14]}} , in162[14:3] };

   // m162_4 = W*in
   wire signed [14:0] m162_4;
   assign m162_4 ={ {4{in162[14]}} , in162[14:4] };

   // m162_5 = W*in
   wire signed [14:0] m162_5;
   assign m162_5 =15'b0;

   // m162_6 = W*in
   wire signed [14:0] m162_6;
   assign m162_6 =15'b0;

   // m162_7 = W*in
   wire signed [14:0] m162_7;
   assign m162_7 =15'b0;

   // m162_8 = W*in
   wire signed [14:0] m162_8;
   assign m162_8 =15'b0;

   // m162_9 = W*in
   wire signed [14:0] m162_9;
   assign m162_9 =15'b0;

   // m162_10 = W*in
   wire signed [14:0] m162_10;
   assign m162_10 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_11 = W*in
   wire signed [14:0] m162_11;
   assign m162_11 =15'b0;

   // m162_12 = W*in
   wire signed [14:0] m162_12;
   assign m162_12 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_13 = W*in
   wire signed [14:0] m162_13;
   assign m162_13 ={ {3{in162[14]}} , in162[14:3] };

   // m162_14 = W*in
   wire signed [14:0] m162_14;
   assign m162_14 =15'b0;

   // m162_15 = W*in
   wire signed [14:0] m162_15;
   assign m162_15 =15'b0;

   // m162_16 = W*in
   wire signed [14:0] m162_16;
   assign m162_16 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_17 = W*in
   wire signed [14:0] m162_17;
   assign m162_17 ={ {3{in162[14]}} , in162[14:3] };

   // m162_18 = W*in
   wire signed [14:0] m162_18;
   assign m162_18 ={ {3{in162[14]}} , in162[14:3] };

   // m162_19 = W*in
   wire signed [14:0] m162_19;
   assign m162_19 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_20 = W*in
   wire signed [14:0] m162_20;
   assign m162_20 ={ {3{in162[14]}} , in162[14:3] };

   // m162_21 = W*in
   wire signed [14:0] m162_21;
   assign m162_21 =15'b0;

   // m162_22 = W*in
   wire signed [14:0] m162_22;
   assign m162_22 =15'b0;

   // m162_23 = W*in
   wire signed [14:0] m162_23;
   assign m162_23 ={ {3{in162[14]}} , in162[14:3] };

   // m162_24 = W*in
   wire signed [14:0] m162_24;
   assign m162_24 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_25 = W*in
   wire signed [14:0] m162_25;
   assign m162_25 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_26 = W*in
   wire signed [14:0] m162_26;
   assign m162_26 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_27 = W*in
   wire signed [14:0] m162_27;
   assign m162_27 ={ {3{in162[14]}} , in162[14:3] };

   // m162_28 = W*in
   wire signed [14:0] m162_28;
   assign m162_28 ={ {3{in162[14]}} , in162[14:3] };

   // m162_29 = W*in
   wire signed [14:0] m162_29;
   assign m162_29 =15'b0;

   // m162_30 = W*in
   wire signed [14:0] m162_30;
   assign m162_30 =15'b0;

   // m162_31 = W*in
   wire signed [14:0] m162_31;
   assign m162_31 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_32 = W*in
   wire signed [14:0] m162_32;
   assign m162_32 =15'b0;

   // m162_33 = W*in
   wire signed [14:0] m162_33;
   assign m162_33 ={ {3{in162[14]}} , in162[14:3] };

   // m162_34 = W*in
   wire signed [14:0] m162_34;
   assign m162_34 =15'b0;

   // m162_35 = W*in
   wire signed [14:0] m162_35;
   assign m162_35 ={ {3{in162[14]}} , in162[14:3] };

   // m162_36 = W*in
   wire signed [14:0] m162_36;
   assign m162_36 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_37 = W*in
   wire signed [14:0] m162_37;
   assign m162_37 =15'b0;

   // m162_38 = W*in
   wire signed [14:0] m162_38;
   assign m162_38 ={ {3{in162[14]}} , in162[14:3] };

   // m162_39 = W*in
   wire signed [14:0] m162_39;
   assign m162_39 ={ {3{in162[14]}} , in162[14:3] };

   // m162_40 = W*in
   wire signed [14:0] m162_40;
   assign m162_40 =15'b0;

   // m162_41 = W*in
   wire signed [14:0] m162_41;
   assign m162_41 =15'b0;

   // m162_42 = W*in
   wire signed [14:0] m162_42;
   assign m162_42 =15'b0;

   // m162_43 = W*in
   wire signed [14:0] m162_43;
   assign m162_43 =15'b0;

   // m162_44 = W*in
   wire signed [14:0] m162_44;
   assign m162_44 =15'b0;

   // m162_45 = W*in
   wire signed [14:0] m162_45;
   assign m162_45 ={ {3{in162[14]}} , in162[14:3] };

   // m162_46 = W*in
   wire signed [14:0] m162_46;
   assign m162_46 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_47 = W*in
   wire signed [14:0] m162_47;
   assign m162_47 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_48 = W*in
   wire signed [14:0] m162_48;
   assign m162_48 ={ {4{neg162[14]}} , neg162[14:4] };

   // m162_49 = W*in
   wire signed [14:0] m162_49;
   assign m162_49 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_50 = W*in
   wire signed [14:0] m162_50;
   assign m162_50 ={ {3{in162[14]}} , in162[14:3] };

   // m162_51 = W*in
   wire signed [14:0] m162_51;
   assign m162_51 =15'b0;

   // m162_52 = W*in
   wire signed [14:0] m162_52;
   assign m162_52 =15'b0;

   // m162_53 = W*in
   wire signed [14:0] m162_53;
   assign m162_53 =15'b0;

   // m162_54 = W*in
   wire signed [14:0] m162_54;
   assign m162_54 =15'b0;

   // m162_55 = W*in
   wire signed [14:0] m162_55;
   assign m162_55 ={ {3{in162[14]}} , in162[14:3] };

   // m162_56 = W*in
   wire signed [14:0] m162_56;
   assign m162_56 =15'b0;

   // m162_57 = W*in
   wire signed [14:0] m162_57;
   assign m162_57 =15'b0;

   // m162_58 = W*in
   wire signed [14:0] m162_58;
   assign m162_58 =15'b0;

   // m162_59 = W*in
   wire signed [14:0] m162_59;
   assign m162_59 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_60 = W*in
   wire signed [14:0] m162_60;
   assign m162_60 =15'b0;

   // m162_61 = W*in
   wire signed [14:0] m162_61;
   assign m162_61 =15'b0;

   // m162_62 = W*in
   wire signed [14:0] m162_62;
   assign m162_62 =15'b0;

   // m162_63 = W*in
   wire signed [14:0] m162_63;
   assign m162_63 =15'b0;

   // m162_64 = W*in
   wire signed [14:0] m162_64;
   assign m162_64 =15'b0;

   // m162_65 = W*in
   wire signed [14:0] m162_65;
   assign m162_65 ={ {4{neg162[14]}} , neg162[14:4] };

   // m162_66 = W*in
   wire signed [14:0] m162_66;
   assign m162_66 ={ {4{neg162[14]}} , neg162[14:4] };

   // m162_67 = W*in
   wire signed [14:0] m162_67;
   assign m162_67 ={ {4{neg162[14]}} , neg162[14:4] };

   // m162_68 = W*in
   wire signed [14:0] m162_68;
   assign m162_68 ={ {3{in162[14]}} , in162[14:3] };

   // m162_69 = W*in
   wire signed [14:0] m162_69;
   assign m162_69 =15'b0;

   // m162_70 = W*in
   wire signed [14:0] m162_70;
   assign m162_70 ={ {3{in162[14]}} , in162[14:3] };

   // m162_71 = W*in
   wire signed [14:0] m162_71;
   assign m162_71 =15'b0;

   // m162_72 = W*in
   wire signed [14:0] m162_72;
   assign m162_72 =15'b0;

   // m162_73 = W*in
   wire signed [14:0] m162_73;
   assign m162_73 =15'b0;

   // m162_74 = W*in
   wire signed [14:0] m162_74;
   assign m162_74 ={ {3{in162[14]}} , in162[14:3] };

   // m162_75 = W*in
   wire signed [14:0] m162_75;
   assign m162_75 =15'b0;

   // m162_76 = W*in
   wire signed [14:0] m162_76;
   assign m162_76 =15'b0;

   // m162_77 = W*in
   wire signed [14:0] m162_77;
   assign m162_77 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_78 = W*in
   wire signed [14:0] m162_78;
   assign m162_78 ={ {3{in162[14]}} , in162[14:3] };

   // m162_79 = W*in
   wire signed [14:0] m162_79;
   assign m162_79 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_80 = W*in
   wire signed [14:0] m162_80;
   assign m162_80 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_81 = W*in
   wire signed [14:0] m162_81;
   assign m162_81 =15'b0;

   // m162_82 = W*in
   wire signed [14:0] m162_82;
   assign m162_82 =15'b0;

   // m162_83 = W*in
   wire signed [14:0] m162_83;
   assign m162_83 =15'b0;

   // m162_84 = W*in
   wire signed [14:0] m162_84;
   assign m162_84 ={ {3{in162[14]}} , in162[14:3] };

   // m162_85 = W*in
   wire signed [14:0] m162_85;
   assign m162_85 =15'b0;

   // m162_86 = W*in
   wire signed [14:0] m162_86;
   assign m162_86 =15'b0;

   // m162_87 = W*in
   wire signed [14:0] m162_87;
   assign m162_87 =15'b0;

   // m162_88 = W*in
   wire signed [14:0] m162_88;
   assign m162_88 =15'b0;

   // m162_89 = W*in
   wire signed [14:0] m162_89;
   assign m162_89 =15'b0;

   // m162_90 = W*in
   wire signed [14:0] m162_90;
   assign m162_90 =15'b0;

   // m162_91 = W*in
   wire signed [14:0] m162_91;
   assign m162_91 =15'b0;

   // m162_92 = W*in
   wire signed [14:0] m162_92;
   assign m162_92 =15'b0;

   // m162_93 = W*in
   wire signed [14:0] m162_93;
   assign m162_93 ={ {3{neg162[14]}} , neg162[14:3] };

   // m162_94 = W*in
   wire signed [14:0] m162_94;
   assign m162_94 ={ {4{in162[14]}} , in162[14:4] };

   // m162_95 = W*in
   wire signed [14:0] m162_95;
   assign m162_95 =15'b0;

   // m162_96 = W*in
   wire signed [14:0] m162_96;
   assign m162_96 =15'b0;

   // m162_97 = W*in
   wire signed [14:0] m162_97;
   assign m162_97 =15'b0;

   // m162_98 = W*in
   wire signed [14:0] m162_98;
   assign m162_98 =15'b0;

   // m162_99 = W*in
   wire signed [14:0] m162_99;
   assign m162_99 =15'b0;

   // m162_100 = W*in
   wire signed [14:0] m162_100;
   assign m162_100 ={ {3{neg162[14]}} , neg162[14:3] };

   // m163_1 = W*in
   wire signed [14:0] m163_1;
   assign m163_1 =15'b0;

   // m163_2 = W*in
   wire signed [14:0] m163_2;
   assign m163_2 =15'b0;

   // m163_3 = W*in
   wire signed [14:0] m163_3;
   assign m163_3 =15'b0;

   // m163_4 = W*in
   wire signed [14:0] m163_4;
   assign m163_4 =15'b0;

   // m163_5 = W*in
   wire signed [14:0] m163_5;
   assign m163_5 =15'b0;

   // m163_6 = W*in
   wire signed [14:0] m163_6;
   assign m163_6 =15'b0;

   // m163_7 = W*in
   wire signed [14:0] m163_7;
   assign m163_7 =15'b0;

   // m163_8 = W*in
   wire signed [14:0] m163_8;
   assign m163_8 =15'b0;

   // m163_9 = W*in
   wire signed [14:0] m163_9;
   assign m163_9 =15'b0;

   // m163_10 = W*in
   wire signed [14:0] m163_10;
   assign m163_10 =15'b0;

   // m163_11 = W*in
   wire signed [14:0] m163_11;
   assign m163_11 =15'b0;

   // m163_12 = W*in
   wire signed [14:0] m163_12;
   assign m163_12 =15'b0;

   // m163_13 = W*in
   wire signed [14:0] m163_13;
   assign m163_13 =15'b0;

   // m163_14 = W*in
   wire signed [14:0] m163_14;
   assign m163_14 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_15 = W*in
   wire signed [14:0] m163_15;
   assign m163_15 =15'b0;

   // m163_16 = W*in
   wire signed [14:0] m163_16;
   assign m163_16 =15'b0;

   // m163_17 = W*in
   wire signed [14:0] m163_17;
   assign m163_17 =15'b0;

   // m163_18 = W*in
   wire signed [14:0] m163_18;
   assign m163_18 =15'b0;

   // m163_19 = W*in
   wire signed [14:0] m163_19;
   assign m163_19 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_20 = W*in
   wire signed [14:0] m163_20;
   assign m163_20 =15'b0;

   // m163_21 = W*in
   wire signed [14:0] m163_21;
   assign m163_21 =15'b0;

   // m163_22 = W*in
   wire signed [14:0] m163_22;
   assign m163_22 ={ {3{in163[14]}} , in163[14:3] };

   // m163_23 = W*in
   wire signed [14:0] m163_23;
   assign m163_23 =15'b0;

   // m163_24 = W*in
   wire signed [14:0] m163_24;
   assign m163_24 =15'b0;

   // m163_25 = W*in
   wire signed [14:0] m163_25;
   assign m163_25 ={ {4{neg163[14]}} , neg163[14:4] };

   // m163_26 = W*in
   wire signed [14:0] m163_26;
   assign m163_26 =15'b0;

   // m163_27 = W*in
   wire signed [14:0] m163_27;
   assign m163_27 ={ {3{in163[14]}} , in163[14:3] };

   // m163_28 = W*in
   wire signed [14:0] m163_28;
   assign m163_28 =15'b0;

   // m163_29 = W*in
   wire signed [14:0] m163_29;
   assign m163_29 =15'b0;

   // m163_30 = W*in
   wire signed [14:0] m163_30;
   assign m163_30 =15'b0;

   // m163_31 = W*in
   wire signed [14:0] m163_31;
   assign m163_31 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_32 = W*in
   wire signed [14:0] m163_32;
   assign m163_32 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_33 = W*in
   wire signed [14:0] m163_33;
   assign m163_33 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_34 = W*in
   wire signed [14:0] m163_34;
   assign m163_34 =15'b0;

   // m163_35 = W*in
   wire signed [14:0] m163_35;
   assign m163_35 =15'b0;

   // m163_36 = W*in
   wire signed [14:0] m163_36;
   assign m163_36 =15'b0;

   // m163_37 = W*in
   wire signed [14:0] m163_37;
   assign m163_37 =15'b0;

   // m163_38 = W*in
   wire signed [14:0] m163_38;
   assign m163_38 =15'b0;

   // m163_39 = W*in
   wire signed [14:0] m163_39;
   assign m163_39 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_40 = W*in
   wire signed [14:0] m163_40;
   assign m163_40 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_41 = W*in
   wire signed [14:0] m163_41;
   assign m163_41 =15'b0;

   // m163_42 = W*in
   wire signed [14:0] m163_42;
   assign m163_42 =15'b0;

   // m163_43 = W*in
   wire signed [14:0] m163_43;
   assign m163_43 =15'b0;

   // m163_44 = W*in
   wire signed [14:0] m163_44;
   assign m163_44 =15'b0;

   // m163_45 = W*in
   wire signed [14:0] m163_45;
   assign m163_45 =15'b0;

   // m163_46 = W*in
   wire signed [14:0] m163_46;
   assign m163_46 =15'b0;

   // m163_47 = W*in
   wire signed [14:0] m163_47;
   assign m163_47 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_48 = W*in
   wire signed [14:0] m163_48;
   assign m163_48 =15'b0;

   // m163_49 = W*in
   wire signed [14:0] m163_49;
   assign m163_49 =15'b0;

   // m163_50 = W*in
   wire signed [14:0] m163_50;
   assign m163_50 =15'b0;

   // m163_51 = W*in
   wire signed [14:0] m163_51;
   assign m163_51 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_52 = W*in
   wire signed [14:0] m163_52;
   assign m163_52 =15'b0;

   // m163_53 = W*in
   wire signed [14:0] m163_53;
   assign m163_53 =15'b0;

   // m163_54 = W*in
   wire signed [14:0] m163_54;
   assign m163_54 =15'b0;

   // m163_55 = W*in
   wire signed [14:0] m163_55;
   assign m163_55 =15'b0;

   // m163_56 = W*in
   wire signed [14:0] m163_56;
   assign m163_56 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_57 = W*in
   wire signed [14:0] m163_57;
   assign m163_57 =15'b0;

   // m163_58 = W*in
   wire signed [14:0] m163_58;
   assign m163_58 =15'b0;

   // m163_59 = W*in
   wire signed [14:0] m163_59;
   assign m163_59 =15'b0;

   // m163_60 = W*in
   wire signed [14:0] m163_60;
   assign m163_60 =15'b0;

   // m163_61 = W*in
   wire signed [14:0] m163_61;
   assign m163_61 =15'b0;

   // m163_62 = W*in
   wire signed [14:0] m163_62;
   assign m163_62 =15'b0;

   // m163_63 = W*in
   wire signed [14:0] m163_63;
   assign m163_63 =15'b0;

   // m163_64 = W*in
   wire signed [14:0] m163_64;
   assign m163_64 =15'b0;

   // m163_65 = W*in
   wire signed [14:0] m163_65;
   assign m163_65 =15'b0;

   // m163_66 = W*in
   wire signed [14:0] m163_66;
   assign m163_66 =15'b0;

   // m163_67 = W*in
   wire signed [14:0] m163_67;
   assign m163_67 =15'b0;

   // m163_68 = W*in
   wire signed [14:0] m163_68;
   assign m163_68 =15'b0;

   // m163_69 = W*in
   wire signed [14:0] m163_69;
   assign m163_69 =15'b0;

   // m163_70 = W*in
   wire signed [14:0] m163_70;
   assign m163_70 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_71 = W*in
   wire signed [14:0] m163_71;
   assign m163_71 =15'b0;

   // m163_72 = W*in
   wire signed [14:0] m163_72;
   assign m163_72 =15'b0;

   // m163_73 = W*in
   wire signed [14:0] m163_73;
   assign m163_73 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_74 = W*in
   wire signed [14:0] m163_74;
   assign m163_74 =15'b0;

   // m163_75 = W*in
   wire signed [14:0] m163_75;
   assign m163_75 =15'b0;

   // m163_76 = W*in
   wire signed [14:0] m163_76;
   assign m163_76 =15'b0;

   // m163_77 = W*in
   wire signed [14:0] m163_77;
   assign m163_77 ={ {3{in163[14]}} , in163[14:3] };

   // m163_78 = W*in
   wire signed [14:0] m163_78;
   assign m163_78 =15'b0;

   // m163_79 = W*in
   wire signed [14:0] m163_79;
   assign m163_79 ={ {4{neg163[14]}} , neg163[14:4] };

   // m163_80 = W*in
   wire signed [14:0] m163_80;
   assign m163_80 =15'b0;

   // m163_81 = W*in
   wire signed [14:0] m163_81;
   assign m163_81 =15'b0;

   // m163_82 = W*in
   wire signed [14:0] m163_82;
   assign m163_82 =15'b0;

   // m163_83 = W*in
   wire signed [14:0] m163_83;
   assign m163_83 =15'b0;

   // m163_84 = W*in
   wire signed [14:0] m163_84;
   assign m163_84 =15'b0;

   // m163_85 = W*in
   wire signed [14:0] m163_85;
   assign m163_85 =15'b0;

   // m163_86 = W*in
   wire signed [14:0] m163_86;
   assign m163_86 =15'b0;

   // m163_87 = W*in
   wire signed [14:0] m163_87;
   assign m163_87 =15'b0;

   // m163_88 = W*in
   wire signed [14:0] m163_88;
   assign m163_88 =15'b0;

   // m163_89 = W*in
   wire signed [14:0] m163_89;
   assign m163_89 =15'b0;

   // m163_90 = W*in
   wire signed [14:0] m163_90;
   assign m163_90 =15'b0;

   // m163_91 = W*in
   wire signed [14:0] m163_91;
   assign m163_91 =15'b0;

   // m163_92 = W*in
   wire signed [14:0] m163_92;
   assign m163_92 =15'b0;

   // m163_93 = W*in
   wire signed [14:0] m163_93;
   assign m163_93 =15'b0;

   // m163_94 = W*in
   wire signed [14:0] m163_94;
   assign m163_94 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_95 = W*in
   wire signed [14:0] m163_95;
   assign m163_95 ={ {3{in163[14]}} , in163[14:3] };

   // m163_96 = W*in
   wire signed [14:0] m163_96;
   assign m163_96 ={ {3{in163[14]}} , in163[14:3] };

   // m163_97 = W*in
   wire signed [14:0] m163_97;
   assign m163_97 =15'b0;

   // m163_98 = W*in
   wire signed [14:0] m163_98;
   assign m163_98 ={ {3{neg163[14]}} , neg163[14:3] };

   // m163_99 = W*in
   wire signed [14:0] m163_99;
   assign m163_99 =15'b0;

   // m163_100 = W*in
   wire signed [14:0] m163_100;
   assign m163_100 =15'b0;

   // m164_1 = W*in
   wire signed [14:0] m164_1;
   assign m164_1 ={ {4{in164[14]}} , in164[14:4] };

   // m164_2 = W*in
   wire signed [14:0] m164_2;
   assign m164_2 =15'b0;

   // m164_3 = W*in
   wire signed [14:0] m164_3;
   assign m164_3 =15'b0;

   // m164_4 = W*in
   wire signed [14:0] m164_4;
   assign m164_4 ={ {4{neg164[14]}} , neg164[14:4] };

   // m164_5 = W*in
   wire signed [14:0] m164_5;
   assign m164_5 =15'b0;

   // m164_6 = W*in
   wire signed [14:0] m164_6;
   assign m164_6 =15'b0;

   // m164_7 = W*in
   wire signed [14:0] m164_7;
   assign m164_7 ={ {2{in164[14]}} , in164[14:2] };

   // m164_8 = W*in
   wire signed [14:0] m164_8;
   assign m164_8 ={ {3{in164[14]}} , in164[14:3] };

   // m164_9 = W*in
   wire signed [14:0] m164_9;
   assign m164_9 =15'b0;

   // m164_10 = W*in
   wire signed [14:0] m164_10;
   assign m164_10 ={ {3{in164[14]}} , in164[14:3] };

   // m164_11 = W*in
   wire signed [14:0] m164_11;
   assign m164_11 =15'b0;

   // m164_12 = W*in
   wire signed [14:0] m164_12;
   assign m164_12 =15'b0;

   // m164_13 = W*in
   wire signed [14:0] m164_13;
   assign m164_13 =15'b0;

   // m164_14 = W*in
   wire signed [14:0] m164_14;
   assign m164_14 =15'b0;

   // m164_15 = W*in
   wire signed [14:0] m164_15;
   assign m164_15 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_16 = W*in
   wire signed [14:0] m164_16;
   assign m164_16 ={ {4{in164[14]}} , in164[14:4] };

   // m164_17 = W*in
   wire signed [14:0] m164_17;
   assign m164_17 =15'b0;

   // m164_18 = W*in
   wire signed [14:0] m164_18;
   assign m164_18 ={ {3{in164[14]}} , in164[14:3] };

   // m164_19 = W*in
   wire signed [14:0] m164_19;
   assign m164_19 ={ {4{neg164[14]}} , neg164[14:4] };

   // m164_20 = W*in
   wire signed [14:0] m164_20;
   assign m164_20 =15'b0;

   // m164_21 = W*in
   wire signed [14:0] m164_21;
   assign m164_21 =15'b0;

   // m164_22 = W*in
   wire signed [14:0] m164_22;
   assign m164_22 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_23 = W*in
   wire signed [14:0] m164_23;
   assign m164_23 ={ {3{in164[14]}} , in164[14:3] };

   // m164_24 = W*in
   wire signed [14:0] m164_24;
   assign m164_24 =15'b0;

   // m164_25 = W*in
   wire signed [14:0] m164_25;
   assign m164_25 =15'b0;

   // m164_26 = W*in
   wire signed [14:0] m164_26;
   assign m164_26 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_27 = W*in
   wire signed [14:0] m164_27;
   assign m164_27 =15'b0;

   // m164_28 = W*in
   wire signed [14:0] m164_28;
   assign m164_28 ={ {3{in164[14]}} , in164[14:3] };

   // m164_29 = W*in
   wire signed [14:0] m164_29;
   assign m164_29 ={ {4{in164[14]}} , in164[14:4] };

   // m164_30 = W*in
   wire signed [14:0] m164_30;
   assign m164_30 ={ {3{in164[14]}} , in164[14:3] };

   // m164_31 = W*in
   wire signed [14:0] m164_31;
   assign m164_31 =15'b0;

   // m164_32 = W*in
   wire signed [14:0] m164_32;
   assign m164_32 ={ {3{in164[14]}} , in164[14:3] };

   // m164_33 = W*in
   wire signed [14:0] m164_33;
   assign m164_33 ={ {4{in164[14]}} , in164[14:4] };

   // m164_34 = W*in
   wire signed [14:0] m164_34;
   assign m164_34 ={ {3{in164[14]}} , in164[14:3] };

   // m164_35 = W*in
   wire signed [14:0] m164_35;
   assign m164_35 =15'b0;

   // m164_36 = W*in
   wire signed [14:0] m164_36;
   assign m164_36 =15'b0;

   // m164_37 = W*in
   wire signed [14:0] m164_37;
   assign m164_37 ={ {3{in164[14]}} , in164[14:3] };

   // m164_38 = W*in
   wire signed [14:0] m164_38;
   assign m164_38 =15'b0;

   // m164_39 = W*in
   wire signed [14:0] m164_39;
   assign m164_39 =15'b0;

   // m164_40 = W*in
   wire signed [14:0] m164_40;
   assign m164_40 =15'b0;

   // m164_41 = W*in
   wire signed [14:0] m164_41;
   assign m164_41 =15'b0;

   // m164_42 = W*in
   wire signed [14:0] m164_42;
   assign m164_42 =15'b0;

   // m164_43 = W*in
   wire signed [14:0] m164_43;
   assign m164_43 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_44 = W*in
   wire signed [14:0] m164_44;
   assign m164_44 ={ {3{in164[14]}} , in164[14:3] };

   // m164_45 = W*in
   wire signed [14:0] m164_45;
   assign m164_45 ={ {3{in164[14]}} , in164[14:3] };

   // m164_46 = W*in
   wire signed [14:0] m164_46;
   assign m164_46 =15'b0;

   // m164_47 = W*in
   wire signed [14:0] m164_47;
   assign m164_47 =15'b0;

   // m164_48 = W*in
   wire signed [14:0] m164_48;
   assign m164_48 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_49 = W*in
   wire signed [14:0] m164_49;
   assign m164_49 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_50 = W*in
   wire signed [14:0] m164_50;
   assign m164_50 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_51 = W*in
   wire signed [14:0] m164_51;
   assign m164_51 ={ {3{in164[14]}} , in164[14:3] };

   // m164_52 = W*in
   wire signed [14:0] m164_52;
   assign m164_52 =15'b0;

   // m164_53 = W*in
   wire signed [14:0] m164_53;
   assign m164_53 =15'b0;

   // m164_54 = W*in
   wire signed [14:0] m164_54;
   assign m164_54 =15'b0;

   // m164_55 = W*in
   wire signed [14:0] m164_55;
   assign m164_55 =15'b0;

   // m164_56 = W*in
   wire signed [14:0] m164_56;
   assign m164_56 =15'b0;

   // m164_57 = W*in
   wire signed [14:0] m164_57;
   assign m164_57 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_58 = W*in
   wire signed [14:0] m164_58;
   assign m164_58 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_59 = W*in
   wire signed [14:0] m164_59;
   assign m164_59 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_60 = W*in
   wire signed [14:0] m164_60;
   assign m164_60 =15'b0;

   // m164_61 = W*in
   wire signed [14:0] m164_61;
   assign m164_61 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_62 = W*in
   wire signed [14:0] m164_62;
   assign m164_62 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_63 = W*in
   wire signed [14:0] m164_63;
   assign m164_63 =15'b0;

   // m164_64 = W*in
   wire signed [14:0] m164_64;
   assign m164_64 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_65 = W*in
   wire signed [14:0] m164_65;
   assign m164_65 ={ {4{in164[14]}} , in164[14:4] };

   // m164_66 = W*in
   wire signed [14:0] m164_66;
   assign m164_66 =15'b0;

   // m164_67 = W*in
   wire signed [14:0] m164_67;
   assign m164_67 =15'b0;

   // m164_68 = W*in
   wire signed [14:0] m164_68;
   assign m164_68 =15'b0;

   // m164_69 = W*in
   wire signed [14:0] m164_69;
   assign m164_69 =15'b0;

   // m164_70 = W*in
   wire signed [14:0] m164_70;
   assign m164_70 =15'b0;

   // m164_71 = W*in
   wire signed [14:0] m164_71;
   assign m164_71 =15'b0;

   // m164_72 = W*in
   wire signed [14:0] m164_72;
   assign m164_72 =15'b0;

   // m164_73 = W*in
   wire signed [14:0] m164_73;
   assign m164_73 =15'b0;

   // m164_74 = W*in
   wire signed [14:0] m164_74;
   assign m164_74 =15'b0;

   // m164_75 = W*in
   wire signed [14:0] m164_75;
   assign m164_75 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_76 = W*in
   wire signed [14:0] m164_76;
   assign m164_76 =15'b0;

   // m164_77 = W*in
   wire signed [14:0] m164_77;
   assign m164_77 ={ {3{in164[14]}} , in164[14:3] };

   // m164_78 = W*in
   wire signed [14:0] m164_78;
   assign m164_78 =15'b0;

   // m164_79 = W*in
   wire signed [14:0] m164_79;
   assign m164_79 =15'b0;

   // m164_80 = W*in
   wire signed [14:0] m164_80;
   assign m164_80 =15'b0;

   // m164_81 = W*in
   wire signed [14:0] m164_81;
   assign m164_81 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_82 = W*in
   wire signed [14:0] m164_82;
   assign m164_82 =15'b0;

   // m164_83 = W*in
   wire signed [14:0] m164_83;
   assign m164_83 ={ {3{in164[14]}} , in164[14:3] };

   // m164_84 = W*in
   wire signed [14:0] m164_84;
   assign m164_84 =15'b0;

   // m164_85 = W*in
   wire signed [14:0] m164_85;
   assign m164_85 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_86 = W*in
   wire signed [14:0] m164_86;
   assign m164_86 =15'b0;

   // m164_87 = W*in
   wire signed [14:0] m164_87;
   assign m164_87 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_88 = W*in
   wire signed [14:0] m164_88;
   assign m164_88 =15'b0;

   // m164_89 = W*in
   wire signed [14:0] m164_89;
   assign m164_89 =15'b0;

   // m164_90 = W*in
   wire signed [14:0] m164_90;
   assign m164_90 =15'b0;

   // m164_91 = W*in
   wire signed [14:0] m164_91;
   assign m164_91 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_92 = W*in
   wire signed [14:0] m164_92;
   assign m164_92 ={ {3{neg164[14]}} , neg164[14:3] };

   // m164_93 = W*in
   wire signed [14:0] m164_93;
   assign m164_93 =15'b0;

   // m164_94 = W*in
   wire signed [14:0] m164_94;
   assign m164_94 ={ {3{in164[14]}} , in164[14:3] };

   // m164_95 = W*in
   wire signed [14:0] m164_95;
   assign m164_95 ={ {3{in164[14]}} , in164[14:3] };

   // m164_96 = W*in
   wire signed [14:0] m164_96;
   assign m164_96 =15'b0;

   // m164_97 = W*in
   wire signed [14:0] m164_97;
   assign m164_97 =15'b0;

   // m164_98 = W*in
   wire signed [14:0] m164_98;
   assign m164_98 =15'b0;

   // m164_99 = W*in
   wire signed [14:0] m164_99;
   assign m164_99 =15'b0;

   // m164_100 = W*in
   wire signed [14:0] m164_100;
   assign m164_100 =15'b0;

   // m165_1 = W*in
   wire signed [14:0] m165_1;
   assign m165_1 =15'b0;

   // m165_2 = W*in
   wire signed [14:0] m165_2;
   assign m165_2 =15'b0;

   // m165_3 = W*in
   wire signed [14:0] m165_3;
   assign m165_3 =15'b0;

   // m165_4 = W*in
   wire signed [14:0] m165_4;
   assign m165_4 ={ {4{in165[14]}} , in165[14:4] };

   // m165_5 = W*in
   wire signed [14:0] m165_5;
   assign m165_5 =15'b0;

   // m165_6 = W*in
   wire signed [14:0] m165_6;
   assign m165_6 =15'b0;

   // m165_7 = W*in
   wire signed [14:0] m165_7;
   assign m165_7 =15'b0;

   // m165_8 = W*in
   wire signed [14:0] m165_8;
   assign m165_8 =15'b0;

   // m165_9 = W*in
   wire signed [14:0] m165_9;
   assign m165_9 =15'b0;

   // m165_10 = W*in
   wire signed [14:0] m165_10;
   assign m165_10 =15'b0;

   // m165_11 = W*in
   wire signed [14:0] m165_11;
   assign m165_11 =15'b0;

   // m165_12 = W*in
   wire signed [14:0] m165_12;
   assign m165_12 =15'b0;

   // m165_13 = W*in
   wire signed [14:0] m165_13;
   assign m165_13 =15'b0;

   // m165_14 = W*in
   wire signed [14:0] m165_14;
   assign m165_14 ={ {3{neg165[14]}} , neg165[14:3] };

   // m165_15 = W*in
   wire signed [14:0] m165_15;
   assign m165_15 =15'b0;

   // m165_16 = W*in
   wire signed [14:0] m165_16;
   assign m165_16 =15'b0;

   // m165_17 = W*in
   wire signed [14:0] m165_17;
   assign m165_17 =15'b0;

   // m165_18 = W*in
   wire signed [14:0] m165_18;
   assign m165_18 =15'b0;

   // m165_19 = W*in
   wire signed [14:0] m165_19;
   assign m165_19 =15'b0;

   // m165_20 = W*in
   wire signed [14:0] m165_20;
   assign m165_20 ={ {3{neg165[14]}} , neg165[14:3] };

   // m165_21 = W*in
   wire signed [14:0] m165_21;
   assign m165_21 =15'b0;

   // m165_22 = W*in
   wire signed [14:0] m165_22;
   assign m165_22 =15'b0;

   // m165_23 = W*in
   wire signed [14:0] m165_23;
   assign m165_23 =15'b0;

   // m165_24 = W*in
   wire signed [14:0] m165_24;
   assign m165_24 =15'b0;

   // m165_25 = W*in
   wire signed [14:0] m165_25;
   assign m165_25 =15'b0;

   // m165_26 = W*in
   wire signed [14:0] m165_26;
   assign m165_26 =15'b0;

   // m165_27 = W*in
   wire signed [14:0] m165_27;
   assign m165_27 =15'b0;

   // m165_28 = W*in
   wire signed [14:0] m165_28;
   assign m165_28 =15'b0;

   // m165_29 = W*in
   wire signed [14:0] m165_29;
   assign m165_29 =15'b0;

   // m165_30 = W*in
   wire signed [14:0] m165_30;
   assign m165_30 =15'b0;

   // m165_31 = W*in
   wire signed [14:0] m165_31;
   assign m165_31 =15'b0;

   // m165_32 = W*in
   wire signed [14:0] m165_32;
   assign m165_32 =15'b0;

   // m165_33 = W*in
   wire signed [14:0] m165_33;
   assign m165_33 =15'b0;

   // m165_34 = W*in
   wire signed [14:0] m165_34;
   assign m165_34 =15'b0;

   // m165_35 = W*in
   wire signed [14:0] m165_35;
   assign m165_35 =15'b0;

   // m165_36 = W*in
   wire signed [14:0] m165_36;
   assign m165_36 =15'b0;

   // m165_37 = W*in
   wire signed [14:0] m165_37;
   assign m165_37 ={ {3{neg165[14]}} , neg165[14:3] };

   // m165_38 = W*in
   wire signed [14:0] m165_38;
   assign m165_38 =15'b0;

   // m165_39 = W*in
   wire signed [14:0] m165_39;
   assign m165_39 =15'b0;

   // m165_40 = W*in
   wire signed [14:0] m165_40;
   assign m165_40 =15'b0;

   // m165_41 = W*in
   wire signed [14:0] m165_41;
   assign m165_41 =15'b0;

   // m165_42 = W*in
   wire signed [14:0] m165_42;
   assign m165_42 =15'b0;

   // m165_43 = W*in
   wire signed [14:0] m165_43;
   assign m165_43 =15'b0;

   // m165_44 = W*in
   wire signed [14:0] m165_44;
   assign m165_44 =15'b0;

   // m165_45 = W*in
   wire signed [14:0] m165_45;
   assign m165_45 ={ {4{in165[14]}} , in165[14:4] };

   // m165_46 = W*in
   wire signed [14:0] m165_46;
   assign m165_46 =15'b0;

   // m165_47 = W*in
   wire signed [14:0] m165_47;
   assign m165_47 =15'b0;

   // m165_48 = W*in
   wire signed [14:0] m165_48;
   assign m165_48 =15'b0;

   // m165_49 = W*in
   wire signed [14:0] m165_49;
   assign m165_49 =15'b0;

   // m165_50 = W*in
   wire signed [14:0] m165_50;
   assign m165_50 =15'b0;

   // m165_51 = W*in
   wire signed [14:0] m165_51;
   assign m165_51 ={ {4{neg165[14]}} , neg165[14:4] };

   // m165_52 = W*in
   wire signed [14:0] m165_52;
   assign m165_52 =15'b0;

   // m165_53 = W*in
   wire signed [14:0] m165_53;
   assign m165_53 =15'b0;

   // m165_54 = W*in
   wire signed [14:0] m165_54;
   assign m165_54 =15'b0;

   // m165_55 = W*in
   wire signed [14:0] m165_55;
   assign m165_55 =15'b0;

   // m165_56 = W*in
   wire signed [14:0] m165_56;
   assign m165_56 =15'b0;

   // m165_57 = W*in
   wire signed [14:0] m165_57;
   assign m165_57 ={ {4{in165[14]}} , in165[14:4] };

   // m165_58 = W*in
   wire signed [14:0] m165_58;
   assign m165_58 =15'b0;

   // m165_59 = W*in
   wire signed [14:0] m165_59;
   assign m165_59 =15'b0;

   // m165_60 = W*in
   wire signed [14:0] m165_60;
   assign m165_60 =15'b0;

   // m165_61 = W*in
   wire signed [14:0] m165_61;
   assign m165_61 =15'b0;

   // m165_62 = W*in
   wire signed [14:0] m165_62;
   assign m165_62 =15'b0;

   // m165_63 = W*in
   wire signed [14:0] m165_63;
   assign m165_63 =15'b0;

   // m165_64 = W*in
   wire signed [14:0] m165_64;
   assign m165_64 =15'b0;

   // m165_65 = W*in
   wire signed [14:0] m165_65;
   assign m165_65 =15'b0;

   // m165_66 = W*in
   wire signed [14:0] m165_66;
   assign m165_66 =15'b0;

   // m165_67 = W*in
   wire signed [14:0] m165_67;
   assign m165_67 =15'b0;

   // m165_68 = W*in
   wire signed [14:0] m165_68;
   assign m165_68 =15'b0;

   // m165_69 = W*in
   wire signed [14:0] m165_69;
   assign m165_69 =15'b0;

   // m165_70 = W*in
   wire signed [14:0] m165_70;
   assign m165_70 =15'b0;

   // m165_71 = W*in
   wire signed [14:0] m165_71;
   assign m165_71 =15'b0;

   // m165_72 = W*in
   wire signed [14:0] m165_72;
   assign m165_72 ={ {3{neg165[14]}} , neg165[14:3] };

   // m165_73 = W*in
   wire signed [14:0] m165_73;
   assign m165_73 =15'b0;

   // m165_74 = W*in
   wire signed [14:0] m165_74;
   assign m165_74 =15'b0;

   // m165_75 = W*in
   wire signed [14:0] m165_75;
   assign m165_75 =15'b0;

   // m165_76 = W*in
   wire signed [14:0] m165_76;
   assign m165_76 =15'b0;

   // m165_77 = W*in
   wire signed [14:0] m165_77;
   assign m165_77 =15'b0;

   // m165_78 = W*in
   wire signed [14:0] m165_78;
   assign m165_78 =15'b0;

   // m165_79 = W*in
   wire signed [14:0] m165_79;
   assign m165_79 =15'b0;

   // m165_80 = W*in
   wire signed [14:0] m165_80;
   assign m165_80 =15'b0;

   // m165_81 = W*in
   wire signed [14:0] m165_81;
   assign m165_81 =15'b0;

   // m165_82 = W*in
   wire signed [14:0] m165_82;
   assign m165_82 =15'b0;

   // m165_83 = W*in
   wire signed [14:0] m165_83;
   assign m165_83 ={ {4{neg165[14]}} , neg165[14:4] };

   // m165_84 = W*in
   wire signed [14:0] m165_84;
   assign m165_84 =15'b0;

   // m165_85 = W*in
   wire signed [14:0] m165_85;
   assign m165_85 =15'b0;

   // m165_86 = W*in
   wire signed [14:0] m165_86;
   assign m165_86 =15'b0;

   // m165_87 = W*in
   wire signed [14:0] m165_87;
   assign m165_87 =15'b0;

   // m165_88 = W*in
   wire signed [14:0] m165_88;
   assign m165_88 =15'b0;

   // m165_89 = W*in
   wire signed [14:0] m165_89;
   assign m165_89 =15'b0;

   // m165_90 = W*in
   wire signed [14:0] m165_90;
   assign m165_90 =15'b0;

   // m165_91 = W*in
   wire signed [14:0] m165_91;
   assign m165_91 =15'b0;

   // m165_92 = W*in
   wire signed [14:0] m165_92;
   assign m165_92 ={ {4{in165[14]}} , in165[14:4] };

   // m165_93 = W*in
   wire signed [14:0] m165_93;
   assign m165_93 =15'b0;

   // m165_94 = W*in
   wire signed [14:0] m165_94;
   assign m165_94 =15'b0;

   // m165_95 = W*in
   wire signed [14:0] m165_95;
   assign m165_95 =15'b0;

   // m165_96 = W*in
   wire signed [14:0] m165_96;
   assign m165_96 =15'b0;

   // m165_97 = W*in
   wire signed [14:0] m165_97;
   assign m165_97 =15'b0;

   // m165_98 = W*in
   wire signed [14:0] m165_98;
   assign m165_98 =15'b0;

   // m165_99 = W*in
   wire signed [14:0] m165_99;
   assign m165_99 =15'b0;

   // m165_100 = W*in
   wire signed [14:0] m165_100;
   assign m165_100 =15'b0;

   // m166_1 = W*in
   wire signed [14:0] m166_1;
   assign m166_1 =15'b0;

   // m166_2 = W*in
   wire signed [14:0] m166_2;
   assign m166_2 =15'b0;

   // m166_3 = W*in
   wire signed [14:0] m166_3;
   assign m166_3 =15'b0;

   // m166_4 = W*in
   wire signed [14:0] m166_4;
   assign m166_4 =15'b0;

   // m166_5 = W*in
   wire signed [14:0] m166_5;
   assign m166_5 =15'b0;

   // m166_6 = W*in
   wire signed [14:0] m166_6;
   assign m166_6 =15'b0;

   // m166_7 = W*in
   wire signed [14:0] m166_7;
   assign m166_7 =15'b0;

   // m166_8 = W*in
   wire signed [14:0] m166_8;
   assign m166_8 =15'b0;

   // m166_9 = W*in
   wire signed [14:0] m166_9;
   assign m166_9 =15'b0;

   // m166_10 = W*in
   wire signed [14:0] m166_10;
   assign m166_10 =15'b0;

   // m166_11 = W*in
   wire signed [14:0] m166_11;
   assign m166_11 =15'b0;

   // m166_12 = W*in
   wire signed [14:0] m166_12;
   assign m166_12 =15'b0;

   // m166_13 = W*in
   wire signed [14:0] m166_13;
   assign m166_13 =15'b0;

   // m166_14 = W*in
   wire signed [14:0] m166_14;
   assign m166_14 =15'b0;

   // m166_15 = W*in
   wire signed [14:0] m166_15;
   assign m166_15 =15'b0;

   // m166_16 = W*in
   wire signed [14:0] m166_16;
   assign m166_16 =15'b0;

   // m166_17 = W*in
   wire signed [14:0] m166_17;
   assign m166_17 =15'b0;

   // m166_18 = W*in
   wire signed [14:0] m166_18;
   assign m166_18 ={ {4{in166[14]}} , in166[14:4] };

   // m166_19 = W*in
   wire signed [14:0] m166_19;
   assign m166_19 =15'b0;

   // m166_20 = W*in
   wire signed [14:0] m166_20;
   assign m166_20 =15'b0;

   // m166_21 = W*in
   wire signed [14:0] m166_21;
   assign m166_21 =15'b0;

   // m166_22 = W*in
   wire signed [14:0] m166_22;
   assign m166_22 ={ {4{neg166[14]}} , neg166[14:4] };

   // m166_23 = W*in
   wire signed [14:0] m166_23;
   assign m166_23 =15'b0;

   // m166_24 = W*in
   wire signed [14:0] m166_24;
   assign m166_24 =15'b0;

   // m166_25 = W*in
   wire signed [14:0] m166_25;
   assign m166_25 =15'b0;

   // m166_26 = W*in
   wire signed [14:0] m166_26;
   assign m166_26 =15'b0;

   // m166_27 = W*in
   wire signed [14:0] m166_27;
   assign m166_27 =15'b0;

   // m166_28 = W*in
   wire signed [14:0] m166_28;
   assign m166_28 =15'b0;

   // m166_29 = W*in
   wire signed [14:0] m166_29;
   assign m166_29 =15'b0;

   // m166_30 = W*in
   wire signed [14:0] m166_30;
   assign m166_30 =15'b0;

   // m166_31 = W*in
   wire signed [14:0] m166_31;
   assign m166_31 =15'b0;

   // m166_32 = W*in
   wire signed [14:0] m166_32;
   assign m166_32 =15'b0;

   // m166_33 = W*in
   wire signed [14:0] m166_33;
   assign m166_33 =15'b0;

   // m166_34 = W*in
   wire signed [14:0] m166_34;
   assign m166_34 =15'b0;

   // m166_35 = W*in
   wire signed [14:0] m166_35;
   assign m166_35 =15'b0;

   // m166_36 = W*in
   wire signed [14:0] m166_36;
   assign m166_36 =15'b0;

   // m166_37 = W*in
   wire signed [14:0] m166_37;
   assign m166_37 =15'b0;

   // m166_38 = W*in
   wire signed [14:0] m166_38;
   assign m166_38 =15'b0;

   // m166_39 = W*in
   wire signed [14:0] m166_39;
   assign m166_39 ={ {3{neg166[14]}} , neg166[14:3] };

   // m166_40 = W*in
   wire signed [14:0] m166_40;
   assign m166_40 =15'b0;

   // m166_41 = W*in
   wire signed [14:0] m166_41;
   assign m166_41 =15'b0;

   // m166_42 = W*in
   wire signed [14:0] m166_42;
   assign m166_42 =15'b0;

   // m166_43 = W*in
   wire signed [14:0] m166_43;
   assign m166_43 =15'b0;

   // m166_44 = W*in
   wire signed [14:0] m166_44;
   assign m166_44 =15'b0;

   // m166_45 = W*in
   wire signed [14:0] m166_45;
   assign m166_45 ={ {4{in166[14]}} , in166[14:4] };

   // m166_46 = W*in
   wire signed [14:0] m166_46;
   assign m166_46 ={ {4{neg166[14]}} , neg166[14:4] };

   // m166_47 = W*in
   wire signed [14:0] m166_47;
   assign m166_47 =15'b0;

   // m166_48 = W*in
   wire signed [14:0] m166_48;
   assign m166_48 =15'b0;

   // m166_49 = W*in
   wire signed [14:0] m166_49;
   assign m166_49 =15'b0;

   // m166_50 = W*in
   wire signed [14:0] m166_50;
   assign m166_50 =15'b0;

   // m166_51 = W*in
   wire signed [14:0] m166_51;
   assign m166_51 =15'b0;

   // m166_52 = W*in
   wire signed [14:0] m166_52;
   assign m166_52 =15'b0;

   // m166_53 = W*in
   wire signed [14:0] m166_53;
   assign m166_53 =15'b0;

   // m166_54 = W*in
   wire signed [14:0] m166_54;
   assign m166_54 =15'b0;

   // m166_55 = W*in
   wire signed [14:0] m166_55;
   assign m166_55 =15'b0;

   // m166_56 = W*in
   wire signed [14:0] m166_56;
   assign m166_56 ={ {4{neg166[14]}} , neg166[14:4] };

   // m166_57 = W*in
   wire signed [14:0] m166_57;
   assign m166_57 =15'b0;

   // m166_58 = W*in
   wire signed [14:0] m166_58;
   assign m166_58 =15'b0;

   // m166_59 = W*in
   wire signed [14:0] m166_59;
   assign m166_59 =15'b0;

   // m166_60 = W*in
   wire signed [14:0] m166_60;
   assign m166_60 =15'b0;

   // m166_61 = W*in
   wire signed [14:0] m166_61;
   assign m166_61 =15'b0;

   // m166_62 = W*in
   wire signed [14:0] m166_62;
   assign m166_62 =15'b0;

   // m166_63 = W*in
   wire signed [14:0] m166_63;
   assign m166_63 =15'b0;

   // m166_64 = W*in
   wire signed [14:0] m166_64;
   assign m166_64 =15'b0;

   // m166_65 = W*in
   wire signed [14:0] m166_65;
   assign m166_65 ={ {4{neg166[14]}} , neg166[14:4] };

   // m166_66 = W*in
   wire signed [14:0] m166_66;
   assign m166_66 =15'b0;

   // m166_67 = W*in
   wire signed [14:0] m166_67;
   assign m166_67 =15'b0;

   // m166_68 = W*in
   wire signed [14:0] m166_68;
   assign m166_68 ={ {4{in166[14]}} , in166[14:4] };

   // m166_69 = W*in
   wire signed [14:0] m166_69;
   assign m166_69 =15'b0;

   // m166_70 = W*in
   wire signed [14:0] m166_70;
   assign m166_70 =15'b0;

   // m166_71 = W*in
   wire signed [14:0] m166_71;
   assign m166_71 =15'b0;

   // m166_72 = W*in
   wire signed [14:0] m166_72;
   assign m166_72 =15'b0;

   // m166_73 = W*in
   wire signed [14:0] m166_73;
   assign m166_73 =15'b0;

   // m166_74 = W*in
   wire signed [14:0] m166_74;
   assign m166_74 ={ {4{neg166[14]}} , neg166[14:4] };

   // m166_75 = W*in
   wire signed [14:0] m166_75;
   assign m166_75 =15'b0;

   // m166_76 = W*in
   wire signed [14:0] m166_76;
   assign m166_76 =15'b0;

   // m166_77 = W*in
   wire signed [14:0] m166_77;
   assign m166_77 =15'b0;

   // m166_78 = W*in
   wire signed [14:0] m166_78;
   assign m166_78 =15'b0;

   // m166_79 = W*in
   wire signed [14:0] m166_79;
   assign m166_79 =15'b0;

   // m166_80 = W*in
   wire signed [14:0] m166_80;
   assign m166_80 =15'b0;

   // m166_81 = W*in
   wire signed [14:0] m166_81;
   assign m166_81 =15'b0;

   // m166_82 = W*in
   wire signed [14:0] m166_82;
   assign m166_82 =15'b0;

   // m166_83 = W*in
   wire signed [14:0] m166_83;
   assign m166_83 =15'b0;

   // m166_84 = W*in
   wire signed [14:0] m166_84;
   assign m166_84 =15'b0;

   // m166_85 = W*in
   wire signed [14:0] m166_85;
   assign m166_85 =15'b0;

   // m166_86 = W*in
   wire signed [14:0] m166_86;
   assign m166_86 =15'b0;

   // m166_87 = W*in
   wire signed [14:0] m166_87;
   assign m166_87 =15'b0;

   // m166_88 = W*in
   wire signed [14:0] m166_88;
   assign m166_88 =15'b0;

   // m166_89 = W*in
   wire signed [14:0] m166_89;
   assign m166_89 =15'b0;

   // m166_90 = W*in
   wire signed [14:0] m166_90;
   assign m166_90 =15'b0;

   // m166_91 = W*in
   wire signed [14:0] m166_91;
   assign m166_91 =15'b0;

   // m166_92 = W*in
   wire signed [14:0] m166_92;
   assign m166_92 =15'b0;

   // m166_93 = W*in
   wire signed [14:0] m166_93;
   assign m166_93 =15'b0;

   // m166_94 = W*in
   wire signed [14:0] m166_94;
   assign m166_94 =15'b0;

   // m166_95 = W*in
   wire signed [14:0] m166_95;
   assign m166_95 =15'b0;

   // m166_96 = W*in
   wire signed [14:0] m166_96;
   assign m166_96 =15'b0;

   // m166_97 = W*in
   wire signed [14:0] m166_97;
   assign m166_97 =15'b0;

   // m166_98 = W*in
   wire signed [14:0] m166_98;
   assign m166_98 =15'b0;

   // m166_99 = W*in
   wire signed [14:0] m166_99;
   assign m166_99 =15'b0;

   // m166_100 = W*in
   wire signed [14:0] m166_100;
   assign m166_100 =15'b0;

   // m167_1 = W*in
   wire signed [14:0] m167_1;
   assign m167_1 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_2 = W*in
   wire signed [14:0] m167_2;
   assign m167_2 =15'b0;

   // m167_3 = W*in
   wire signed [14:0] m167_3;
   assign m167_3 =15'b0;

   // m167_4 = W*in
   wire signed [14:0] m167_4;
   assign m167_4 =15'b0;

   // m167_5 = W*in
   wire signed [14:0] m167_5;
   assign m167_5 =15'b0;

   // m167_6 = W*in
   wire signed [14:0] m167_6;
   assign m167_6 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_7 = W*in
   wire signed [14:0] m167_7;
   assign m167_7 =15'b0;

   // m167_8 = W*in
   wire signed [14:0] m167_8;
   assign m167_8 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_9 = W*in
   wire signed [14:0] m167_9;
   assign m167_9 =15'b0;

   // m167_10 = W*in
   wire signed [14:0] m167_10;
   assign m167_10 =15'b0;

   // m167_11 = W*in
   wire signed [14:0] m167_11;
   assign m167_11 =15'b0;

   // m167_12 = W*in
   wire signed [14:0] m167_12;
   assign m167_12 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_13 = W*in
   wire signed [14:0] m167_13;
   assign m167_13 =15'b0;

   // m167_14 = W*in
   wire signed [14:0] m167_14;
   assign m167_14 =15'b0;

   // m167_15 = W*in
   wire signed [14:0] m167_15;
   assign m167_15 =15'b0;

   // m167_16 = W*in
   wire signed [14:0] m167_16;
   assign m167_16 =15'b0;

   // m167_17 = W*in
   wire signed [14:0] m167_17;
   assign m167_17 ={ {3{in167[14]}} , in167[14:3] };

   // m167_18 = W*in
   wire signed [14:0] m167_18;
   assign m167_18 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_19 = W*in
   wire signed [14:0] m167_19;
   assign m167_19 =15'b0;

   // m167_20 = W*in
   wire signed [14:0] m167_20;
   assign m167_20 =15'b0;

   // m167_21 = W*in
   wire signed [14:0] m167_21;
   assign m167_21 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_22 = W*in
   wire signed [14:0] m167_22;
   assign m167_22 =15'b0;

   // m167_23 = W*in
   wire signed [14:0] m167_23;
   assign m167_23 =15'b0;

   // m167_24 = W*in
   wire signed [14:0] m167_24;
   assign m167_24 =15'b0;

   // m167_25 = W*in
   wire signed [14:0] m167_25;
   assign m167_25 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_26 = W*in
   wire signed [14:0] m167_26;
   assign m167_26 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_27 = W*in
   wire signed [14:0] m167_27;
   assign m167_27 =15'b0;

   // m167_28 = W*in
   wire signed [14:0] m167_28;
   assign m167_28 =15'b0;

   // m167_29 = W*in
   wire signed [14:0] m167_29;
   assign m167_29 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_30 = W*in
   wire signed [14:0] m167_30;
   assign m167_30 =15'b0;

   // m167_31 = W*in
   wire signed [14:0] m167_31;
   assign m167_31 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_32 = W*in
   wire signed [14:0] m167_32;
   assign m167_32 =15'b0;

   // m167_33 = W*in
   wire signed [14:0] m167_33;
   assign m167_33 ={ {4{in167[14]}} , in167[14:4] };

   // m167_34 = W*in
   wire signed [14:0] m167_34;
   assign m167_34 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_35 = W*in
   wire signed [14:0] m167_35;
   assign m167_35 =15'b0;

   // m167_36 = W*in
   wire signed [14:0] m167_36;
   assign m167_36 =15'b0;

   // m167_37 = W*in
   wire signed [14:0] m167_37;
   assign m167_37 =15'b0;

   // m167_38 = W*in
   wire signed [14:0] m167_38;
   assign m167_38 =15'b0;

   // m167_39 = W*in
   wire signed [14:0] m167_39;
   assign m167_39 =15'b0;

   // m167_40 = W*in
   wire signed [14:0] m167_40;
   assign m167_40 =15'b0;

   // m167_41 = W*in
   wire signed [14:0] m167_41;
   assign m167_41 =15'b0;

   // m167_42 = W*in
   wire signed [14:0] m167_42;
   assign m167_42 =15'b0;

   // m167_43 = W*in
   wire signed [14:0] m167_43;
   assign m167_43 =15'b0;

   // m167_44 = W*in
   wire signed [14:0] m167_44;
   assign m167_44 =15'b0;

   // m167_45 = W*in
   wire signed [14:0] m167_45;
   assign m167_45 =15'b0;

   // m167_46 = W*in
   wire signed [14:0] m167_46;
   assign m167_46 =15'b0;

   // m167_47 = W*in
   wire signed [14:0] m167_47;
   assign m167_47 =15'b0;

   // m167_48 = W*in
   wire signed [14:0] m167_48;
   assign m167_48 =15'b0;

   // m167_49 = W*in
   wire signed [14:0] m167_49;
   assign m167_49 =15'b0;

   // m167_50 = W*in
   wire signed [14:0] m167_50;
   assign m167_50 =15'b0;

   // m167_51 = W*in
   wire signed [14:0] m167_51;
   assign m167_51 =15'b0;

   // m167_52 = W*in
   wire signed [14:0] m167_52;
   assign m167_52 =15'b0;

   // m167_53 = W*in
   wire signed [14:0] m167_53;
   assign m167_53 =15'b0;

   // m167_54 = W*in
   wire signed [14:0] m167_54;
   assign m167_54 =15'b0;

   // m167_55 = W*in
   wire signed [14:0] m167_55;
   assign m167_55 =15'b0;

   // m167_56 = W*in
   wire signed [14:0] m167_56;
   assign m167_56 ={ {2{in167[14]}} , in167[14:2] };

   // m167_57 = W*in
   wire signed [14:0] m167_57;
   assign m167_57 =15'b0;

   // m167_58 = W*in
   wire signed [14:0] m167_58;
   assign m167_58 =15'b0;

   // m167_59 = W*in
   wire signed [14:0] m167_59;
   assign m167_59 ={ {4{in167[14]}} , in167[14:4] };

   // m167_60 = W*in
   wire signed [14:0] m167_60;
   assign m167_60 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_61 = W*in
   wire signed [14:0] m167_61;
   assign m167_61 =15'b0;

   // m167_62 = W*in
   wire signed [14:0] m167_62;
   assign m167_62 =15'b0;

   // m167_63 = W*in
   wire signed [14:0] m167_63;
   assign m167_63 =15'b0;

   // m167_64 = W*in
   wire signed [14:0] m167_64;
   assign m167_64 =15'b0;

   // m167_65 = W*in
   wire signed [14:0] m167_65;
   assign m167_65 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_66 = W*in
   wire signed [14:0] m167_66;
   assign m167_66 =15'b0;

   // m167_67 = W*in
   wire signed [14:0] m167_67;
   assign m167_67 =15'b0;

   // m167_68 = W*in
   wire signed [14:0] m167_68;
   assign m167_68 =15'b0;

   // m167_69 = W*in
   wire signed [14:0] m167_69;
   assign m167_69 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_70 = W*in
   wire signed [14:0] m167_70;
   assign m167_70 ={ {3{in167[14]}} , in167[14:3] };

   // m167_71 = W*in
   wire signed [14:0] m167_71;
   assign m167_71 =15'b0;

   // m167_72 = W*in
   wire signed [14:0] m167_72;
   assign m167_72 =15'b0;

   // m167_73 = W*in
   wire signed [14:0] m167_73;
   assign m167_73 =15'b0;

   // m167_74 = W*in
   wire signed [14:0] m167_74;
   assign m167_74 ={ {4{in167[14]}} , in167[14:4] };

   // m167_75 = W*in
   wire signed [14:0] m167_75;
   assign m167_75 =15'b0;

   // m167_76 = W*in
   wire signed [14:0] m167_76;
   assign m167_76 ={ {4{neg167[14]}} , neg167[14:4] };

   // m167_77 = W*in
   wire signed [14:0] m167_77;
   assign m167_77 =15'b0;

   // m167_78 = W*in
   wire signed [14:0] m167_78;
   assign m167_78 =15'b0;

   // m167_79 = W*in
   wire signed [14:0] m167_79;
   assign m167_79 =15'b0;

   // m167_80 = W*in
   wire signed [14:0] m167_80;
   assign m167_80 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_81 = W*in
   wire signed [14:0] m167_81;
   assign m167_81 =15'b0;

   // m167_82 = W*in
   wire signed [14:0] m167_82;
   assign m167_82 =15'b0;

   // m167_83 = W*in
   wire signed [14:0] m167_83;
   assign m167_83 =15'b0;

   // m167_84 = W*in
   wire signed [14:0] m167_84;
   assign m167_84 =15'b0;

   // m167_85 = W*in
   wire signed [14:0] m167_85;
   assign m167_85 =15'b0;

   // m167_86 = W*in
   wire signed [14:0] m167_86;
   assign m167_86 =15'b0;

   // m167_87 = W*in
   wire signed [14:0] m167_87;
   assign m167_87 =15'b0;

   // m167_88 = W*in
   wire signed [14:0] m167_88;
   assign m167_88 =15'b0;

   // m167_89 = W*in
   wire signed [14:0] m167_89;
   assign m167_89 =15'b0;

   // m167_90 = W*in
   wire signed [14:0] m167_90;
   assign m167_90 =15'b0;

   // m167_91 = W*in
   wire signed [14:0] m167_91;
   assign m167_91 =15'b0;

   // m167_92 = W*in
   wire signed [14:0] m167_92;
   assign m167_92 =15'b0;

   // m167_93 = W*in
   wire signed [14:0] m167_93;
   assign m167_93 =15'b0;

   // m167_94 = W*in
   wire signed [14:0] m167_94;
   assign m167_94 ={ {4{in167[14]}} , in167[14:4] };

   // m167_95 = W*in
   wire signed [14:0] m167_95;
   assign m167_95 =15'b0;

   // m167_96 = W*in
   wire signed [14:0] m167_96;
   assign m167_96 ={ {3{neg167[14]}} , neg167[14:3] };

   // m167_97 = W*in
   wire signed [14:0] m167_97;
   assign m167_97 =15'b0;

   // m167_98 = W*in
   wire signed [14:0] m167_98;
   assign m167_98 =15'b0;

   // m167_99 = W*in
   wire signed [14:0] m167_99;
   assign m167_99 ={ {3{in167[14]}} , in167[14:3] };

   // m167_100 = W*in
   wire signed [14:0] m167_100;
   assign m167_100 =15'b0;

   // m168_1 = W*in
   wire signed [14:0] m168_1;
   assign m168_1 ={ {3{in168[14]}} , in168[14:3] };

   // m168_2 = W*in
   wire signed [14:0] m168_2;
   assign m168_2 ={ {3{in168[14]}} , in168[14:3] };

   // m168_3 = W*in
   wire signed [14:0] m168_3;
   assign m168_3 =15'b0;

   // m168_4 = W*in
   wire signed [14:0] m168_4;
   assign m168_4 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_5 = W*in
   wire signed [14:0] m168_5;
   assign m168_5 =15'b0;

   // m168_6 = W*in
   wire signed [14:0] m168_6;
   assign m168_6 =15'b0;

   // m168_7 = W*in
   wire signed [14:0] m168_7;
   assign m168_7 =15'b0;

   // m168_8 = W*in
   wire signed [14:0] m168_8;
   assign m168_8 =15'b0;

   // m168_9 = W*in
   wire signed [14:0] m168_9;
   assign m168_9 =15'b0;

   // m168_10 = W*in
   wire signed [14:0] m168_10;
   assign m168_10 ={ {3{in168[14]}} , in168[14:3] };

   // m168_11 = W*in
   wire signed [14:0] m168_11;
   assign m168_11 =15'b0;

   // m168_12 = W*in
   wire signed [14:0] m168_12;
   assign m168_12 =15'b0;

   // m168_13 = W*in
   wire signed [14:0] m168_13;
   assign m168_13 =15'b0;

   // m168_14 = W*in
   wire signed [14:0] m168_14;
   assign m168_14 =15'b0;

   // m168_15 = W*in
   wire signed [14:0] m168_15;
   assign m168_15 =15'b0;

   // m168_16 = W*in
   wire signed [14:0] m168_16;
   assign m168_16 ={ {3{in168[14]}} , in168[14:3] };

   // m168_17 = W*in
   wire signed [14:0] m168_17;
   assign m168_17 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_18 = W*in
   wire signed [14:0] m168_18;
   assign m168_18 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_19 = W*in
   wire signed [14:0] m168_19;
   assign m168_19 ={ {3{in168[14]}} , in168[14:3] };

   // m168_20 = W*in
   wire signed [14:0] m168_20;
   assign m168_20 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_21 = W*in
   wire signed [14:0] m168_21;
   assign m168_21 =15'b0;

   // m168_22 = W*in
   wire signed [14:0] m168_22;
   assign m168_22 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_23 = W*in
   wire signed [14:0] m168_23;
   assign m168_23 =15'b0;

   // m168_24 = W*in
   wire signed [14:0] m168_24;
   assign m168_24 ={ {3{in168[14]}} , in168[14:3] };

   // m168_25 = W*in
   wire signed [14:0] m168_25;
   assign m168_25 =15'b0;

   // m168_26 = W*in
   wire signed [14:0] m168_26;
   assign m168_26 ={ {3{in168[14]}} , in168[14:3] };

   // m168_27 = W*in
   wire signed [14:0] m168_27;
   assign m168_27 =15'b0;

   // m168_28 = W*in
   wire signed [14:0] m168_28;
   assign m168_28 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_29 = W*in
   wire signed [14:0] m168_29;
   assign m168_29 =15'b0;

   // m168_30 = W*in
   wire signed [14:0] m168_30;
   assign m168_30 =15'b0;

   // m168_31 = W*in
   wire signed [14:0] m168_31;
   assign m168_31 =15'b0;

   // m168_32 = W*in
   wire signed [14:0] m168_32;
   assign m168_32 ={ {3{in168[14]}} , in168[14:3] };

   // m168_33 = W*in
   wire signed [14:0] m168_33;
   assign m168_33 =15'b0;

   // m168_34 = W*in
   wire signed [14:0] m168_34;
   assign m168_34 =15'b0;

   // m168_35 = W*in
   wire signed [14:0] m168_35;
   assign m168_35 =15'b0;

   // m168_36 = W*in
   wire signed [14:0] m168_36;
   assign m168_36 =15'b0;

   // m168_37 = W*in
   wire signed [14:0] m168_37;
   assign m168_37 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_38 = W*in
   wire signed [14:0] m168_38;
   assign m168_38 =15'b0;

   // m168_39 = W*in
   wire signed [14:0] m168_39;
   assign m168_39 =15'b0;

   // m168_40 = W*in
   wire signed [14:0] m168_40;
   assign m168_40 =15'b0;

   // m168_41 = W*in
   wire signed [14:0] m168_41;
   assign m168_41 =15'b0;

   // m168_42 = W*in
   wire signed [14:0] m168_42;
   assign m168_42 ={ {3{in168[14]}} , in168[14:3] };

   // m168_43 = W*in
   wire signed [14:0] m168_43;
   assign m168_43 =15'b0;

   // m168_44 = W*in
   wire signed [14:0] m168_44;
   assign m168_44 =15'b0;

   // m168_45 = W*in
   wire signed [14:0] m168_45;
   assign m168_45 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_46 = W*in
   wire signed [14:0] m168_46;
   assign m168_46 ={ {4{in168[14]}} , in168[14:4] };

   // m168_47 = W*in
   wire signed [14:0] m168_47;
   assign m168_47 ={ {3{in168[14]}} , in168[14:3] };

   // m168_48 = W*in
   wire signed [14:0] m168_48;
   assign m168_48 =15'b0;

   // m168_49 = W*in
   wire signed [14:0] m168_49;
   assign m168_49 =15'b0;

   // m168_50 = W*in
   wire signed [14:0] m168_50;
   assign m168_50 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_51 = W*in
   wire signed [14:0] m168_51;
   assign m168_51 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_52 = W*in
   wire signed [14:0] m168_52;
   assign m168_52 =15'b0;

   // m168_53 = W*in
   wire signed [14:0] m168_53;
   assign m168_53 =15'b0;

   // m168_54 = W*in
   wire signed [14:0] m168_54;
   assign m168_54 =15'b0;

   // m168_55 = W*in
   wire signed [14:0] m168_55;
   assign m168_55 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_56 = W*in
   wire signed [14:0] m168_56;
   assign m168_56 =15'b0;

   // m168_57 = W*in
   wire signed [14:0] m168_57;
   assign m168_57 =15'b0;

   // m168_58 = W*in
   wire signed [14:0] m168_58;
   assign m168_58 =15'b0;

   // m168_59 = W*in
   wire signed [14:0] m168_59;
   assign m168_59 =15'b0;

   // m168_60 = W*in
   wire signed [14:0] m168_60;
   assign m168_60 =15'b0;

   // m168_61 = W*in
   wire signed [14:0] m168_61;
   assign m168_61 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_62 = W*in
   wire signed [14:0] m168_62;
   assign m168_62 =15'b0;

   // m168_63 = W*in
   wire signed [14:0] m168_63;
   assign m168_63 ={ {4{in168[14]}} , in168[14:4] };

   // m168_64 = W*in
   wire signed [14:0] m168_64;
   assign m168_64 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_65 = W*in
   wire signed [14:0] m168_65;
   assign m168_65 ={ {3{in168[14]}} , in168[14:3] };

   // m168_66 = W*in
   wire signed [14:0] m168_66;
   assign m168_66 =15'b0;

   // m168_67 = W*in
   wire signed [14:0] m168_67;
   assign m168_67 =15'b0;

   // m168_68 = W*in
   wire signed [14:0] m168_68;
   assign m168_68 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_69 = W*in
   wire signed [14:0] m168_69;
   assign m168_69 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_70 = W*in
   wire signed [14:0] m168_70;
   assign m168_70 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_71 = W*in
   wire signed [14:0] m168_71;
   assign m168_71 =15'b0;

   // m168_72 = W*in
   wire signed [14:0] m168_72;
   assign m168_72 =15'b0;

   // m168_73 = W*in
   wire signed [14:0] m168_73;
   assign m168_73 =15'b0;

   // m168_74 = W*in
   wire signed [14:0] m168_74;
   assign m168_74 ={ {4{neg168[14]}} , neg168[14:4] };

   // m168_75 = W*in
   wire signed [14:0] m168_75;
   assign m168_75 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_76 = W*in
   wire signed [14:0] m168_76;
   assign m168_76 =15'b0;

   // m168_77 = W*in
   wire signed [14:0] m168_77;
   assign m168_77 =15'b0;

   // m168_78 = W*in
   wire signed [14:0] m168_78;
   assign m168_78 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_79 = W*in
   wire signed [14:0] m168_79;
   assign m168_79 ={ {3{in168[14]}} , in168[14:3] };

   // m168_80 = W*in
   wire signed [14:0] m168_80;
   assign m168_80 =15'b0;

   // m168_81 = W*in
   wire signed [14:0] m168_81;
   assign m168_81 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_82 = W*in
   wire signed [14:0] m168_82;
   assign m168_82 =15'b0;

   // m168_83 = W*in
   wire signed [14:0] m168_83;
   assign m168_83 =15'b0;

   // m168_84 = W*in
   wire signed [14:0] m168_84;
   assign m168_84 =15'b0;

   // m168_85 = W*in
   wire signed [14:0] m168_85;
   assign m168_85 =15'b0;

   // m168_86 = W*in
   wire signed [14:0] m168_86;
   assign m168_86 =15'b0;

   // m168_87 = W*in
   wire signed [14:0] m168_87;
   assign m168_87 =15'b0;

   // m168_88 = W*in
   wire signed [14:0] m168_88;
   assign m168_88 =15'b0;

   // m168_89 = W*in
   wire signed [14:0] m168_89;
   assign m168_89 ={ {3{neg168[14]}} , neg168[14:3] };

   // m168_90 = W*in
   wire signed [14:0] m168_90;
   assign m168_90 =15'b0;

   // m168_91 = W*in
   wire signed [14:0] m168_91;
   assign m168_91 =15'b0;

   // m168_92 = W*in
   wire signed [14:0] m168_92;
   assign m168_92 =15'b0;

   // m168_93 = W*in
   wire signed [14:0] m168_93;
   assign m168_93 =15'b0;

   // m168_94 = W*in
   wire signed [14:0] m168_94;
   assign m168_94 =15'b0;

   // m168_95 = W*in
   wire signed [14:0] m168_95;
   assign m168_95 =15'b0;

   // m168_96 = W*in
   wire signed [14:0] m168_96;
   assign m168_96 =15'b0;

   // m168_97 = W*in
   wire signed [14:0] m168_97;
   assign m168_97 =15'b0;

   // m168_98 = W*in
   wire signed [14:0] m168_98;
   assign m168_98 =15'b0;

   // m168_99 = W*in
   wire signed [14:0] m168_99;
   assign m168_99 =15'b0;

   // m168_100 = W*in
   wire signed [14:0] m168_100;
   assign m168_100 =15'b0;

   // m169_1 = W*in
   wire signed [14:0] m169_1;
   assign m169_1 =15'b0;

   // m169_2 = W*in
   wire signed [14:0] m169_2;
   assign m169_2 =15'b0;

   // m169_3 = W*in
   wire signed [14:0] m169_3;
   assign m169_3 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_4 = W*in
   wire signed [14:0] m169_4;
   assign m169_4 =15'b0;

   // m169_5 = W*in
   wire signed [14:0] m169_5;
   assign m169_5 =15'b0;

   // m169_6 = W*in
   wire signed [14:0] m169_6;
   assign m169_6 =15'b0;

   // m169_7 = W*in
   wire signed [14:0] m169_7;
   assign m169_7 =15'b0;

   // m169_8 = W*in
   wire signed [14:0] m169_8;
   assign m169_8 =15'b0;

   // m169_9 = W*in
   wire signed [14:0] m169_9;
   assign m169_9 =15'b0;

   // m169_10 = W*in
   wire signed [14:0] m169_10;
   assign m169_10 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_11 = W*in
   wire signed [14:0] m169_11;
   assign m169_11 =15'b0;

   // m169_12 = W*in
   wire signed [14:0] m169_12;
   assign m169_12 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_13 = W*in
   wire signed [14:0] m169_13;
   assign m169_13 =15'b0;

   // m169_14 = W*in
   wire signed [14:0] m169_14;
   assign m169_14 =15'b0;

   // m169_15 = W*in
   wire signed [14:0] m169_15;
   assign m169_15 =15'b0;

   // m169_16 = W*in
   wire signed [14:0] m169_16;
   assign m169_16 =15'b0;

   // m169_17 = W*in
   wire signed [14:0] m169_17;
   assign m169_17 =15'b0;

   // m169_18 = W*in
   wire signed [14:0] m169_18;
   assign m169_18 =15'b0;

   // m169_19 = W*in
   wire signed [14:0] m169_19;
   assign m169_19 =15'b0;

   // m169_20 = W*in
   wire signed [14:0] m169_20;
   assign m169_20 =15'b0;

   // m169_21 = W*in
   wire signed [14:0] m169_21;
   assign m169_21 =15'b0;

   // m169_22 = W*in
   wire signed [14:0] m169_22;
   assign m169_22 =15'b0;

   // m169_23 = W*in
   wire signed [14:0] m169_23;
   assign m169_23 =15'b0;

   // m169_24 = W*in
   wire signed [14:0] m169_24;
   assign m169_24 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_25 = W*in
   wire signed [14:0] m169_25;
   assign m169_25 =15'b0;

   // m169_26 = W*in
   wire signed [14:0] m169_26;
   assign m169_26 =15'b0;

   // m169_27 = W*in
   wire signed [14:0] m169_27;
   assign m169_27 =15'b0;

   // m169_28 = W*in
   wire signed [14:0] m169_28;
   assign m169_28 =15'b0;

   // m169_29 = W*in
   wire signed [14:0] m169_29;
   assign m169_29 =15'b0;

   // m169_30 = W*in
   wire signed [14:0] m169_30;
   assign m169_30 ={ {3{in169[14]}} , in169[14:3] };

   // m169_31 = W*in
   wire signed [14:0] m169_31;
   assign m169_31 =15'b0;

   // m169_32 = W*in
   wire signed [14:0] m169_32;
   assign m169_32 ={ {3{in169[14]}} , in169[14:3] };

   // m169_33 = W*in
   wire signed [14:0] m169_33;
   assign m169_33 ={ {4{in169[14]}} , in169[14:4] };

   // m169_34 = W*in
   wire signed [14:0] m169_34;
   assign m169_34 =15'b0;

   // m169_35 = W*in
   wire signed [14:0] m169_35;
   assign m169_35 =15'b0;

   // m169_36 = W*in
   wire signed [14:0] m169_36;
   assign m169_36 =15'b0;

   // m169_37 = W*in
   wire signed [14:0] m169_37;
   assign m169_37 =15'b0;

   // m169_38 = W*in
   wire signed [14:0] m169_38;
   assign m169_38 =15'b0;

   // m169_39 = W*in
   wire signed [14:0] m169_39;
   assign m169_39 =15'b0;

   // m169_40 = W*in
   wire signed [14:0] m169_40;
   assign m169_40 =15'b0;

   // m169_41 = W*in
   wire signed [14:0] m169_41;
   assign m169_41 =15'b0;

   // m169_42 = W*in
   wire signed [14:0] m169_42;
   assign m169_42 =15'b0;

   // m169_43 = W*in
   wire signed [14:0] m169_43;
   assign m169_43 =15'b0;

   // m169_44 = W*in
   wire signed [14:0] m169_44;
   assign m169_44 =15'b0;

   // m169_45 = W*in
   wire signed [14:0] m169_45;
   assign m169_45 =15'b0;

   // m169_46 = W*in
   wire signed [14:0] m169_46;
   assign m169_46 =15'b0;

   // m169_47 = W*in
   wire signed [14:0] m169_47;
   assign m169_47 =15'b0;

   // m169_48 = W*in
   wire signed [14:0] m169_48;
   assign m169_48 =15'b0;

   // m169_49 = W*in
   wire signed [14:0] m169_49;
   assign m169_49 =15'b0;

   // m169_50 = W*in
   wire signed [14:0] m169_50;
   assign m169_50 =15'b0;

   // m169_51 = W*in
   wire signed [14:0] m169_51;
   assign m169_51 =15'b0;

   // m169_52 = W*in
   wire signed [14:0] m169_52;
   assign m169_52 =15'b0;

   // m169_53 = W*in
   wire signed [14:0] m169_53;
   assign m169_53 =15'b0;

   // m169_54 = W*in
   wire signed [14:0] m169_54;
   assign m169_54 =15'b0;

   // m169_55 = W*in
   wire signed [14:0] m169_55;
   assign m169_55 ={ {3{in169[14]}} , in169[14:3] };

   // m169_56 = W*in
   wire signed [14:0] m169_56;
   assign m169_56 =15'b0;

   // m169_57 = W*in
   wire signed [14:0] m169_57;
   assign m169_57 =15'b0;

   // m169_58 = W*in
   wire signed [14:0] m169_58;
   assign m169_58 =15'b0;

   // m169_59 = W*in
   wire signed [14:0] m169_59;
   assign m169_59 ={ {4{neg169[14]}} , neg169[14:4] };

   // m169_60 = W*in
   wire signed [14:0] m169_60;
   assign m169_60 =15'b0;

   // m169_61 = W*in
   wire signed [14:0] m169_61;
   assign m169_61 =15'b0;

   // m169_62 = W*in
   wire signed [14:0] m169_62;
   assign m169_62 =15'b0;

   // m169_63 = W*in
   wire signed [14:0] m169_63;
   assign m169_63 =15'b0;

   // m169_64 = W*in
   wire signed [14:0] m169_64;
   assign m169_64 =15'b0;

   // m169_65 = W*in
   wire signed [14:0] m169_65;
   assign m169_65 =15'b0;

   // m169_66 = W*in
   wire signed [14:0] m169_66;
   assign m169_66 =15'b0;

   // m169_67 = W*in
   wire signed [14:0] m169_67;
   assign m169_67 =15'b0;

   // m169_68 = W*in
   wire signed [14:0] m169_68;
   assign m169_68 ={ {3{in169[14]}} , in169[14:3] };

   // m169_69 = W*in
   wire signed [14:0] m169_69;
   assign m169_69 =15'b0;

   // m169_70 = W*in
   wire signed [14:0] m169_70;
   assign m169_70 =15'b0;

   // m169_71 = W*in
   wire signed [14:0] m169_71;
   assign m169_71 =15'b0;

   // m169_72 = W*in
   wire signed [14:0] m169_72;
   assign m169_72 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_73 = W*in
   wire signed [14:0] m169_73;
   assign m169_73 =15'b0;

   // m169_74 = W*in
   wire signed [14:0] m169_74;
   assign m169_74 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_75 = W*in
   wire signed [14:0] m169_75;
   assign m169_75 =15'b0;

   // m169_76 = W*in
   wire signed [14:0] m169_76;
   assign m169_76 =15'b0;

   // m169_77 = W*in
   wire signed [14:0] m169_77;
   assign m169_77 =15'b0;

   // m169_78 = W*in
   wire signed [14:0] m169_78;
   assign m169_78 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_79 = W*in
   wire signed [14:0] m169_79;
   assign m169_79 =15'b0;

   // m169_80 = W*in
   wire signed [14:0] m169_80;
   assign m169_80 =15'b0;

   // m169_81 = W*in
   wire signed [14:0] m169_81;
   assign m169_81 =15'b0;

   // m169_82 = W*in
   wire signed [14:0] m169_82;
   assign m169_82 =15'b0;

   // m169_83 = W*in
   wire signed [14:0] m169_83;
   assign m169_83 =15'b0;

   // m169_84 = W*in
   wire signed [14:0] m169_84;
   assign m169_84 =15'b0;

   // m169_85 = W*in
   wire signed [14:0] m169_85;
   assign m169_85 =15'b0;

   // m169_86 = W*in
   wire signed [14:0] m169_86;
   assign m169_86 =15'b0;

   // m169_87 = W*in
   wire signed [14:0] m169_87;
   assign m169_87 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_88 = W*in
   wire signed [14:0] m169_88;
   assign m169_88 =15'b0;

   // m169_89 = W*in
   wire signed [14:0] m169_89;
   assign m169_89 =15'b0;

   // m169_90 = W*in
   wire signed [14:0] m169_90;
   assign m169_90 =15'b0;

   // m169_91 = W*in
   wire signed [14:0] m169_91;
   assign m169_91 =15'b0;

   // m169_92 = W*in
   wire signed [14:0] m169_92;
   assign m169_92 =15'b0;

   // m169_93 = W*in
   wire signed [14:0] m169_93;
   assign m169_93 ={ {3{neg169[14]}} , neg169[14:3] };

   // m169_94 = W*in
   wire signed [14:0] m169_94;
   assign m169_94 ={ {3{in169[14]}} , in169[14:3] };

   // m169_95 = W*in
   wire signed [14:0] m169_95;
   assign m169_95 =15'b0;

   // m169_96 = W*in
   wire signed [14:0] m169_96;
   assign m169_96 =15'b0;

   // m169_97 = W*in
   wire signed [14:0] m169_97;
   assign m169_97 =15'b0;

   // m169_98 = W*in
   wire signed [14:0] m169_98;
   assign m169_98 =15'b0;

   // m169_99 = W*in
   wire signed [14:0] m169_99;
   assign m169_99 =15'b0;

   // m169_100 = W*in
   wire signed [14:0] m169_100;
   assign m169_100 =15'b0;

   // m170_1 = W*in
   wire signed [14:0] m170_1;
   assign m170_1 =15'b0;

   // m170_2 = W*in
   wire signed [14:0] m170_2;
   assign m170_2 =15'b0;

   // m170_3 = W*in
   wire signed [14:0] m170_3;
   assign m170_3 =15'b0;

   // m170_4 = W*in
   wire signed [14:0] m170_4;
   assign m170_4 =15'b0;

   // m170_5 = W*in
   wire signed [14:0] m170_5;
   assign m170_5 =15'b0;

   // m170_6 = W*in
   wire signed [14:0] m170_6;
   assign m170_6 =15'b0;

   // m170_7 = W*in
   wire signed [14:0] m170_7;
   assign m170_7 =15'b0;

   // m170_8 = W*in
   wire signed [14:0] m170_8;
   assign m170_8 =15'b0;

   // m170_9 = W*in
   wire signed [14:0] m170_9;
   assign m170_9 =15'b0;

   // m170_10 = W*in
   wire signed [14:0] m170_10;
   assign m170_10 =15'b0;

   // m170_11 = W*in
   wire signed [14:0] m170_11;
   assign m170_11 ={ {3{neg170[14]}} , neg170[14:3] };

   // m170_12 = W*in
   wire signed [14:0] m170_12;
   assign m170_12 =15'b0;

   // m170_13 = W*in
   wire signed [14:0] m170_13;
   assign m170_13 =15'b0;

   // m170_14 = W*in
   wire signed [14:0] m170_14;
   assign m170_14 =15'b0;

   // m170_15 = W*in
   wire signed [14:0] m170_15;
   assign m170_15 =15'b0;

   // m170_16 = W*in
   wire signed [14:0] m170_16;
   assign m170_16 =15'b0;

   // m170_17 = W*in
   wire signed [14:0] m170_17;
   assign m170_17 =15'b0;

   // m170_18 = W*in
   wire signed [14:0] m170_18;
   assign m170_18 =15'b0;

   // m170_19 = W*in
   wire signed [14:0] m170_19;
   assign m170_19 =15'b0;

   // m170_20 = W*in
   wire signed [14:0] m170_20;
   assign m170_20 =15'b0;

   // m170_21 = W*in
   wire signed [14:0] m170_21;
   assign m170_21 =15'b0;

   // m170_22 = W*in
   wire signed [14:0] m170_22;
   assign m170_22 =15'b0;

   // m170_23 = W*in
   wire signed [14:0] m170_23;
   assign m170_23 =15'b0;

   // m170_24 = W*in
   wire signed [14:0] m170_24;
   assign m170_24 =15'b0;

   // m170_25 = W*in
   wire signed [14:0] m170_25;
   assign m170_25 =15'b0;

   // m170_26 = W*in
   wire signed [14:0] m170_26;
   assign m170_26 =15'b0;

   // m170_27 = W*in
   wire signed [14:0] m170_27;
   assign m170_27 =15'b0;

   // m170_28 = W*in
   wire signed [14:0] m170_28;
   assign m170_28 =15'b0;

   // m170_29 = W*in
   wire signed [14:0] m170_29;
   assign m170_29 =15'b0;

   // m170_30 = W*in
   wire signed [14:0] m170_30;
   assign m170_30 ={ {3{neg170[14]}} , neg170[14:3] };

   // m170_31 = W*in
   wire signed [14:0] m170_31;
   assign m170_31 =15'b0;

   // m170_32 = W*in
   wire signed [14:0] m170_32;
   assign m170_32 =15'b0;

   // m170_33 = W*in
   wire signed [14:0] m170_33;
   assign m170_33 ={ {4{neg170[14]}} , neg170[14:4] };

   // m170_34 = W*in
   wire signed [14:0] m170_34;
   assign m170_34 =15'b0;

   // m170_35 = W*in
   wire signed [14:0] m170_35;
   assign m170_35 =15'b0;

   // m170_36 = W*in
   wire signed [14:0] m170_36;
   assign m170_36 =15'b0;

   // m170_37 = W*in
   wire signed [14:0] m170_37;
   assign m170_37 =15'b0;

   // m170_38 = W*in
   wire signed [14:0] m170_38;
   assign m170_38 =15'b0;

   // m170_39 = W*in
   wire signed [14:0] m170_39;
   assign m170_39 =15'b0;

   // m170_40 = W*in
   wire signed [14:0] m170_40;
   assign m170_40 =15'b0;

   // m170_41 = W*in
   wire signed [14:0] m170_41;
   assign m170_41 =15'b0;

   // m170_42 = W*in
   wire signed [14:0] m170_42;
   assign m170_42 =15'b0;

   // m170_43 = W*in
   wire signed [14:0] m170_43;
   assign m170_43 =15'b0;

   // m170_44 = W*in
   wire signed [14:0] m170_44;
   assign m170_44 =15'b0;

   // m170_45 = W*in
   wire signed [14:0] m170_45;
   assign m170_45 =15'b0;

   // m170_46 = W*in
   wire signed [14:0] m170_46;
   assign m170_46 =15'b0;

   // m170_47 = W*in
   wire signed [14:0] m170_47;
   assign m170_47 =15'b0;

   // m170_48 = W*in
   wire signed [14:0] m170_48;
   assign m170_48 =15'b0;

   // m170_49 = W*in
   wire signed [14:0] m170_49;
   assign m170_49 =15'b0;

   // m170_50 = W*in
   wire signed [14:0] m170_50;
   assign m170_50 =15'b0;

   // m170_51 = W*in
   wire signed [14:0] m170_51;
   assign m170_51 ={ {4{in170[14]}} , in170[14:4] };

   // m170_52 = W*in
   wire signed [14:0] m170_52;
   assign m170_52 =15'b0;

   // m170_53 = W*in
   wire signed [14:0] m170_53;
   assign m170_53 ={ {3{neg170[14]}} , neg170[14:3] };

   // m170_54 = W*in
   wire signed [14:0] m170_54;
   assign m170_54 =15'b0;

   // m170_55 = W*in
   wire signed [14:0] m170_55;
   assign m170_55 =15'b0;

   // m170_56 = W*in
   wire signed [14:0] m170_56;
   assign m170_56 =15'b0;

   // m170_57 = W*in
   wire signed [14:0] m170_57;
   assign m170_57 =15'b0;

   // m170_58 = W*in
   wire signed [14:0] m170_58;
   assign m170_58 =15'b0;

   // m170_59 = W*in
   wire signed [14:0] m170_59;
   assign m170_59 ={ {4{in170[14]}} , in170[14:4] };

   // m170_60 = W*in
   wire signed [14:0] m170_60;
   assign m170_60 =15'b0;

   // m170_61 = W*in
   wire signed [14:0] m170_61;
   assign m170_61 =15'b0;

   // m170_62 = W*in
   wire signed [14:0] m170_62;
   assign m170_62 =15'b0;

   // m170_63 = W*in
   wire signed [14:0] m170_63;
   assign m170_63 =15'b0;

   // m170_64 = W*in
   wire signed [14:0] m170_64;
   assign m170_64 =15'b0;

   // m170_65 = W*in
   wire signed [14:0] m170_65;
   assign m170_65 =15'b0;

   // m170_66 = W*in
   wire signed [14:0] m170_66;
   assign m170_66 =15'b0;

   // m170_67 = W*in
   wire signed [14:0] m170_67;
   assign m170_67 ={ {3{neg170[14]}} , neg170[14:3] };

   // m170_68 = W*in
   wire signed [14:0] m170_68;
   assign m170_68 =15'b0;

   // m170_69 = W*in
   wire signed [14:0] m170_69;
   assign m170_69 =15'b0;

   // m170_70 = W*in
   wire signed [14:0] m170_70;
   assign m170_70 =15'b0;

   // m170_71 = W*in
   wire signed [14:0] m170_71;
   assign m170_71 ={ {3{in170[14]}} , in170[14:3] };

   // m170_72 = W*in
   wire signed [14:0] m170_72;
   assign m170_72 =15'b0;

   // m170_73 = W*in
   wire signed [14:0] m170_73;
   assign m170_73 =15'b0;

   // m170_74 = W*in
   wire signed [14:0] m170_74;
   assign m170_74 =15'b0;

   // m170_75 = W*in
   wire signed [14:0] m170_75;
   assign m170_75 =15'b0;

   // m170_76 = W*in
   wire signed [14:0] m170_76;
   assign m170_76 ={ {4{neg170[14]}} , neg170[14:4] };

   // m170_77 = W*in
   wire signed [14:0] m170_77;
   assign m170_77 =15'b0;

   // m170_78 = W*in
   wire signed [14:0] m170_78;
   assign m170_78 =15'b0;

   // m170_79 = W*in
   wire signed [14:0] m170_79;
   assign m170_79 =15'b0;

   // m170_80 = W*in
   wire signed [14:0] m170_80;
   assign m170_80 =15'b0;

   // m170_81 = W*in
   wire signed [14:0] m170_81;
   assign m170_81 ={ {4{neg170[14]}} , neg170[14:4] };

   // m170_82 = W*in
   wire signed [14:0] m170_82;
   assign m170_82 =15'b0;

   // m170_83 = W*in
   wire signed [14:0] m170_83;
   assign m170_83 ={ {3{in170[14]}} , in170[14:3] };

   // m170_84 = W*in
   wire signed [14:0] m170_84;
   assign m170_84 =15'b0;

   // m170_85 = W*in
   wire signed [14:0] m170_85;
   assign m170_85 =15'b0;

   // m170_86 = W*in
   wire signed [14:0] m170_86;
   assign m170_86 =15'b0;

   // m170_87 = W*in
   wire signed [14:0] m170_87;
   assign m170_87 =15'b0;

   // m170_88 = W*in
   wire signed [14:0] m170_88;
   assign m170_88 =15'b0;

   // m170_89 = W*in
   wire signed [14:0] m170_89;
   assign m170_89 =15'b0;

   // m170_90 = W*in
   wire signed [14:0] m170_90;
   assign m170_90 =15'b0;

   // m170_91 = W*in
   wire signed [14:0] m170_91;
   assign m170_91 =15'b0;

   // m170_92 = W*in
   wire signed [14:0] m170_92;
   assign m170_92 =15'b0;

   // m170_93 = W*in
   wire signed [14:0] m170_93;
   assign m170_93 =15'b0;

   // m170_94 = W*in
   wire signed [14:0] m170_94;
   assign m170_94 =15'b0;

   // m170_95 = W*in
   wire signed [14:0] m170_95;
   assign m170_95 =15'b0;

   // m170_96 = W*in
   wire signed [14:0] m170_96;
   assign m170_96 =15'b0;

   // m170_97 = W*in
   wire signed [14:0] m170_97;
   assign m170_97 =15'b0;

   // m170_98 = W*in
   wire signed [14:0] m170_98;
   assign m170_98 =15'b0;

   // m170_99 = W*in
   wire signed [14:0] m170_99;
   assign m170_99 =15'b0;

   // m170_100 = W*in
   wire signed [14:0] m170_100;
   assign m170_100 =15'b0;

   // m171_1 = W*in
   wire signed [14:0] m171_1;
   assign m171_1 =15'b0;

   // m171_2 = W*in
   wire signed [14:0] m171_2;
   assign m171_2 =15'b0;

   // m171_3 = W*in
   wire signed [14:0] m171_3;
   assign m171_3 =15'b0;

   // m171_4 = W*in
   wire signed [14:0] m171_4;
   assign m171_4 ={ {3{in171[14]}} , in171[14:3] };

   // m171_5 = W*in
   wire signed [14:0] m171_5;
   assign m171_5 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_6 = W*in
   wire signed [14:0] m171_6;
   assign m171_6 =15'b0;

   // m171_7 = W*in
   wire signed [14:0] m171_7;
   assign m171_7 =15'b0;

   // m171_8 = W*in
   wire signed [14:0] m171_8;
   assign m171_8 =15'b0;

   // m171_9 = W*in
   wire signed [14:0] m171_9;
   assign m171_9 =15'b0;

   // m171_10 = W*in
   wire signed [14:0] m171_10;
   assign m171_10 =15'b0;

   // m171_11 = W*in
   wire signed [14:0] m171_11;
   assign m171_11 =15'b0;

   // m171_12 = W*in
   wire signed [14:0] m171_12;
   assign m171_12 =15'b0;

   // m171_13 = W*in
   wire signed [14:0] m171_13;
   assign m171_13 =15'b0;

   // m171_14 = W*in
   wire signed [14:0] m171_14;
   assign m171_14 =15'b0;

   // m171_15 = W*in
   wire signed [14:0] m171_15;
   assign m171_15 =15'b0;

   // m171_16 = W*in
   wire signed [14:0] m171_16;
   assign m171_16 =15'b0;

   // m171_17 = W*in
   wire signed [14:0] m171_17;
   assign m171_17 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_18 = W*in
   wire signed [14:0] m171_18;
   assign m171_18 =15'b0;

   // m171_19 = W*in
   wire signed [14:0] m171_19;
   assign m171_19 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_20 = W*in
   wire signed [14:0] m171_20;
   assign m171_20 =15'b0;

   // m171_21 = W*in
   wire signed [14:0] m171_21;
   assign m171_21 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_22 = W*in
   wire signed [14:0] m171_22;
   assign m171_22 =15'b0;

   // m171_23 = W*in
   wire signed [14:0] m171_23;
   assign m171_23 =15'b0;

   // m171_24 = W*in
   wire signed [14:0] m171_24;
   assign m171_24 =15'b0;

   // m171_25 = W*in
   wire signed [14:0] m171_25;
   assign m171_25 =15'b0;

   // m171_26 = W*in
   wire signed [14:0] m171_26;
   assign m171_26 ={ {3{in171[14]}} , in171[14:3] };

   // m171_27 = W*in
   wire signed [14:0] m171_27;
   assign m171_27 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_28 = W*in
   wire signed [14:0] m171_28;
   assign m171_28 ={ {4{neg171[14]}} , neg171[14:4] };

   // m171_29 = W*in
   wire signed [14:0] m171_29;
   assign m171_29 ={ {3{in171[14]}} , in171[14:3] };

   // m171_30 = W*in
   wire signed [14:0] m171_30;
   assign m171_30 =15'b0;

   // m171_31 = W*in
   wire signed [14:0] m171_31;
   assign m171_31 ={ {3{in171[14]}} , in171[14:3] };

   // m171_32 = W*in
   wire signed [14:0] m171_32;
   assign m171_32 =15'b0;

   // m171_33 = W*in
   wire signed [14:0] m171_33;
   assign m171_33 =15'b0;

   // m171_34 = W*in
   wire signed [14:0] m171_34;
   assign m171_34 =15'b0;

   // m171_35 = W*in
   wire signed [14:0] m171_35;
   assign m171_35 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_36 = W*in
   wire signed [14:0] m171_36;
   assign m171_36 =15'b0;

   // m171_37 = W*in
   wire signed [14:0] m171_37;
   assign m171_37 =15'b0;

   // m171_38 = W*in
   wire signed [14:0] m171_38;
   assign m171_38 =15'b0;

   // m171_39 = W*in
   wire signed [14:0] m171_39;
   assign m171_39 =15'b0;

   // m171_40 = W*in
   wire signed [14:0] m171_40;
   assign m171_40 =15'b0;

   // m171_41 = W*in
   wire signed [14:0] m171_41;
   assign m171_41 =15'b0;

   // m171_42 = W*in
   wire signed [14:0] m171_42;
   assign m171_42 =15'b0;

   // m171_43 = W*in
   wire signed [14:0] m171_43;
   assign m171_43 =15'b0;

   // m171_44 = W*in
   wire signed [14:0] m171_44;
   assign m171_44 =15'b0;

   // m171_45 = W*in
   wire signed [14:0] m171_45;
   assign m171_45 =15'b0;

   // m171_46 = W*in
   wire signed [14:0] m171_46;
   assign m171_46 =15'b0;

   // m171_47 = W*in
   wire signed [14:0] m171_47;
   assign m171_47 =15'b0;

   // m171_48 = W*in
   wire signed [14:0] m171_48;
   assign m171_48 =15'b0;

   // m171_49 = W*in
   wire signed [14:0] m171_49;
   assign m171_49 =15'b0;

   // m171_50 = W*in
   wire signed [14:0] m171_50;
   assign m171_50 ={ {3{in171[14]}} , in171[14:3] };

   // m171_51 = W*in
   wire signed [14:0] m171_51;
   assign m171_51 =15'b0;

   // m171_52 = W*in
   wire signed [14:0] m171_52;
   assign m171_52 =15'b0;

   // m171_53 = W*in
   wire signed [14:0] m171_53;
   assign m171_53 =15'b0;

   // m171_54 = W*in
   wire signed [14:0] m171_54;
   assign m171_54 =15'b0;

   // m171_55 = W*in
   wire signed [14:0] m171_55;
   assign m171_55 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_56 = W*in
   wire signed [14:0] m171_56;
   assign m171_56 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_57 = W*in
   wire signed [14:0] m171_57;
   assign m171_57 =15'b0;

   // m171_58 = W*in
   wire signed [14:0] m171_58;
   assign m171_58 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_59 = W*in
   wire signed [14:0] m171_59;
   assign m171_59 =15'b0;

   // m171_60 = W*in
   wire signed [14:0] m171_60;
   assign m171_60 =15'b0;

   // m171_61 = W*in
   wire signed [14:0] m171_61;
   assign m171_61 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_62 = W*in
   wire signed [14:0] m171_62;
   assign m171_62 =15'b0;

   // m171_63 = W*in
   wire signed [14:0] m171_63;
   assign m171_63 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_64 = W*in
   wire signed [14:0] m171_64;
   assign m171_64 =15'b0;

   // m171_65 = W*in
   wire signed [14:0] m171_65;
   assign m171_65 ={ {4{neg171[14]}} , neg171[14:4] };

   // m171_66 = W*in
   wire signed [14:0] m171_66;
   assign m171_66 =15'b0;

   // m171_67 = W*in
   wire signed [14:0] m171_67;
   assign m171_67 =15'b0;

   // m171_68 = W*in
   wire signed [14:0] m171_68;
   assign m171_68 =15'b0;

   // m171_69 = W*in
   wire signed [14:0] m171_69;
   assign m171_69 =15'b0;

   // m171_70 = W*in
   wire signed [14:0] m171_70;
   assign m171_70 =15'b0;

   // m171_71 = W*in
   wire signed [14:0] m171_71;
   assign m171_71 =15'b0;

   // m171_72 = W*in
   wire signed [14:0] m171_72;
   assign m171_72 =15'b0;

   // m171_73 = W*in
   wire signed [14:0] m171_73;
   assign m171_73 =15'b0;

   // m171_74 = W*in
   wire signed [14:0] m171_74;
   assign m171_74 =15'b0;

   // m171_75 = W*in
   wire signed [14:0] m171_75;
   assign m171_75 =15'b0;

   // m171_76 = W*in
   wire signed [14:0] m171_76;
   assign m171_76 ={ {4{neg171[14]}} , neg171[14:4] };

   // m171_77 = W*in
   wire signed [14:0] m171_77;
   assign m171_77 =15'b0;

   // m171_78 = W*in
   wire signed [14:0] m171_78;
   assign m171_78 =15'b0;

   // m171_79 = W*in
   wire signed [14:0] m171_79;
   assign m171_79 =15'b0;

   // m171_80 = W*in
   wire signed [14:0] m171_80;
   assign m171_80 ={ {2{in171[14]}} , in171[14:2] };

   // m171_81 = W*in
   wire signed [14:0] m171_81;
   assign m171_81 =15'b0;

   // m171_82 = W*in
   wire signed [14:0] m171_82;
   assign m171_82 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_83 = W*in
   wire signed [14:0] m171_83;
   assign m171_83 =15'b0;

   // m171_84 = W*in
   wire signed [14:0] m171_84;
   assign m171_84 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_85 = W*in
   wire signed [14:0] m171_85;
   assign m171_85 =15'b0;

   // m171_86 = W*in
   wire signed [14:0] m171_86;
   assign m171_86 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_87 = W*in
   wire signed [14:0] m171_87;
   assign m171_87 =15'b0;

   // m171_88 = W*in
   wire signed [14:0] m171_88;
   assign m171_88 =15'b0;

   // m171_89 = W*in
   wire signed [14:0] m171_89;
   assign m171_89 =15'b0;

   // m171_90 = W*in
   wire signed [14:0] m171_90;
   assign m171_90 =15'b0;

   // m171_91 = W*in
   wire signed [14:0] m171_91;
   assign m171_91 ={ {3{in171[14]}} , in171[14:3] };

   // m171_92 = W*in
   wire signed [14:0] m171_92;
   assign m171_92 =15'b0;

   // m171_93 = W*in
   wire signed [14:0] m171_93;
   assign m171_93 =15'b0;

   // m171_94 = W*in
   wire signed [14:0] m171_94;
   assign m171_94 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_95 = W*in
   wire signed [14:0] m171_95;
   assign m171_95 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_96 = W*in
   wire signed [14:0] m171_96;
   assign m171_96 ={ {3{in171[14]}} , in171[14:3] };

   // m171_97 = W*in
   wire signed [14:0] m171_97;
   assign m171_97 ={ {3{neg171[14]}} , neg171[14:3] };

   // m171_98 = W*in
   wire signed [14:0] m171_98;
   assign m171_98 =15'b0;

   // m171_99 = W*in
   wire signed [14:0] m171_99;
   assign m171_99 =15'b0;

   // m171_100 = W*in
   wire signed [14:0] m171_100;
   assign m171_100 =15'b0;

   // m172_1 = W*in
   wire signed [14:0] m172_1;
   assign m172_1 =15'b0;

   // m172_2 = W*in
   wire signed [14:0] m172_2;
   assign m172_2 =15'b0;

   // m172_3 = W*in
   wire signed [14:0] m172_3;
   assign m172_3 =15'b0;

   // m172_4 = W*in
   wire signed [14:0] m172_4;
   assign m172_4 =15'b0;

   // m172_5 = W*in
   wire signed [14:0] m172_5;
   assign m172_5 ={ {3{in172[14]}} , in172[14:3] };

   // m172_6 = W*in
   wire signed [14:0] m172_6;
   assign m172_6 =15'b0;

   // m172_7 = W*in
   wire signed [14:0] m172_7;
   assign m172_7 =15'b0;

   // m172_8 = W*in
   wire signed [14:0] m172_8;
   assign m172_8 =15'b0;

   // m172_9 = W*in
   wire signed [14:0] m172_9;
   assign m172_9 =15'b0;

   // m172_10 = W*in
   wire signed [14:0] m172_10;
   assign m172_10 =15'b0;

   // m172_11 = W*in
   wire signed [14:0] m172_11;
   assign m172_11 =15'b0;

   // m172_12 = W*in
   wire signed [14:0] m172_12;
   assign m172_12 =15'b0;

   // m172_13 = W*in
   wire signed [14:0] m172_13;
   assign m172_13 =15'b0;

   // m172_14 = W*in
   wire signed [14:0] m172_14;
   assign m172_14 =15'b0;

   // m172_15 = W*in
   wire signed [14:0] m172_15;
   assign m172_15 =15'b0;

   // m172_16 = W*in
   wire signed [14:0] m172_16;
   assign m172_16 =15'b0;

   // m172_17 = W*in
   wire signed [14:0] m172_17;
   assign m172_17 =15'b0;

   // m172_18 = W*in
   wire signed [14:0] m172_18;
   assign m172_18 ={ {4{in172[14]}} , in172[14:4] };

   // m172_19 = W*in
   wire signed [14:0] m172_19;
   assign m172_19 =15'b0;

   // m172_20 = W*in
   wire signed [14:0] m172_20;
   assign m172_20 =15'b0;

   // m172_21 = W*in
   wire signed [14:0] m172_21;
   assign m172_21 =15'b0;

   // m172_22 = W*in
   wire signed [14:0] m172_22;
   assign m172_22 =15'b0;

   // m172_23 = W*in
   wire signed [14:0] m172_23;
   assign m172_23 =15'b0;

   // m172_24 = W*in
   wire signed [14:0] m172_24;
   assign m172_24 =15'b0;

   // m172_25 = W*in
   wire signed [14:0] m172_25;
   assign m172_25 ={ {4{neg172[14]}} , neg172[14:4] };

   // m172_26 = W*in
   wire signed [14:0] m172_26;
   assign m172_26 ={ {4{in172[14]}} , in172[14:4] };

   // m172_27 = W*in
   wire signed [14:0] m172_27;
   assign m172_27 =15'b0;

   // m172_28 = W*in
   wire signed [14:0] m172_28;
   assign m172_28 =15'b0;

   // m172_29 = W*in
   wire signed [14:0] m172_29;
   assign m172_29 =15'b0;

   // m172_30 = W*in
   wire signed [14:0] m172_30;
   assign m172_30 =15'b0;

   // m172_31 = W*in
   wire signed [14:0] m172_31;
   assign m172_31 =15'b0;

   // m172_32 = W*in
   wire signed [14:0] m172_32;
   assign m172_32 =15'b0;

   // m172_33 = W*in
   wire signed [14:0] m172_33;
   assign m172_33 =15'b0;

   // m172_34 = W*in
   wire signed [14:0] m172_34;
   assign m172_34 =15'b0;

   // m172_35 = W*in
   wire signed [14:0] m172_35;
   assign m172_35 =15'b0;

   // m172_36 = W*in
   wire signed [14:0] m172_36;
   assign m172_36 =15'b0;

   // m172_37 = W*in
   wire signed [14:0] m172_37;
   assign m172_37 =15'b0;

   // m172_38 = W*in
   wire signed [14:0] m172_38;
   assign m172_38 =15'b0;

   // m172_39 = W*in
   wire signed [14:0] m172_39;
   assign m172_39 ={ {3{neg172[14]}} , neg172[14:3] };

   // m172_40 = W*in
   wire signed [14:0] m172_40;
   assign m172_40 =15'b0;

   // m172_41 = W*in
   wire signed [14:0] m172_41;
   assign m172_41 =15'b0;

   // m172_42 = W*in
   wire signed [14:0] m172_42;
   assign m172_42 =15'b0;

   // m172_43 = W*in
   wire signed [14:0] m172_43;
   assign m172_43 =15'b0;

   // m172_44 = W*in
   wire signed [14:0] m172_44;
   assign m172_44 =15'b0;

   // m172_45 = W*in
   wire signed [14:0] m172_45;
   assign m172_45 =15'b0;

   // m172_46 = W*in
   wire signed [14:0] m172_46;
   assign m172_46 =15'b0;

   // m172_47 = W*in
   wire signed [14:0] m172_47;
   assign m172_47 ={ {4{in172[14]}} , in172[14:4] };

   // m172_48 = W*in
   wire signed [14:0] m172_48;
   assign m172_48 =15'b0;

   // m172_49 = W*in
   wire signed [14:0] m172_49;
   assign m172_49 =15'b0;

   // m172_50 = W*in
   wire signed [14:0] m172_50;
   assign m172_50 =15'b0;

   // m172_51 = W*in
   wire signed [14:0] m172_51;
   assign m172_51 =15'b0;

   // m172_52 = W*in
   wire signed [14:0] m172_52;
   assign m172_52 =15'b0;

   // m172_53 = W*in
   wire signed [14:0] m172_53;
   assign m172_53 ={ {4{in172[14]}} , in172[14:4] };

   // m172_54 = W*in
   wire signed [14:0] m172_54;
   assign m172_54 =15'b0;

   // m172_55 = W*in
   wire signed [14:0] m172_55;
   assign m172_55 =15'b0;

   // m172_56 = W*in
   wire signed [14:0] m172_56;
   assign m172_56 =15'b0;

   // m172_57 = W*in
   wire signed [14:0] m172_57;
   assign m172_57 =15'b0;

   // m172_58 = W*in
   wire signed [14:0] m172_58;
   assign m172_58 =15'b0;

   // m172_59 = W*in
   wire signed [14:0] m172_59;
   assign m172_59 =15'b0;

   // m172_60 = W*in
   wire signed [14:0] m172_60;
   assign m172_60 =15'b0;

   // m172_61 = W*in
   wire signed [14:0] m172_61;
   assign m172_61 =15'b0;

   // m172_62 = W*in
   wire signed [14:0] m172_62;
   assign m172_62 =15'b0;

   // m172_63 = W*in
   wire signed [14:0] m172_63;
   assign m172_63 =15'b0;

   // m172_64 = W*in
   wire signed [14:0] m172_64;
   assign m172_64 =15'b0;

   // m172_65 = W*in
   wire signed [14:0] m172_65;
   assign m172_65 =15'b0;

   // m172_66 = W*in
   wire signed [14:0] m172_66;
   assign m172_66 ={ {3{neg172[14]}} , neg172[14:3] };

   // m172_67 = W*in
   wire signed [14:0] m172_67;
   assign m172_67 =15'b0;

   // m172_68 = W*in
   wire signed [14:0] m172_68;
   assign m172_68 =15'b0;

   // m172_69 = W*in
   wire signed [14:0] m172_69;
   assign m172_69 =15'b0;

   // m172_70 = W*in
   wire signed [14:0] m172_70;
   assign m172_70 =15'b0;

   // m172_71 = W*in
   wire signed [14:0] m172_71;
   assign m172_71 =15'b0;

   // m172_72 = W*in
   wire signed [14:0] m172_72;
   assign m172_72 ={ {3{neg172[14]}} , neg172[14:3] };

   // m172_73 = W*in
   wire signed [14:0] m172_73;
   assign m172_73 =15'b0;

   // m172_74 = W*in
   wire signed [14:0] m172_74;
   assign m172_74 =15'b0;

   // m172_75 = W*in
   wire signed [14:0] m172_75;
   assign m172_75 =15'b0;

   // m172_76 = W*in
   wire signed [14:0] m172_76;
   assign m172_76 =15'b0;

   // m172_77 = W*in
   wire signed [14:0] m172_77;
   assign m172_77 =15'b0;

   // m172_78 = W*in
   wire signed [14:0] m172_78;
   assign m172_78 =15'b0;

   // m172_79 = W*in
   wire signed [14:0] m172_79;
   assign m172_79 =15'b0;

   // m172_80 = W*in
   wire signed [14:0] m172_80;
   assign m172_80 =15'b0;

   // m172_81 = W*in
   wire signed [14:0] m172_81;
   assign m172_81 =15'b0;

   // m172_82 = W*in
   wire signed [14:0] m172_82;
   assign m172_82 =15'b0;

   // m172_83 = W*in
   wire signed [14:0] m172_83;
   assign m172_83 =15'b0;

   // m172_84 = W*in
   wire signed [14:0] m172_84;
   assign m172_84 =15'b0;

   // m172_85 = W*in
   wire signed [14:0] m172_85;
   assign m172_85 =15'b0;

   // m172_86 = W*in
   wire signed [14:0] m172_86;
   assign m172_86 =15'b0;

   // m172_87 = W*in
   wire signed [14:0] m172_87;
   assign m172_87 =15'b0;

   // m172_88 = W*in
   wire signed [14:0] m172_88;
   assign m172_88 =15'b0;

   // m172_89 = W*in
   wire signed [14:0] m172_89;
   assign m172_89 ={ {4{in172[14]}} , in172[14:4] };

   // m172_90 = W*in
   wire signed [14:0] m172_90;
   assign m172_90 =15'b0;

   // m172_91 = W*in
   wire signed [14:0] m172_91;
   assign m172_91 =15'b0;

   // m172_92 = W*in
   wire signed [14:0] m172_92;
   assign m172_92 =15'b0;

   // m172_93 = W*in
   wire signed [14:0] m172_93;
   assign m172_93 =15'b0;

   // m172_94 = W*in
   wire signed [14:0] m172_94;
   assign m172_94 =15'b0;

   // m172_95 = W*in
   wire signed [14:0] m172_95;
   assign m172_95 =15'b0;

   // m172_96 = W*in
   wire signed [14:0] m172_96;
   assign m172_96 ={ {4{in172[14]}} , in172[14:4] };

   // m172_97 = W*in
   wire signed [14:0] m172_97;
   assign m172_97 =15'b0;

   // m172_98 = W*in
   wire signed [14:0] m172_98;
   assign m172_98 =15'b0;

   // m172_99 = W*in
   wire signed [14:0] m172_99;
   assign m172_99 =15'b0;

   // m172_100 = W*in
   wire signed [14:0] m172_100;
   assign m172_100 =15'b0;

   // m173_1 = W*in
   wire signed [14:0] m173_1;
   assign m173_1 =15'b0;

   // m173_2 = W*in
   wire signed [14:0] m173_2;
   assign m173_2 =15'b0;

   // m173_3 = W*in
   wire signed [14:0] m173_3;
   assign m173_3 =15'b0;

   // m173_4 = W*in
   wire signed [14:0] m173_4;
   assign m173_4 =15'b0;

   // m173_5 = W*in
   wire signed [14:0] m173_5;
   assign m173_5 =15'b0;

   // m173_6 = W*in
   wire signed [14:0] m173_6;
   assign m173_6 =15'b0;

   // m173_7 = W*in
   wire signed [14:0] m173_7;
   assign m173_7 =15'b0;

   // m173_8 = W*in
   wire signed [14:0] m173_8;
   assign m173_8 =15'b0;

   // m173_9 = W*in
   wire signed [14:0] m173_9;
   assign m173_9 =15'b0;

   // m173_10 = W*in
   wire signed [14:0] m173_10;
   assign m173_10 =15'b0;

   // m173_11 = W*in
   wire signed [14:0] m173_11;
   assign m173_11 =15'b0;

   // m173_12 = W*in
   wire signed [14:0] m173_12;
   assign m173_12 =15'b0;

   // m173_13 = W*in
   wire signed [14:0] m173_13;
   assign m173_13 =15'b0;

   // m173_14 = W*in
   wire signed [14:0] m173_14;
   assign m173_14 =15'b0;

   // m173_15 = W*in
   wire signed [14:0] m173_15;
   assign m173_15 =15'b0;

   // m173_16 = W*in
   wire signed [14:0] m173_16;
   assign m173_16 =15'b0;

   // m173_17 = W*in
   wire signed [14:0] m173_17;
   assign m173_17 =15'b0;

   // m173_18 = W*in
   wire signed [14:0] m173_18;
   assign m173_18 =15'b0;

   // m173_19 = W*in
   wire signed [14:0] m173_19;
   assign m173_19 =15'b0;

   // m173_20 = W*in
   wire signed [14:0] m173_20;
   assign m173_20 =15'b0;

   // m173_21 = W*in
   wire signed [14:0] m173_21;
   assign m173_21 =15'b0;

   // m173_22 = W*in
   wire signed [14:0] m173_22;
   assign m173_22 =15'b0;

   // m173_23 = W*in
   wire signed [14:0] m173_23;
   assign m173_23 =15'b0;

   // m173_24 = W*in
   wire signed [14:0] m173_24;
   assign m173_24 =15'b0;

   // m173_25 = W*in
   wire signed [14:0] m173_25;
   assign m173_25 =15'b0;

   // m173_26 = W*in
   wire signed [14:0] m173_26;
   assign m173_26 =15'b0;

   // m173_27 = W*in
   wire signed [14:0] m173_27;
   assign m173_27 =15'b0;

   // m173_28 = W*in
   wire signed [14:0] m173_28;
   assign m173_28 =15'b0;

   // m173_29 = W*in
   wire signed [14:0] m173_29;
   assign m173_29 =15'b0;

   // m173_30 = W*in
   wire signed [14:0] m173_30;
   assign m173_30 =15'b0;

   // m173_31 = W*in
   wire signed [14:0] m173_31;
   assign m173_31 =15'b0;

   // m173_32 = W*in
   wire signed [14:0] m173_32;
   assign m173_32 =15'b0;

   // m173_33 = W*in
   wire signed [14:0] m173_33;
   assign m173_33 =15'b0;

   // m173_34 = W*in
   wire signed [14:0] m173_34;
   assign m173_34 ={ {4{neg173[14]}} , neg173[14:4] };

   // m173_35 = W*in
   wire signed [14:0] m173_35;
   assign m173_35 =15'b0;

   // m173_36 = W*in
   wire signed [14:0] m173_36;
   assign m173_36 =15'b0;

   // m173_37 = W*in
   wire signed [14:0] m173_37;
   assign m173_37 ={ {4{neg173[14]}} , neg173[14:4] };

   // m173_38 = W*in
   wire signed [14:0] m173_38;
   assign m173_38 =15'b0;

   // m173_39 = W*in
   wire signed [14:0] m173_39;
   assign m173_39 =15'b0;

   // m173_40 = W*in
   wire signed [14:0] m173_40;
   assign m173_40 ={ {2{in173[14]}} , in173[14:2] };

   // m173_41 = W*in
   wire signed [14:0] m173_41;
   assign m173_41 =15'b0;

   // m173_42 = W*in
   wire signed [14:0] m173_42;
   assign m173_42 =15'b0;

   // m173_43 = W*in
   wire signed [14:0] m173_43;
   assign m173_43 =15'b0;

   // m173_44 = W*in
   wire signed [14:0] m173_44;
   assign m173_44 =15'b0;

   // m173_45 = W*in
   wire signed [14:0] m173_45;
   assign m173_45 =15'b0;

   // m173_46 = W*in
   wire signed [14:0] m173_46;
   assign m173_46 =15'b0;

   // m173_47 = W*in
   wire signed [14:0] m173_47;
   assign m173_47 =15'b0;

   // m173_48 = W*in
   wire signed [14:0] m173_48;
   assign m173_48 =15'b0;

   // m173_49 = W*in
   wire signed [14:0] m173_49;
   assign m173_49 =15'b0;

   // m173_50 = W*in
   wire signed [14:0] m173_50;
   assign m173_50 =15'b0;

   // m173_51 = W*in
   wire signed [14:0] m173_51;
   assign m173_51 =15'b0;

   // m173_52 = W*in
   wire signed [14:0] m173_52;
   assign m173_52 =15'b0;

   // m173_53 = W*in
   wire signed [14:0] m173_53;
   assign m173_53 ={ {4{in173[14]}} , in173[14:4] };

   // m173_54 = W*in
   wire signed [14:0] m173_54;
   assign m173_54 ={ {3{in173[14]}} , in173[14:3] };

   // m173_55 = W*in
   wire signed [14:0] m173_55;
   assign m173_55 =15'b0;

   // m173_56 = W*in
   wire signed [14:0] m173_56;
   assign m173_56 =15'b0;

   // m173_57 = W*in
   wire signed [14:0] m173_57;
   assign m173_57 ={ {3{in173[14]}} , in173[14:3] };

   // m173_58 = W*in
   wire signed [14:0] m173_58;
   assign m173_58 =15'b0;

   // m173_59 = W*in
   wire signed [14:0] m173_59;
   assign m173_59 ={ {4{in173[14]}} , in173[14:4] };

   // m173_60 = W*in
   wire signed [14:0] m173_60;
   assign m173_60 =15'b0;

   // m173_61 = W*in
   wire signed [14:0] m173_61;
   assign m173_61 =15'b0;

   // m173_62 = W*in
   wire signed [14:0] m173_62;
   assign m173_62 =15'b0;

   // m173_63 = W*in
   wire signed [14:0] m173_63;
   assign m173_63 =15'b0;

   // m173_64 = W*in
   wire signed [14:0] m173_64;
   assign m173_64 =15'b0;

   // m173_65 = W*in
   wire signed [14:0] m173_65;
   assign m173_65 =15'b0;

   // m173_66 = W*in
   wire signed [14:0] m173_66;
   assign m173_66 =15'b0;

   // m173_67 = W*in
   wire signed [14:0] m173_67;
   assign m173_67 =15'b0;

   // m173_68 = W*in
   wire signed [14:0] m173_68;
   assign m173_68 =15'b0;

   // m173_69 = W*in
   wire signed [14:0] m173_69;
   assign m173_69 ={ {4{neg173[14]}} , neg173[14:4] };

   // m173_70 = W*in
   wire signed [14:0] m173_70;
   assign m173_70 =15'b0;

   // m173_71 = W*in
   wire signed [14:0] m173_71;
   assign m173_71 =15'b0;

   // m173_72 = W*in
   wire signed [14:0] m173_72;
   assign m173_72 =15'b0;

   // m173_73 = W*in
   wire signed [14:0] m173_73;
   assign m173_73 =15'b0;

   // m173_74 = W*in
   wire signed [14:0] m173_74;
   assign m173_74 ={ {4{in173[14]}} , in173[14:4] };

   // m173_75 = W*in
   wire signed [14:0] m173_75;
   assign m173_75 =15'b0;

   // m173_76 = W*in
   wire signed [14:0] m173_76;
   assign m173_76 =15'b0;

   // m173_77 = W*in
   wire signed [14:0] m173_77;
   assign m173_77 =15'b0;

   // m173_78 = W*in
   wire signed [14:0] m173_78;
   assign m173_78 =15'b0;

   // m173_79 = W*in
   wire signed [14:0] m173_79;
   assign m173_79 =15'b0;

   // m173_80 = W*in
   wire signed [14:0] m173_80;
   assign m173_80 ={ {4{in173[14]}} , in173[14:4] };

   // m173_81 = W*in
   wire signed [14:0] m173_81;
   assign m173_81 =15'b0;

   // m173_82 = W*in
   wire signed [14:0] m173_82;
   assign m173_82 =15'b0;

   // m173_83 = W*in
   wire signed [14:0] m173_83;
   assign m173_83 =15'b0;

   // m173_84 = W*in
   wire signed [14:0] m173_84;
   assign m173_84 ={ {3{neg173[14]}} , neg173[14:3] };

   // m173_85 = W*in
   wire signed [14:0] m173_85;
   assign m173_85 =15'b0;

   // m173_86 = W*in
   wire signed [14:0] m173_86;
   assign m173_86 =15'b0;

   // m173_87 = W*in
   wire signed [14:0] m173_87;
   assign m173_87 =15'b0;

   // m173_88 = W*in
   wire signed [14:0] m173_88;
   assign m173_88 =15'b0;

   // m173_89 = W*in
   wire signed [14:0] m173_89;
   assign m173_89 =15'b0;

   // m173_90 = W*in
   wire signed [14:0] m173_90;
   assign m173_90 =15'b0;

   // m173_91 = W*in
   wire signed [14:0] m173_91;
   assign m173_91 =15'b0;

   // m173_92 = W*in
   wire signed [14:0] m173_92;
   assign m173_92 =15'b0;

   // m173_93 = W*in
   wire signed [14:0] m173_93;
   assign m173_93 =15'b0;

   // m173_94 = W*in
   wire signed [14:0] m173_94;
   assign m173_94 =15'b0;

   // m173_95 = W*in
   wire signed [14:0] m173_95;
   assign m173_95 =15'b0;

   // m173_96 = W*in
   wire signed [14:0] m173_96;
   assign m173_96 =15'b0;

   // m173_97 = W*in
   wire signed [14:0] m173_97;
   assign m173_97 =15'b0;

   // m173_98 = W*in
   wire signed [14:0] m173_98;
   assign m173_98 =15'b0;

   // m173_99 = W*in
   wire signed [14:0] m173_99;
   assign m173_99 ={ {4{in173[14]}} , in173[14:4] };

   // m173_100 = W*in
   wire signed [14:0] m173_100;
   assign m173_100 ={ {3{in173[14]}} , in173[14:3] };

   // m174_1 = W*in
   wire signed [14:0] m174_1;
   assign m174_1 =15'b0;

   // m174_2 = W*in
   wire signed [14:0] m174_2;
   assign m174_2 =15'b0;

   // m174_3 = W*in
   wire signed [14:0] m174_3;
   assign m174_3 =15'b0;

   // m174_4 = W*in
   wire signed [14:0] m174_4;
   assign m174_4 =15'b0;

   // m174_5 = W*in
   wire signed [14:0] m174_5;
   assign m174_5 =15'b0;

   // m174_6 = W*in
   wire signed [14:0] m174_6;
   assign m174_6 =15'b0;

   // m174_7 = W*in
   wire signed [14:0] m174_7;
   assign m174_7 ={ {3{in174[14]}} , in174[14:3] };

   // m174_8 = W*in
   wire signed [14:0] m174_8;
   assign m174_8 ={ {3{in174[14]}} , in174[14:3] };

   // m174_9 = W*in
   wire signed [14:0] m174_9;
   assign m174_9 =15'b0;

   // m174_10 = W*in
   wire signed [14:0] m174_10;
   assign m174_10 =15'b0;

   // m174_11 = W*in
   wire signed [14:0] m174_11;
   assign m174_11 =15'b0;

   // m174_12 = W*in
   wire signed [14:0] m174_12;
   assign m174_12 =15'b0;

   // m174_13 = W*in
   wire signed [14:0] m174_13;
   assign m174_13 =15'b0;

   // m174_14 = W*in
   wire signed [14:0] m174_14;
   assign m174_14 =15'b0;

   // m174_15 = W*in
   wire signed [14:0] m174_15;
   assign m174_15 =15'b0;

   // m174_16 = W*in
   wire signed [14:0] m174_16;
   assign m174_16 =15'b0;

   // m174_17 = W*in
   wire signed [14:0] m174_17;
   assign m174_17 =15'b0;

   // m174_18 = W*in
   wire signed [14:0] m174_18;
   assign m174_18 ={ {4{in174[14]}} , in174[14:4] };

   // m174_19 = W*in
   wire signed [14:0] m174_19;
   assign m174_19 =15'b0;

   // m174_20 = W*in
   wire signed [14:0] m174_20;
   assign m174_20 =15'b0;

   // m174_21 = W*in
   wire signed [14:0] m174_21;
   assign m174_21 ={ {3{in174[14]}} , in174[14:3] };

   // m174_22 = W*in
   wire signed [14:0] m174_22;
   assign m174_22 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_23 = W*in
   wire signed [14:0] m174_23;
   assign m174_23 =15'b0;

   // m174_24 = W*in
   wire signed [14:0] m174_24;
   assign m174_24 =15'b0;

   // m174_25 = W*in
   wire signed [14:0] m174_25;
   assign m174_25 =15'b0;

   // m174_26 = W*in
   wire signed [14:0] m174_26;
   assign m174_26 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_27 = W*in
   wire signed [14:0] m174_27;
   assign m174_27 =15'b0;

   // m174_28 = W*in
   wire signed [14:0] m174_28;
   assign m174_28 =15'b0;

   // m174_29 = W*in
   wire signed [14:0] m174_29;
   assign m174_29 =15'b0;

   // m174_30 = W*in
   wire signed [14:0] m174_30;
   assign m174_30 =15'b0;

   // m174_31 = W*in
   wire signed [14:0] m174_31;
   assign m174_31 =15'b0;

   // m174_32 = W*in
   wire signed [14:0] m174_32;
   assign m174_32 ={ {3{in174[14]}} , in174[14:3] };

   // m174_33 = W*in
   wire signed [14:0] m174_33;
   assign m174_33 ={ {3{in174[14]}} , in174[14:3] };

   // m174_34 = W*in
   wire signed [14:0] m174_34;
   assign m174_34 =15'b0;

   // m174_35 = W*in
   wire signed [14:0] m174_35;
   assign m174_35 ={ {3{in174[14]}} , in174[14:3] };

   // m174_36 = W*in
   wire signed [14:0] m174_36;
   assign m174_36 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_37 = W*in
   wire signed [14:0] m174_37;
   assign m174_37 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_38 = W*in
   wire signed [14:0] m174_38;
   assign m174_38 =15'b0;

   // m174_39 = W*in
   wire signed [14:0] m174_39;
   assign m174_39 =15'b0;

   // m174_40 = W*in
   wire signed [14:0] m174_40;
   assign m174_40 =15'b0;

   // m174_41 = W*in
   wire signed [14:0] m174_41;
   assign m174_41 =15'b0;

   // m174_42 = W*in
   wire signed [14:0] m174_42;
   assign m174_42 =15'b0;

   // m174_43 = W*in
   wire signed [14:0] m174_43;
   assign m174_43 =15'b0;

   // m174_44 = W*in
   wire signed [14:0] m174_44;
   assign m174_44 ={ {2{in174[14]}} , in174[14:2] };

   // m174_45 = W*in
   wire signed [14:0] m174_45;
   assign m174_45 =15'b0;

   // m174_46 = W*in
   wire signed [14:0] m174_46;
   assign m174_46 ={ {4{neg174[14]}} , neg174[14:4] };

   // m174_47 = W*in
   wire signed [14:0] m174_47;
   assign m174_47 =15'b0;

   // m174_48 = W*in
   wire signed [14:0] m174_48;
   assign m174_48 ={ {4{in174[14]}} , in174[14:4] };

   // m174_49 = W*in
   wire signed [14:0] m174_49;
   assign m174_49 =15'b0;

   // m174_50 = W*in
   wire signed [14:0] m174_50;
   assign m174_50 =15'b0;

   // m174_51 = W*in
   wire signed [14:0] m174_51;
   assign m174_51 =15'b0;

   // m174_52 = W*in
   wire signed [14:0] m174_52;
   assign m174_52 =15'b0;

   // m174_53 = W*in
   wire signed [14:0] m174_53;
   assign m174_53 =15'b0;

   // m174_54 = W*in
   wire signed [14:0] m174_54;
   assign m174_54 =15'b0;

   // m174_55 = W*in
   wire signed [14:0] m174_55;
   assign m174_55 =15'b0;

   // m174_56 = W*in
   wire signed [14:0] m174_56;
   assign m174_56 =15'b0;

   // m174_57 = W*in
   wire signed [14:0] m174_57;
   assign m174_57 ={ {4{neg174[14]}} , neg174[14:4] };

   // m174_58 = W*in
   wire signed [14:0] m174_58;
   assign m174_58 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_59 = W*in
   wire signed [14:0] m174_59;
   assign m174_59 =15'b0;

   // m174_60 = W*in
   wire signed [14:0] m174_60;
   assign m174_60 =15'b0;

   // m174_61 = W*in
   wire signed [14:0] m174_61;
   assign m174_61 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_62 = W*in
   wire signed [14:0] m174_62;
   assign m174_62 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_63 = W*in
   wire signed [14:0] m174_63;
   assign m174_63 =15'b0;

   // m174_64 = W*in
   wire signed [14:0] m174_64;
   assign m174_64 ={ {4{neg174[14]}} , neg174[14:4] };

   // m174_65 = W*in
   wire signed [14:0] m174_65;
   assign m174_65 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_66 = W*in
   wire signed [14:0] m174_66;
   assign m174_66 =15'b0;

   // m174_67 = W*in
   wire signed [14:0] m174_67;
   assign m174_67 =15'b0;

   // m174_68 = W*in
   wire signed [14:0] m174_68;
   assign m174_68 ={ {4{neg174[14]}} , neg174[14:4] };

   // m174_69 = W*in
   wire signed [14:0] m174_69;
   assign m174_69 =15'b0;

   // m174_70 = W*in
   wire signed [14:0] m174_70;
   assign m174_70 ={ {3{in174[14]}} , in174[14:3] };

   // m174_71 = W*in
   wire signed [14:0] m174_71;
   assign m174_71 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_72 = W*in
   wire signed [14:0] m174_72;
   assign m174_72 =15'b0;

   // m174_73 = W*in
   wire signed [14:0] m174_73;
   assign m174_73 =15'b0;

   // m174_74 = W*in
   wire signed [14:0] m174_74;
   assign m174_74 ={ {4{in174[14]}} , in174[14:4] };

   // m174_75 = W*in
   wire signed [14:0] m174_75;
   assign m174_75 =15'b0;

   // m174_76 = W*in
   wire signed [14:0] m174_76;
   assign m174_76 =15'b0;

   // m174_77 = W*in
   wire signed [14:0] m174_77;
   assign m174_77 =15'b0;

   // m174_78 = W*in
   wire signed [14:0] m174_78;
   assign m174_78 =15'b0;

   // m174_79 = W*in
   wire signed [14:0] m174_79;
   assign m174_79 =15'b0;

   // m174_80 = W*in
   wire signed [14:0] m174_80;
   assign m174_80 =15'b0;

   // m174_81 = W*in
   wire signed [14:0] m174_81;
   assign m174_81 =15'b0;

   // m174_82 = W*in
   wire signed [14:0] m174_82;
   assign m174_82 =15'b0;

   // m174_83 = W*in
   wire signed [14:0] m174_83;
   assign m174_83 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_84 = W*in
   wire signed [14:0] m174_84;
   assign m174_84 =15'b0;

   // m174_85 = W*in
   wire signed [14:0] m174_85;
   assign m174_85 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_86 = W*in
   wire signed [14:0] m174_86;
   assign m174_86 =15'b0;

   // m174_87 = W*in
   wire signed [14:0] m174_87;
   assign m174_87 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_88 = W*in
   wire signed [14:0] m174_88;
   assign m174_88 =15'b0;

   // m174_89 = W*in
   wire signed [14:0] m174_89;
   assign m174_89 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_90 = W*in
   wire signed [14:0] m174_90;
   assign m174_90 ={ {3{in174[14]}} , in174[14:3] };

   // m174_91 = W*in
   wire signed [14:0] m174_91;
   assign m174_91 =15'b0;

   // m174_92 = W*in
   wire signed [14:0] m174_92;
   assign m174_92 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_93 = W*in
   wire signed [14:0] m174_93;
   assign m174_93 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_94 = W*in
   wire signed [14:0] m174_94;
   assign m174_94 ={ {3{in174[14]}} , in174[14:3] };

   // m174_95 = W*in
   wire signed [14:0] m174_95;
   assign m174_95 ={ {3{in174[14]}} , in174[14:3] };

   // m174_96 = W*in
   wire signed [14:0] m174_96;
   assign m174_96 =15'b0;

   // m174_97 = W*in
   wire signed [14:0] m174_97;
   assign m174_97 ={ {3{neg174[14]}} , neg174[14:3] };

   // m174_98 = W*in
   wire signed [14:0] m174_98;
   assign m174_98 ={ {3{in174[14]}} , in174[14:3] };

   // m174_99 = W*in
   wire signed [14:0] m174_99;
   assign m174_99 =15'b0;

   // m174_100 = W*in
   wire signed [14:0] m174_100;
   assign m174_100 =15'b0;

   // m175_1 = W*in
   wire signed [14:0] m175_1;
   assign m175_1 =15'b0;

   // m175_2 = W*in
   wire signed [14:0] m175_2;
   assign m175_2 =15'b0;

   // m175_3 = W*in
   wire signed [14:0] m175_3;
   assign m175_3 =15'b0;

   // m175_4 = W*in
   wire signed [14:0] m175_4;
   assign m175_4 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_5 = W*in
   wire signed [14:0] m175_5;
   assign m175_5 =15'b0;

   // m175_6 = W*in
   wire signed [14:0] m175_6;
   assign m175_6 =15'b0;

   // m175_7 = W*in
   wire signed [14:0] m175_7;
   assign m175_7 =15'b0;

   // m175_8 = W*in
   wire signed [14:0] m175_8;
   assign m175_8 =15'b0;

   // m175_9 = W*in
   wire signed [14:0] m175_9;
   assign m175_9 =15'b0;

   // m175_10 = W*in
   wire signed [14:0] m175_10;
   assign m175_10 =15'b0;

   // m175_11 = W*in
   wire signed [14:0] m175_11;
   assign m175_11 =15'b0;

   // m175_12 = W*in
   wire signed [14:0] m175_12;
   assign m175_12 =15'b0;

   // m175_13 = W*in
   wire signed [14:0] m175_13;
   assign m175_13 =15'b0;

   // m175_14 = W*in
   wire signed [14:0] m175_14;
   assign m175_14 =15'b0;

   // m175_15 = W*in
   wire signed [14:0] m175_15;
   assign m175_15 =15'b0;

   // m175_16 = W*in
   wire signed [14:0] m175_16;
   assign m175_16 =15'b0;

   // m175_17 = W*in
   wire signed [14:0] m175_17;
   assign m175_17 =15'b0;

   // m175_18 = W*in
   wire signed [14:0] m175_18;
   assign m175_18 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_19 = W*in
   wire signed [14:0] m175_19;
   assign m175_19 ={ {4{in175[14]}} , in175[14:4] };

   // m175_20 = W*in
   wire signed [14:0] m175_20;
   assign m175_20 =15'b0;

   // m175_21 = W*in
   wire signed [14:0] m175_21;
   assign m175_21 =15'b0;

   // m175_22 = W*in
   wire signed [14:0] m175_22;
   assign m175_22 ={ {4{in175[14]}} , in175[14:4] };

   // m175_23 = W*in
   wire signed [14:0] m175_23;
   assign m175_23 =15'b0;

   // m175_24 = W*in
   wire signed [14:0] m175_24;
   assign m175_24 =15'b0;

   // m175_25 = W*in
   wire signed [14:0] m175_25;
   assign m175_25 ={ {4{in175[14]}} , in175[14:4] };

   // m175_26 = W*in
   wire signed [14:0] m175_26;
   assign m175_26 =15'b0;

   // m175_27 = W*in
   wire signed [14:0] m175_27;
   assign m175_27 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_28 = W*in
   wire signed [14:0] m175_28;
   assign m175_28 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_29 = W*in
   wire signed [14:0] m175_29;
   assign m175_29 =15'b0;

   // m175_30 = W*in
   wire signed [14:0] m175_30;
   assign m175_30 =15'b0;

   // m175_31 = W*in
   wire signed [14:0] m175_31;
   assign m175_31 =15'b0;

   // m175_32 = W*in
   wire signed [14:0] m175_32;
   assign m175_32 =15'b0;

   // m175_33 = W*in
   wire signed [14:0] m175_33;
   assign m175_33 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_34 = W*in
   wire signed [14:0] m175_34;
   assign m175_34 =15'b0;

   // m175_35 = W*in
   wire signed [14:0] m175_35;
   assign m175_35 =15'b0;

   // m175_36 = W*in
   wire signed [14:0] m175_36;
   assign m175_36 =15'b0;

   // m175_37 = W*in
   wire signed [14:0] m175_37;
   assign m175_37 =15'b0;

   // m175_38 = W*in
   wire signed [14:0] m175_38;
   assign m175_38 =15'b0;

   // m175_39 = W*in
   wire signed [14:0] m175_39;
   assign m175_39 =15'b0;

   // m175_40 = W*in
   wire signed [14:0] m175_40;
   assign m175_40 =15'b0;

   // m175_41 = W*in
   wire signed [14:0] m175_41;
   assign m175_41 =15'b0;

   // m175_42 = W*in
   wire signed [14:0] m175_42;
   assign m175_42 =15'b0;

   // m175_43 = W*in
   wire signed [14:0] m175_43;
   assign m175_43 =15'b0;

   // m175_44 = W*in
   wire signed [14:0] m175_44;
   assign m175_44 =15'b0;

   // m175_45 = W*in
   wire signed [14:0] m175_45;
   assign m175_45 =15'b0;

   // m175_46 = W*in
   wire signed [14:0] m175_46;
   assign m175_46 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_47 = W*in
   wire signed [14:0] m175_47;
   assign m175_47 =15'b0;

   // m175_48 = W*in
   wire signed [14:0] m175_48;
   assign m175_48 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_49 = W*in
   wire signed [14:0] m175_49;
   assign m175_49 =15'b0;

   // m175_50 = W*in
   wire signed [14:0] m175_50;
   assign m175_50 =15'b0;

   // m175_51 = W*in
   wire signed [14:0] m175_51;
   assign m175_51 =15'b0;

   // m175_52 = W*in
   wire signed [14:0] m175_52;
   assign m175_52 =15'b0;

   // m175_53 = W*in
   wire signed [14:0] m175_53;
   assign m175_53 =15'b0;

   // m175_54 = W*in
   wire signed [14:0] m175_54;
   assign m175_54 =15'b0;

   // m175_55 = W*in
   wire signed [14:0] m175_55;
   assign m175_55 =15'b0;

   // m175_56 = W*in
   wire signed [14:0] m175_56;
   assign m175_56 =15'b0;

   // m175_57 = W*in
   wire signed [14:0] m175_57;
   assign m175_57 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_58 = W*in
   wire signed [14:0] m175_58;
   assign m175_58 =15'b0;

   // m175_59 = W*in
   wire signed [14:0] m175_59;
   assign m175_59 ={ {3{in175[14]}} , in175[14:3] };

   // m175_60 = W*in
   wire signed [14:0] m175_60;
   assign m175_60 =15'b0;

   // m175_61 = W*in
   wire signed [14:0] m175_61;
   assign m175_61 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_62 = W*in
   wire signed [14:0] m175_62;
   assign m175_62 =15'b0;

   // m175_63 = W*in
   wire signed [14:0] m175_63;
   assign m175_63 ={ {3{neg175[14]}} , neg175[14:3] };

   // m175_64 = W*in
   wire signed [14:0] m175_64;
   assign m175_64 ={ {4{in175[14]}} , in175[14:4] };

   // m175_65 = W*in
   wire signed [14:0] m175_65;
   assign m175_65 =15'b0;

   // m175_66 = W*in
   wire signed [14:0] m175_66;
   assign m175_66 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_67 = W*in
   wire signed [14:0] m175_67;
   assign m175_67 =15'b0;

   // m175_68 = W*in
   wire signed [14:0] m175_68;
   assign m175_68 ={ {4{neg175[14]}} , neg175[14:4] };

   // m175_69 = W*in
   wire signed [14:0] m175_69;
   assign m175_69 ={ {4{in175[14]}} , in175[14:4] };

   // m175_70 = W*in
   wire signed [14:0] m175_70;
   assign m175_70 ={ {3{in175[14]}} , in175[14:3] };

   // m175_71 = W*in
   wire signed [14:0] m175_71;
   assign m175_71 =15'b0;

   // m175_72 = W*in
   wire signed [14:0] m175_72;
   assign m175_72 =15'b0;

   // m175_73 = W*in
   wire signed [14:0] m175_73;
   assign m175_73 =15'b0;

   // m175_74 = W*in
   wire signed [14:0] m175_74;
   assign m175_74 =15'b0;

   // m175_75 = W*in
   wire signed [14:0] m175_75;
   assign m175_75 ={ {3{in175[14]}} , in175[14:3] };

   // m175_76 = W*in
   wire signed [14:0] m175_76;
   assign m175_76 =15'b0;

   // m175_77 = W*in
   wire signed [14:0] m175_77;
   assign m175_77 =15'b0;

   // m175_78 = W*in
   wire signed [14:0] m175_78;
   assign m175_78 =15'b0;

   // m175_79 = W*in
   wire signed [14:0] m175_79;
   assign m175_79 =15'b0;

   // m175_80 = W*in
   wire signed [14:0] m175_80;
   assign m175_80 =15'b0;

   // m175_81 = W*in
   wire signed [14:0] m175_81;
   assign m175_81 =15'b0;

   // m175_82 = W*in
   wire signed [14:0] m175_82;
   assign m175_82 =15'b0;

   // m175_83 = W*in
   wire signed [14:0] m175_83;
   assign m175_83 =15'b0;

   // m175_84 = W*in
   wire signed [14:0] m175_84;
   assign m175_84 =15'b0;

   // m175_85 = W*in
   wire signed [14:0] m175_85;
   assign m175_85 =15'b0;

   // m175_86 = W*in
   wire signed [14:0] m175_86;
   assign m175_86 =15'b0;

   // m175_87 = W*in
   wire signed [14:0] m175_87;
   assign m175_87 =15'b0;

   // m175_88 = W*in
   wire signed [14:0] m175_88;
   assign m175_88 ={ {3{in175[14]}} , in175[14:3] };

   // m175_89 = W*in
   wire signed [14:0] m175_89;
   assign m175_89 =15'b0;

   // m175_90 = W*in
   wire signed [14:0] m175_90;
   assign m175_90 =15'b0;

   // m175_91 = W*in
   wire signed [14:0] m175_91;
   assign m175_91 =15'b0;

   // m175_92 = W*in
   wire signed [14:0] m175_92;
   assign m175_92 =15'b0;

   // m175_93 = W*in
   wire signed [14:0] m175_93;
   assign m175_93 =15'b0;

   // m175_94 = W*in
   wire signed [14:0] m175_94;
   assign m175_94 =15'b0;

   // m175_95 = W*in
   wire signed [14:0] m175_95;
   assign m175_95 =15'b0;

   // m175_96 = W*in
   wire signed [14:0] m175_96;
   assign m175_96 =15'b0;

   // m175_97 = W*in
   wire signed [14:0] m175_97;
   assign m175_97 =15'b0;

   // m175_98 = W*in
   wire signed [14:0] m175_98;
   assign m175_98 =15'b0;

   // m175_99 = W*in
   wire signed [14:0] m175_99;
   assign m175_99 =15'b0;

   // m175_100 = W*in
   wire signed [14:0] m175_100;
   assign m175_100 =15'b0;

   // m176_1 = W*in
   wire signed [14:0] m176_1;
   assign m176_1 ={ {3{in176[14]}} , in176[14:3] };

   // m176_2 = W*in
   wire signed [14:0] m176_2;
   assign m176_2 =15'b0;

   // m176_3 = W*in
   wire signed [14:0] m176_3;
   assign m176_3 =15'b0;

   // m176_4 = W*in
   wire signed [14:0] m176_4;
   assign m176_4 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_5 = W*in
   wire signed [14:0] m176_5;
   assign m176_5 =15'b0;

   // m176_6 = W*in
   wire signed [14:0] m176_6;
   assign m176_6 =15'b0;

   // m176_7 = W*in
   wire signed [14:0] m176_7;
   assign m176_7 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_8 = W*in
   wire signed [14:0] m176_8;
   assign m176_8 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_9 = W*in
   wire signed [14:0] m176_9;
   assign m176_9 =15'b0;

   // m176_10 = W*in
   wire signed [14:0] m176_10;
   assign m176_10 =15'b0;

   // m176_11 = W*in
   wire signed [14:0] m176_11;
   assign m176_11 =15'b0;

   // m176_12 = W*in
   wire signed [14:0] m176_12;
   assign m176_12 =15'b0;

   // m176_13 = W*in
   wire signed [14:0] m176_13;
   assign m176_13 =15'b0;

   // m176_14 = W*in
   wire signed [14:0] m176_14;
   assign m176_14 =15'b0;

   // m176_15 = W*in
   wire signed [14:0] m176_15;
   assign m176_15 =15'b0;

   // m176_16 = W*in
   wire signed [14:0] m176_16;
   assign m176_16 =15'b0;

   // m176_17 = W*in
   wire signed [14:0] m176_17;
   assign m176_17 =15'b0;

   // m176_18 = W*in
   wire signed [14:0] m176_18;
   assign m176_18 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_19 = W*in
   wire signed [14:0] m176_19;
   assign m176_19 ={ {4{in176[14]}} , in176[14:4] };

   // m176_20 = W*in
   wire signed [14:0] m176_20;
   assign m176_20 =15'b0;

   // m176_21 = W*in
   wire signed [14:0] m176_21;
   assign m176_21 ={ {3{in176[14]}} , in176[14:3] };

   // m176_22 = W*in
   wire signed [14:0] m176_22;
   assign m176_22 =15'b0;

   // m176_23 = W*in
   wire signed [14:0] m176_23;
   assign m176_23 =15'b0;

   // m176_24 = W*in
   wire signed [14:0] m176_24;
   assign m176_24 =15'b0;

   // m176_25 = W*in
   wire signed [14:0] m176_25;
   assign m176_25 ={ {3{in176[14]}} , in176[14:3] };

   // m176_26 = W*in
   wire signed [14:0] m176_26;
   assign m176_26 =15'b0;

   // m176_27 = W*in
   wire signed [14:0] m176_27;
   assign m176_27 =15'b0;

   // m176_28 = W*in
   wire signed [14:0] m176_28;
   assign m176_28 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_29 = W*in
   wire signed [14:0] m176_29;
   assign m176_29 =15'b0;

   // m176_30 = W*in
   wire signed [14:0] m176_30;
   assign m176_30 =15'b0;

   // m176_31 = W*in
   wire signed [14:0] m176_31;
   assign m176_31 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_32 = W*in
   wire signed [14:0] m176_32;
   assign m176_32 =15'b0;

   // m176_33 = W*in
   wire signed [14:0] m176_33;
   assign m176_33 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_34 = W*in
   wire signed [14:0] m176_34;
   assign m176_34 =15'b0;

   // m176_35 = W*in
   wire signed [14:0] m176_35;
   assign m176_35 =15'b0;

   // m176_36 = W*in
   wire signed [14:0] m176_36;
   assign m176_36 =15'b0;

   // m176_37 = W*in
   wire signed [14:0] m176_37;
   assign m176_37 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_38 = W*in
   wire signed [14:0] m176_38;
   assign m176_38 =15'b0;

   // m176_39 = W*in
   wire signed [14:0] m176_39;
   assign m176_39 =15'b0;

   // m176_40 = W*in
   wire signed [14:0] m176_40;
   assign m176_40 =15'b0;

   // m176_41 = W*in
   wire signed [14:0] m176_41;
   assign m176_41 =15'b0;

   // m176_42 = W*in
   wire signed [14:0] m176_42;
   assign m176_42 =15'b0;

   // m176_43 = W*in
   wire signed [14:0] m176_43;
   assign m176_43 =15'b0;

   // m176_44 = W*in
   wire signed [14:0] m176_44;
   assign m176_44 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_45 = W*in
   wire signed [14:0] m176_45;
   assign m176_45 =15'b0;

   // m176_46 = W*in
   wire signed [14:0] m176_46;
   assign m176_46 =15'b0;

   // m176_47 = W*in
   wire signed [14:0] m176_47;
   assign m176_47 =15'b0;

   // m176_48 = W*in
   wire signed [14:0] m176_48;
   assign m176_48 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_49 = W*in
   wire signed [14:0] m176_49;
   assign m176_49 =15'b0;

   // m176_50 = W*in
   wire signed [14:0] m176_50;
   assign m176_50 =15'b0;

   // m176_51 = W*in
   wire signed [14:0] m176_51;
   assign m176_51 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_52 = W*in
   wire signed [14:0] m176_52;
   assign m176_52 =15'b0;

   // m176_53 = W*in
   wire signed [14:0] m176_53;
   assign m176_53 =15'b0;

   // m176_54 = W*in
   wire signed [14:0] m176_54;
   assign m176_54 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_55 = W*in
   wire signed [14:0] m176_55;
   assign m176_55 =15'b0;

   // m176_56 = W*in
   wire signed [14:0] m176_56;
   assign m176_56 =15'b0;

   // m176_57 = W*in
   wire signed [14:0] m176_57;
   assign m176_57 =15'b0;

   // m176_58 = W*in
   wire signed [14:0] m176_58;
   assign m176_58 =15'b0;

   // m176_59 = W*in
   wire signed [14:0] m176_59;
   assign m176_59 ={ {4{in176[14]}} , in176[14:4] };

   // m176_60 = W*in
   wire signed [14:0] m176_60;
   assign m176_60 =15'b0;

   // m176_61 = W*in
   wire signed [14:0] m176_61;
   assign m176_61 ={ {4{in176[14]}} , in176[14:4] };

   // m176_62 = W*in
   wire signed [14:0] m176_62;
   assign m176_62 =15'b0;

   // m176_63 = W*in
   wire signed [14:0] m176_63;
   assign m176_63 =15'b0;

   // m176_64 = W*in
   wire signed [14:0] m176_64;
   assign m176_64 ={ {4{in176[14]}} , in176[14:4] };

   // m176_65 = W*in
   wire signed [14:0] m176_65;
   assign m176_65 ={ {4{in176[14]}} , in176[14:4] };

   // m176_66 = W*in
   wire signed [14:0] m176_66;
   assign m176_66 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_67 = W*in
   wire signed [14:0] m176_67;
   assign m176_67 =15'b0;

   // m176_68 = W*in
   wire signed [14:0] m176_68;
   assign m176_68 =15'b0;

   // m176_69 = W*in
   wire signed [14:0] m176_69;
   assign m176_69 ={ {3{in176[14]}} , in176[14:3] };

   // m176_70 = W*in
   wire signed [14:0] m176_70;
   assign m176_70 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_71 = W*in
   wire signed [14:0] m176_71;
   assign m176_71 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_72 = W*in
   wire signed [14:0] m176_72;
   assign m176_72 =15'b0;

   // m176_73 = W*in
   wire signed [14:0] m176_73;
   assign m176_73 =15'b0;

   // m176_74 = W*in
   wire signed [14:0] m176_74;
   assign m176_74 ={ {4{neg176[14]}} , neg176[14:4] };

   // m176_75 = W*in
   wire signed [14:0] m176_75;
   assign m176_75 ={ {3{in176[14]}} , in176[14:3] };

   // m176_76 = W*in
   wire signed [14:0] m176_76;
   assign m176_76 =15'b0;

   // m176_77 = W*in
   wire signed [14:0] m176_77;
   assign m176_77 =15'b0;

   // m176_78 = W*in
   wire signed [14:0] m176_78;
   assign m176_78 =15'b0;

   // m176_79 = W*in
   wire signed [14:0] m176_79;
   assign m176_79 =15'b0;

   // m176_80 = W*in
   wire signed [14:0] m176_80;
   assign m176_80 =15'b0;

   // m176_81 = W*in
   wire signed [14:0] m176_81;
   assign m176_81 =15'b0;

   // m176_82 = W*in
   wire signed [14:0] m176_82;
   assign m176_82 =15'b0;

   // m176_83 = W*in
   wire signed [14:0] m176_83;
   assign m176_83 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_84 = W*in
   wire signed [14:0] m176_84;
   assign m176_84 =15'b0;

   // m176_85 = W*in
   wire signed [14:0] m176_85;
   assign m176_85 =15'b0;

   // m176_86 = W*in
   wire signed [14:0] m176_86;
   assign m176_86 =15'b0;

   // m176_87 = W*in
   wire signed [14:0] m176_87;
   assign m176_87 =15'b0;

   // m176_88 = W*in
   wire signed [14:0] m176_88;
   assign m176_88 =15'b0;

   // m176_89 = W*in
   wire signed [14:0] m176_89;
   assign m176_89 =15'b0;

   // m176_90 = W*in
   wire signed [14:0] m176_90;
   assign m176_90 =15'b0;

   // m176_91 = W*in
   wire signed [14:0] m176_91;
   assign m176_91 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_92 = W*in
   wire signed [14:0] m176_92;
   assign m176_92 ={ {3{in176[14]}} , in176[14:3] };

   // m176_93 = W*in
   wire signed [14:0] m176_93;
   assign m176_93 =15'b0;

   // m176_94 = W*in
   wire signed [14:0] m176_94;
   assign m176_94 ={ {3{neg176[14]}} , neg176[14:3] };

   // m176_95 = W*in
   wire signed [14:0] m176_95;
   assign m176_95 =15'b0;

   // m176_96 = W*in
   wire signed [14:0] m176_96;
   assign m176_96 =15'b0;

   // m176_97 = W*in
   wire signed [14:0] m176_97;
   assign m176_97 =15'b0;

   // m176_98 = W*in
   wire signed [14:0] m176_98;
   assign m176_98 =15'b0;

   // m176_99 = W*in
   wire signed [14:0] m176_99;
   assign m176_99 =15'b0;

   // m176_100 = W*in
   wire signed [14:0] m176_100;
   assign m176_100 =15'b0;

   // m177_1 = W*in
   wire signed [14:0] m177_1;
   assign m177_1 =15'b0;

   // m177_2 = W*in
   wire signed [14:0] m177_2;
   assign m177_2 =15'b0;

   // m177_3 = W*in
   wire signed [14:0] m177_3;
   assign m177_3 =15'b0;

   // m177_4 = W*in
   wire signed [14:0] m177_4;
   assign m177_4 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_5 = W*in
   wire signed [14:0] m177_5;
   assign m177_5 =15'b0;

   // m177_6 = W*in
   wire signed [14:0] m177_6;
   assign m177_6 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_7 = W*in
   wire signed [14:0] m177_7;
   assign m177_7 =15'b0;

   // m177_8 = W*in
   wire signed [14:0] m177_8;
   assign m177_8 =15'b0;

   // m177_9 = W*in
   wire signed [14:0] m177_9;
   assign m177_9 =15'b0;

   // m177_10 = W*in
   wire signed [14:0] m177_10;
   assign m177_10 =15'b0;

   // m177_11 = W*in
   wire signed [14:0] m177_11;
   assign m177_11 =15'b0;

   // m177_12 = W*in
   wire signed [14:0] m177_12;
   assign m177_12 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_13 = W*in
   wire signed [14:0] m177_13;
   assign m177_13 ={ {3{in177[14]}} , in177[14:3] };

   // m177_14 = W*in
   wire signed [14:0] m177_14;
   assign m177_14 =15'b0;

   // m177_15 = W*in
   wire signed [14:0] m177_15;
   assign m177_15 =15'b0;

   // m177_16 = W*in
   wire signed [14:0] m177_16;
   assign m177_16 =15'b0;

   // m177_17 = W*in
   wire signed [14:0] m177_17;
   assign m177_17 =15'b0;

   // m177_18 = W*in
   wire signed [14:0] m177_18;
   assign m177_18 ={ {3{in177[14]}} , in177[14:3] };

   // m177_19 = W*in
   wire signed [14:0] m177_19;
   assign m177_19 =15'b0;

   // m177_20 = W*in
   wire signed [14:0] m177_20;
   assign m177_20 =15'b0;

   // m177_21 = W*in
   wire signed [14:0] m177_21;
   assign m177_21 =15'b0;

   // m177_22 = W*in
   wire signed [14:0] m177_22;
   assign m177_22 =15'b0;

   // m177_23 = W*in
   wire signed [14:0] m177_23;
   assign m177_23 =15'b0;

   // m177_24 = W*in
   wire signed [14:0] m177_24;
   assign m177_24 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_25 = W*in
   wire signed [14:0] m177_25;
   assign m177_25 =15'b0;

   // m177_26 = W*in
   wire signed [14:0] m177_26;
   assign m177_26 ={ {4{neg177[14]}} , neg177[14:4] };

   // m177_27 = W*in
   wire signed [14:0] m177_27;
   assign m177_27 =15'b0;

   // m177_28 = W*in
   wire signed [14:0] m177_28;
   assign m177_28 ={ {4{in177[14]}} , in177[14:4] };

   // m177_29 = W*in
   wire signed [14:0] m177_29;
   assign m177_29 =15'b0;

   // m177_30 = W*in
   wire signed [14:0] m177_30;
   assign m177_30 =15'b0;

   // m177_31 = W*in
   wire signed [14:0] m177_31;
   assign m177_31 =15'b0;

   // m177_32 = W*in
   wire signed [14:0] m177_32;
   assign m177_32 =15'b0;

   // m177_33 = W*in
   wire signed [14:0] m177_33;
   assign m177_33 =15'b0;

   // m177_34 = W*in
   wire signed [14:0] m177_34;
   assign m177_34 =15'b0;

   // m177_35 = W*in
   wire signed [14:0] m177_35;
   assign m177_35 =15'b0;

   // m177_36 = W*in
   wire signed [14:0] m177_36;
   assign m177_36 =15'b0;

   // m177_37 = W*in
   wire signed [14:0] m177_37;
   assign m177_37 =15'b0;

   // m177_38 = W*in
   wire signed [14:0] m177_38;
   assign m177_38 ={ {3{in177[14]}} , in177[14:3] };

   // m177_39 = W*in
   wire signed [14:0] m177_39;
   assign m177_39 =15'b0;

   // m177_40 = W*in
   wire signed [14:0] m177_40;
   assign m177_40 ={ {3{in177[14]}} , in177[14:3] };

   // m177_41 = W*in
   wire signed [14:0] m177_41;
   assign m177_41 =15'b0;

   // m177_42 = W*in
   wire signed [14:0] m177_42;
   assign m177_42 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_43 = W*in
   wire signed [14:0] m177_43;
   assign m177_43 =15'b0;

   // m177_44 = W*in
   wire signed [14:0] m177_44;
   assign m177_44 =15'b0;

   // m177_45 = W*in
   wire signed [14:0] m177_45;
   assign m177_45 =15'b0;

   // m177_46 = W*in
   wire signed [14:0] m177_46;
   assign m177_46 =15'b0;

   // m177_47 = W*in
   wire signed [14:0] m177_47;
   assign m177_47 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_48 = W*in
   wire signed [14:0] m177_48;
   assign m177_48 =15'b0;

   // m177_49 = W*in
   wire signed [14:0] m177_49;
   assign m177_49 =15'b0;

   // m177_50 = W*in
   wire signed [14:0] m177_50;
   assign m177_50 =15'b0;

   // m177_51 = W*in
   wire signed [14:0] m177_51;
   assign m177_51 =15'b0;

   // m177_52 = W*in
   wire signed [14:0] m177_52;
   assign m177_52 =15'b0;

   // m177_53 = W*in
   wire signed [14:0] m177_53;
   assign m177_53 =15'b0;

   // m177_54 = W*in
   wire signed [14:0] m177_54;
   assign m177_54 =15'b0;

   // m177_55 = W*in
   wire signed [14:0] m177_55;
   assign m177_55 ={ {3{in177[14]}} , in177[14:3] };

   // m177_56 = W*in
   wire signed [14:0] m177_56;
   assign m177_56 ={ {3{in177[14]}} , in177[14:3] };

   // m177_57 = W*in
   wire signed [14:0] m177_57;
   assign m177_57 =15'b0;

   // m177_58 = W*in
   wire signed [14:0] m177_58;
   assign m177_58 =15'b0;

   // m177_59 = W*in
   wire signed [14:0] m177_59;
   assign m177_59 =15'b0;

   // m177_60 = W*in
   wire signed [14:0] m177_60;
   assign m177_60 =15'b0;

   // m177_61 = W*in
   wire signed [14:0] m177_61;
   assign m177_61 =15'b0;

   // m177_62 = W*in
   wire signed [14:0] m177_62;
   assign m177_62 =15'b0;

   // m177_63 = W*in
   wire signed [14:0] m177_63;
   assign m177_63 =15'b0;

   // m177_64 = W*in
   wire signed [14:0] m177_64;
   assign m177_64 =15'b0;

   // m177_65 = W*in
   wire signed [14:0] m177_65;
   assign m177_65 =15'b0;

   // m177_66 = W*in
   wire signed [14:0] m177_66;
   assign m177_66 =15'b0;

   // m177_67 = W*in
   wire signed [14:0] m177_67;
   assign m177_67 =15'b0;

   // m177_68 = W*in
   wire signed [14:0] m177_68;
   assign m177_68 ={ {3{in177[14]}} , in177[14:3] };

   // m177_69 = W*in
   wire signed [14:0] m177_69;
   assign m177_69 =15'b0;

   // m177_70 = W*in
   wire signed [14:0] m177_70;
   assign m177_70 =15'b0;

   // m177_71 = W*in
   wire signed [14:0] m177_71;
   assign m177_71 =15'b0;

   // m177_72 = W*in
   wire signed [14:0] m177_72;
   assign m177_72 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_73 = W*in
   wire signed [14:0] m177_73;
   assign m177_73 =15'b0;

   // m177_74 = W*in
   wire signed [14:0] m177_74;
   assign m177_74 =15'b0;

   // m177_75 = W*in
   wire signed [14:0] m177_75;
   assign m177_75 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_76 = W*in
   wire signed [14:0] m177_76;
   assign m177_76 =15'b0;

   // m177_77 = W*in
   wire signed [14:0] m177_77;
   assign m177_77 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_78 = W*in
   wire signed [14:0] m177_78;
   assign m177_78 =15'b0;

   // m177_79 = W*in
   wire signed [14:0] m177_79;
   assign m177_79 =15'b0;

   // m177_80 = W*in
   wire signed [14:0] m177_80;
   assign m177_80 =15'b0;

   // m177_81 = W*in
   wire signed [14:0] m177_81;
   assign m177_81 =15'b0;

   // m177_82 = W*in
   wire signed [14:0] m177_82;
   assign m177_82 =15'b0;

   // m177_83 = W*in
   wire signed [14:0] m177_83;
   assign m177_83 =15'b0;

   // m177_84 = W*in
   wire signed [14:0] m177_84;
   assign m177_84 =15'b0;

   // m177_85 = W*in
   wire signed [14:0] m177_85;
   assign m177_85 =15'b0;

   // m177_86 = W*in
   wire signed [14:0] m177_86;
   assign m177_86 =15'b0;

   // m177_87 = W*in
   wire signed [14:0] m177_87;
   assign m177_87 =15'b0;

   // m177_88 = W*in
   wire signed [14:0] m177_88;
   assign m177_88 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_89 = W*in
   wire signed [14:0] m177_89;
   assign m177_89 =15'b0;

   // m177_90 = W*in
   wire signed [14:0] m177_90;
   assign m177_90 =15'b0;

   // m177_91 = W*in
   wire signed [14:0] m177_91;
   assign m177_91 =15'b0;

   // m177_92 = W*in
   wire signed [14:0] m177_92;
   assign m177_92 =15'b0;

   // m177_93 = W*in
   wire signed [14:0] m177_93;
   assign m177_93 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_94 = W*in
   wire signed [14:0] m177_94;
   assign m177_94 =15'b0;

   // m177_95 = W*in
   wire signed [14:0] m177_95;
   assign m177_95 =15'b0;

   // m177_96 = W*in
   wire signed [14:0] m177_96;
   assign m177_96 ={ {3{neg177[14]}} , neg177[14:3] };

   // m177_97 = W*in
   wire signed [14:0] m177_97;
   assign m177_97 =15'b0;

   // m177_98 = W*in
   wire signed [14:0] m177_98;
   assign m177_98 =15'b0;

   // m177_99 = W*in
   wire signed [14:0] m177_99;
   assign m177_99 =15'b0;

   // m177_100 = W*in
   wire signed [14:0] m177_100;
   assign m177_100 =15'b0;

   // m178_1 = W*in
   wire signed [14:0] m178_1;
   assign m178_1 =15'b0;

   // m178_2 = W*in
   wire signed [14:0] m178_2;
   assign m178_2 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_3 = W*in
   wire signed [14:0] m178_3;
   assign m178_3 ={ {3{in178[14]}} , in178[14:3] };

   // m178_4 = W*in
   wire signed [14:0] m178_4;
   assign m178_4 =15'b0;

   // m178_5 = W*in
   wire signed [14:0] m178_5;
   assign m178_5 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_6 = W*in
   wire signed [14:0] m178_6;
   assign m178_6 =15'b0;

   // m178_7 = W*in
   wire signed [14:0] m178_7;
   assign m178_7 ={ {3{in178[14]}} , in178[14:3] };

   // m178_8 = W*in
   wire signed [14:0] m178_8;
   assign m178_8 ={ {3{in178[14]}} , in178[14:3] };

   // m178_9 = W*in
   wire signed [14:0] m178_9;
   assign m178_9 =15'b0;

   // m178_10 = W*in
   wire signed [14:0] m178_10;
   assign m178_10 =15'b0;

   // m178_11 = W*in
   wire signed [14:0] m178_11;
   assign m178_11 =15'b0;

   // m178_12 = W*in
   wire signed [14:0] m178_12;
   assign m178_12 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_13 = W*in
   wire signed [14:0] m178_13;
   assign m178_13 =15'b0;

   // m178_14 = W*in
   wire signed [14:0] m178_14;
   assign m178_14 =15'b0;

   // m178_15 = W*in
   wire signed [14:0] m178_15;
   assign m178_15 =15'b0;

   // m178_16 = W*in
   wire signed [14:0] m178_16;
   assign m178_16 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_17 = W*in
   wire signed [14:0] m178_17;
   assign m178_17 =15'b0;

   // m178_18 = W*in
   wire signed [14:0] m178_18;
   assign m178_18 ={ {3{in178[14]}} , in178[14:3] };

   // m178_19 = W*in
   wire signed [14:0] m178_19;
   assign m178_19 =15'b0;

   // m178_20 = W*in
   wire signed [14:0] m178_20;
   assign m178_20 =15'b0;

   // m178_21 = W*in
   wire signed [14:0] m178_21;
   assign m178_21 ={ {3{in178[14]}} , in178[14:3] };

   // m178_22 = W*in
   wire signed [14:0] m178_22;
   assign m178_22 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_23 = W*in
   wire signed [14:0] m178_23;
   assign m178_23 =15'b0;

   // m178_24 = W*in
   wire signed [14:0] m178_24;
   assign m178_24 =15'b0;

   // m178_25 = W*in
   wire signed [14:0] m178_25;
   assign m178_25 =15'b0;

   // m178_26 = W*in
   wire signed [14:0] m178_26;
   assign m178_26 ={ {4{neg178[14]}} , neg178[14:4] };

   // m178_27 = W*in
   wire signed [14:0] m178_27;
   assign m178_27 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_28 = W*in
   wire signed [14:0] m178_28;
   assign m178_28 ={ {3{in178[14]}} , in178[14:3] };

   // m178_29 = W*in
   wire signed [14:0] m178_29;
   assign m178_29 =15'b0;

   // m178_30 = W*in
   wire signed [14:0] m178_30;
   assign m178_30 =15'b0;

   // m178_31 = W*in
   wire signed [14:0] m178_31;
   assign m178_31 =15'b0;

   // m178_32 = W*in
   wire signed [14:0] m178_32;
   assign m178_32 =15'b0;

   // m178_33 = W*in
   wire signed [14:0] m178_33;
   assign m178_33 =15'b0;

   // m178_34 = W*in
   wire signed [14:0] m178_34;
   assign m178_34 =15'b0;

   // m178_35 = W*in
   wire signed [14:0] m178_35;
   assign m178_35 =15'b0;

   // m178_36 = W*in
   wire signed [14:0] m178_36;
   assign m178_36 =15'b0;

   // m178_37 = W*in
   wire signed [14:0] m178_37;
   assign m178_37 ={ {3{in178[14]}} , in178[14:3] };

   // m178_38 = W*in
   wire signed [14:0] m178_38;
   assign m178_38 =15'b0;

   // m178_39 = W*in
   wire signed [14:0] m178_39;
   assign m178_39 =15'b0;

   // m178_40 = W*in
   wire signed [14:0] m178_40;
   assign m178_40 =15'b0;

   // m178_41 = W*in
   wire signed [14:0] m178_41;
   assign m178_41 =15'b0;

   // m178_42 = W*in
   wire signed [14:0] m178_42;
   assign m178_42 =15'b0;

   // m178_43 = W*in
   wire signed [14:0] m178_43;
   assign m178_43 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_44 = W*in
   wire signed [14:0] m178_44;
   assign m178_44 ={ {3{in178[14]}} , in178[14:3] };

   // m178_45 = W*in
   wire signed [14:0] m178_45;
   assign m178_45 =15'b0;

   // m178_46 = W*in
   wire signed [14:0] m178_46;
   assign m178_46 =15'b0;

   // m178_47 = W*in
   wire signed [14:0] m178_47;
   assign m178_47 =15'b0;

   // m178_48 = W*in
   wire signed [14:0] m178_48;
   assign m178_48 ={ {4{in178[14]}} , in178[14:4] };

   // m178_49 = W*in
   wire signed [14:0] m178_49;
   assign m178_49 =15'b0;

   // m178_50 = W*in
   wire signed [14:0] m178_50;
   assign m178_50 =15'b0;

   // m178_51 = W*in
   wire signed [14:0] m178_51;
   assign m178_51 ={ {3{in178[14]}} , in178[14:3] };

   // m178_52 = W*in
   wire signed [14:0] m178_52;
   assign m178_52 =15'b0;

   // m178_53 = W*in
   wire signed [14:0] m178_53;
   assign m178_53 =15'b0;

   // m178_54 = W*in
   wire signed [14:0] m178_54;
   assign m178_54 =15'b0;

   // m178_55 = W*in
   wire signed [14:0] m178_55;
   assign m178_55 =15'b0;

   // m178_56 = W*in
   wire signed [14:0] m178_56;
   assign m178_56 ={ {3{in178[14]}} , in178[14:3] };

   // m178_57 = W*in
   wire signed [14:0] m178_57;
   assign m178_57 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_58 = W*in
   wire signed [14:0] m178_58;
   assign m178_58 ={ {4{neg178[14]}} , neg178[14:4] };

   // m178_59 = W*in
   wire signed [14:0] m178_59;
   assign m178_59 =15'b0;

   // m178_60 = W*in
   wire signed [14:0] m178_60;
   assign m178_60 =15'b0;

   // m178_61 = W*in
   wire signed [14:0] m178_61;
   assign m178_61 ={ {4{neg178[14]}} , neg178[14:4] };

   // m178_62 = W*in
   wire signed [14:0] m178_62;
   assign m178_62 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_63 = W*in
   wire signed [14:0] m178_63;
   assign m178_63 =15'b0;

   // m178_64 = W*in
   wire signed [14:0] m178_64;
   assign m178_64 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_65 = W*in
   wire signed [14:0] m178_65;
   assign m178_65 =15'b0;

   // m178_66 = W*in
   wire signed [14:0] m178_66;
   assign m178_66 =15'b0;

   // m178_67 = W*in
   wire signed [14:0] m178_67;
   assign m178_67 =15'b0;

   // m178_68 = W*in
   wire signed [14:0] m178_68;
   assign m178_68 =15'b0;

   // m178_69 = W*in
   wire signed [14:0] m178_69;
   assign m178_69 ={ {3{in178[14]}} , in178[14:3] };

   // m178_70 = W*in
   wire signed [14:0] m178_70;
   assign m178_70 ={ {3{in178[14]}} , in178[14:3] };

   // m178_71 = W*in
   wire signed [14:0] m178_71;
   assign m178_71 ={ {3{in178[14]}} , in178[14:3] };

   // m178_72 = W*in
   wire signed [14:0] m178_72;
   assign m178_72 =15'b0;

   // m178_73 = W*in
   wire signed [14:0] m178_73;
   assign m178_73 =15'b0;

   // m178_74 = W*in
   wire signed [14:0] m178_74;
   assign m178_74 ={ {4{in178[14]}} , in178[14:4] };

   // m178_75 = W*in
   wire signed [14:0] m178_75;
   assign m178_75 ={ {4{neg178[14]}} , neg178[14:4] };

   // m178_76 = W*in
   wire signed [14:0] m178_76;
   assign m178_76 ={ {4{neg178[14]}} , neg178[14:4] };

   // m178_77 = W*in
   wire signed [14:0] m178_77;
   assign m178_77 ={ {3{in178[14]}} , in178[14:3] };

   // m178_78 = W*in
   wire signed [14:0] m178_78;
   assign m178_78 =15'b0;

   // m178_79 = W*in
   wire signed [14:0] m178_79;
   assign m178_79 =15'b0;

   // m178_80 = W*in
   wire signed [14:0] m178_80;
   assign m178_80 =15'b0;

   // m178_81 = W*in
   wire signed [14:0] m178_81;
   assign m178_81 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_82 = W*in
   wire signed [14:0] m178_82;
   assign m178_82 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_83 = W*in
   wire signed [14:0] m178_83;
   assign m178_83 =15'b0;

   // m178_84 = W*in
   wire signed [14:0] m178_84;
   assign m178_84 =15'b0;

   // m178_85 = W*in
   wire signed [14:0] m178_85;
   assign m178_85 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_86 = W*in
   wire signed [14:0] m178_86;
   assign m178_86 =15'b0;

   // m178_87 = W*in
   wire signed [14:0] m178_87;
   assign m178_87 =15'b0;

   // m178_88 = W*in
   wire signed [14:0] m178_88;
   assign m178_88 ={ {3{in178[14]}} , in178[14:3] };

   // m178_89 = W*in
   wire signed [14:0] m178_89;
   assign m178_89 ={ {3{in178[14]}} , in178[14:3] };

   // m178_90 = W*in
   wire signed [14:0] m178_90;
   assign m178_90 =15'b0;

   // m178_91 = W*in
   wire signed [14:0] m178_91;
   assign m178_91 =15'b0;

   // m178_92 = W*in
   wire signed [14:0] m178_92;
   assign m178_92 =15'b0;

   // m178_93 = W*in
   wire signed [14:0] m178_93;
   assign m178_93 =15'b0;

   // m178_94 = W*in
   wire signed [14:0] m178_94;
   assign m178_94 =15'b0;

   // m178_95 = W*in
   wire signed [14:0] m178_95;
   assign m178_95 =15'b0;

   // m178_96 = W*in
   wire signed [14:0] m178_96;
   assign m178_96 =15'b0;

   // m178_97 = W*in
   wire signed [14:0] m178_97;
   assign m178_97 ={ {3{neg178[14]}} , neg178[14:3] };

   // m178_98 = W*in
   wire signed [14:0] m178_98;
   assign m178_98 ={ {3{in178[14]}} , in178[14:3] };

   // m178_99 = W*in
   wire signed [14:0] m178_99;
   assign m178_99 =15'b0;

   // m178_100 = W*in
   wire signed [14:0] m178_100;
   assign m178_100 =15'b0;

   // m179_1 = W*in
   wire signed [14:0] m179_1;
   assign m179_1 =15'b0;

   // m179_2 = W*in
   wire signed [14:0] m179_2;
   assign m179_2 =15'b0;

   // m179_3 = W*in
   wire signed [14:0] m179_3;
   assign m179_3 =15'b0;

   // m179_4 = W*in
   wire signed [14:0] m179_4;
   assign m179_4 =15'b0;

   // m179_5 = W*in
   wire signed [14:0] m179_5;
   assign m179_5 =15'b0;

   // m179_6 = W*in
   wire signed [14:0] m179_6;
   assign m179_6 =15'b0;

   // m179_7 = W*in
   wire signed [14:0] m179_7;
   assign m179_7 =15'b0;

   // m179_8 = W*in
   wire signed [14:0] m179_8;
   assign m179_8 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_9 = W*in
   wire signed [14:0] m179_9;
   assign m179_9 =15'b0;

   // m179_10 = W*in
   wire signed [14:0] m179_10;
   assign m179_10 =15'b0;

   // m179_11 = W*in
   wire signed [14:0] m179_11;
   assign m179_11 =15'b0;

   // m179_12 = W*in
   wire signed [14:0] m179_12;
   assign m179_12 =15'b0;

   // m179_13 = W*in
   wire signed [14:0] m179_13;
   assign m179_13 =15'b0;

   // m179_14 = W*in
   wire signed [14:0] m179_14;
   assign m179_14 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_15 = W*in
   wire signed [14:0] m179_15;
   assign m179_15 ={ {3{in179[14]}} , in179[14:3] };

   // m179_16 = W*in
   wire signed [14:0] m179_16;
   assign m179_16 =15'b0;

   // m179_17 = W*in
   wire signed [14:0] m179_17;
   assign m179_17 =15'b0;

   // m179_18 = W*in
   wire signed [14:0] m179_18;
   assign m179_18 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_19 = W*in
   wire signed [14:0] m179_19;
   assign m179_19 ={ {3{in179[14]}} , in179[14:3] };

   // m179_20 = W*in
   wire signed [14:0] m179_20;
   assign m179_20 =15'b0;

   // m179_21 = W*in
   wire signed [14:0] m179_21;
   assign m179_21 ={ {4{neg179[14]}} , neg179[14:4] };

   // m179_22 = W*in
   wire signed [14:0] m179_22;
   assign m179_22 =15'b0;

   // m179_23 = W*in
   wire signed [14:0] m179_23;
   assign m179_23 =15'b0;

   // m179_24 = W*in
   wire signed [14:0] m179_24;
   assign m179_24 =15'b0;

   // m179_25 = W*in
   wire signed [14:0] m179_25;
   assign m179_25 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_26 = W*in
   wire signed [14:0] m179_26;
   assign m179_26 =15'b0;

   // m179_27 = W*in
   wire signed [14:0] m179_27;
   assign m179_27 =15'b0;

   // m179_28 = W*in
   wire signed [14:0] m179_28;
   assign m179_28 =15'b0;

   // m179_29 = W*in
   wire signed [14:0] m179_29;
   assign m179_29 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_30 = W*in
   wire signed [14:0] m179_30;
   assign m179_30 =15'b0;

   // m179_31 = W*in
   wire signed [14:0] m179_31;
   assign m179_31 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_32 = W*in
   wire signed [14:0] m179_32;
   assign m179_32 =15'b0;

   // m179_33 = W*in
   wire signed [14:0] m179_33;
   assign m179_33 =15'b0;

   // m179_34 = W*in
   wire signed [14:0] m179_34;
   assign m179_34 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_35 = W*in
   wire signed [14:0] m179_35;
   assign m179_35 ={ {3{in179[14]}} , in179[14:3] };

   // m179_36 = W*in
   wire signed [14:0] m179_36;
   assign m179_36 =15'b0;

   // m179_37 = W*in
   wire signed [14:0] m179_37;
   assign m179_37 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_38 = W*in
   wire signed [14:0] m179_38;
   assign m179_38 ={ {3{in179[14]}} , in179[14:3] };

   // m179_39 = W*in
   wire signed [14:0] m179_39;
   assign m179_39 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_40 = W*in
   wire signed [14:0] m179_40;
   assign m179_40 =15'b0;

   // m179_41 = W*in
   wire signed [14:0] m179_41;
   assign m179_41 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_42 = W*in
   wire signed [14:0] m179_42;
   assign m179_42 ={ {3{in179[14]}} , in179[14:3] };

   // m179_43 = W*in
   wire signed [14:0] m179_43;
   assign m179_43 =15'b0;

   // m179_44 = W*in
   wire signed [14:0] m179_44;
   assign m179_44 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_45 = W*in
   wire signed [14:0] m179_45;
   assign m179_45 =15'b0;

   // m179_46 = W*in
   wire signed [14:0] m179_46;
   assign m179_46 ={ {3{in179[14]}} , in179[14:3] };

   // m179_47 = W*in
   wire signed [14:0] m179_47;
   assign m179_47 =15'b0;

   // m179_48 = W*in
   wire signed [14:0] m179_48;
   assign m179_48 =15'b0;

   // m179_49 = W*in
   wire signed [14:0] m179_49;
   assign m179_49 ={ {3{in179[14]}} , in179[14:3] };

   // m179_50 = W*in
   wire signed [14:0] m179_50;
   assign m179_50 ={ {3{in179[14]}} , in179[14:3] };

   // m179_51 = W*in
   wire signed [14:0] m179_51;
   assign m179_51 =15'b0;

   // m179_52 = W*in
   wire signed [14:0] m179_52;
   assign m179_52 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_53 = W*in
   wire signed [14:0] m179_53;
   assign m179_53 =15'b0;

   // m179_54 = W*in
   wire signed [14:0] m179_54;
   assign m179_54 =15'b0;

   // m179_55 = W*in
   wire signed [14:0] m179_55;
   assign m179_55 =15'b0;

   // m179_56 = W*in
   wire signed [14:0] m179_56;
   assign m179_56 ={ {3{in179[14]}} , in179[14:3] };

   // m179_57 = W*in
   wire signed [14:0] m179_57;
   assign m179_57 =15'b0;

   // m179_58 = W*in
   wire signed [14:0] m179_58;
   assign m179_58 =15'b0;

   // m179_59 = W*in
   wire signed [14:0] m179_59;
   assign m179_59 ={ {4{in179[14]}} , in179[14:4] };

   // m179_60 = W*in
   wire signed [14:0] m179_60;
   assign m179_60 ={ {4{neg179[14]}} , neg179[14:4] };

   // m179_61 = W*in
   wire signed [14:0] m179_61;
   assign m179_61 =15'b0;

   // m179_62 = W*in
   wire signed [14:0] m179_62;
   assign m179_62 =15'b0;

   // m179_63 = W*in
   wire signed [14:0] m179_63;
   assign m179_63 =15'b0;

   // m179_64 = W*in
   wire signed [14:0] m179_64;
   assign m179_64 =15'b0;

   // m179_65 = W*in
   wire signed [14:0] m179_65;
   assign m179_65 =15'b0;

   // m179_66 = W*in
   wire signed [14:0] m179_66;
   assign m179_66 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_67 = W*in
   wire signed [14:0] m179_67;
   assign m179_67 ={ {3{in179[14]}} , in179[14:3] };

   // m179_68 = W*in
   wire signed [14:0] m179_68;
   assign m179_68 =15'b0;

   // m179_69 = W*in
   wire signed [14:0] m179_69;
   assign m179_69 =15'b0;

   // m179_70 = W*in
   wire signed [14:0] m179_70;
   assign m179_70 ={ {3{in179[14]}} , in179[14:3] };

   // m179_71 = W*in
   wire signed [14:0] m179_71;
   assign m179_71 =15'b0;

   // m179_72 = W*in
   wire signed [14:0] m179_72;
   assign m179_72 =15'b0;

   // m179_73 = W*in
   wire signed [14:0] m179_73;
   assign m179_73 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_74 = W*in
   wire signed [14:0] m179_74;
   assign m179_74 =15'b0;

   // m179_75 = W*in
   wire signed [14:0] m179_75;
   assign m179_75 ={ {3{in179[14]}} , in179[14:3] };

   // m179_76 = W*in
   wire signed [14:0] m179_76;
   assign m179_76 ={ {4{neg179[14]}} , neg179[14:4] };

   // m179_77 = W*in
   wire signed [14:0] m179_77;
   assign m179_77 =15'b0;

   // m179_78 = W*in
   wire signed [14:0] m179_78;
   assign m179_78 =15'b0;

   // m179_79 = W*in
   wire signed [14:0] m179_79;
   assign m179_79 =15'b0;

   // m179_80 = W*in
   wire signed [14:0] m179_80;
   assign m179_80 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_81 = W*in
   wire signed [14:0] m179_81;
   assign m179_81 ={ {3{in179[14]}} , in179[14:3] };

   // m179_82 = W*in
   wire signed [14:0] m179_82;
   assign m179_82 =15'b0;

   // m179_83 = W*in
   wire signed [14:0] m179_83;
   assign m179_83 =15'b0;

   // m179_84 = W*in
   wire signed [14:0] m179_84;
   assign m179_84 ={ {4{in179[14]}} , in179[14:4] };

   // m179_85 = W*in
   wire signed [14:0] m179_85;
   assign m179_85 ={ {3{in179[14]}} , in179[14:3] };

   // m179_86 = W*in
   wire signed [14:0] m179_86;
   assign m179_86 ={ {3{in179[14]}} , in179[14:3] };

   // m179_87 = W*in
   wire signed [14:0] m179_87;
   assign m179_87 ={ {3{in179[14]}} , in179[14:3] };

   // m179_88 = W*in
   wire signed [14:0] m179_88;
   assign m179_88 =15'b0;

   // m179_89 = W*in
   wire signed [14:0] m179_89;
   assign m179_89 =15'b0;

   // m179_90 = W*in
   wire signed [14:0] m179_90;
   assign m179_90 =15'b0;

   // m179_91 = W*in
   wire signed [14:0] m179_91;
   assign m179_91 =15'b0;

   // m179_92 = W*in
   wire signed [14:0] m179_92;
   assign m179_92 =15'b0;

   // m179_93 = W*in
   wire signed [14:0] m179_93;
   assign m179_93 ={ {3{in179[14]}} , in179[14:3] };

   // m179_94 = W*in
   wire signed [14:0] m179_94;
   assign m179_94 =15'b0;

   // m179_95 = W*in
   wire signed [14:0] m179_95;
   assign m179_95 ={ {3{in179[14]}} , in179[14:3] };

   // m179_96 = W*in
   wire signed [14:0] m179_96;
   assign m179_96 ={ {3{neg179[14]}} , neg179[14:3] };

   // m179_97 = W*in
   wire signed [14:0] m179_97;
   assign m179_97 =15'b0;

   // m179_98 = W*in
   wire signed [14:0] m179_98;
   assign m179_98 =15'b0;

   // m179_99 = W*in
   wire signed [14:0] m179_99;
   assign m179_99 =15'b0;

   // m179_100 = W*in
   wire signed [14:0] m179_100;
   assign m179_100 =15'b0;

   // m180_1 = W*in
   wire signed [14:0] m180_1;
   assign m180_1 =15'b0;

   // m180_2 = W*in
   wire signed [14:0] m180_2;
   assign m180_2 =15'b0;

   // m180_3 = W*in
   wire signed [14:0] m180_3;
   assign m180_3 =15'b0;

   // m180_4 = W*in
   wire signed [14:0] m180_4;
   assign m180_4 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_5 = W*in
   wire signed [14:0] m180_5;
   assign m180_5 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_6 = W*in
   wire signed [14:0] m180_6;
   assign m180_6 ={ {3{in180[14]}} , in180[14:3] };

   // m180_7 = W*in
   wire signed [14:0] m180_7;
   assign m180_7 ={ {3{in180[14]}} , in180[14:3] };

   // m180_8 = W*in
   wire signed [14:0] m180_8;
   assign m180_8 ={ {3{in180[14]}} , in180[14:3] };

   // m180_9 = W*in
   wire signed [14:0] m180_9;
   assign m180_9 =15'b0;

   // m180_10 = W*in
   wire signed [14:0] m180_10;
   assign m180_10 =15'b0;

   // m180_11 = W*in
   wire signed [14:0] m180_11;
   assign m180_11 =15'b0;

   // m180_12 = W*in
   wire signed [14:0] m180_12;
   assign m180_12 =15'b0;

   // m180_13 = W*in
   wire signed [14:0] m180_13;
   assign m180_13 =15'b0;

   // m180_14 = W*in
   wire signed [14:0] m180_14;
   assign m180_14 ={ {3{in180[14]}} , in180[14:3] };

   // m180_15 = W*in
   wire signed [14:0] m180_15;
   assign m180_15 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_16 = W*in
   wire signed [14:0] m180_16;
   assign m180_16 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_17 = W*in
   wire signed [14:0] m180_17;
   assign m180_17 =15'b0;

   // m180_18 = W*in
   wire signed [14:0] m180_18;
   assign m180_18 ={ {3{in180[14]}} , in180[14:3] };

   // m180_19 = W*in
   wire signed [14:0] m180_19;
   assign m180_19 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_20 = W*in
   wire signed [14:0] m180_20;
   assign m180_20 =15'b0;

   // m180_21 = W*in
   wire signed [14:0] m180_21;
   assign m180_21 ={ {4{in180[14]}} , in180[14:4] };

   // m180_22 = W*in
   wire signed [14:0] m180_22;
   assign m180_22 =15'b0;

   // m180_23 = W*in
   wire signed [14:0] m180_23;
   assign m180_23 ={ {3{in180[14]}} , in180[14:3] };

   // m180_24 = W*in
   wire signed [14:0] m180_24;
   assign m180_24 =15'b0;

   // m180_25 = W*in
   wire signed [14:0] m180_25;
   assign m180_25 =15'b0;

   // m180_26 = W*in
   wire signed [14:0] m180_26;
   assign m180_26 =15'b0;

   // m180_27 = W*in
   wire signed [14:0] m180_27;
   assign m180_27 =15'b0;

   // m180_28 = W*in
   wire signed [14:0] m180_28;
   assign m180_28 =15'b0;

   // m180_29 = W*in
   wire signed [14:0] m180_29;
   assign m180_29 =15'b0;

   // m180_30 = W*in
   wire signed [14:0] m180_30;
   assign m180_30 =15'b0;

   // m180_31 = W*in
   wire signed [14:0] m180_31;
   assign m180_31 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_32 = W*in
   wire signed [14:0] m180_32;
   assign m180_32 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_33 = W*in
   wire signed [14:0] m180_33;
   assign m180_33 =15'b0;

   // m180_34 = W*in
   wire signed [14:0] m180_34;
   assign m180_34 =15'b0;

   // m180_35 = W*in
   wire signed [14:0] m180_35;
   assign m180_35 =15'b0;

   // m180_36 = W*in
   wire signed [14:0] m180_36;
   assign m180_36 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_37 = W*in
   wire signed [14:0] m180_37;
   assign m180_37 =15'b0;

   // m180_38 = W*in
   wire signed [14:0] m180_38;
   assign m180_38 =15'b0;

   // m180_39 = W*in
   wire signed [14:0] m180_39;
   assign m180_39 =15'b0;

   // m180_40 = W*in
   wire signed [14:0] m180_40;
   assign m180_40 =15'b0;

   // m180_41 = W*in
   wire signed [14:0] m180_41;
   assign m180_41 ={ {2{in180[14]}} , in180[14:2] };

   // m180_42 = W*in
   wire signed [14:0] m180_42;
   assign m180_42 =15'b0;

   // m180_43 = W*in
   wire signed [14:0] m180_43;
   assign m180_43 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_44 = W*in
   wire signed [14:0] m180_44;
   assign m180_44 =15'b0;

   // m180_45 = W*in
   wire signed [14:0] m180_45;
   assign m180_45 =15'b0;

   // m180_46 = W*in
   wire signed [14:0] m180_46;
   assign m180_46 =15'b0;

   // m180_47 = W*in
   wire signed [14:0] m180_47;
   assign m180_47 ={ {4{neg180[14]}} , neg180[14:4] };

   // m180_48 = W*in
   wire signed [14:0] m180_48;
   assign m180_48 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_49 = W*in
   wire signed [14:0] m180_49;
   assign m180_49 =15'b0;

   // m180_50 = W*in
   wire signed [14:0] m180_50;
   assign m180_50 =15'b0;

   // m180_51 = W*in
   wire signed [14:0] m180_51;
   assign m180_51 =15'b0;

   // m180_52 = W*in
   wire signed [14:0] m180_52;
   assign m180_52 =15'b0;

   // m180_53 = W*in
   wire signed [14:0] m180_53;
   assign m180_53 =15'b0;

   // m180_54 = W*in
   wire signed [14:0] m180_54;
   assign m180_54 =15'b0;

   // m180_55 = W*in
   wire signed [14:0] m180_55;
   assign m180_55 =15'b0;

   // m180_56 = W*in
   wire signed [14:0] m180_56;
   assign m180_56 =15'b0;

   // m180_57 = W*in
   wire signed [14:0] m180_57;
   assign m180_57 =15'b0;

   // m180_58 = W*in
   wire signed [14:0] m180_58;
   assign m180_58 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_59 = W*in
   wire signed [14:0] m180_59;
   assign m180_59 ={ {4{neg180[14]}} , neg180[14:4] };

   // m180_60 = W*in
   wire signed [14:0] m180_60;
   assign m180_60 =15'b0;

   // m180_61 = W*in
   wire signed [14:0] m180_61;
   assign m180_61 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_62 = W*in
   wire signed [14:0] m180_62;
   assign m180_62 =15'b0;

   // m180_63 = W*in
   wire signed [14:0] m180_63;
   assign m180_63 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_64 = W*in
   wire signed [14:0] m180_64;
   assign m180_64 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_65 = W*in
   wire signed [14:0] m180_65;
   assign m180_65 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_66 = W*in
   wire signed [14:0] m180_66;
   assign m180_66 =15'b0;

   // m180_67 = W*in
   wire signed [14:0] m180_67;
   assign m180_67 =15'b0;

   // m180_68 = W*in
   wire signed [14:0] m180_68;
   assign m180_68 ={ {4{neg180[14]}} , neg180[14:4] };

   // m180_69 = W*in
   wire signed [14:0] m180_69;
   assign m180_69 =15'b0;

   // m180_70 = W*in
   wire signed [14:0] m180_70;
   assign m180_70 =15'b0;

   // m180_71 = W*in
   wire signed [14:0] m180_71;
   assign m180_71 =15'b0;

   // m180_72 = W*in
   wire signed [14:0] m180_72;
   assign m180_72 =15'b0;

   // m180_73 = W*in
   wire signed [14:0] m180_73;
   assign m180_73 =15'b0;

   // m180_74 = W*in
   wire signed [14:0] m180_74;
   assign m180_74 =15'b0;

   // m180_75 = W*in
   wire signed [14:0] m180_75;
   assign m180_75 =15'b0;

   // m180_76 = W*in
   wire signed [14:0] m180_76;
   assign m180_76 =15'b0;

   // m180_77 = W*in
   wire signed [14:0] m180_77;
   assign m180_77 =15'b0;

   // m180_78 = W*in
   wire signed [14:0] m180_78;
   assign m180_78 ={ {3{in180[14]}} , in180[14:3] };

   // m180_79 = W*in
   wire signed [14:0] m180_79;
   assign m180_79 =15'b0;

   // m180_80 = W*in
   wire signed [14:0] m180_80;
   assign m180_80 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_81 = W*in
   wire signed [14:0] m180_81;
   assign m180_81 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_82 = W*in
   wire signed [14:0] m180_82;
   assign m180_82 =15'b0;

   // m180_83 = W*in
   wire signed [14:0] m180_83;
   assign m180_83 =15'b0;

   // m180_84 = W*in
   wire signed [14:0] m180_84;
   assign m180_84 =15'b0;

   // m180_85 = W*in
   wire signed [14:0] m180_85;
   assign m180_85 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_86 = W*in
   wire signed [14:0] m180_86;
   assign m180_86 =15'b0;

   // m180_87 = W*in
   wire signed [14:0] m180_87;
   assign m180_87 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_88 = W*in
   wire signed [14:0] m180_88;
   assign m180_88 ={ {3{in180[14]}} , in180[14:3] };

   // m180_89 = W*in
   wire signed [14:0] m180_89;
   assign m180_89 =15'b0;

   // m180_90 = W*in
   wire signed [14:0] m180_90;
   assign m180_90 =15'b0;

   // m180_91 = W*in
   wire signed [14:0] m180_91;
   assign m180_91 =15'b0;

   // m180_92 = W*in
   wire signed [14:0] m180_92;
   assign m180_92 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_93 = W*in
   wire signed [14:0] m180_93;
   assign m180_93 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_94 = W*in
   wire signed [14:0] m180_94;
   assign m180_94 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_95 = W*in
   wire signed [14:0] m180_95;
   assign m180_95 ={ {3{neg180[14]}} , neg180[14:3] };

   // m180_96 = W*in
   wire signed [14:0] m180_96;
   assign m180_96 ={ {3{in180[14]}} , in180[14:3] };

   // m180_97 = W*in
   wire signed [14:0] m180_97;
   assign m180_97 =15'b0;

   // m180_98 = W*in
   wire signed [14:0] m180_98;
   assign m180_98 =15'b0;

   // m180_99 = W*in
   wire signed [14:0] m180_99;
   assign m180_99 =15'b0;

   // m180_100 = W*in
   wire signed [14:0] m180_100;
   assign m180_100 =15'b0;

   // m181_1 = W*in
   wire signed [14:0] m181_1;
   assign m181_1 =15'b0;

   // m181_2 = W*in
   wire signed [14:0] m181_2;
   assign m181_2 =15'b0;

   // m181_3 = W*in
   wire signed [14:0] m181_3;
   assign m181_3 =15'b0;

   // m181_4 = W*in
   wire signed [14:0] m181_4;
   assign m181_4 =15'b0;

   // m181_5 = W*in
   wire signed [14:0] m181_5;
   assign m181_5 =15'b0;

   // m181_6 = W*in
   wire signed [14:0] m181_6;
   assign m181_6 =15'b0;

   // m181_7 = W*in
   wire signed [14:0] m181_7;
   assign m181_7 =15'b0;

   // m181_8 = W*in
   wire signed [14:0] m181_8;
   assign m181_8 ={ {3{in181[14]}} , in181[14:3] };

   // m181_9 = W*in
   wire signed [14:0] m181_9;
   assign m181_9 =15'b0;

   // m181_10 = W*in
   wire signed [14:0] m181_10;
   assign m181_10 =15'b0;

   // m181_11 = W*in
   wire signed [14:0] m181_11;
   assign m181_11 =15'b0;

   // m181_12 = W*in
   wire signed [14:0] m181_12;
   assign m181_12 =15'b0;

   // m181_13 = W*in
   wire signed [14:0] m181_13;
   assign m181_13 =15'b0;

   // m181_14 = W*in
   wire signed [14:0] m181_14;
   assign m181_14 =15'b0;

   // m181_15 = W*in
   wire signed [14:0] m181_15;
   assign m181_15 =15'b0;

   // m181_16 = W*in
   wire signed [14:0] m181_16;
   assign m181_16 =15'b0;

   // m181_17 = W*in
   wire signed [14:0] m181_17;
   assign m181_17 =15'b0;

   // m181_18 = W*in
   wire signed [14:0] m181_18;
   assign m181_18 ={ {4{in181[14]}} , in181[14:4] };

   // m181_19 = W*in
   wire signed [14:0] m181_19;
   assign m181_19 =15'b0;

   // m181_20 = W*in
   wire signed [14:0] m181_20;
   assign m181_20 =15'b0;

   // m181_21 = W*in
   wire signed [14:0] m181_21;
   assign m181_21 =15'b0;

   // m181_22 = W*in
   wire signed [14:0] m181_22;
   assign m181_22 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_23 = W*in
   wire signed [14:0] m181_23;
   assign m181_23 =15'b0;

   // m181_24 = W*in
   wire signed [14:0] m181_24;
   assign m181_24 =15'b0;

   // m181_25 = W*in
   wire signed [14:0] m181_25;
   assign m181_25 =15'b0;

   // m181_26 = W*in
   wire signed [14:0] m181_26;
   assign m181_26 =15'b0;

   // m181_27 = W*in
   wire signed [14:0] m181_27;
   assign m181_27 ={ {4{neg181[14]}} , neg181[14:4] };

   // m181_28 = W*in
   wire signed [14:0] m181_28;
   assign m181_28 =15'b0;

   // m181_29 = W*in
   wire signed [14:0] m181_29;
   assign m181_29 ={ {4{in181[14]}} , in181[14:4] };

   // m181_30 = W*in
   wire signed [14:0] m181_30;
   assign m181_30 =15'b0;

   // m181_31 = W*in
   wire signed [14:0] m181_31;
   assign m181_31 ={ {3{in181[14]}} , in181[14:3] };

   // m181_32 = W*in
   wire signed [14:0] m181_32;
   assign m181_32 ={ {4{in181[14]}} , in181[14:4] };

   // m181_33 = W*in
   wire signed [14:0] m181_33;
   assign m181_33 =15'b0;

   // m181_34 = W*in
   wire signed [14:0] m181_34;
   assign m181_34 =15'b0;

   // m181_35 = W*in
   wire signed [14:0] m181_35;
   assign m181_35 =15'b0;

   // m181_36 = W*in
   wire signed [14:0] m181_36;
   assign m181_36 =15'b0;

   // m181_37 = W*in
   wire signed [14:0] m181_37;
   assign m181_37 =15'b0;

   // m181_38 = W*in
   wire signed [14:0] m181_38;
   assign m181_38 =15'b0;

   // m181_39 = W*in
   wire signed [14:0] m181_39;
   assign m181_39 =15'b0;

   // m181_40 = W*in
   wire signed [14:0] m181_40;
   assign m181_40 =15'b0;

   // m181_41 = W*in
   wire signed [14:0] m181_41;
   assign m181_41 =15'b0;

   // m181_42 = W*in
   wire signed [14:0] m181_42;
   assign m181_42 =15'b0;

   // m181_43 = W*in
   wire signed [14:0] m181_43;
   assign m181_43 =15'b0;

   // m181_44 = W*in
   wire signed [14:0] m181_44;
   assign m181_44 ={ {3{in181[14]}} , in181[14:3] };

   // m181_45 = W*in
   wire signed [14:0] m181_45;
   assign m181_45 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_46 = W*in
   wire signed [14:0] m181_46;
   assign m181_46 =15'b0;

   // m181_47 = W*in
   wire signed [14:0] m181_47;
   assign m181_47 =15'b0;

   // m181_48 = W*in
   wire signed [14:0] m181_48;
   assign m181_48 =15'b0;

   // m181_49 = W*in
   wire signed [14:0] m181_49;
   assign m181_49 =15'b0;

   // m181_50 = W*in
   wire signed [14:0] m181_50;
   assign m181_50 =15'b0;

   // m181_51 = W*in
   wire signed [14:0] m181_51;
   assign m181_51 =15'b0;

   // m181_52 = W*in
   wire signed [14:0] m181_52;
   assign m181_52 =15'b0;

   // m181_53 = W*in
   wire signed [14:0] m181_53;
   assign m181_53 =15'b0;

   // m181_54 = W*in
   wire signed [14:0] m181_54;
   assign m181_54 ={ {3{in181[14]}} , in181[14:3] };

   // m181_55 = W*in
   wire signed [14:0] m181_55;
   assign m181_55 =15'b0;

   // m181_56 = W*in
   wire signed [14:0] m181_56;
   assign m181_56 =15'b0;

   // m181_57 = W*in
   wire signed [14:0] m181_57;
   assign m181_57 =15'b0;

   // m181_58 = W*in
   wire signed [14:0] m181_58;
   assign m181_58 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_59 = W*in
   wire signed [14:0] m181_59;
   assign m181_59 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_60 = W*in
   wire signed [14:0] m181_60;
   assign m181_60 ={ {4{in181[14]}} , in181[14:4] };

   // m181_61 = W*in
   wire signed [14:0] m181_61;
   assign m181_61 ={ {4{neg181[14]}} , neg181[14:4] };

   // m181_62 = W*in
   wire signed [14:0] m181_62;
   assign m181_62 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_63 = W*in
   wire signed [14:0] m181_63;
   assign m181_63 =15'b0;

   // m181_64 = W*in
   wire signed [14:0] m181_64;
   assign m181_64 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_65 = W*in
   wire signed [14:0] m181_65;
   assign m181_65 ={ {4{in181[14]}} , in181[14:4] };

   // m181_66 = W*in
   wire signed [14:0] m181_66;
   assign m181_66 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_67 = W*in
   wire signed [14:0] m181_67;
   assign m181_67 =15'b0;

   // m181_68 = W*in
   wire signed [14:0] m181_68;
   assign m181_68 =15'b0;

   // m181_69 = W*in
   wire signed [14:0] m181_69;
   assign m181_69 ={ {4{in181[14]}} , in181[14:4] };

   // m181_70 = W*in
   wire signed [14:0] m181_70;
   assign m181_70 =15'b0;

   // m181_71 = W*in
   wire signed [14:0] m181_71;
   assign m181_71 =15'b0;

   // m181_72 = W*in
   wire signed [14:0] m181_72;
   assign m181_72 =15'b0;

   // m181_73 = W*in
   wire signed [14:0] m181_73;
   assign m181_73 =15'b0;

   // m181_74 = W*in
   wire signed [14:0] m181_74;
   assign m181_74 ={ {4{neg181[14]}} , neg181[14:4] };

   // m181_75 = W*in
   wire signed [14:0] m181_75;
   assign m181_75 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_76 = W*in
   wire signed [14:0] m181_76;
   assign m181_76 ={ {4{neg181[14]}} , neg181[14:4] };

   // m181_77 = W*in
   wire signed [14:0] m181_77;
   assign m181_77 =15'b0;

   // m181_78 = W*in
   wire signed [14:0] m181_78;
   assign m181_78 =15'b0;

   // m181_79 = W*in
   wire signed [14:0] m181_79;
   assign m181_79 =15'b0;

   // m181_80 = W*in
   wire signed [14:0] m181_80;
   assign m181_80 =15'b0;

   // m181_81 = W*in
   wire signed [14:0] m181_81;
   assign m181_81 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_82 = W*in
   wire signed [14:0] m181_82;
   assign m181_82 =15'b0;

   // m181_83 = W*in
   wire signed [14:0] m181_83;
   assign m181_83 =15'b0;

   // m181_84 = W*in
   wire signed [14:0] m181_84;
   assign m181_84 =15'b0;

   // m181_85 = W*in
   wire signed [14:0] m181_85;
   assign m181_85 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_86 = W*in
   wire signed [14:0] m181_86;
   assign m181_86 =15'b0;

   // m181_87 = W*in
   wire signed [14:0] m181_87;
   assign m181_87 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_88 = W*in
   wire signed [14:0] m181_88;
   assign m181_88 =15'b0;

   // m181_89 = W*in
   wire signed [14:0] m181_89;
   assign m181_89 =15'b0;

   // m181_90 = W*in
   wire signed [14:0] m181_90;
   assign m181_90 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_91 = W*in
   wire signed [14:0] m181_91;
   assign m181_91 =15'b0;

   // m181_92 = W*in
   wire signed [14:0] m181_92;
   assign m181_92 =15'b0;

   // m181_93 = W*in
   wire signed [14:0] m181_93;
   assign m181_93 ={ {3{neg181[14]}} , neg181[14:3] };

   // m181_94 = W*in
   wire signed [14:0] m181_94;
   assign m181_94 ={ {4{neg181[14]}} , neg181[14:4] };

   // m181_95 = W*in
   wire signed [14:0] m181_95;
   assign m181_95 =15'b0;

   // m181_96 = W*in
   wire signed [14:0] m181_96;
   assign m181_96 ={ {4{in181[14]}} , in181[14:4] };

   // m181_97 = W*in
   wire signed [14:0] m181_97;
   assign m181_97 =15'b0;

   // m181_98 = W*in
   wire signed [14:0] m181_98;
   assign m181_98 =15'b0;

   // m181_99 = W*in
   wire signed [14:0] m181_99;
   assign m181_99 =15'b0;

   // m181_100 = W*in
   wire signed [14:0] m181_100;
   assign m181_100 =15'b0;

   // m182_1 = W*in
   wire signed [14:0] m182_1;
   assign m182_1 ={ {4{neg182[14]}} , neg182[14:4] };

   // m182_2 = W*in
   wire signed [14:0] m182_2;
   assign m182_2 =15'b0;

   // m182_3 = W*in
   wire signed [14:0] m182_3;
   assign m182_3 ={ {4{in182[14]}} , in182[14:4] };

   // m182_4 = W*in
   wire signed [14:0] m182_4;
   assign m182_4 =15'b0;

   // m182_5 = W*in
   wire signed [14:0] m182_5;
   assign m182_5 =15'b0;

   // m182_6 = W*in
   wire signed [14:0] m182_6;
   assign m182_6 =15'b0;

   // m182_7 = W*in
   wire signed [14:0] m182_7;
   assign m182_7 =15'b0;

   // m182_8 = W*in
   wire signed [14:0] m182_8;
   assign m182_8 =15'b0;

   // m182_9 = W*in
   wire signed [14:0] m182_9;
   assign m182_9 =15'b0;

   // m182_10 = W*in
   wire signed [14:0] m182_10;
   assign m182_10 =15'b0;

   // m182_11 = W*in
   wire signed [14:0] m182_11;
   assign m182_11 =15'b0;

   // m182_12 = W*in
   wire signed [14:0] m182_12;
   assign m182_12 =15'b0;

   // m182_13 = W*in
   wire signed [14:0] m182_13;
   assign m182_13 =15'b0;

   // m182_14 = W*in
   wire signed [14:0] m182_14;
   assign m182_14 =15'b0;

   // m182_15 = W*in
   wire signed [14:0] m182_15;
   assign m182_15 =15'b0;

   // m182_16 = W*in
   wire signed [14:0] m182_16;
   assign m182_16 =15'b0;

   // m182_17 = W*in
   wire signed [14:0] m182_17;
   assign m182_17 =15'b0;

   // m182_18 = W*in
   wire signed [14:0] m182_18;
   assign m182_18 =15'b0;

   // m182_19 = W*in
   wire signed [14:0] m182_19;
   assign m182_19 =15'b0;

   // m182_20 = W*in
   wire signed [14:0] m182_20;
   assign m182_20 ={ {3{in182[14]}} , in182[14:3] };

   // m182_21 = W*in
   wire signed [14:0] m182_21;
   assign m182_21 =15'b0;

   // m182_22 = W*in
   wire signed [14:0] m182_22;
   assign m182_22 =15'b0;

   // m182_23 = W*in
   wire signed [14:0] m182_23;
   assign m182_23 =15'b0;

   // m182_24 = W*in
   wire signed [14:0] m182_24;
   assign m182_24 =15'b0;

   // m182_25 = W*in
   wire signed [14:0] m182_25;
   assign m182_25 =15'b0;

   // m182_26 = W*in
   wire signed [14:0] m182_26;
   assign m182_26 =15'b0;

   // m182_27 = W*in
   wire signed [14:0] m182_27;
   assign m182_27 ={ {4{in182[14]}} , in182[14:4] };

   // m182_28 = W*in
   wire signed [14:0] m182_28;
   assign m182_28 =15'b0;

   // m182_29 = W*in
   wire signed [14:0] m182_29;
   assign m182_29 =15'b0;

   // m182_30 = W*in
   wire signed [14:0] m182_30;
   assign m182_30 =15'b0;

   // m182_31 = W*in
   wire signed [14:0] m182_31;
   assign m182_31 =15'b0;

   // m182_32 = W*in
   wire signed [14:0] m182_32;
   assign m182_32 =15'b0;

   // m182_33 = W*in
   wire signed [14:0] m182_33;
   assign m182_33 =15'b0;

   // m182_34 = W*in
   wire signed [14:0] m182_34;
   assign m182_34 =15'b0;

   // m182_35 = W*in
   wire signed [14:0] m182_35;
   assign m182_35 =15'b0;

   // m182_36 = W*in
   wire signed [14:0] m182_36;
   assign m182_36 =15'b0;

   // m182_37 = W*in
   wire signed [14:0] m182_37;
   assign m182_37 =15'b0;

   // m182_38 = W*in
   wire signed [14:0] m182_38;
   assign m182_38 =15'b0;

   // m182_39 = W*in
   wire signed [14:0] m182_39;
   assign m182_39 =15'b0;

   // m182_40 = W*in
   wire signed [14:0] m182_40;
   assign m182_40 =15'b0;

   // m182_41 = W*in
   wire signed [14:0] m182_41;
   assign m182_41 =15'b0;

   // m182_42 = W*in
   wire signed [14:0] m182_42;
   assign m182_42 =15'b0;

   // m182_43 = W*in
   wire signed [14:0] m182_43;
   assign m182_43 =15'b0;

   // m182_44 = W*in
   wire signed [14:0] m182_44;
   assign m182_44 =15'b0;

   // m182_45 = W*in
   wire signed [14:0] m182_45;
   assign m182_45 ={ {3{neg182[14]}} , neg182[14:3] };

   // m182_46 = W*in
   wire signed [14:0] m182_46;
   assign m182_46 =15'b0;

   // m182_47 = W*in
   wire signed [14:0] m182_47;
   assign m182_47 =15'b0;

   // m182_48 = W*in
   wire signed [14:0] m182_48;
   assign m182_48 =15'b0;

   // m182_49 = W*in
   wire signed [14:0] m182_49;
   assign m182_49 =15'b0;

   // m182_50 = W*in
   wire signed [14:0] m182_50;
   assign m182_50 =15'b0;

   // m182_51 = W*in
   wire signed [14:0] m182_51;
   assign m182_51 =15'b0;

   // m182_52 = W*in
   wire signed [14:0] m182_52;
   assign m182_52 =15'b0;

   // m182_53 = W*in
   wire signed [14:0] m182_53;
   assign m182_53 =15'b0;

   // m182_54 = W*in
   wire signed [14:0] m182_54;
   assign m182_54 =15'b0;

   // m182_55 = W*in
   wire signed [14:0] m182_55;
   assign m182_55 =15'b0;

   // m182_56 = W*in
   wire signed [14:0] m182_56;
   assign m182_56 =15'b0;

   // m182_57 = W*in
   wire signed [14:0] m182_57;
   assign m182_57 =15'b0;

   // m182_58 = W*in
   wire signed [14:0] m182_58;
   assign m182_58 =15'b0;

   // m182_59 = W*in
   wire signed [14:0] m182_59;
   assign m182_59 =15'b0;

   // m182_60 = W*in
   wire signed [14:0] m182_60;
   assign m182_60 =15'b0;

   // m182_61 = W*in
   wire signed [14:0] m182_61;
   assign m182_61 =15'b0;

   // m182_62 = W*in
   wire signed [14:0] m182_62;
   assign m182_62 =15'b0;

   // m182_63 = W*in
   wire signed [14:0] m182_63;
   assign m182_63 =15'b0;

   // m182_64 = W*in
   wire signed [14:0] m182_64;
   assign m182_64 =15'b0;

   // m182_65 = W*in
   wire signed [14:0] m182_65;
   assign m182_65 =15'b0;

   // m182_66 = W*in
   wire signed [14:0] m182_66;
   assign m182_66 =15'b0;

   // m182_67 = W*in
   wire signed [14:0] m182_67;
   assign m182_67 =15'b0;

   // m182_68 = W*in
   wire signed [14:0] m182_68;
   assign m182_68 =15'b0;

   // m182_69 = W*in
   wire signed [14:0] m182_69;
   assign m182_69 =15'b0;

   // m182_70 = W*in
   wire signed [14:0] m182_70;
   assign m182_70 =15'b0;

   // m182_71 = W*in
   wire signed [14:0] m182_71;
   assign m182_71 =15'b0;

   // m182_72 = W*in
   wire signed [14:0] m182_72;
   assign m182_72 =15'b0;

   // m182_73 = W*in
   wire signed [14:0] m182_73;
   assign m182_73 =15'b0;

   // m182_74 = W*in
   wire signed [14:0] m182_74;
   assign m182_74 ={ {3{in182[14]}} , in182[14:3] };

   // m182_75 = W*in
   wire signed [14:0] m182_75;
   assign m182_75 ={ {3{in182[14]}} , in182[14:3] };

   // m182_76 = W*in
   wire signed [14:0] m182_76;
   assign m182_76 ={ {4{neg182[14]}} , neg182[14:4] };

   // m182_77 = W*in
   wire signed [14:0] m182_77;
   assign m182_77 =15'b0;

   // m182_78 = W*in
   wire signed [14:0] m182_78;
   assign m182_78 =15'b0;

   // m182_79 = W*in
   wire signed [14:0] m182_79;
   assign m182_79 =15'b0;

   // m182_80 = W*in
   wire signed [14:0] m182_80;
   assign m182_80 ={ {4{neg182[14]}} , neg182[14:4] };

   // m182_81 = W*in
   wire signed [14:0] m182_81;
   assign m182_81 =15'b0;

   // m182_82 = W*in
   wire signed [14:0] m182_82;
   assign m182_82 =15'b0;

   // m182_83 = W*in
   wire signed [14:0] m182_83;
   assign m182_83 =15'b0;

   // m182_84 = W*in
   wire signed [14:0] m182_84;
   assign m182_84 =15'b0;

   // m182_85 = W*in
   wire signed [14:0] m182_85;
   assign m182_85 =15'b0;

   // m182_86 = W*in
   wire signed [14:0] m182_86;
   assign m182_86 =15'b0;

   // m182_87 = W*in
   wire signed [14:0] m182_87;
   assign m182_87 =15'b0;

   // m182_88 = W*in
   wire signed [14:0] m182_88;
   assign m182_88 =15'b0;

   // m182_89 = W*in
   wire signed [14:0] m182_89;
   assign m182_89 ={ {4{neg182[14]}} , neg182[14:4] };

   // m182_90 = W*in
   wire signed [14:0] m182_90;
   assign m182_90 =15'b0;

   // m182_91 = W*in
   wire signed [14:0] m182_91;
   assign m182_91 =15'b0;

   // m182_92 = W*in
   wire signed [14:0] m182_92;
   assign m182_92 =15'b0;

   // m182_93 = W*in
   wire signed [14:0] m182_93;
   assign m182_93 =15'b0;

   // m182_94 = W*in
   wire signed [14:0] m182_94;
   assign m182_94 =15'b0;

   // m182_95 = W*in
   wire signed [14:0] m182_95;
   assign m182_95 =15'b0;

   // m182_96 = W*in
   wire signed [14:0] m182_96;
   assign m182_96 =15'b0;

   // m182_97 = W*in
   wire signed [14:0] m182_97;
   assign m182_97 =15'b0;

   // m182_98 = W*in
   wire signed [14:0] m182_98;
   assign m182_98 =15'b0;

   // m182_99 = W*in
   wire signed [14:0] m182_99;
   assign m182_99 =15'b0;

   // m182_100 = W*in
   wire signed [14:0] m182_100;
   assign m182_100 =15'b0;

   // m183_1 = W*in
   wire signed [14:0] m183_1;
   assign m183_1 =15'b0;

   // m183_2 = W*in
   wire signed [14:0] m183_2;
   assign m183_2 =15'b0;

   // m183_3 = W*in
   wire signed [14:0] m183_3;
   assign m183_3 =15'b0;

   // m183_4 = W*in
   wire signed [14:0] m183_4;
   assign m183_4 =15'b0;

   // m183_5 = W*in
   wire signed [14:0] m183_5;
   assign m183_5 =15'b0;

   // m183_6 = W*in
   wire signed [14:0] m183_6;
   assign m183_6 =15'b0;

   // m183_7 = W*in
   wire signed [14:0] m183_7;
   assign m183_7 =15'b0;

   // m183_8 = W*in
   wire signed [14:0] m183_8;
   assign m183_8 =15'b0;

   // m183_9 = W*in
   wire signed [14:0] m183_9;
   assign m183_9 ={ {4{neg183[14]}} , neg183[14:4] };

   // m183_10 = W*in
   wire signed [14:0] m183_10;
   assign m183_10 =15'b0;

   // m183_11 = W*in
   wire signed [14:0] m183_11;
   assign m183_11 =15'b0;

   // m183_12 = W*in
   wire signed [14:0] m183_12;
   assign m183_12 =15'b0;

   // m183_13 = W*in
   wire signed [14:0] m183_13;
   assign m183_13 =15'b0;

   // m183_14 = W*in
   wire signed [14:0] m183_14;
   assign m183_14 ={ {3{neg183[14]}} , neg183[14:3] };

   // m183_15 = W*in
   wire signed [14:0] m183_15;
   assign m183_15 =15'b0;

   // m183_16 = W*in
   wire signed [14:0] m183_16;
   assign m183_16 ={ {3{neg183[14]}} , neg183[14:3] };

   // m183_17 = W*in
   wire signed [14:0] m183_17;
   assign m183_17 =15'b0;

   // m183_18 = W*in
   wire signed [14:0] m183_18;
   assign m183_18 =15'b0;

   // m183_19 = W*in
   wire signed [14:0] m183_19;
   assign m183_19 =15'b0;

   // m183_20 = W*in
   wire signed [14:0] m183_20;
   assign m183_20 =15'b0;

   // m183_21 = W*in
   wire signed [14:0] m183_21;
   assign m183_21 =15'b0;

   // m183_22 = W*in
   wire signed [14:0] m183_22;
   assign m183_22 =15'b0;

   // m183_23 = W*in
   wire signed [14:0] m183_23;
   assign m183_23 =15'b0;

   // m183_24 = W*in
   wire signed [14:0] m183_24;
   assign m183_24 ={ {3{in183[14]}} , in183[14:3] };

   // m183_25 = W*in
   wire signed [14:0] m183_25;
   assign m183_25 ={ {4{in183[14]}} , in183[14:4] };

   // m183_26 = W*in
   wire signed [14:0] m183_26;
   assign m183_26 =15'b0;

   // m183_27 = W*in
   wire signed [14:0] m183_27;
   assign m183_27 =15'b0;

   // m183_28 = W*in
   wire signed [14:0] m183_28;
   assign m183_28 =15'b0;

   // m183_29 = W*in
   wire signed [14:0] m183_29;
   assign m183_29 ={ {4{neg183[14]}} , neg183[14:4] };

   // m183_30 = W*in
   wire signed [14:0] m183_30;
   assign m183_30 =15'b0;

   // m183_31 = W*in
   wire signed [14:0] m183_31;
   assign m183_31 =15'b0;

   // m183_32 = W*in
   wire signed [14:0] m183_32;
   assign m183_32 =15'b0;

   // m183_33 = W*in
   wire signed [14:0] m183_33;
   assign m183_33 =15'b0;

   // m183_34 = W*in
   wire signed [14:0] m183_34;
   assign m183_34 =15'b0;

   // m183_35 = W*in
   wire signed [14:0] m183_35;
   assign m183_35 ={ {3{neg183[14]}} , neg183[14:3] };

   // m183_36 = W*in
   wire signed [14:0] m183_36;
   assign m183_36 ={ {3{in183[14]}} , in183[14:3] };

   // m183_37 = W*in
   wire signed [14:0] m183_37;
   assign m183_37 =15'b0;

   // m183_38 = W*in
   wire signed [14:0] m183_38;
   assign m183_38 =15'b0;

   // m183_39 = W*in
   wire signed [14:0] m183_39;
   assign m183_39 =15'b0;

   // m183_40 = W*in
   wire signed [14:0] m183_40;
   assign m183_40 =15'b0;

   // m183_41 = W*in
   wire signed [14:0] m183_41;
   assign m183_41 =15'b0;

   // m183_42 = W*in
   wire signed [14:0] m183_42;
   assign m183_42 ={ {3{neg183[14]}} , neg183[14:3] };

   // m183_43 = W*in
   wire signed [14:0] m183_43;
   assign m183_43 ={ {3{in183[14]}} , in183[14:3] };

   // m183_44 = W*in
   wire signed [14:0] m183_44;
   assign m183_44 =15'b0;

   // m183_45 = W*in
   wire signed [14:0] m183_45;
   assign m183_45 =15'b0;

   // m183_46 = W*in
   wire signed [14:0] m183_46;
   assign m183_46 =15'b0;

   // m183_47 = W*in
   wire signed [14:0] m183_47;
   assign m183_47 =15'b0;

   // m183_48 = W*in
   wire signed [14:0] m183_48;
   assign m183_48 =15'b0;

   // m183_49 = W*in
   wire signed [14:0] m183_49;
   assign m183_49 =15'b0;

   // m183_50 = W*in
   wire signed [14:0] m183_50;
   assign m183_50 ={ {3{in183[14]}} , in183[14:3] };

   // m183_51 = W*in
   wire signed [14:0] m183_51;
   assign m183_51 =15'b0;

   // m183_52 = W*in
   wire signed [14:0] m183_52;
   assign m183_52 =15'b0;

   // m183_53 = W*in
   wire signed [14:0] m183_53;
   assign m183_53 =15'b0;

   // m183_54 = W*in
   wire signed [14:0] m183_54;
   assign m183_54 =15'b0;

   // m183_55 = W*in
   wire signed [14:0] m183_55;
   assign m183_55 =15'b0;

   // m183_56 = W*in
   wire signed [14:0] m183_56;
   assign m183_56 =15'b0;

   // m183_57 = W*in
   wire signed [14:0] m183_57;
   assign m183_57 =15'b0;

   // m183_58 = W*in
   wire signed [14:0] m183_58;
   assign m183_58 =15'b0;

   // m183_59 = W*in
   wire signed [14:0] m183_59;
   assign m183_59 =15'b0;

   // m183_60 = W*in
   wire signed [14:0] m183_60;
   assign m183_60 =15'b0;

   // m183_61 = W*in
   wire signed [14:0] m183_61;
   assign m183_61 =15'b0;

   // m183_62 = W*in
   wire signed [14:0] m183_62;
   assign m183_62 ={ {4{neg183[14]}} , neg183[14:4] };

   // m183_63 = W*in
   wire signed [14:0] m183_63;
   assign m183_63 =15'b0;

   // m183_64 = W*in
   wire signed [14:0] m183_64;
   assign m183_64 =15'b0;

   // m183_65 = W*in
   wire signed [14:0] m183_65;
   assign m183_65 =15'b0;

   // m183_66 = W*in
   wire signed [14:0] m183_66;
   assign m183_66 =15'b0;

   // m183_67 = W*in
   wire signed [14:0] m183_67;
   assign m183_67 =15'b0;

   // m183_68 = W*in
   wire signed [14:0] m183_68;
   assign m183_68 ={ {3{neg183[14]}} , neg183[14:3] };

   // m183_69 = W*in
   wire signed [14:0] m183_69;
   assign m183_69 ={ {3{in183[14]}} , in183[14:3] };

   // m183_70 = W*in
   wire signed [14:0] m183_70;
   assign m183_70 =15'b0;

   // m183_71 = W*in
   wire signed [14:0] m183_71;
   assign m183_71 =15'b0;

   // m183_72 = W*in
   wire signed [14:0] m183_72;
   assign m183_72 =15'b0;

   // m183_73 = W*in
   wire signed [14:0] m183_73;
   assign m183_73 =15'b0;

   // m183_74 = W*in
   wire signed [14:0] m183_74;
   assign m183_74 ={ {4{neg183[14]}} , neg183[14:4] };

   // m183_75 = W*in
   wire signed [14:0] m183_75;
   assign m183_75 =15'b0;

   // m183_76 = W*in
   wire signed [14:0] m183_76;
   assign m183_76 ={ {4{neg183[14]}} , neg183[14:4] };

   // m183_77 = W*in
   wire signed [14:0] m183_77;
   assign m183_77 ={ {2{in183[14]}} , in183[14:2] };

   // m183_78 = W*in
   wire signed [14:0] m183_78;
   assign m183_78 =15'b0;

   // m183_79 = W*in
   wire signed [14:0] m183_79;
   assign m183_79 ={ {3{in183[14]}} , in183[14:3] };

   // m183_80 = W*in
   wire signed [14:0] m183_80;
   assign m183_80 =15'b0;

   // m183_81 = W*in
   wire signed [14:0] m183_81;
   assign m183_81 =15'b0;

   // m183_82 = W*in
   wire signed [14:0] m183_82;
   assign m183_82 =15'b0;

   // m183_83 = W*in
   wire signed [14:0] m183_83;
   assign m183_83 =15'b0;

   // m183_84 = W*in
   wire signed [14:0] m183_84;
   assign m183_84 =15'b0;

   // m183_85 = W*in
   wire signed [14:0] m183_85;
   assign m183_85 =15'b0;

   // m183_86 = W*in
   wire signed [14:0] m183_86;
   assign m183_86 =15'b0;

   // m183_87 = W*in
   wire signed [14:0] m183_87;
   assign m183_87 =15'b0;

   // m183_88 = W*in
   wire signed [14:0] m183_88;
   assign m183_88 =15'b0;

   // m183_89 = W*in
   wire signed [14:0] m183_89;
   assign m183_89 =15'b0;

   // m183_90 = W*in
   wire signed [14:0] m183_90;
   assign m183_90 =15'b0;

   // m183_91 = W*in
   wire signed [14:0] m183_91;
   assign m183_91 =15'b0;

   // m183_92 = W*in
   wire signed [14:0] m183_92;
   assign m183_92 =15'b0;

   // m183_93 = W*in
   wire signed [14:0] m183_93;
   assign m183_93 =15'b0;

   // m183_94 = W*in
   wire signed [14:0] m183_94;
   assign m183_94 ={ {4{neg183[14]}} , neg183[14:4] };

   // m183_95 = W*in
   wire signed [14:0] m183_95;
   assign m183_95 =15'b0;

   // m183_96 = W*in
   wire signed [14:0] m183_96;
   assign m183_96 =15'b0;

   // m183_97 = W*in
   wire signed [14:0] m183_97;
   assign m183_97 =15'b0;

   // m183_98 = W*in
   wire signed [14:0] m183_98;
   assign m183_98 =15'b0;

   // m183_99 = W*in
   wire signed [14:0] m183_99;
   assign m183_99 =15'b0;

   // m183_100 = W*in
   wire signed [14:0] m183_100;
   assign m183_100 =15'b0;

   // m184_1 = W*in
   wire signed [14:0] m184_1;
   assign m184_1 =15'b0;

   // m184_2 = W*in
   wire signed [14:0] m184_2;
   assign m184_2 ={ {3{in184[14]}} , in184[14:3] };

   // m184_3 = W*in
   wire signed [14:0] m184_3;
   assign m184_3 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_4 = W*in
   wire signed [14:0] m184_4;
   assign m184_4 =15'b0;

   // m184_5 = W*in
   wire signed [14:0] m184_5;
   assign m184_5 =15'b0;

   // m184_6 = W*in
   wire signed [14:0] m184_6;
   assign m184_6 =15'b0;

   // m184_7 = W*in
   wire signed [14:0] m184_7;
   assign m184_7 =15'b0;

   // m184_8 = W*in
   wire signed [14:0] m184_8;
   assign m184_8 ={ {3{in184[14]}} , in184[14:3] };

   // m184_9 = W*in
   wire signed [14:0] m184_9;
   assign m184_9 =15'b0;

   // m184_10 = W*in
   wire signed [14:0] m184_10;
   assign m184_10 =15'b0;

   // m184_11 = W*in
   wire signed [14:0] m184_11;
   assign m184_11 =15'b0;

   // m184_12 = W*in
   wire signed [14:0] m184_12;
   assign m184_12 =15'b0;

   // m184_13 = W*in
   wire signed [14:0] m184_13;
   assign m184_13 ={ {3{in184[14]}} , in184[14:3] };

   // m184_14 = W*in
   wire signed [14:0] m184_14;
   assign m184_14 =15'b0;

   // m184_15 = W*in
   wire signed [14:0] m184_15;
   assign m184_15 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_16 = W*in
   wire signed [14:0] m184_16;
   assign m184_16 =15'b0;

   // m184_17 = W*in
   wire signed [14:0] m184_17;
   assign m184_17 =15'b0;

   // m184_18 = W*in
   wire signed [14:0] m184_18;
   assign m184_18 ={ {3{in184[14]}} , in184[14:3] };

   // m184_19 = W*in
   wire signed [14:0] m184_19;
   assign m184_19 ={ {3{in184[14]}} , in184[14:3] };

   // m184_20 = W*in
   wire signed [14:0] m184_20;
   assign m184_20 =15'b0;

   // m184_21 = W*in
   wire signed [14:0] m184_21;
   assign m184_21 =15'b0;

   // m184_22 = W*in
   wire signed [14:0] m184_22;
   assign m184_22 =15'b0;

   // m184_23 = W*in
   wire signed [14:0] m184_23;
   assign m184_23 =15'b0;

   // m184_24 = W*in
   wire signed [14:0] m184_24;
   assign m184_24 =15'b0;

   // m184_25 = W*in
   wire signed [14:0] m184_25;
   assign m184_25 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_26 = W*in
   wire signed [14:0] m184_26;
   assign m184_26 ={ {4{in184[14]}} , in184[14:4] };

   // m184_27 = W*in
   wire signed [14:0] m184_27;
   assign m184_27 ={ {3{in184[14]}} , in184[14:3] };

   // m184_28 = W*in
   wire signed [14:0] m184_28;
   assign m184_28 ={ {3{in184[14]}} , in184[14:3] };

   // m184_29 = W*in
   wire signed [14:0] m184_29;
   assign m184_29 ={ {3{in184[14]}} , in184[14:3] };

   // m184_30 = W*in
   wire signed [14:0] m184_30;
   assign m184_30 =15'b0;

   // m184_31 = W*in
   wire signed [14:0] m184_31;
   assign m184_31 ={ {3{in184[14]}} , in184[14:3] };

   // m184_32 = W*in
   wire signed [14:0] m184_32;
   assign m184_32 =15'b0;

   // m184_33 = W*in
   wire signed [14:0] m184_33;
   assign m184_33 ={ {4{in184[14]}} , in184[14:4] };

   // m184_34 = W*in
   wire signed [14:0] m184_34;
   assign m184_34 =15'b0;

   // m184_35 = W*in
   wire signed [14:0] m184_35;
   assign m184_35 =15'b0;

   // m184_36 = W*in
   wire signed [14:0] m184_36;
   assign m184_36 =15'b0;

   // m184_37 = W*in
   wire signed [14:0] m184_37;
   assign m184_37 =15'b0;

   // m184_38 = W*in
   wire signed [14:0] m184_38;
   assign m184_38 =15'b0;

   // m184_39 = W*in
   wire signed [14:0] m184_39;
   assign m184_39 =15'b0;

   // m184_40 = W*in
   wire signed [14:0] m184_40;
   assign m184_40 =15'b0;

   // m184_41 = W*in
   wire signed [14:0] m184_41;
   assign m184_41 =15'b0;

   // m184_42 = W*in
   wire signed [14:0] m184_42;
   assign m184_42 =15'b0;

   // m184_43 = W*in
   wire signed [14:0] m184_43;
   assign m184_43 =15'b0;

   // m184_44 = W*in
   wire signed [14:0] m184_44;
   assign m184_44 =15'b0;

   // m184_45 = W*in
   wire signed [14:0] m184_45;
   assign m184_45 =15'b0;

   // m184_46 = W*in
   wire signed [14:0] m184_46;
   assign m184_46 =15'b0;

   // m184_47 = W*in
   wire signed [14:0] m184_47;
   assign m184_47 =15'b0;

   // m184_48 = W*in
   wire signed [14:0] m184_48;
   assign m184_48 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_49 = W*in
   wire signed [14:0] m184_49;
   assign m184_49 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_50 = W*in
   wire signed [14:0] m184_50;
   assign m184_50 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_51 = W*in
   wire signed [14:0] m184_51;
   assign m184_51 =15'b0;

   // m184_52 = W*in
   wire signed [14:0] m184_52;
   assign m184_52 =15'b0;

   // m184_53 = W*in
   wire signed [14:0] m184_53;
   assign m184_53 =15'b0;

   // m184_54 = W*in
   wire signed [14:0] m184_54;
   assign m184_54 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_55 = W*in
   wire signed [14:0] m184_55;
   assign m184_55 =15'b0;

   // m184_56 = W*in
   wire signed [14:0] m184_56;
   assign m184_56 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_57 = W*in
   wire signed [14:0] m184_57;
   assign m184_57 =15'b0;

   // m184_58 = W*in
   wire signed [14:0] m184_58;
   assign m184_58 ={ {4{neg184[14]}} , neg184[14:4] };

   // m184_59 = W*in
   wire signed [14:0] m184_59;
   assign m184_59 =15'b0;

   // m184_60 = W*in
   wire signed [14:0] m184_60;
   assign m184_60 ={ {4{neg184[14]}} , neg184[14:4] };

   // m184_61 = W*in
   wire signed [14:0] m184_61;
   assign m184_61 =15'b0;

   // m184_62 = W*in
   wire signed [14:0] m184_62;
   assign m184_62 =15'b0;

   // m184_63 = W*in
   wire signed [14:0] m184_63;
   assign m184_63 =15'b0;

   // m184_64 = W*in
   wire signed [14:0] m184_64;
   assign m184_64 =15'b0;

   // m184_65 = W*in
   wire signed [14:0] m184_65;
   assign m184_65 =15'b0;

   // m184_66 = W*in
   wire signed [14:0] m184_66;
   assign m184_66 ={ {4{neg184[14]}} , neg184[14:4] };

   // m184_67 = W*in
   wire signed [14:0] m184_67;
   assign m184_67 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_68 = W*in
   wire signed [14:0] m184_68;
   assign m184_68 ={ {4{in184[14]}} , in184[14:4] };

   // m184_69 = W*in
   wire signed [14:0] m184_69;
   assign m184_69 ={ {4{neg184[14]}} , neg184[14:4] };

   // m184_70 = W*in
   wire signed [14:0] m184_70;
   assign m184_70 =15'b0;

   // m184_71 = W*in
   wire signed [14:0] m184_71;
   assign m184_71 =15'b0;

   // m184_72 = W*in
   wire signed [14:0] m184_72;
   assign m184_72 =15'b0;

   // m184_73 = W*in
   wire signed [14:0] m184_73;
   assign m184_73 =15'b0;

   // m184_74 = W*in
   wire signed [14:0] m184_74;
   assign m184_74 =15'b0;

   // m184_75 = W*in
   wire signed [14:0] m184_75;
   assign m184_75 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_76 = W*in
   wire signed [14:0] m184_76;
   assign m184_76 =15'b0;

   // m184_77 = W*in
   wire signed [14:0] m184_77;
   assign m184_77 =15'b0;

   // m184_78 = W*in
   wire signed [14:0] m184_78;
   assign m184_78 =15'b0;

   // m184_79 = W*in
   wire signed [14:0] m184_79;
   assign m184_79 =15'b0;

   // m184_80 = W*in
   wire signed [14:0] m184_80;
   assign m184_80 =15'b0;

   // m184_81 = W*in
   wire signed [14:0] m184_81;
   assign m184_81 =15'b0;

   // m184_82 = W*in
   wire signed [14:0] m184_82;
   assign m184_82 =15'b0;

   // m184_83 = W*in
   wire signed [14:0] m184_83;
   assign m184_83 =15'b0;

   // m184_84 = W*in
   wire signed [14:0] m184_84;
   assign m184_84 =15'b0;

   // m184_85 = W*in
   wire signed [14:0] m184_85;
   assign m184_85 =15'b0;

   // m184_86 = W*in
   wire signed [14:0] m184_86;
   assign m184_86 =15'b0;

   // m184_87 = W*in
   wire signed [14:0] m184_87;
   assign m184_87 =15'b0;

   // m184_88 = W*in
   wire signed [14:0] m184_88;
   assign m184_88 =15'b0;

   // m184_89 = W*in
   wire signed [14:0] m184_89;
   assign m184_89 =15'b0;

   // m184_90 = W*in
   wire signed [14:0] m184_90;
   assign m184_90 ={ {3{in184[14]}} , in184[14:3] };

   // m184_91 = W*in
   wire signed [14:0] m184_91;
   assign m184_91 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_92 = W*in
   wire signed [14:0] m184_92;
   assign m184_92 =15'b0;

   // m184_93 = W*in
   wire signed [14:0] m184_93;
   assign m184_93 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_94 = W*in
   wire signed [14:0] m184_94;
   assign m184_94 ={ {4{in184[14]}} , in184[14:4] };

   // m184_95 = W*in
   wire signed [14:0] m184_95;
   assign m184_95 ={ {3{neg184[14]}} , neg184[14:3] };

   // m184_96 = W*in
   wire signed [14:0] m184_96;
   assign m184_96 =15'b0;

   // m184_97 = W*in
   wire signed [14:0] m184_97;
   assign m184_97 ={ {3{in184[14]}} , in184[14:3] };

   // m184_98 = W*in
   wire signed [14:0] m184_98;
   assign m184_98 =15'b0;

   // m184_99 = W*in
   wire signed [14:0] m184_99;
   assign m184_99 =15'b0;

   // m184_100 = W*in
   wire signed [14:0] m184_100;
   assign m184_100 =15'b0;

   // m185_1 = W*in
   wire signed [14:0] m185_1;
   assign m185_1 =15'b0;

   // m185_2 = W*in
   wire signed [14:0] m185_2;
   assign m185_2 =15'b0;

   // m185_3 = W*in
   wire signed [14:0] m185_3;
   assign m185_3 =15'b0;

   // m185_4 = W*in
   wire signed [14:0] m185_4;
   assign m185_4 =15'b0;

   // m185_5 = W*in
   wire signed [14:0] m185_5;
   assign m185_5 =15'b0;

   // m185_6 = W*in
   wire signed [14:0] m185_6;
   assign m185_6 =15'b0;

   // m185_7 = W*in
   wire signed [14:0] m185_7;
   assign m185_7 ={ {3{neg185[14]}} , neg185[14:3] };

   // m185_8 = W*in
   wire signed [14:0] m185_8;
   assign m185_8 =15'b0;

   // m185_9 = W*in
   wire signed [14:0] m185_9;
   assign m185_9 =15'b0;

   // m185_10 = W*in
   wire signed [14:0] m185_10;
   assign m185_10 =15'b0;

   // m185_11 = W*in
   wire signed [14:0] m185_11;
   assign m185_11 ={ {3{in185[14]}} , in185[14:3] };

   // m185_12 = W*in
   wire signed [14:0] m185_12;
   assign m185_12 =15'b0;

   // m185_13 = W*in
   wire signed [14:0] m185_13;
   assign m185_13 =15'b0;

   // m185_14 = W*in
   wire signed [14:0] m185_14;
   assign m185_14 =15'b0;

   // m185_15 = W*in
   wire signed [14:0] m185_15;
   assign m185_15 =15'b0;

   // m185_16 = W*in
   wire signed [14:0] m185_16;
   assign m185_16 =15'b0;

   // m185_17 = W*in
   wire signed [14:0] m185_17;
   assign m185_17 =15'b0;

   // m185_18 = W*in
   wire signed [14:0] m185_18;
   assign m185_18 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_19 = W*in
   wire signed [14:0] m185_19;
   assign m185_19 =15'b0;

   // m185_20 = W*in
   wire signed [14:0] m185_20;
   assign m185_20 =15'b0;

   // m185_21 = W*in
   wire signed [14:0] m185_21;
   assign m185_21 ={ {3{in185[14]}} , in185[14:3] };

   // m185_22 = W*in
   wire signed [14:0] m185_22;
   assign m185_22 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_23 = W*in
   wire signed [14:0] m185_23;
   assign m185_23 =15'b0;

   // m185_24 = W*in
   wire signed [14:0] m185_24;
   assign m185_24 =15'b0;

   // m185_25 = W*in
   wire signed [14:0] m185_25;
   assign m185_25 ={ {3{in185[14]}} , in185[14:3] };

   // m185_26 = W*in
   wire signed [14:0] m185_26;
   assign m185_26 =15'b0;

   // m185_27 = W*in
   wire signed [14:0] m185_27;
   assign m185_27 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_28 = W*in
   wire signed [14:0] m185_28;
   assign m185_28 ={ {3{neg185[14]}} , neg185[14:3] };

   // m185_29 = W*in
   wire signed [14:0] m185_29;
   assign m185_29 =15'b0;

   // m185_30 = W*in
   wire signed [14:0] m185_30;
   assign m185_30 =15'b0;

   // m185_31 = W*in
   wire signed [14:0] m185_31;
   assign m185_31 =15'b0;

   // m185_32 = W*in
   wire signed [14:0] m185_32;
   assign m185_32 ={ {4{in185[14]}} , in185[14:4] };

   // m185_33 = W*in
   wire signed [14:0] m185_33;
   assign m185_33 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_34 = W*in
   wire signed [14:0] m185_34;
   assign m185_34 =15'b0;

   // m185_35 = W*in
   wire signed [14:0] m185_35;
   assign m185_35 =15'b0;

   // m185_36 = W*in
   wire signed [14:0] m185_36;
   assign m185_36 =15'b0;

   // m185_37 = W*in
   wire signed [14:0] m185_37;
   assign m185_37 ={ {3{neg185[14]}} , neg185[14:3] };

   // m185_38 = W*in
   wire signed [14:0] m185_38;
   assign m185_38 =15'b0;

   // m185_39 = W*in
   wire signed [14:0] m185_39;
   assign m185_39 =15'b0;

   // m185_40 = W*in
   wire signed [14:0] m185_40;
   assign m185_40 ={ {3{neg185[14]}} , neg185[14:3] };

   // m185_41 = W*in
   wire signed [14:0] m185_41;
   assign m185_41 =15'b0;

   // m185_42 = W*in
   wire signed [14:0] m185_42;
   assign m185_42 =15'b0;

   // m185_43 = W*in
   wire signed [14:0] m185_43;
   assign m185_43 =15'b0;

   // m185_44 = W*in
   wire signed [14:0] m185_44;
   assign m185_44 =15'b0;

   // m185_45 = W*in
   wire signed [14:0] m185_45;
   assign m185_45 =15'b0;

   // m185_46 = W*in
   wire signed [14:0] m185_46;
   assign m185_46 =15'b0;

   // m185_47 = W*in
   wire signed [14:0] m185_47;
   assign m185_47 =15'b0;

   // m185_48 = W*in
   wire signed [14:0] m185_48;
   assign m185_48 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_49 = W*in
   wire signed [14:0] m185_49;
   assign m185_49 ={ {3{in185[14]}} , in185[14:3] };

   // m185_50 = W*in
   wire signed [14:0] m185_50;
   assign m185_50 ={ {3{in185[14]}} , in185[14:3] };

   // m185_51 = W*in
   wire signed [14:0] m185_51;
   assign m185_51 =15'b0;

   // m185_52 = W*in
   wire signed [14:0] m185_52;
   assign m185_52 =15'b0;

   // m185_53 = W*in
   wire signed [14:0] m185_53;
   assign m185_53 =15'b0;

   // m185_54 = W*in
   wire signed [14:0] m185_54;
   assign m185_54 =15'b0;

   // m185_55 = W*in
   wire signed [14:0] m185_55;
   assign m185_55 =15'b0;

   // m185_56 = W*in
   wire signed [14:0] m185_56;
   assign m185_56 =15'b0;

   // m185_57 = W*in
   wire signed [14:0] m185_57;
   assign m185_57 ={ {3{neg185[14]}} , neg185[14:3] };

   // m185_58 = W*in
   wire signed [14:0] m185_58;
   assign m185_58 =15'b0;

   // m185_59 = W*in
   wire signed [14:0] m185_59;
   assign m185_59 ={ {4{in185[14]}} , in185[14:4] };

   // m185_60 = W*in
   wire signed [14:0] m185_60;
   assign m185_60 =15'b0;

   // m185_61 = W*in
   wire signed [14:0] m185_61;
   assign m185_61 =15'b0;

   // m185_62 = W*in
   wire signed [14:0] m185_62;
   assign m185_62 =15'b0;

   // m185_63 = W*in
   wire signed [14:0] m185_63;
   assign m185_63 =15'b0;

   // m185_64 = W*in
   wire signed [14:0] m185_64;
   assign m185_64 =15'b0;

   // m185_65 = W*in
   wire signed [14:0] m185_65;
   assign m185_65 ={ {3{in185[14]}} , in185[14:3] };

   // m185_66 = W*in
   wire signed [14:0] m185_66;
   assign m185_66 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_67 = W*in
   wire signed [14:0] m185_67;
   assign m185_67 ={ {4{in185[14]}} , in185[14:4] };

   // m185_68 = W*in
   wire signed [14:0] m185_68;
   assign m185_68 =15'b0;

   // m185_69 = W*in
   wire signed [14:0] m185_69;
   assign m185_69 ={ {3{in185[14]}} , in185[14:3] };

   // m185_70 = W*in
   wire signed [14:0] m185_70;
   assign m185_70 =15'b0;

   // m185_71 = W*in
   wire signed [14:0] m185_71;
   assign m185_71 =15'b0;

   // m185_72 = W*in
   wire signed [14:0] m185_72;
   assign m185_72 =15'b0;

   // m185_73 = W*in
   wire signed [14:0] m185_73;
   assign m185_73 ={ {3{in185[14]}} , in185[14:3] };

   // m185_74 = W*in
   wire signed [14:0] m185_74;
   assign m185_74 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_75 = W*in
   wire signed [14:0] m185_75;
   assign m185_75 ={ {3{in185[14]}} , in185[14:3] };

   // m185_76 = W*in
   wire signed [14:0] m185_76;
   assign m185_76 =15'b0;

   // m185_77 = W*in
   wire signed [14:0] m185_77;
   assign m185_77 ={ {3{in185[14]}} , in185[14:3] };

   // m185_78 = W*in
   wire signed [14:0] m185_78;
   assign m185_78 =15'b0;

   // m185_79 = W*in
   wire signed [14:0] m185_79;
   assign m185_79 =15'b0;

   // m185_80 = W*in
   wire signed [14:0] m185_80;
   assign m185_80 =15'b0;

   // m185_81 = W*in
   wire signed [14:0] m185_81;
   assign m185_81 =15'b0;

   // m185_82 = W*in
   wire signed [14:0] m185_82;
   assign m185_82 =15'b0;

   // m185_83 = W*in
   wire signed [14:0] m185_83;
   assign m185_83 =15'b0;

   // m185_84 = W*in
   wire signed [14:0] m185_84;
   assign m185_84 =15'b0;

   // m185_85 = W*in
   wire signed [14:0] m185_85;
   assign m185_85 =15'b0;

   // m185_86 = W*in
   wire signed [14:0] m185_86;
   assign m185_86 ={ {3{in185[14]}} , in185[14:3] };

   // m185_87 = W*in
   wire signed [14:0] m185_87;
   assign m185_87 =15'b0;

   // m185_88 = W*in
   wire signed [14:0] m185_88;
   assign m185_88 =15'b0;

   // m185_89 = W*in
   wire signed [14:0] m185_89;
   assign m185_89 =15'b0;

   // m185_90 = W*in
   wire signed [14:0] m185_90;
   assign m185_90 =15'b0;

   // m185_91 = W*in
   wire signed [14:0] m185_91;
   assign m185_91 =15'b0;

   // m185_92 = W*in
   wire signed [14:0] m185_92;
   assign m185_92 =15'b0;

   // m185_93 = W*in
   wire signed [14:0] m185_93;
   assign m185_93 =15'b0;

   // m185_94 = W*in
   wire signed [14:0] m185_94;
   assign m185_94 ={ {4{neg185[14]}} , neg185[14:4] };

   // m185_95 = W*in
   wire signed [14:0] m185_95;
   assign m185_95 ={ {3{in185[14]}} , in185[14:3] };

   // m185_96 = W*in
   wire signed [14:0] m185_96;
   assign m185_96 =15'b0;

   // m185_97 = W*in
   wire signed [14:0] m185_97;
   assign m185_97 =15'b0;

   // m185_98 = W*in
   wire signed [14:0] m185_98;
   assign m185_98 =15'b0;

   // m185_99 = W*in
   wire signed [14:0] m185_99;
   assign m185_99 =15'b0;

   // m185_100 = W*in
   wire signed [14:0] m185_100;
   assign m185_100 =15'b0;

   // m186_1 = W*in
   wire signed [14:0] m186_1;
   assign m186_1 =15'b0;

   // m186_2 = W*in
   wire signed [14:0] m186_2;
   assign m186_2 =15'b0;

   // m186_3 = W*in
   wire signed [14:0] m186_3;
   assign m186_3 =15'b0;

   // m186_4 = W*in
   wire signed [14:0] m186_4;
   assign m186_4 ={ {4{in186[14]}} , in186[14:4] };

   // m186_5 = W*in
   wire signed [14:0] m186_5;
   assign m186_5 ={ {4{neg186[14]}} , neg186[14:4] };

   // m186_6 = W*in
   wire signed [14:0] m186_6;
   assign m186_6 ={ {3{in186[14]}} , in186[14:3] };

   // m186_7 = W*in
   wire signed [14:0] m186_7;
   assign m186_7 ={ {3{in186[14]}} , in186[14:3] };

   // m186_8 = W*in
   wire signed [14:0] m186_8;
   assign m186_8 ={ {3{in186[14]}} , in186[14:3] };

   // m186_9 = W*in
   wire signed [14:0] m186_9;
   assign m186_9 =15'b0;

   // m186_10 = W*in
   wire signed [14:0] m186_10;
   assign m186_10 =15'b0;

   // m186_11 = W*in
   wire signed [14:0] m186_11;
   assign m186_11 =15'b0;

   // m186_12 = W*in
   wire signed [14:0] m186_12;
   assign m186_12 =15'b0;

   // m186_13 = W*in
   wire signed [14:0] m186_13;
   assign m186_13 =15'b0;

   // m186_14 = W*in
   wire signed [14:0] m186_14;
   assign m186_14 =15'b0;

   // m186_15 = W*in
   wire signed [14:0] m186_15;
   assign m186_15 =15'b0;

   // m186_16 = W*in
   wire signed [14:0] m186_16;
   assign m186_16 =15'b0;

   // m186_17 = W*in
   wire signed [14:0] m186_17;
   assign m186_17 =15'b0;

   // m186_18 = W*in
   wire signed [14:0] m186_18;
   assign m186_18 ={ {3{in186[14]}} , in186[14:3] };

   // m186_19 = W*in
   wire signed [14:0] m186_19;
   assign m186_19 =15'b0;

   // m186_20 = W*in
   wire signed [14:0] m186_20;
   assign m186_20 =15'b0;

   // m186_21 = W*in
   wire signed [14:0] m186_21;
   assign m186_21 ={ {4{in186[14]}} , in186[14:4] };

   // m186_22 = W*in
   wire signed [14:0] m186_22;
   assign m186_22 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_23 = W*in
   wire signed [14:0] m186_23;
   assign m186_23 =15'b0;

   // m186_24 = W*in
   wire signed [14:0] m186_24;
   assign m186_24 =15'b0;

   // m186_25 = W*in
   wire signed [14:0] m186_25;
   assign m186_25 =15'b0;

   // m186_26 = W*in
   wire signed [14:0] m186_26;
   assign m186_26 =15'b0;

   // m186_27 = W*in
   wire signed [14:0] m186_27;
   assign m186_27 ={ {4{neg186[14]}} , neg186[14:4] };

   // m186_28 = W*in
   wire signed [14:0] m186_28;
   assign m186_28 =15'b0;

   // m186_29 = W*in
   wire signed [14:0] m186_29;
   assign m186_29 =15'b0;

   // m186_30 = W*in
   wire signed [14:0] m186_30;
   assign m186_30 =15'b0;

   // m186_31 = W*in
   wire signed [14:0] m186_31;
   assign m186_31 ={ {4{in186[14]}} , in186[14:4] };

   // m186_32 = W*in
   wire signed [14:0] m186_32;
   assign m186_32 =15'b0;

   // m186_33 = W*in
   wire signed [14:0] m186_33;
   assign m186_33 =15'b0;

   // m186_34 = W*in
   wire signed [14:0] m186_34;
   assign m186_34 =15'b0;

   // m186_35 = W*in
   wire signed [14:0] m186_35;
   assign m186_35 =15'b0;

   // m186_36 = W*in
   wire signed [14:0] m186_36;
   assign m186_36 =15'b0;

   // m186_37 = W*in
   wire signed [14:0] m186_37;
   assign m186_37 =15'b0;

   // m186_38 = W*in
   wire signed [14:0] m186_38;
   assign m186_38 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_39 = W*in
   wire signed [14:0] m186_39;
   assign m186_39 =15'b0;

   // m186_40 = W*in
   wire signed [14:0] m186_40;
   assign m186_40 =15'b0;

   // m186_41 = W*in
   wire signed [14:0] m186_41;
   assign m186_41 ={ {3{in186[14]}} , in186[14:3] };

   // m186_42 = W*in
   wire signed [14:0] m186_42;
   assign m186_42 =15'b0;

   // m186_43 = W*in
   wire signed [14:0] m186_43;
   assign m186_43 =15'b0;

   // m186_44 = W*in
   wire signed [14:0] m186_44;
   assign m186_44 =15'b0;

   // m186_45 = W*in
   wire signed [14:0] m186_45;
   assign m186_45 =15'b0;

   // m186_46 = W*in
   wire signed [14:0] m186_46;
   assign m186_46 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_47 = W*in
   wire signed [14:0] m186_47;
   assign m186_47 =15'b0;

   // m186_48 = W*in
   wire signed [14:0] m186_48;
   assign m186_48 ={ {3{in186[14]}} , in186[14:3] };

   // m186_49 = W*in
   wire signed [14:0] m186_49;
   assign m186_49 =15'b0;

   // m186_50 = W*in
   wire signed [14:0] m186_50;
   assign m186_50 =15'b0;

   // m186_51 = W*in
   wire signed [14:0] m186_51;
   assign m186_51 =15'b0;

   // m186_52 = W*in
   wire signed [14:0] m186_52;
   assign m186_52 ={ {3{in186[14]}} , in186[14:3] };

   // m186_53 = W*in
   wire signed [14:0] m186_53;
   assign m186_53 =15'b0;

   // m186_54 = W*in
   wire signed [14:0] m186_54;
   assign m186_54 =15'b0;

   // m186_55 = W*in
   wire signed [14:0] m186_55;
   assign m186_55 =15'b0;

   // m186_56 = W*in
   wire signed [14:0] m186_56;
   assign m186_56 =15'b0;

   // m186_57 = W*in
   wire signed [14:0] m186_57;
   assign m186_57 =15'b0;

   // m186_58 = W*in
   wire signed [14:0] m186_58;
   assign m186_58 ={ {4{neg186[14]}} , neg186[14:4] };

   // m186_59 = W*in
   wire signed [14:0] m186_59;
   assign m186_59 =15'b0;

   // m186_60 = W*in
   wire signed [14:0] m186_60;
   assign m186_60 ={ {4{in186[14]}} , in186[14:4] };

   // m186_61 = W*in
   wire signed [14:0] m186_61;
   assign m186_61 ={ {4{neg186[14]}} , neg186[14:4] };

   // m186_62 = W*in
   wire signed [14:0] m186_62;
   assign m186_62 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_63 = W*in
   wire signed [14:0] m186_63;
   assign m186_63 =15'b0;

   // m186_64 = W*in
   wire signed [14:0] m186_64;
   assign m186_64 ={ {4{neg186[14]}} , neg186[14:4] };

   // m186_65 = W*in
   wire signed [14:0] m186_65;
   assign m186_65 =15'b0;

   // m186_66 = W*in
   wire signed [14:0] m186_66;
   assign m186_66 =15'b0;

   // m186_67 = W*in
   wire signed [14:0] m186_67;
   assign m186_67 =15'b0;

   // m186_68 = W*in
   wire signed [14:0] m186_68;
   assign m186_68 ={ {3{in186[14]}} , in186[14:3] };

   // m186_69 = W*in
   wire signed [14:0] m186_69;
   assign m186_69 ={ {4{in186[14]}} , in186[14:4] };

   // m186_70 = W*in
   wire signed [14:0] m186_70;
   assign m186_70 ={ {4{in186[14]}} , in186[14:4] };

   // m186_71 = W*in
   wire signed [14:0] m186_71;
   assign m186_71 =15'b0;

   // m186_72 = W*in
   wire signed [14:0] m186_72;
   assign m186_72 =15'b0;

   // m186_73 = W*in
   wire signed [14:0] m186_73;
   assign m186_73 ={ {3{in186[14]}} , in186[14:3] };

   // m186_74 = W*in
   wire signed [14:0] m186_74;
   assign m186_74 =15'b0;

   // m186_75 = W*in
   wire signed [14:0] m186_75;
   assign m186_75 =15'b0;

   // m186_76 = W*in
   wire signed [14:0] m186_76;
   assign m186_76 ={ {4{neg186[14]}} , neg186[14:4] };

   // m186_77 = W*in
   wire signed [14:0] m186_77;
   assign m186_77 =15'b0;

   // m186_78 = W*in
   wire signed [14:0] m186_78;
   assign m186_78 ={ {3{in186[14]}} , in186[14:3] };

   // m186_79 = W*in
   wire signed [14:0] m186_79;
   assign m186_79 =15'b0;

   // m186_80 = W*in
   wire signed [14:0] m186_80;
   assign m186_80 =15'b0;

   // m186_81 = W*in
   wire signed [14:0] m186_81;
   assign m186_81 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_82 = W*in
   wire signed [14:0] m186_82;
   assign m186_82 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_83 = W*in
   wire signed [14:0] m186_83;
   assign m186_83 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_84 = W*in
   wire signed [14:0] m186_84;
   assign m186_84 =15'b0;

   // m186_85 = W*in
   wire signed [14:0] m186_85;
   assign m186_85 =15'b0;

   // m186_86 = W*in
   wire signed [14:0] m186_86;
   assign m186_86 =15'b0;

   // m186_87 = W*in
   wire signed [14:0] m186_87;
   assign m186_87 =15'b0;

   // m186_88 = W*in
   wire signed [14:0] m186_88;
   assign m186_88 ={ {3{in186[14]}} , in186[14:3] };

   // m186_89 = W*in
   wire signed [14:0] m186_89;
   assign m186_89 =15'b0;

   // m186_90 = W*in
   wire signed [14:0] m186_90;
   assign m186_90 =15'b0;

   // m186_91 = W*in
   wire signed [14:0] m186_91;
   assign m186_91 =15'b0;

   // m186_92 = W*in
   wire signed [14:0] m186_92;
   assign m186_92 =15'b0;

   // m186_93 = W*in
   wire signed [14:0] m186_93;
   assign m186_93 =15'b0;

   // m186_94 = W*in
   wire signed [14:0] m186_94;
   assign m186_94 ={ {3{neg186[14]}} , neg186[14:3] };

   // m186_95 = W*in
   wire signed [14:0] m186_95;
   assign m186_95 =15'b0;

   // m186_96 = W*in
   wire signed [14:0] m186_96;
   assign m186_96 ={ {3{in186[14]}} , in186[14:3] };

   // m186_97 = W*in
   wire signed [14:0] m186_97;
   assign m186_97 =15'b0;

   // m186_98 = W*in
   wire signed [14:0] m186_98;
   assign m186_98 ={ {3{in186[14]}} , in186[14:3] };

   // m186_99 = W*in
   wire signed [14:0] m186_99;
   assign m186_99 =15'b0;

   // m186_100 = W*in
   wire signed [14:0] m186_100;
   assign m186_100 =15'b0;

   // m187_1 = W*in
   wire signed [14:0] m187_1;
   assign m187_1 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_2 = W*in
   wire signed [14:0] m187_2;
   assign m187_2 =15'b0;

   // m187_3 = W*in
   wire signed [14:0] m187_3;
   assign m187_3 =15'b0;

   // m187_4 = W*in
   wire signed [14:0] m187_4;
   assign m187_4 =15'b0;

   // m187_5 = W*in
   wire signed [14:0] m187_5;
   assign m187_5 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_6 = W*in
   wire signed [14:0] m187_6;
   assign m187_6 ={ {3{in187[14]}} , in187[14:3] };

   // m187_7 = W*in
   wire signed [14:0] m187_7;
   assign m187_7 =15'b0;

   // m187_8 = W*in
   wire signed [14:0] m187_8;
   assign m187_8 =15'b0;

   // m187_9 = W*in
   wire signed [14:0] m187_9;
   assign m187_9 ={ {3{in187[14]}} , in187[14:3] };

   // m187_10 = W*in
   wire signed [14:0] m187_10;
   assign m187_10 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_11 = W*in
   wire signed [14:0] m187_11;
   assign m187_11 =15'b0;

   // m187_12 = W*in
   wire signed [14:0] m187_12;
   assign m187_12 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_13 = W*in
   wire signed [14:0] m187_13;
   assign m187_13 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_14 = W*in
   wire signed [14:0] m187_14;
   assign m187_14 =15'b0;

   // m187_15 = W*in
   wire signed [14:0] m187_15;
   assign m187_15 =15'b0;

   // m187_16 = W*in
   wire signed [14:0] m187_16;
   assign m187_16 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_17 = W*in
   wire signed [14:0] m187_17;
   assign m187_17 ={ {3{in187[14]}} , in187[14:3] };

   // m187_18 = W*in
   wire signed [14:0] m187_18;
   assign m187_18 =15'b0;

   // m187_19 = W*in
   wire signed [14:0] m187_19;
   assign m187_19 =15'b0;

   // m187_20 = W*in
   wire signed [14:0] m187_20;
   assign m187_20 =15'b0;

   // m187_21 = W*in
   wire signed [14:0] m187_21;
   assign m187_21 =15'b0;

   // m187_22 = W*in
   wire signed [14:0] m187_22;
   assign m187_22 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_23 = W*in
   wire signed [14:0] m187_23;
   assign m187_23 =15'b0;

   // m187_24 = W*in
   wire signed [14:0] m187_24;
   assign m187_24 =15'b0;

   // m187_25 = W*in
   wire signed [14:0] m187_25;
   assign m187_25 =15'b0;

   // m187_26 = W*in
   wire signed [14:0] m187_26;
   assign m187_26 =15'b0;

   // m187_27 = W*in
   wire signed [14:0] m187_27;
   assign m187_27 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_28 = W*in
   wire signed [14:0] m187_28;
   assign m187_28 =15'b0;

   // m187_29 = W*in
   wire signed [14:0] m187_29;
   assign m187_29 =15'b0;

   // m187_30 = W*in
   wire signed [14:0] m187_30;
   assign m187_30 =15'b0;

   // m187_31 = W*in
   wire signed [14:0] m187_31;
   assign m187_31 =15'b0;

   // m187_32 = W*in
   wire signed [14:0] m187_32;
   assign m187_32 =15'b0;

   // m187_33 = W*in
   wire signed [14:0] m187_33;
   assign m187_33 =15'b0;

   // m187_34 = W*in
   wire signed [14:0] m187_34;
   assign m187_34 =15'b0;

   // m187_35 = W*in
   wire signed [14:0] m187_35;
   assign m187_35 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_36 = W*in
   wire signed [14:0] m187_36;
   assign m187_36 =15'b0;

   // m187_37 = W*in
   wire signed [14:0] m187_37;
   assign m187_37 =15'b0;

   // m187_38 = W*in
   wire signed [14:0] m187_38;
   assign m187_38 =15'b0;

   // m187_39 = W*in
   wire signed [14:0] m187_39;
   assign m187_39 =15'b0;

   // m187_40 = W*in
   wire signed [14:0] m187_40;
   assign m187_40 =15'b0;

   // m187_41 = W*in
   wire signed [14:0] m187_41;
   assign m187_41 =15'b0;

   // m187_42 = W*in
   wire signed [14:0] m187_42;
   assign m187_42 =15'b0;

   // m187_43 = W*in
   wire signed [14:0] m187_43;
   assign m187_43 =15'b0;

   // m187_44 = W*in
   wire signed [14:0] m187_44;
   assign m187_44 =15'b0;

   // m187_45 = W*in
   wire signed [14:0] m187_45;
   assign m187_45 =15'b0;

   // m187_46 = W*in
   wire signed [14:0] m187_46;
   assign m187_46 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_47 = W*in
   wire signed [14:0] m187_47;
   assign m187_47 ={ {3{in187[14]}} , in187[14:3] };

   // m187_48 = W*in
   wire signed [14:0] m187_48;
   assign m187_48 =15'b0;

   // m187_49 = W*in
   wire signed [14:0] m187_49;
   assign m187_49 ={ {3{in187[14]}} , in187[14:3] };

   // m187_50 = W*in
   wire signed [14:0] m187_50;
   assign m187_50 =15'b0;

   // m187_51 = W*in
   wire signed [14:0] m187_51;
   assign m187_51 =15'b0;

   // m187_52 = W*in
   wire signed [14:0] m187_52;
   assign m187_52 ={ {3{in187[14]}} , in187[14:3] };

   // m187_53 = W*in
   wire signed [14:0] m187_53;
   assign m187_53 =15'b0;

   // m187_54 = W*in
   wire signed [14:0] m187_54;
   assign m187_54 =15'b0;

   // m187_55 = W*in
   wire signed [14:0] m187_55;
   assign m187_55 =15'b0;

   // m187_56 = W*in
   wire signed [14:0] m187_56;
   assign m187_56 =15'b0;

   // m187_57 = W*in
   wire signed [14:0] m187_57;
   assign m187_57 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_58 = W*in
   wire signed [14:0] m187_58;
   assign m187_58 =15'b0;

   // m187_59 = W*in
   wire signed [14:0] m187_59;
   assign m187_59 ={ {3{in187[14]}} , in187[14:3] };

   // m187_60 = W*in
   wire signed [14:0] m187_60;
   assign m187_60 =15'b0;

   // m187_61 = W*in
   wire signed [14:0] m187_61;
   assign m187_61 ={ {4{neg187[14]}} , neg187[14:4] };

   // m187_62 = W*in
   wire signed [14:0] m187_62;
   assign m187_62 =15'b0;

   // m187_63 = W*in
   wire signed [14:0] m187_63;
   assign m187_63 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_64 = W*in
   wire signed [14:0] m187_64;
   assign m187_64 =15'b0;

   // m187_65 = W*in
   wire signed [14:0] m187_65;
   assign m187_65 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_66 = W*in
   wire signed [14:0] m187_66;
   assign m187_66 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_67 = W*in
   wire signed [14:0] m187_67;
   assign m187_67 =15'b0;

   // m187_68 = W*in
   wire signed [14:0] m187_68;
   assign m187_68 ={ {2{neg187[14]}} , neg187[14:2] };

   // m187_69 = W*in
   wire signed [14:0] m187_69;
   assign m187_69 =15'b0;

   // m187_70 = W*in
   wire signed [14:0] m187_70;
   assign m187_70 ={ {3{in187[14]}} , in187[14:3] };

   // m187_71 = W*in
   wire signed [14:0] m187_71;
   assign m187_71 =15'b0;

   // m187_72 = W*in
   wire signed [14:0] m187_72;
   assign m187_72 =15'b0;

   // m187_73 = W*in
   wire signed [14:0] m187_73;
   assign m187_73 =15'b0;

   // m187_74 = W*in
   wire signed [14:0] m187_74;
   assign m187_74 =15'b0;

   // m187_75 = W*in
   wire signed [14:0] m187_75;
   assign m187_75 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_76 = W*in
   wire signed [14:0] m187_76;
   assign m187_76 =15'b0;

   // m187_77 = W*in
   wire signed [14:0] m187_77;
   assign m187_77 =15'b0;

   // m187_78 = W*in
   wire signed [14:0] m187_78;
   assign m187_78 =15'b0;

   // m187_79 = W*in
   wire signed [14:0] m187_79;
   assign m187_79 =15'b0;

   // m187_80 = W*in
   wire signed [14:0] m187_80;
   assign m187_80 =15'b0;

   // m187_81 = W*in
   wire signed [14:0] m187_81;
   assign m187_81 =15'b0;

   // m187_82 = W*in
   wire signed [14:0] m187_82;
   assign m187_82 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_83 = W*in
   wire signed [14:0] m187_83;
   assign m187_83 =15'b0;

   // m187_84 = W*in
   wire signed [14:0] m187_84;
   assign m187_84 =15'b0;

   // m187_85 = W*in
   wire signed [14:0] m187_85;
   assign m187_85 =15'b0;

   // m187_86 = W*in
   wire signed [14:0] m187_86;
   assign m187_86 =15'b0;

   // m187_87 = W*in
   wire signed [14:0] m187_87;
   assign m187_87 =15'b0;

   // m187_88 = W*in
   wire signed [14:0] m187_88;
   assign m187_88 =15'b0;

   // m187_89 = W*in
   wire signed [14:0] m187_89;
   assign m187_89 =15'b0;

   // m187_90 = W*in
   wire signed [14:0] m187_90;
   assign m187_90 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_91 = W*in
   wire signed [14:0] m187_91;
   assign m187_91 =15'b0;

   // m187_92 = W*in
   wire signed [14:0] m187_92;
   assign m187_92 ={ {3{neg187[14]}} , neg187[14:3] };

   // m187_93 = W*in
   wire signed [14:0] m187_93;
   assign m187_93 =15'b0;

   // m187_94 = W*in
   wire signed [14:0] m187_94;
   assign m187_94 ={ {4{neg187[14]}} , neg187[14:4] };

   // m187_95 = W*in
   wire signed [14:0] m187_95;
   assign m187_95 ={ {3{in187[14]}} , in187[14:3] };

   // m187_96 = W*in
   wire signed [14:0] m187_96;
   assign m187_96 =15'b0;

   // m187_97 = W*in
   wire signed [14:0] m187_97;
   assign m187_97 ={ {2{neg187[14]}} , neg187[14:2] };

   // m187_98 = W*in
   wire signed [14:0] m187_98;
   assign m187_98 ={ {3{in187[14]}} , in187[14:3] };

   // m187_99 = W*in
   wire signed [14:0] m187_99;
   assign m187_99 =15'b0;

   // m187_100 = W*in
   wire signed [14:0] m187_100;
   assign m187_100 =15'b0;

   // m188_1 = W*in
   wire signed [14:0] m188_1;
   assign m188_1 =15'b0;

   // m188_2 = W*in
   wire signed [14:0] m188_2;
   assign m188_2 =15'b0;

   // m188_3 = W*in
   wire signed [14:0] m188_3;
   assign m188_3 =15'b0;

   // m188_4 = W*in
   wire signed [14:0] m188_4;
   assign m188_4 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_5 = W*in
   wire signed [14:0] m188_5;
   assign m188_5 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_6 = W*in
   wire signed [14:0] m188_6;
   assign m188_6 ={ {3{in188[14]}} , in188[14:3] };

   // m188_7 = W*in
   wire signed [14:0] m188_7;
   assign m188_7 =15'b0;

   // m188_8 = W*in
   wire signed [14:0] m188_8;
   assign m188_8 ={ {3{in188[14]}} , in188[14:3] };

   // m188_9 = W*in
   wire signed [14:0] m188_9;
   assign m188_9 =15'b0;

   // m188_10 = W*in
   wire signed [14:0] m188_10;
   assign m188_10 =15'b0;

   // m188_11 = W*in
   wire signed [14:0] m188_11;
   assign m188_11 =15'b0;

   // m188_12 = W*in
   wire signed [14:0] m188_12;
   assign m188_12 ={ {3{in188[14]}} , in188[14:3] };

   // m188_13 = W*in
   wire signed [14:0] m188_13;
   assign m188_13 =15'b0;

   // m188_14 = W*in
   wire signed [14:0] m188_14;
   assign m188_14 =15'b0;

   // m188_15 = W*in
   wire signed [14:0] m188_15;
   assign m188_15 =15'b0;

   // m188_16 = W*in
   wire signed [14:0] m188_16;
   assign m188_16 =15'b0;

   // m188_17 = W*in
   wire signed [14:0] m188_17;
   assign m188_17 =15'b0;

   // m188_18 = W*in
   wire signed [14:0] m188_18;
   assign m188_18 =15'b0;

   // m188_19 = W*in
   wire signed [14:0] m188_19;
   assign m188_19 ={ {4{neg188[14]}} , neg188[14:4] };

   // m188_20 = W*in
   wire signed [14:0] m188_20;
   assign m188_20 =15'b0;

   // m188_21 = W*in
   wire signed [14:0] m188_21;
   assign m188_21 =15'b0;

   // m188_22 = W*in
   wire signed [14:0] m188_22;
   assign m188_22 =15'b0;

   // m188_23 = W*in
   wire signed [14:0] m188_23;
   assign m188_23 =15'b0;

   // m188_24 = W*in
   wire signed [14:0] m188_24;
   assign m188_24 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_25 = W*in
   wire signed [14:0] m188_25;
   assign m188_25 =15'b0;

   // m188_26 = W*in
   wire signed [14:0] m188_26;
   assign m188_26 =15'b0;

   // m188_27 = W*in
   wire signed [14:0] m188_27;
   assign m188_27 =15'b0;

   // m188_28 = W*in
   wire signed [14:0] m188_28;
   assign m188_28 ={ {4{neg188[14]}} , neg188[14:4] };

   // m188_29 = W*in
   wire signed [14:0] m188_29;
   assign m188_29 ={ {3{in188[14]}} , in188[14:3] };

   // m188_30 = W*in
   wire signed [14:0] m188_30;
   assign m188_30 =15'b0;

   // m188_31 = W*in
   wire signed [14:0] m188_31;
   assign m188_31 =15'b0;

   // m188_32 = W*in
   wire signed [14:0] m188_32;
   assign m188_32 ={ {3{in188[14]}} , in188[14:3] };

   // m188_33 = W*in
   wire signed [14:0] m188_33;
   assign m188_33 =15'b0;

   // m188_34 = W*in
   wire signed [14:0] m188_34;
   assign m188_34 ={ {3{in188[14]}} , in188[14:3] };

   // m188_35 = W*in
   wire signed [14:0] m188_35;
   assign m188_35 =15'b0;

   // m188_36 = W*in
   wire signed [14:0] m188_36;
   assign m188_36 =15'b0;

   // m188_37 = W*in
   wire signed [14:0] m188_37;
   assign m188_37 =15'b0;

   // m188_38 = W*in
   wire signed [14:0] m188_38;
   assign m188_38 =15'b0;

   // m188_39 = W*in
   wire signed [14:0] m188_39;
   assign m188_39 =15'b0;

   // m188_40 = W*in
   wire signed [14:0] m188_40;
   assign m188_40 =15'b0;

   // m188_41 = W*in
   wire signed [14:0] m188_41;
   assign m188_41 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_42 = W*in
   wire signed [14:0] m188_42;
   assign m188_42 =15'b0;

   // m188_43 = W*in
   wire signed [14:0] m188_43;
   assign m188_43 =15'b0;

   // m188_44 = W*in
   wire signed [14:0] m188_44;
   assign m188_44 =15'b0;

   // m188_45 = W*in
   wire signed [14:0] m188_45;
   assign m188_45 =15'b0;

   // m188_46 = W*in
   wire signed [14:0] m188_46;
   assign m188_46 =15'b0;

   // m188_47 = W*in
   wire signed [14:0] m188_47;
   assign m188_47 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_48 = W*in
   wire signed [14:0] m188_48;
   assign m188_48 ={ {4{neg188[14]}} , neg188[14:4] };

   // m188_49 = W*in
   wire signed [14:0] m188_49;
   assign m188_49 =15'b0;

   // m188_50 = W*in
   wire signed [14:0] m188_50;
   assign m188_50 =15'b0;

   // m188_51 = W*in
   wire signed [14:0] m188_51;
   assign m188_51 =15'b0;

   // m188_52 = W*in
   wire signed [14:0] m188_52;
   assign m188_52 =15'b0;

   // m188_53 = W*in
   wire signed [14:0] m188_53;
   assign m188_53 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_54 = W*in
   wire signed [14:0] m188_54;
   assign m188_54 =15'b0;

   // m188_55 = W*in
   wire signed [14:0] m188_55;
   assign m188_55 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_56 = W*in
   wire signed [14:0] m188_56;
   assign m188_56 =15'b0;

   // m188_57 = W*in
   wire signed [14:0] m188_57;
   assign m188_57 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_58 = W*in
   wire signed [14:0] m188_58;
   assign m188_58 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_59 = W*in
   wire signed [14:0] m188_59;
   assign m188_59 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_60 = W*in
   wire signed [14:0] m188_60;
   assign m188_60 =15'b0;

   // m188_61 = W*in
   wire signed [14:0] m188_61;
   assign m188_61 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_62 = W*in
   wire signed [14:0] m188_62;
   assign m188_62 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_63 = W*in
   wire signed [14:0] m188_63;
   assign m188_63 ={ {3{in188[14]}} , in188[14:3] };

   // m188_64 = W*in
   wire signed [14:0] m188_64;
   assign m188_64 =15'b0;

   // m188_65 = W*in
   wire signed [14:0] m188_65;
   assign m188_65 =15'b0;

   // m188_66 = W*in
   wire signed [14:0] m188_66;
   assign m188_66 ={ {3{in188[14]}} , in188[14:3] };

   // m188_67 = W*in
   wire signed [14:0] m188_67;
   assign m188_67 =15'b0;

   // m188_68 = W*in
   wire signed [14:0] m188_68;
   assign m188_68 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_69 = W*in
   wire signed [14:0] m188_69;
   assign m188_69 ={ {4{in188[14]}} , in188[14:4] };

   // m188_70 = W*in
   wire signed [14:0] m188_70;
   assign m188_70 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_71 = W*in
   wire signed [14:0] m188_71;
   assign m188_71 =15'b0;

   // m188_72 = W*in
   wire signed [14:0] m188_72;
   assign m188_72 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_73 = W*in
   wire signed [14:0] m188_73;
   assign m188_73 =15'b0;

   // m188_74 = W*in
   wire signed [14:0] m188_74;
   assign m188_74 =15'b0;

   // m188_75 = W*in
   wire signed [14:0] m188_75;
   assign m188_75 =15'b0;

   // m188_76 = W*in
   wire signed [14:0] m188_76;
   assign m188_76 =15'b0;

   // m188_77 = W*in
   wire signed [14:0] m188_77;
   assign m188_77 ={ {4{in188[14]}} , in188[14:4] };

   // m188_78 = W*in
   wire signed [14:0] m188_78;
   assign m188_78 =15'b0;

   // m188_79 = W*in
   wire signed [14:0] m188_79;
   assign m188_79 =15'b0;

   // m188_80 = W*in
   wire signed [14:0] m188_80;
   assign m188_80 =15'b0;

   // m188_81 = W*in
   wire signed [14:0] m188_81;
   assign m188_81 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_82 = W*in
   wire signed [14:0] m188_82;
   assign m188_82 =15'b0;

   // m188_83 = W*in
   wire signed [14:0] m188_83;
   assign m188_83 =15'b0;

   // m188_84 = W*in
   wire signed [14:0] m188_84;
   assign m188_84 =15'b0;

   // m188_85 = W*in
   wire signed [14:0] m188_85;
   assign m188_85 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_86 = W*in
   wire signed [14:0] m188_86;
   assign m188_86 =15'b0;

   // m188_87 = W*in
   wire signed [14:0] m188_87;
   assign m188_87 =15'b0;

   // m188_88 = W*in
   wire signed [14:0] m188_88;
   assign m188_88 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_89 = W*in
   wire signed [14:0] m188_89;
   assign m188_89 =15'b0;

   // m188_90 = W*in
   wire signed [14:0] m188_90;
   assign m188_90 ={ {3{in188[14]}} , in188[14:3] };

   // m188_91 = W*in
   wire signed [14:0] m188_91;
   assign m188_91 =15'b0;

   // m188_92 = W*in
   wire signed [14:0] m188_92;
   assign m188_92 ={ {3{neg188[14]}} , neg188[14:3] };

   // m188_93 = W*in
   wire signed [14:0] m188_93;
   assign m188_93 =15'b0;

   // m188_94 = W*in
   wire signed [14:0] m188_94;
   assign m188_94 =15'b0;

   // m188_95 = W*in
   wire signed [14:0] m188_95;
   assign m188_95 =15'b0;

   // m188_96 = W*in
   wire signed [14:0] m188_96;
   assign m188_96 ={ {3{in188[14]}} , in188[14:3] };

   // m188_97 = W*in
   wire signed [14:0] m188_97;
   assign m188_97 =15'b0;

   // m188_98 = W*in
   wire signed [14:0] m188_98;
   assign m188_98 =15'b0;

   // m188_99 = W*in
   wire signed [14:0] m188_99;
   assign m188_99 =15'b0;

   // m188_100 = W*in
   wire signed [14:0] m188_100;
   assign m188_100 =15'b0;

   // m189_1 = W*in
   wire signed [14:0] m189_1;
   assign m189_1 =15'b0;

   // m189_2 = W*in
   wire signed [14:0] m189_2;
   assign m189_2 =15'b0;

   // m189_3 = W*in
   wire signed [14:0] m189_3;
   assign m189_3 =15'b0;

   // m189_4 = W*in
   wire signed [14:0] m189_4;
   assign m189_4 =15'b0;

   // m189_5 = W*in
   wire signed [14:0] m189_5;
   assign m189_5 =15'b0;

   // m189_6 = W*in
   wire signed [14:0] m189_6;
   assign m189_6 =15'b0;

   // m189_7 = W*in
   wire signed [14:0] m189_7;
   assign m189_7 =15'b0;

   // m189_8 = W*in
   wire signed [14:0] m189_8;
   assign m189_8 =15'b0;

   // m189_9 = W*in
   wire signed [14:0] m189_9;
   assign m189_9 =15'b0;

   // m189_10 = W*in
   wire signed [14:0] m189_10;
   assign m189_10 =15'b0;

   // m189_11 = W*in
   wire signed [14:0] m189_11;
   assign m189_11 =15'b0;

   // m189_12 = W*in
   wire signed [14:0] m189_12;
   assign m189_12 =15'b0;

   // m189_13 = W*in
   wire signed [14:0] m189_13;
   assign m189_13 =15'b0;

   // m189_14 = W*in
   wire signed [14:0] m189_14;
   assign m189_14 =15'b0;

   // m189_15 = W*in
   wire signed [14:0] m189_15;
   assign m189_15 =15'b0;

   // m189_16 = W*in
   wire signed [14:0] m189_16;
   assign m189_16 =15'b0;

   // m189_17 = W*in
   wire signed [14:0] m189_17;
   assign m189_17 =15'b0;

   // m189_18 = W*in
   wire signed [14:0] m189_18;
   assign m189_18 =15'b0;

   // m189_19 = W*in
   wire signed [14:0] m189_19;
   assign m189_19 =15'b0;

   // m189_20 = W*in
   wire signed [14:0] m189_20;
   assign m189_20 =15'b0;

   // m189_21 = W*in
   wire signed [14:0] m189_21;
   assign m189_21 =15'b0;

   // m189_22 = W*in
   wire signed [14:0] m189_22;
   assign m189_22 ={ {4{in189[14]}} , in189[14:4] };

   // m189_23 = W*in
   wire signed [14:0] m189_23;
   assign m189_23 =15'b0;

   // m189_24 = W*in
   wire signed [14:0] m189_24;
   assign m189_24 =15'b0;

   // m189_25 = W*in
   wire signed [14:0] m189_25;
   assign m189_25 =15'b0;

   // m189_26 = W*in
   wire signed [14:0] m189_26;
   assign m189_26 =15'b0;

   // m189_27 = W*in
   wire signed [14:0] m189_27;
   assign m189_27 ={ {4{in189[14]}} , in189[14:4] };

   // m189_28 = W*in
   wire signed [14:0] m189_28;
   assign m189_28 =15'b0;

   // m189_29 = W*in
   wire signed [14:0] m189_29;
   assign m189_29 ={ {4{in189[14]}} , in189[14:4] };

   // m189_30 = W*in
   wire signed [14:0] m189_30;
   assign m189_30 =15'b0;

   // m189_31 = W*in
   wire signed [14:0] m189_31;
   assign m189_31 =15'b0;

   // m189_32 = W*in
   wire signed [14:0] m189_32;
   assign m189_32 =15'b0;

   // m189_33 = W*in
   wire signed [14:0] m189_33;
   assign m189_33 =15'b0;

   // m189_34 = W*in
   wire signed [14:0] m189_34;
   assign m189_34 =15'b0;

   // m189_35 = W*in
   wire signed [14:0] m189_35;
   assign m189_35 =15'b0;

   // m189_36 = W*in
   wire signed [14:0] m189_36;
   assign m189_36 =15'b0;

   // m189_37 = W*in
   wire signed [14:0] m189_37;
   assign m189_37 =15'b0;

   // m189_38 = W*in
   wire signed [14:0] m189_38;
   assign m189_38 =15'b0;

   // m189_39 = W*in
   wire signed [14:0] m189_39;
   assign m189_39 =15'b0;

   // m189_40 = W*in
   wire signed [14:0] m189_40;
   assign m189_40 =15'b0;

   // m189_41 = W*in
   wire signed [14:0] m189_41;
   assign m189_41 =15'b0;

   // m189_42 = W*in
   wire signed [14:0] m189_42;
   assign m189_42 =15'b0;

   // m189_43 = W*in
   wire signed [14:0] m189_43;
   assign m189_43 =15'b0;

   // m189_44 = W*in
   wire signed [14:0] m189_44;
   assign m189_44 =15'b0;

   // m189_45 = W*in
   wire signed [14:0] m189_45;
   assign m189_45 =15'b0;

   // m189_46 = W*in
   wire signed [14:0] m189_46;
   assign m189_46 ={ {4{in189[14]}} , in189[14:4] };

   // m189_47 = W*in
   wire signed [14:0] m189_47;
   assign m189_47 =15'b0;

   // m189_48 = W*in
   wire signed [14:0] m189_48;
   assign m189_48 =15'b0;

   // m189_49 = W*in
   wire signed [14:0] m189_49;
   assign m189_49 =15'b0;

   // m189_50 = W*in
   wire signed [14:0] m189_50;
   assign m189_50 =15'b0;

   // m189_51 = W*in
   wire signed [14:0] m189_51;
   assign m189_51 =15'b0;

   // m189_52 = W*in
   wire signed [14:0] m189_52;
   assign m189_52 =15'b0;

   // m189_53 = W*in
   wire signed [14:0] m189_53;
   assign m189_53 =15'b0;

   // m189_54 = W*in
   wire signed [14:0] m189_54;
   assign m189_54 =15'b0;

   // m189_55 = W*in
   wire signed [14:0] m189_55;
   assign m189_55 =15'b0;

   // m189_56 = W*in
   wire signed [14:0] m189_56;
   assign m189_56 =15'b0;

   // m189_57 = W*in
   wire signed [14:0] m189_57;
   assign m189_57 =15'b0;

   // m189_58 = W*in
   wire signed [14:0] m189_58;
   assign m189_58 =15'b0;

   // m189_59 = W*in
   wire signed [14:0] m189_59;
   assign m189_59 =15'b0;

   // m189_60 = W*in
   wire signed [14:0] m189_60;
   assign m189_60 =15'b0;

   // m189_61 = W*in
   wire signed [14:0] m189_61;
   assign m189_61 =15'b0;

   // m189_62 = W*in
   wire signed [14:0] m189_62;
   assign m189_62 =15'b0;

   // m189_63 = W*in
   wire signed [14:0] m189_63;
   assign m189_63 =15'b0;

   // m189_64 = W*in
   wire signed [14:0] m189_64;
   assign m189_64 =15'b0;

   // m189_65 = W*in
   wire signed [14:0] m189_65;
   assign m189_65 =15'b0;

   // m189_66 = W*in
   wire signed [14:0] m189_66;
   assign m189_66 =15'b0;

   // m189_67 = W*in
   wire signed [14:0] m189_67;
   assign m189_67 =15'b0;

   // m189_68 = W*in
   wire signed [14:0] m189_68;
   assign m189_68 ={ {4{in189[14]}} , in189[14:4] };

   // m189_69 = W*in
   wire signed [14:0] m189_69;
   assign m189_69 =15'b0;

   // m189_70 = W*in
   wire signed [14:0] m189_70;
   assign m189_70 =15'b0;

   // m189_71 = W*in
   wire signed [14:0] m189_71;
   assign m189_71 =15'b0;

   // m189_72 = W*in
   wire signed [14:0] m189_72;
   assign m189_72 =15'b0;

   // m189_73 = W*in
   wire signed [14:0] m189_73;
   assign m189_73 =15'b0;

   // m189_74 = W*in
   wire signed [14:0] m189_74;
   assign m189_74 =15'b0;

   // m189_75 = W*in
   wire signed [14:0] m189_75;
   assign m189_75 =15'b0;

   // m189_76 = W*in
   wire signed [14:0] m189_76;
   assign m189_76 =15'b0;

   // m189_77 = W*in
   wire signed [14:0] m189_77;
   assign m189_77 =15'b0;

   // m189_78 = W*in
   wire signed [14:0] m189_78;
   assign m189_78 =15'b0;

   // m189_79 = W*in
   wire signed [14:0] m189_79;
   assign m189_79 =15'b0;

   // m189_80 = W*in
   wire signed [14:0] m189_80;
   assign m189_80 =15'b0;

   // m189_81 = W*in
   wire signed [14:0] m189_81;
   assign m189_81 =15'b0;

   // m189_82 = W*in
   wire signed [14:0] m189_82;
   assign m189_82 =15'b0;

   // m189_83 = W*in
   wire signed [14:0] m189_83;
   assign m189_83 =15'b0;

   // m189_84 = W*in
   wire signed [14:0] m189_84;
   assign m189_84 =15'b0;

   // m189_85 = W*in
   wire signed [14:0] m189_85;
   assign m189_85 =15'b0;

   // m189_86 = W*in
   wire signed [14:0] m189_86;
   assign m189_86 =15'b0;

   // m189_87 = W*in
   wire signed [14:0] m189_87;
   assign m189_87 =15'b0;

   // m189_88 = W*in
   wire signed [14:0] m189_88;
   assign m189_88 =15'b0;

   // m189_89 = W*in
   wire signed [14:0] m189_89;
   assign m189_89 =15'b0;

   // m189_90 = W*in
   wire signed [14:0] m189_90;
   assign m189_90 =15'b0;

   // m189_91 = W*in
   wire signed [14:0] m189_91;
   assign m189_91 =15'b0;

   // m189_92 = W*in
   wire signed [14:0] m189_92;
   assign m189_92 =15'b0;

   // m189_93 = W*in
   wire signed [14:0] m189_93;
   assign m189_93 =15'b0;

   // m189_94 = W*in
   wire signed [14:0] m189_94;
   assign m189_94 =15'b0;

   // m189_95 = W*in
   wire signed [14:0] m189_95;
   assign m189_95 =15'b0;

   // m189_96 = W*in
   wire signed [14:0] m189_96;
   assign m189_96 =15'b0;

   // m189_97 = W*in
   wire signed [14:0] m189_97;
   assign m189_97 =15'b0;

   // m189_98 = W*in
   wire signed [14:0] m189_98;
   assign m189_98 =15'b0;

   // m189_99 = W*in
   wire signed [14:0] m189_99;
   assign m189_99 =15'b0;

   // m189_100 = W*in
   wire signed [14:0] m189_100;
   assign m189_100 =15'b0;

   // m190_1 = W*in
   wire signed [14:0] m190_1;
   assign m190_1 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_2 = W*in
   wire signed [14:0] m190_2;
   assign m190_2 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_3 = W*in
   wire signed [14:0] m190_3;
   assign m190_3 =15'b0;

   // m190_4 = W*in
   wire signed [14:0] m190_4;
   assign m190_4 =15'b0;

   // m190_5 = W*in
   wire signed [14:0] m190_5;
   assign m190_5 ={ {4{neg190[14]}} , neg190[14:4] };

   // m190_6 = W*in
   wire signed [14:0] m190_6;
   assign m190_6 =15'b0;

   // m190_7 = W*in
   wire signed [14:0] m190_7;
   assign m190_7 =15'b0;

   // m190_8 = W*in
   wire signed [14:0] m190_8;
   assign m190_8 =15'b0;

   // m190_9 = W*in
   wire signed [14:0] m190_9;
   assign m190_9 =15'b0;

   // m190_10 = W*in
   wire signed [14:0] m190_10;
   assign m190_10 =15'b0;

   // m190_11 = W*in
   wire signed [14:0] m190_11;
   assign m190_11 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_12 = W*in
   wire signed [14:0] m190_12;
   assign m190_12 =15'b0;

   // m190_13 = W*in
   wire signed [14:0] m190_13;
   assign m190_13 =15'b0;

   // m190_14 = W*in
   wire signed [14:0] m190_14;
   assign m190_14 =15'b0;

   // m190_15 = W*in
   wire signed [14:0] m190_15;
   assign m190_15 =15'b0;

   // m190_16 = W*in
   wire signed [14:0] m190_16;
   assign m190_16 =15'b0;

   // m190_17 = W*in
   wire signed [14:0] m190_17;
   assign m190_17 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_18 = W*in
   wire signed [14:0] m190_18;
   assign m190_18 =15'b0;

   // m190_19 = W*in
   wire signed [14:0] m190_19;
   assign m190_19 =15'b0;

   // m190_20 = W*in
   wire signed [14:0] m190_20;
   assign m190_20 =15'b0;

   // m190_21 = W*in
   wire signed [14:0] m190_21;
   assign m190_21 ={ {4{neg190[14]}} , neg190[14:4] };

   // m190_22 = W*in
   wire signed [14:0] m190_22;
   assign m190_22 ={ {4{neg190[14]}} , neg190[14:4] };

   // m190_23 = W*in
   wire signed [14:0] m190_23;
   assign m190_23 =15'b0;

   // m190_24 = W*in
   wire signed [14:0] m190_24;
   assign m190_24 =15'b0;

   // m190_25 = W*in
   wire signed [14:0] m190_25;
   assign m190_25 =15'b0;

   // m190_26 = W*in
   wire signed [14:0] m190_26;
   assign m190_26 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_27 = W*in
   wire signed [14:0] m190_27;
   assign m190_27 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_28 = W*in
   wire signed [14:0] m190_28;
   assign m190_28 =15'b0;

   // m190_29 = W*in
   wire signed [14:0] m190_29;
   assign m190_29 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_30 = W*in
   wire signed [14:0] m190_30;
   assign m190_30 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_31 = W*in
   wire signed [14:0] m190_31;
   assign m190_31 =15'b0;

   // m190_32 = W*in
   wire signed [14:0] m190_32;
   assign m190_32 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_33 = W*in
   wire signed [14:0] m190_33;
   assign m190_33 =15'b0;

   // m190_34 = W*in
   wire signed [14:0] m190_34;
   assign m190_34 =15'b0;

   // m190_35 = W*in
   wire signed [14:0] m190_35;
   assign m190_35 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_36 = W*in
   wire signed [14:0] m190_36;
   assign m190_36 =15'b0;

   // m190_37 = W*in
   wire signed [14:0] m190_37;
   assign m190_37 =15'b0;

   // m190_38 = W*in
   wire signed [14:0] m190_38;
   assign m190_38 =15'b0;

   // m190_39 = W*in
   wire signed [14:0] m190_39;
   assign m190_39 =15'b0;

   // m190_40 = W*in
   wire signed [14:0] m190_40;
   assign m190_40 =15'b0;

   // m190_41 = W*in
   wire signed [14:0] m190_41;
   assign m190_41 =15'b0;

   // m190_42 = W*in
   wire signed [14:0] m190_42;
   assign m190_42 =15'b0;

   // m190_43 = W*in
   wire signed [14:0] m190_43;
   assign m190_43 =15'b0;

   // m190_44 = W*in
   wire signed [14:0] m190_44;
   assign m190_44 =15'b0;

   // m190_45 = W*in
   wire signed [14:0] m190_45;
   assign m190_45 =15'b0;

   // m190_46 = W*in
   wire signed [14:0] m190_46;
   assign m190_46 =15'b0;

   // m190_47 = W*in
   wire signed [14:0] m190_47;
   assign m190_47 =15'b0;

   // m190_48 = W*in
   wire signed [14:0] m190_48;
   assign m190_48 ={ {3{in190[14]}} , in190[14:3] };

   // m190_49 = W*in
   wire signed [14:0] m190_49;
   assign m190_49 =15'b0;

   // m190_50 = W*in
   wire signed [14:0] m190_50;
   assign m190_50 =15'b0;

   // m190_51 = W*in
   wire signed [14:0] m190_51;
   assign m190_51 ={ {3{in190[14]}} , in190[14:3] };

   // m190_52 = W*in
   wire signed [14:0] m190_52;
   assign m190_52 =15'b0;

   // m190_53 = W*in
   wire signed [14:0] m190_53;
   assign m190_53 ={ {3{in190[14]}} , in190[14:3] };

   // m190_54 = W*in
   wire signed [14:0] m190_54;
   assign m190_54 =15'b0;

   // m190_55 = W*in
   wire signed [14:0] m190_55;
   assign m190_55 =15'b0;

   // m190_56 = W*in
   wire signed [14:0] m190_56;
   assign m190_56 ={ {3{in190[14]}} , in190[14:3] };

   // m190_57 = W*in
   wire signed [14:0] m190_57;
   assign m190_57 ={ {3{in190[14]}} , in190[14:3] };

   // m190_58 = W*in
   wire signed [14:0] m190_58;
   assign m190_58 ={ {3{in190[14]}} , in190[14:3] };

   // m190_59 = W*in
   wire signed [14:0] m190_59;
   assign m190_59 =15'b0;

   // m190_60 = W*in
   wire signed [14:0] m190_60;
   assign m190_60 ={ {4{neg190[14]}} , neg190[14:4] };

   // m190_61 = W*in
   wire signed [14:0] m190_61;
   assign m190_61 =15'b0;

   // m190_62 = W*in
   wire signed [14:0] m190_62;
   assign m190_62 =15'b0;

   // m190_63 = W*in
   wire signed [14:0] m190_63;
   assign m190_63 =15'b0;

   // m190_64 = W*in
   wire signed [14:0] m190_64;
   assign m190_64 ={ {3{in190[14]}} , in190[14:3] };

   // m190_65 = W*in
   wire signed [14:0] m190_65;
   assign m190_65 =15'b0;

   // m190_66 = W*in
   wire signed [14:0] m190_66;
   assign m190_66 =15'b0;

   // m190_67 = W*in
   wire signed [14:0] m190_67;
   assign m190_67 =15'b0;

   // m190_68 = W*in
   wire signed [14:0] m190_68;
   assign m190_68 =15'b0;

   // m190_69 = W*in
   wire signed [14:0] m190_69;
   assign m190_69 =15'b0;

   // m190_70 = W*in
   wire signed [14:0] m190_70;
   assign m190_70 =15'b0;

   // m190_71 = W*in
   wire signed [14:0] m190_71;
   assign m190_71 =15'b0;

   // m190_72 = W*in
   wire signed [14:0] m190_72;
   assign m190_72 =15'b0;

   // m190_73 = W*in
   wire signed [14:0] m190_73;
   assign m190_73 =15'b0;

   // m190_74 = W*in
   wire signed [14:0] m190_74;
   assign m190_74 ={ {3{in190[14]}} , in190[14:3] };

   // m190_75 = W*in
   wire signed [14:0] m190_75;
   assign m190_75 =15'b0;

   // m190_76 = W*in
   wire signed [14:0] m190_76;
   assign m190_76 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_77 = W*in
   wire signed [14:0] m190_77;
   assign m190_77 =15'b0;

   // m190_78 = W*in
   wire signed [14:0] m190_78;
   assign m190_78 =15'b0;

   // m190_79 = W*in
   wire signed [14:0] m190_79;
   assign m190_79 =15'b0;

   // m190_80 = W*in
   wire signed [14:0] m190_80;
   assign m190_80 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_81 = W*in
   wire signed [14:0] m190_81;
   assign m190_81 =15'b0;

   // m190_82 = W*in
   wire signed [14:0] m190_82;
   assign m190_82 =15'b0;

   // m190_83 = W*in
   wire signed [14:0] m190_83;
   assign m190_83 =15'b0;

   // m190_84 = W*in
   wire signed [14:0] m190_84;
   assign m190_84 =15'b0;

   // m190_85 = W*in
   wire signed [14:0] m190_85;
   assign m190_85 ={ {3{in190[14]}} , in190[14:3] };

   // m190_86 = W*in
   wire signed [14:0] m190_86;
   assign m190_86 =15'b0;

   // m190_87 = W*in
   wire signed [14:0] m190_87;
   assign m190_87 =15'b0;

   // m190_88 = W*in
   wire signed [14:0] m190_88;
   assign m190_88 =15'b0;

   // m190_89 = W*in
   wire signed [14:0] m190_89;
   assign m190_89 =15'b0;

   // m190_90 = W*in
   wire signed [14:0] m190_90;
   assign m190_90 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_91 = W*in
   wire signed [14:0] m190_91;
   assign m190_91 ={ {3{in190[14]}} , in190[14:3] };

   // m190_92 = W*in
   wire signed [14:0] m190_92;
   assign m190_92 ={ {3{in190[14]}} , in190[14:3] };

   // m190_93 = W*in
   wire signed [14:0] m190_93;
   assign m190_93 =15'b0;

   // m190_94 = W*in
   wire signed [14:0] m190_94;
   assign m190_94 ={ {4{neg190[14]}} , neg190[14:4] };

   // m190_95 = W*in
   wire signed [14:0] m190_95;
   assign m190_95 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_96 = W*in
   wire signed [14:0] m190_96;
   assign m190_96 ={ {3{neg190[14]}} , neg190[14:3] };

   // m190_97 = W*in
   wire signed [14:0] m190_97;
   assign m190_97 =15'b0;

   // m190_98 = W*in
   wire signed [14:0] m190_98;
   assign m190_98 =15'b0;

   // m190_99 = W*in
   wire signed [14:0] m190_99;
   assign m190_99 =15'b0;

   // m190_100 = W*in
   wire signed [14:0] m190_100;
   assign m190_100 =15'b0;

   // m191_1 = W*in
   wire signed [14:0] m191_1;
   assign m191_1 =15'b0;

   // m191_2 = W*in
   wire signed [14:0] m191_2;
   assign m191_2 =15'b0;

   // m191_3 = W*in
   wire signed [14:0] m191_3;
   assign m191_3 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_4 = W*in
   wire signed [14:0] m191_4;
   assign m191_4 =15'b0;

   // m191_5 = W*in
   wire signed [14:0] m191_5;
   assign m191_5 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_6 = W*in
   wire signed [14:0] m191_6;
   assign m191_6 =15'b0;

   // m191_7 = W*in
   wire signed [14:0] m191_7;
   assign m191_7 ={ {2{in191[14]}} , in191[14:2] };

   // m191_8 = W*in
   wire signed [14:0] m191_8;
   assign m191_8 ={ {3{in191[14]}} , in191[14:3] };

   // m191_9 = W*in
   wire signed [14:0] m191_9;
   assign m191_9 =15'b0;

   // m191_10 = W*in
   wire signed [14:0] m191_10;
   assign m191_10 =15'b0;

   // m191_11 = W*in
   wire signed [14:0] m191_11;
   assign m191_11 =15'b0;

   // m191_12 = W*in
   wire signed [14:0] m191_12;
   assign m191_12 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_13 = W*in
   wire signed [14:0] m191_13;
   assign m191_13 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_14 = W*in
   wire signed [14:0] m191_14;
   assign m191_14 ={ {3{in191[14]}} , in191[14:3] };

   // m191_15 = W*in
   wire signed [14:0] m191_15;
   assign m191_15 =15'b0;

   // m191_16 = W*in
   wire signed [14:0] m191_16;
   assign m191_16 =15'b0;

   // m191_17 = W*in
   wire signed [14:0] m191_17;
   assign m191_17 =15'b0;

   // m191_18 = W*in
   wire signed [14:0] m191_18;
   assign m191_18 =15'b0;

   // m191_19 = W*in
   wire signed [14:0] m191_19;
   assign m191_19 ={ {4{in191[14]}} , in191[14:4] };

   // m191_20 = W*in
   wire signed [14:0] m191_20;
   assign m191_20 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_21 = W*in
   wire signed [14:0] m191_21;
   assign m191_21 =15'b0;

   // m191_22 = W*in
   wire signed [14:0] m191_22;
   assign m191_22 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_23 = W*in
   wire signed [14:0] m191_23;
   assign m191_23 =15'b0;

   // m191_24 = W*in
   wire signed [14:0] m191_24;
   assign m191_24 =15'b0;

   // m191_25 = W*in
   wire signed [14:0] m191_25;
   assign m191_25 =15'b0;

   // m191_26 = W*in
   wire signed [14:0] m191_26;
   assign m191_26 =15'b0;

   // m191_27 = W*in
   wire signed [14:0] m191_27;
   assign m191_27 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_28 = W*in
   wire signed [14:0] m191_28;
   assign m191_28 =15'b0;

   // m191_29 = W*in
   wire signed [14:0] m191_29;
   assign m191_29 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_30 = W*in
   wire signed [14:0] m191_30;
   assign m191_30 =15'b0;

   // m191_31 = W*in
   wire signed [14:0] m191_31;
   assign m191_31 ={ {3{in191[14]}} , in191[14:3] };

   // m191_32 = W*in
   wire signed [14:0] m191_32;
   assign m191_32 ={ {3{in191[14]}} , in191[14:3] };

   // m191_33 = W*in
   wire signed [14:0] m191_33;
   assign m191_33 =15'b0;

   // m191_34 = W*in
   wire signed [14:0] m191_34;
   assign m191_34 =15'b0;

   // m191_35 = W*in
   wire signed [14:0] m191_35;
   assign m191_35 =15'b0;

   // m191_36 = W*in
   wire signed [14:0] m191_36;
   assign m191_36 =15'b0;

   // m191_37 = W*in
   wire signed [14:0] m191_37;
   assign m191_37 =15'b0;

   // m191_38 = W*in
   wire signed [14:0] m191_38;
   assign m191_38 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_39 = W*in
   wire signed [14:0] m191_39;
   assign m191_39 =15'b0;

   // m191_40 = W*in
   wire signed [14:0] m191_40;
   assign m191_40 =15'b0;

   // m191_41 = W*in
   wire signed [14:0] m191_41;
   assign m191_41 =15'b0;

   // m191_42 = W*in
   wire signed [14:0] m191_42;
   assign m191_42 ={ {3{in191[14]}} , in191[14:3] };

   // m191_43 = W*in
   wire signed [14:0] m191_43;
   assign m191_43 =15'b0;

   // m191_44 = W*in
   wire signed [14:0] m191_44;
   assign m191_44 ={ {3{in191[14]}} , in191[14:3] };

   // m191_45 = W*in
   wire signed [14:0] m191_45;
   assign m191_45 =15'b0;

   // m191_46 = W*in
   wire signed [14:0] m191_46;
   assign m191_46 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_47 = W*in
   wire signed [14:0] m191_47;
   assign m191_47 ={ {3{in191[14]}} , in191[14:3] };

   // m191_48 = W*in
   wire signed [14:0] m191_48;
   assign m191_48 =15'b0;

   // m191_49 = W*in
   wire signed [14:0] m191_49;
   assign m191_49 =15'b0;

   // m191_50 = W*in
   wire signed [14:0] m191_50;
   assign m191_50 =15'b0;

   // m191_51 = W*in
   wire signed [14:0] m191_51;
   assign m191_51 =15'b0;

   // m191_52 = W*in
   wire signed [14:0] m191_52;
   assign m191_52 =15'b0;

   // m191_53 = W*in
   wire signed [14:0] m191_53;
   assign m191_53 =15'b0;

   // m191_54 = W*in
   wire signed [14:0] m191_54;
   assign m191_54 ={ {3{in191[14]}} , in191[14:3] };

   // m191_55 = W*in
   wire signed [14:0] m191_55;
   assign m191_55 =15'b0;

   // m191_56 = W*in
   wire signed [14:0] m191_56;
   assign m191_56 =15'b0;

   // m191_57 = W*in
   wire signed [14:0] m191_57;
   assign m191_57 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_58 = W*in
   wire signed [14:0] m191_58;
   assign m191_58 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_59 = W*in
   wire signed [14:0] m191_59;
   assign m191_59 =15'b0;

   // m191_60 = W*in
   wire signed [14:0] m191_60;
   assign m191_60 =15'b0;

   // m191_61 = W*in
   wire signed [14:0] m191_61;
   assign m191_61 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_62 = W*in
   wire signed [14:0] m191_62;
   assign m191_62 ={ {2{neg191[14]}} , neg191[14:2] };

   // m191_63 = W*in
   wire signed [14:0] m191_63;
   assign m191_63 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_64 = W*in
   wire signed [14:0] m191_64;
   assign m191_64 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_65 = W*in
   wire signed [14:0] m191_65;
   assign m191_65 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_66 = W*in
   wire signed [14:0] m191_66;
   assign m191_66 =15'b0;

   // m191_67 = W*in
   wire signed [14:0] m191_67;
   assign m191_67 ={ {3{in191[14]}} , in191[14:3] };

   // m191_68 = W*in
   wire signed [14:0] m191_68;
   assign m191_68 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_69 = W*in
   wire signed [14:0] m191_69;
   assign m191_69 =15'b0;

   // m191_70 = W*in
   wire signed [14:0] m191_70;
   assign m191_70 ={ {3{in191[14]}} , in191[14:3] };

   // m191_71 = W*in
   wire signed [14:0] m191_71;
   assign m191_71 =15'b0;

   // m191_72 = W*in
   wire signed [14:0] m191_72;
   assign m191_72 =15'b0;

   // m191_73 = W*in
   wire signed [14:0] m191_73;
   assign m191_73 =15'b0;

   // m191_74 = W*in
   wire signed [14:0] m191_74;
   assign m191_74 ={ {4{neg191[14]}} , neg191[14:4] };

   // m191_75 = W*in
   wire signed [14:0] m191_75;
   assign m191_75 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_76 = W*in
   wire signed [14:0] m191_76;
   assign m191_76 =15'b0;

   // m191_77 = W*in
   wire signed [14:0] m191_77;
   assign m191_77 =15'b0;

   // m191_78 = W*in
   wire signed [14:0] m191_78;
   assign m191_78 =15'b0;

   // m191_79 = W*in
   wire signed [14:0] m191_79;
   assign m191_79 =15'b0;

   // m191_80 = W*in
   wire signed [14:0] m191_80;
   assign m191_80 =15'b0;

   // m191_81 = W*in
   wire signed [14:0] m191_81;
   assign m191_81 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_82 = W*in
   wire signed [14:0] m191_82;
   assign m191_82 =15'b0;

   // m191_83 = W*in
   wire signed [14:0] m191_83;
   assign m191_83 =15'b0;

   // m191_84 = W*in
   wire signed [14:0] m191_84;
   assign m191_84 =15'b0;

   // m191_85 = W*in
   wire signed [14:0] m191_85;
   assign m191_85 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_86 = W*in
   wire signed [14:0] m191_86;
   assign m191_86 =15'b0;

   // m191_87 = W*in
   wire signed [14:0] m191_87;
   assign m191_87 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_88 = W*in
   wire signed [14:0] m191_88;
   assign m191_88 =15'b0;

   // m191_89 = W*in
   wire signed [14:0] m191_89;
   assign m191_89 =15'b0;

   // m191_90 = W*in
   wire signed [14:0] m191_90;
   assign m191_90 =15'b0;

   // m191_91 = W*in
   wire signed [14:0] m191_91;
   assign m191_91 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_92 = W*in
   wire signed [14:0] m191_92;
   assign m191_92 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_93 = W*in
   wire signed [14:0] m191_93;
   assign m191_93 ={ {3{neg191[14]}} , neg191[14:3] };

   // m191_94 = W*in
   wire signed [14:0] m191_94;
   assign m191_94 ={ {4{in191[14]}} , in191[14:4] };

   // m191_95 = W*in
   wire signed [14:0] m191_95;
   assign m191_95 ={ {3{in191[14]}} , in191[14:3] };

   // m191_96 = W*in
   wire signed [14:0] m191_96;
   assign m191_96 =15'b0;

   // m191_97 = W*in
   wire signed [14:0] m191_97;
   assign m191_97 ={ {2{neg191[14]}} , neg191[14:2] };

   // m191_98 = W*in
   wire signed [14:0] m191_98;
   assign m191_98 ={ {3{in191[14]}} , in191[14:3] };

   // m191_99 = W*in
   wire signed [14:0] m191_99;
   assign m191_99 =15'b0;

   // m191_100 = W*in
   wire signed [14:0] m191_100;
   assign m191_100 =15'b0;

   // m192_1 = W*in
   wire signed [14:0] m192_1;
   assign m192_1 =15'b0;

   // m192_2 = W*in
   wire signed [14:0] m192_2;
   assign m192_2 =15'b0;

   // m192_3 = W*in
   wire signed [14:0] m192_3;
   assign m192_3 ={ {4{neg192[14]}} , neg192[14:4] };

   // m192_4 = W*in
   wire signed [14:0] m192_4;
   assign m192_4 =15'b0;

   // m192_5 = W*in
   wire signed [14:0] m192_5;
   assign m192_5 =15'b0;

   // m192_6 = W*in
   wire signed [14:0] m192_6;
   assign m192_6 =15'b0;

   // m192_7 = W*in
   wire signed [14:0] m192_7;
   assign m192_7 =15'b0;

   // m192_8 = W*in
   wire signed [14:0] m192_8;
   assign m192_8 =15'b0;

   // m192_9 = W*in
   wire signed [14:0] m192_9;
   assign m192_9 =15'b0;

   // m192_10 = W*in
   wire signed [14:0] m192_10;
   assign m192_10 ={ {3{in192[14]}} , in192[14:3] };

   // m192_11 = W*in
   wire signed [14:0] m192_11;
   assign m192_11 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_12 = W*in
   wire signed [14:0] m192_12;
   assign m192_12 =15'b0;

   // m192_13 = W*in
   wire signed [14:0] m192_13;
   assign m192_13 =15'b0;

   // m192_14 = W*in
   wire signed [14:0] m192_14;
   assign m192_14 =15'b0;

   // m192_15 = W*in
   wire signed [14:0] m192_15;
   assign m192_15 =15'b0;

   // m192_16 = W*in
   wire signed [14:0] m192_16;
   assign m192_16 ={ {3{in192[14]}} , in192[14:3] };

   // m192_17 = W*in
   wire signed [14:0] m192_17;
   assign m192_17 =15'b0;

   // m192_18 = W*in
   wire signed [14:0] m192_18;
   assign m192_18 =15'b0;

   // m192_19 = W*in
   wire signed [14:0] m192_19;
   assign m192_19 =15'b0;

   // m192_20 = W*in
   wire signed [14:0] m192_20;
   assign m192_20 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_21 = W*in
   wire signed [14:0] m192_21;
   assign m192_21 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_22 = W*in
   wire signed [14:0] m192_22;
   assign m192_22 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_23 = W*in
   wire signed [14:0] m192_23;
   assign m192_23 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_24 = W*in
   wire signed [14:0] m192_24;
   assign m192_24 =15'b0;

   // m192_25 = W*in
   wire signed [14:0] m192_25;
   assign m192_25 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_26 = W*in
   wire signed [14:0] m192_26;
   assign m192_26 =15'b0;

   // m192_27 = W*in
   wire signed [14:0] m192_27;
   assign m192_27 =15'b0;

   // m192_28 = W*in
   wire signed [14:0] m192_28;
   assign m192_28 =15'b0;

   // m192_29 = W*in
   wire signed [14:0] m192_29;
   assign m192_29 =15'b0;

   // m192_30 = W*in
   wire signed [14:0] m192_30;
   assign m192_30 =15'b0;

   // m192_31 = W*in
   wire signed [14:0] m192_31;
   assign m192_31 =15'b0;

   // m192_32 = W*in
   wire signed [14:0] m192_32;
   assign m192_32 =15'b0;

   // m192_33 = W*in
   wire signed [14:0] m192_33;
   assign m192_33 =15'b0;

   // m192_34 = W*in
   wire signed [14:0] m192_34;
   assign m192_34 ={ {4{neg192[14]}} , neg192[14:4] };

   // m192_35 = W*in
   wire signed [14:0] m192_35;
   assign m192_35 =15'b0;

   // m192_36 = W*in
   wire signed [14:0] m192_36;
   assign m192_36 ={ {3{in192[14]}} , in192[14:3] };

   // m192_37 = W*in
   wire signed [14:0] m192_37;
   assign m192_37 =15'b0;

   // m192_38 = W*in
   wire signed [14:0] m192_38;
   assign m192_38 =15'b0;

   // m192_39 = W*in
   wire signed [14:0] m192_39;
   assign m192_39 =15'b0;

   // m192_40 = W*in
   wire signed [14:0] m192_40;
   assign m192_40 =15'b0;

   // m192_41 = W*in
   wire signed [14:0] m192_41;
   assign m192_41 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_42 = W*in
   wire signed [14:0] m192_42;
   assign m192_42 =15'b0;

   // m192_43 = W*in
   wire signed [14:0] m192_43;
   assign m192_43 =15'b0;

   // m192_44 = W*in
   wire signed [14:0] m192_44;
   assign m192_44 =15'b0;

   // m192_45 = W*in
   wire signed [14:0] m192_45;
   assign m192_45 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_46 = W*in
   wire signed [14:0] m192_46;
   assign m192_46 =15'b0;

   // m192_47 = W*in
   wire signed [14:0] m192_47;
   assign m192_47 =15'b0;

   // m192_48 = W*in
   wire signed [14:0] m192_48;
   assign m192_48 ={ {3{in192[14]}} , in192[14:3] };

   // m192_49 = W*in
   wire signed [14:0] m192_49;
   assign m192_49 =15'b0;

   // m192_50 = W*in
   wire signed [14:0] m192_50;
   assign m192_50 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_51 = W*in
   wire signed [14:0] m192_51;
   assign m192_51 =15'b0;

   // m192_52 = W*in
   wire signed [14:0] m192_52;
   assign m192_52 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_53 = W*in
   wire signed [14:0] m192_53;
   assign m192_53 =15'b0;

   // m192_54 = W*in
   wire signed [14:0] m192_54;
   assign m192_54 =15'b0;

   // m192_55 = W*in
   wire signed [14:0] m192_55;
   assign m192_55 ={ {3{in192[14]}} , in192[14:3] };

   // m192_56 = W*in
   wire signed [14:0] m192_56;
   assign m192_56 =15'b0;

   // m192_57 = W*in
   wire signed [14:0] m192_57;
   assign m192_57 =15'b0;

   // m192_58 = W*in
   wire signed [14:0] m192_58;
   assign m192_58 =15'b0;

   // m192_59 = W*in
   wire signed [14:0] m192_59;
   assign m192_59 =15'b0;

   // m192_60 = W*in
   wire signed [14:0] m192_60;
   assign m192_60 =15'b0;

   // m192_61 = W*in
   wire signed [14:0] m192_61;
   assign m192_61 ={ {3{in192[14]}} , in192[14:3] };

   // m192_62 = W*in
   wire signed [14:0] m192_62;
   assign m192_62 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_63 = W*in
   wire signed [14:0] m192_63;
   assign m192_63 ={ {2{in192[14]}} , in192[14:2] };

   // m192_64 = W*in
   wire signed [14:0] m192_64;
   assign m192_64 ={ {4{neg192[14]}} , neg192[14:4] };

   // m192_65 = W*in
   wire signed [14:0] m192_65;
   assign m192_65 =15'b0;

   // m192_66 = W*in
   wire signed [14:0] m192_66;
   assign m192_66 ={ {2{in192[14]}} , in192[14:2] };

   // m192_67 = W*in
   wire signed [14:0] m192_67;
   assign m192_67 ={ {4{neg192[14]}} , neg192[14:4] };

   // m192_68 = W*in
   wire signed [14:0] m192_68;
   assign m192_68 =15'b0;

   // m192_69 = W*in
   wire signed [14:0] m192_69;
   assign m192_69 =15'b0;

   // m192_70 = W*in
   wire signed [14:0] m192_70;
   assign m192_70 =15'b0;

   // m192_71 = W*in
   wire signed [14:0] m192_71;
   assign m192_71 ={ {3{in192[14]}} , in192[14:3] };

   // m192_72 = W*in
   wire signed [14:0] m192_72;
   assign m192_72 =15'b0;

   // m192_73 = W*in
   wire signed [14:0] m192_73;
   assign m192_73 =15'b0;

   // m192_74 = W*in
   wire signed [14:0] m192_74;
   assign m192_74 ={ {4{neg192[14]}} , neg192[14:4] };

   // m192_75 = W*in
   wire signed [14:0] m192_75;
   assign m192_75 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_76 = W*in
   wire signed [14:0] m192_76;
   assign m192_76 =15'b0;

   // m192_77 = W*in
   wire signed [14:0] m192_77;
   assign m192_77 =15'b0;

   // m192_78 = W*in
   wire signed [14:0] m192_78;
   assign m192_78 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_79 = W*in
   wire signed [14:0] m192_79;
   assign m192_79 =15'b0;

   // m192_80 = W*in
   wire signed [14:0] m192_80;
   assign m192_80 =15'b0;

   // m192_81 = W*in
   wire signed [14:0] m192_81;
   assign m192_81 =15'b0;

   // m192_82 = W*in
   wire signed [14:0] m192_82;
   assign m192_82 =15'b0;

   // m192_83 = W*in
   wire signed [14:0] m192_83;
   assign m192_83 ={ {3{in192[14]}} , in192[14:3] };

   // m192_84 = W*in
   wire signed [14:0] m192_84;
   assign m192_84 =15'b0;

   // m192_85 = W*in
   wire signed [14:0] m192_85;
   assign m192_85 =15'b0;

   // m192_86 = W*in
   wire signed [14:0] m192_86;
   assign m192_86 =15'b0;

   // m192_87 = W*in
   wire signed [14:0] m192_87;
   assign m192_87 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_88 = W*in
   wire signed [14:0] m192_88;
   assign m192_88 ={ {3{neg192[14]}} , neg192[14:3] };

   // m192_89 = W*in
   wire signed [14:0] m192_89;
   assign m192_89 ={ {3{in192[14]}} , in192[14:3] };

   // m192_90 = W*in
   wire signed [14:0] m192_90;
   assign m192_90 =15'b0;

   // m192_91 = W*in
   wire signed [14:0] m192_91;
   assign m192_91 =15'b0;

   // m192_92 = W*in
   wire signed [14:0] m192_92;
   assign m192_92 =15'b0;

   // m192_93 = W*in
   wire signed [14:0] m192_93;
   assign m192_93 ={ {3{in192[14]}} , in192[14:3] };

   // m192_94 = W*in
   wire signed [14:0] m192_94;
   assign m192_94 =15'b0;

   // m192_95 = W*in
   wire signed [14:0] m192_95;
   assign m192_95 =15'b0;

   // m192_96 = W*in
   wire signed [14:0] m192_96;
   assign m192_96 ={ {4{neg192[14]}} , neg192[14:4] };

   // m192_97 = W*in
   wire signed [14:0] m192_97;
   assign m192_97 =15'b0;

   // m192_98 = W*in
   wire signed [14:0] m192_98;
   assign m192_98 =15'b0;

   // m192_99 = W*in
   wire signed [14:0] m192_99;
   assign m192_99 =15'b0;

   // m192_100 = W*in
   wire signed [14:0] m192_100;
   assign m192_100 ={ {2{in192[14]}} , in192[14:2] };

   // m193_1 = W*in
   wire signed [14:0] m193_1;
   assign m193_1 =15'b0;

   // m193_2 = W*in
   wire signed [14:0] m193_2;
   assign m193_2 =15'b0;

   // m193_3 = W*in
   wire signed [14:0] m193_3;
   assign m193_3 =15'b0;

   // m193_4 = W*in
   wire signed [14:0] m193_4;
   assign m193_4 =15'b0;

   // m193_5 = W*in
   wire signed [14:0] m193_5;
   assign m193_5 =15'b0;

   // m193_6 = W*in
   wire signed [14:0] m193_6;
   assign m193_6 =15'b0;

   // m193_7 = W*in
   wire signed [14:0] m193_7;
   assign m193_7 =15'b0;

   // m193_8 = W*in
   wire signed [14:0] m193_8;
   assign m193_8 =15'b0;

   // m193_9 = W*in
   wire signed [14:0] m193_9;
   assign m193_9 =15'b0;

   // m193_10 = W*in
   wire signed [14:0] m193_10;
   assign m193_10 =15'b0;

   // m193_11 = W*in
   wire signed [14:0] m193_11;
   assign m193_11 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_12 = W*in
   wire signed [14:0] m193_12;
   assign m193_12 =15'b0;

   // m193_13 = W*in
   wire signed [14:0] m193_13;
   assign m193_13 =15'b0;

   // m193_14 = W*in
   wire signed [14:0] m193_14;
   assign m193_14 =15'b0;

   // m193_15 = W*in
   wire signed [14:0] m193_15;
   assign m193_15 =15'b0;

   // m193_16 = W*in
   wire signed [14:0] m193_16;
   assign m193_16 =15'b0;

   // m193_17 = W*in
   wire signed [14:0] m193_17;
   assign m193_17 =15'b0;

   // m193_18 = W*in
   wire signed [14:0] m193_18;
   assign m193_18 =15'b0;

   // m193_19 = W*in
   wire signed [14:0] m193_19;
   assign m193_19 =15'b0;

   // m193_20 = W*in
   wire signed [14:0] m193_20;
   assign m193_20 =15'b0;

   // m193_21 = W*in
   wire signed [14:0] m193_21;
   assign m193_21 =15'b0;

   // m193_22 = W*in
   wire signed [14:0] m193_22;
   assign m193_22 =15'b0;

   // m193_23 = W*in
   wire signed [14:0] m193_23;
   assign m193_23 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_24 = W*in
   wire signed [14:0] m193_24;
   assign m193_24 =15'b0;

   // m193_25 = W*in
   wire signed [14:0] m193_25;
   assign m193_25 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_26 = W*in
   wire signed [14:0] m193_26;
   assign m193_26 =15'b0;

   // m193_27 = W*in
   wire signed [14:0] m193_27;
   assign m193_27 =15'b0;

   // m193_28 = W*in
   wire signed [14:0] m193_28;
   assign m193_28 =15'b0;

   // m193_29 = W*in
   wire signed [14:0] m193_29;
   assign m193_29 =15'b0;

   // m193_30 = W*in
   wire signed [14:0] m193_30;
   assign m193_30 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_31 = W*in
   wire signed [14:0] m193_31;
   assign m193_31 =15'b0;

   // m193_32 = W*in
   wire signed [14:0] m193_32;
   assign m193_32 =15'b0;

   // m193_33 = W*in
   wire signed [14:0] m193_33;
   assign m193_33 =15'b0;

   // m193_34 = W*in
   wire signed [14:0] m193_34;
   assign m193_34 =15'b0;

   // m193_35 = W*in
   wire signed [14:0] m193_35;
   assign m193_35 =15'b0;

   // m193_36 = W*in
   wire signed [14:0] m193_36;
   assign m193_36 =15'b0;

   // m193_37 = W*in
   wire signed [14:0] m193_37;
   assign m193_37 ={ {3{in193[14]}} , in193[14:3] };

   // m193_38 = W*in
   wire signed [14:0] m193_38;
   assign m193_38 =15'b0;

   // m193_39 = W*in
   wire signed [14:0] m193_39;
   assign m193_39 =15'b0;

   // m193_40 = W*in
   wire signed [14:0] m193_40;
   assign m193_40 =15'b0;

   // m193_41 = W*in
   wire signed [14:0] m193_41;
   assign m193_41 =15'b0;

   // m193_42 = W*in
   wire signed [14:0] m193_42;
   assign m193_42 =15'b0;

   // m193_43 = W*in
   wire signed [14:0] m193_43;
   assign m193_43 =15'b0;

   // m193_44 = W*in
   wire signed [14:0] m193_44;
   assign m193_44 =15'b0;

   // m193_45 = W*in
   wire signed [14:0] m193_45;
   assign m193_45 =15'b0;

   // m193_46 = W*in
   wire signed [14:0] m193_46;
   assign m193_46 =15'b0;

   // m193_47 = W*in
   wire signed [14:0] m193_47;
   assign m193_47 =15'b0;

   // m193_48 = W*in
   wire signed [14:0] m193_48;
   assign m193_48 ={ {3{in193[14]}} , in193[14:3] };

   // m193_49 = W*in
   wire signed [14:0] m193_49;
   assign m193_49 =15'b0;

   // m193_50 = W*in
   wire signed [14:0] m193_50;
   assign m193_50 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_51 = W*in
   wire signed [14:0] m193_51;
   assign m193_51 ={ {3{in193[14]}} , in193[14:3] };

   // m193_52 = W*in
   wire signed [14:0] m193_52;
   assign m193_52 =15'b0;

   // m193_53 = W*in
   wire signed [14:0] m193_53;
   assign m193_53 =15'b0;

   // m193_54 = W*in
   wire signed [14:0] m193_54;
   assign m193_54 =15'b0;

   // m193_55 = W*in
   wire signed [14:0] m193_55;
   assign m193_55 =15'b0;

   // m193_56 = W*in
   wire signed [14:0] m193_56;
   assign m193_56 =15'b0;

   // m193_57 = W*in
   wire signed [14:0] m193_57;
   assign m193_57 ={ {4{in193[14]}} , in193[14:4] };

   // m193_58 = W*in
   wire signed [14:0] m193_58;
   assign m193_58 ={ {3{in193[14]}} , in193[14:3] };

   // m193_59 = W*in
   wire signed [14:0] m193_59;
   assign m193_59 =15'b0;

   // m193_60 = W*in
   wire signed [14:0] m193_60;
   assign m193_60 =15'b0;

   // m193_61 = W*in
   wire signed [14:0] m193_61;
   assign m193_61 ={ {3{in193[14]}} , in193[14:3] };

   // m193_62 = W*in
   wire signed [14:0] m193_62;
   assign m193_62 =15'b0;

   // m193_63 = W*in
   wire signed [14:0] m193_63;
   assign m193_63 ={ {3{in193[14]}} , in193[14:3] };

   // m193_64 = W*in
   wire signed [14:0] m193_64;
   assign m193_64 =15'b0;

   // m193_65 = W*in
   wire signed [14:0] m193_65;
   assign m193_65 =15'b0;

   // m193_66 = W*in
   wire signed [14:0] m193_66;
   assign m193_66 =15'b0;

   // m193_67 = W*in
   wire signed [14:0] m193_67;
   assign m193_67 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_68 = W*in
   wire signed [14:0] m193_68;
   assign m193_68 ={ {3{in193[14]}} , in193[14:3] };

   // m193_69 = W*in
   wire signed [14:0] m193_69;
   assign m193_69 =15'b0;

   // m193_70 = W*in
   wire signed [14:0] m193_70;
   assign m193_70 =15'b0;

   // m193_71 = W*in
   wire signed [14:0] m193_71;
   assign m193_71 ={ {3{in193[14]}} , in193[14:3] };

   // m193_72 = W*in
   wire signed [14:0] m193_72;
   assign m193_72 =15'b0;

   // m193_73 = W*in
   wire signed [14:0] m193_73;
   assign m193_73 =15'b0;

   // m193_74 = W*in
   wire signed [14:0] m193_74;
   assign m193_74 =15'b0;

   // m193_75 = W*in
   wire signed [14:0] m193_75;
   assign m193_75 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_76 = W*in
   wire signed [14:0] m193_76;
   assign m193_76 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_77 = W*in
   wire signed [14:0] m193_77;
   assign m193_77 =15'b0;

   // m193_78 = W*in
   wire signed [14:0] m193_78;
   assign m193_78 =15'b0;

   // m193_79 = W*in
   wire signed [14:0] m193_79;
   assign m193_79 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_80 = W*in
   wire signed [14:0] m193_80;
   assign m193_80 =15'b0;

   // m193_81 = W*in
   wire signed [14:0] m193_81;
   assign m193_81 =15'b0;

   // m193_82 = W*in
   wire signed [14:0] m193_82;
   assign m193_82 =15'b0;

   // m193_83 = W*in
   wire signed [14:0] m193_83;
   assign m193_83 ={ {3{in193[14]}} , in193[14:3] };

   // m193_84 = W*in
   wire signed [14:0] m193_84;
   assign m193_84 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_85 = W*in
   wire signed [14:0] m193_85;
   assign m193_85 =15'b0;

   // m193_86 = W*in
   wire signed [14:0] m193_86;
   assign m193_86 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_87 = W*in
   wire signed [14:0] m193_87;
   assign m193_87 =15'b0;

   // m193_88 = W*in
   wire signed [14:0] m193_88;
   assign m193_88 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_89 = W*in
   wire signed [14:0] m193_89;
   assign m193_89 ={ {2{in193[14]}} , in193[14:2] };

   // m193_90 = W*in
   wire signed [14:0] m193_90;
   assign m193_90 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_91 = W*in
   wire signed [14:0] m193_91;
   assign m193_91 ={ {3{in193[14]}} , in193[14:3] };

   // m193_92 = W*in
   wire signed [14:0] m193_92;
   assign m193_92 =15'b0;

   // m193_93 = W*in
   wire signed [14:0] m193_93;
   assign m193_93 =15'b0;

   // m193_94 = W*in
   wire signed [14:0] m193_94;
   assign m193_94 =15'b0;

   // m193_95 = W*in
   wire signed [14:0] m193_95;
   assign m193_95 ={ {3{neg193[14]}} , neg193[14:3] };

   // m193_96 = W*in
   wire signed [14:0] m193_96;
   assign m193_96 =15'b0;

   // m193_97 = W*in
   wire signed [14:0] m193_97;
   assign m193_97 =15'b0;

   // m193_98 = W*in
   wire signed [14:0] m193_98;
   assign m193_98 =15'b0;

   // m193_99 = W*in
   wire signed [14:0] m193_99;
   assign m193_99 =15'b0;

   // m193_100 = W*in
   wire signed [14:0] m193_100;
   assign m193_100 ={ {3{in193[14]}} , in193[14:3] };

   // m194_1 = W*in
   wire signed [14:0] m194_1;
   assign m194_1 =15'b0;

   // m194_2 = W*in
   wire signed [14:0] m194_2;
   assign m194_2 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_3 = W*in
   wire signed [14:0] m194_3;
   assign m194_3 =15'b0;

   // m194_4 = W*in
   wire signed [14:0] m194_4;
   assign m194_4 =15'b0;

   // m194_5 = W*in
   wire signed [14:0] m194_5;
   assign m194_5 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_6 = W*in
   wire signed [14:0] m194_6;
   assign m194_6 ={ {3{in194[14]}} , in194[14:3] };

   // m194_7 = W*in
   wire signed [14:0] m194_7;
   assign m194_7 =15'b0;

   // m194_8 = W*in
   wire signed [14:0] m194_8;
   assign m194_8 ={ {3{in194[14]}} , in194[14:3] };

   // m194_9 = W*in
   wire signed [14:0] m194_9;
   assign m194_9 ={ {3{in194[14]}} , in194[14:3] };

   // m194_10 = W*in
   wire signed [14:0] m194_10;
   assign m194_10 =15'b0;

   // m194_11 = W*in
   wire signed [14:0] m194_11;
   assign m194_11 =15'b0;

   // m194_12 = W*in
   wire signed [14:0] m194_12;
   assign m194_12 =15'b0;

   // m194_13 = W*in
   wire signed [14:0] m194_13;
   assign m194_13 =15'b0;

   // m194_14 = W*in
   wire signed [14:0] m194_14;
   assign m194_14 =15'b0;

   // m194_15 = W*in
   wire signed [14:0] m194_15;
   assign m194_15 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_16 = W*in
   wire signed [14:0] m194_16;
   assign m194_16 =15'b0;

   // m194_17 = W*in
   wire signed [14:0] m194_17;
   assign m194_17 =15'b0;

   // m194_18 = W*in
   wire signed [14:0] m194_18;
   assign m194_18 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_19 = W*in
   wire signed [14:0] m194_19;
   assign m194_19 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_20 = W*in
   wire signed [14:0] m194_20;
   assign m194_20 =15'b0;

   // m194_21 = W*in
   wire signed [14:0] m194_21;
   assign m194_21 =15'b0;

   // m194_22 = W*in
   wire signed [14:0] m194_22;
   assign m194_22 =15'b0;

   // m194_23 = W*in
   wire signed [14:0] m194_23;
   assign m194_23 =15'b0;

   // m194_24 = W*in
   wire signed [14:0] m194_24;
   assign m194_24 =15'b0;

   // m194_25 = W*in
   wire signed [14:0] m194_25;
   assign m194_25 ={ {3{in194[14]}} , in194[14:3] };

   // m194_26 = W*in
   wire signed [14:0] m194_26;
   assign m194_26 =15'b0;

   // m194_27 = W*in
   wire signed [14:0] m194_27;
   assign m194_27 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_28 = W*in
   wire signed [14:0] m194_28;
   assign m194_28 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_29 = W*in
   wire signed [14:0] m194_29;
   assign m194_29 ={ {3{in194[14]}} , in194[14:3] };

   // m194_30 = W*in
   wire signed [14:0] m194_30;
   assign m194_30 =15'b0;

   // m194_31 = W*in
   wire signed [14:0] m194_31;
   assign m194_31 ={ {3{in194[14]}} , in194[14:3] };

   // m194_32 = W*in
   wire signed [14:0] m194_32;
   assign m194_32 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_33 = W*in
   wire signed [14:0] m194_33;
   assign m194_33 =15'b0;

   // m194_34 = W*in
   wire signed [14:0] m194_34;
   assign m194_34 ={ {3{in194[14]}} , in194[14:3] };

   // m194_35 = W*in
   wire signed [14:0] m194_35;
   assign m194_35 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_36 = W*in
   wire signed [14:0] m194_36;
   assign m194_36 =15'b0;

   // m194_37 = W*in
   wire signed [14:0] m194_37;
   assign m194_37 =15'b0;

   // m194_38 = W*in
   wire signed [14:0] m194_38;
   assign m194_38 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_39 = W*in
   wire signed [14:0] m194_39;
   assign m194_39 =15'b0;

   // m194_40 = W*in
   wire signed [14:0] m194_40;
   assign m194_40 =15'b0;

   // m194_41 = W*in
   wire signed [14:0] m194_41;
   assign m194_41 =15'b0;

   // m194_42 = W*in
   wire signed [14:0] m194_42;
   assign m194_42 =15'b0;

   // m194_43 = W*in
   wire signed [14:0] m194_43;
   assign m194_43 =15'b0;

   // m194_44 = W*in
   wire signed [14:0] m194_44;
   assign m194_44 =15'b0;

   // m194_45 = W*in
   wire signed [14:0] m194_45;
   assign m194_45 =15'b0;

   // m194_46 = W*in
   wire signed [14:0] m194_46;
   assign m194_46 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_47 = W*in
   wire signed [14:0] m194_47;
   assign m194_47 ={ {3{in194[14]}} , in194[14:3] };

   // m194_48 = W*in
   wire signed [14:0] m194_48;
   assign m194_48 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_49 = W*in
   wire signed [14:0] m194_49;
   assign m194_49 =15'b0;

   // m194_50 = W*in
   wire signed [14:0] m194_50;
   assign m194_50 =15'b0;

   // m194_51 = W*in
   wire signed [14:0] m194_51;
   assign m194_51 =15'b0;

   // m194_52 = W*in
   wire signed [14:0] m194_52;
   assign m194_52 ={ {3{in194[14]}} , in194[14:3] };

   // m194_53 = W*in
   wire signed [14:0] m194_53;
   assign m194_53 =15'b0;

   // m194_54 = W*in
   wire signed [14:0] m194_54;
   assign m194_54 =15'b0;

   // m194_55 = W*in
   wire signed [14:0] m194_55;
   assign m194_55 =15'b0;

   // m194_56 = W*in
   wire signed [14:0] m194_56;
   assign m194_56 =15'b0;

   // m194_57 = W*in
   wire signed [14:0] m194_57;
   assign m194_57 =15'b0;

   // m194_58 = W*in
   wire signed [14:0] m194_58;
   assign m194_58 ={ {3{in194[14]}} , in194[14:3] };

   // m194_59 = W*in
   wire signed [14:0] m194_59;
   assign m194_59 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_60 = W*in
   wire signed [14:0] m194_60;
   assign m194_60 ={ {3{in194[14]}} , in194[14:3] };

   // m194_61 = W*in
   wire signed [14:0] m194_61;
   assign m194_61 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_62 = W*in
   wire signed [14:0] m194_62;
   assign m194_62 =15'b0;

   // m194_63 = W*in
   wire signed [14:0] m194_63;
   assign m194_63 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_64 = W*in
   wire signed [14:0] m194_64;
   assign m194_64 =15'b0;

   // m194_65 = W*in
   wire signed [14:0] m194_65;
   assign m194_65 =15'b0;

   // m194_66 = W*in
   wire signed [14:0] m194_66;
   assign m194_66 =15'b0;

   // m194_67 = W*in
   wire signed [14:0] m194_67;
   assign m194_67 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_68 = W*in
   wire signed [14:0] m194_68;
   assign m194_68 ={ {4{neg194[14]}} , neg194[14:4] };

   // m194_69 = W*in
   wire signed [14:0] m194_69;
   assign m194_69 =15'b0;

   // m194_70 = W*in
   wire signed [14:0] m194_70;
   assign m194_70 =15'b0;

   // m194_71 = W*in
   wire signed [14:0] m194_71;
   assign m194_71 =15'b0;

   // m194_72 = W*in
   wire signed [14:0] m194_72;
   assign m194_72 =15'b0;

   // m194_73 = W*in
   wire signed [14:0] m194_73;
   assign m194_73 =15'b0;

   // m194_74 = W*in
   wire signed [14:0] m194_74;
   assign m194_74 =15'b0;

   // m194_75 = W*in
   wire signed [14:0] m194_75;
   assign m194_75 =15'b0;

   // m194_76 = W*in
   wire signed [14:0] m194_76;
   assign m194_76 =15'b0;

   // m194_77 = W*in
   wire signed [14:0] m194_77;
   assign m194_77 =15'b0;

   // m194_78 = W*in
   wire signed [14:0] m194_78;
   assign m194_78 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_79 = W*in
   wire signed [14:0] m194_79;
   assign m194_79 ={ {3{in194[14]}} , in194[14:3] };

   // m194_80 = W*in
   wire signed [14:0] m194_80;
   assign m194_80 ={ {2{in194[14]}} , in194[14:2] };

   // m194_81 = W*in
   wire signed [14:0] m194_81;
   assign m194_81 =15'b0;

   // m194_82 = W*in
   wire signed [14:0] m194_82;
   assign m194_82 =15'b0;

   // m194_83 = W*in
   wire signed [14:0] m194_83;
   assign m194_83 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_84 = W*in
   wire signed [14:0] m194_84;
   assign m194_84 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_85 = W*in
   wire signed [14:0] m194_85;
   assign m194_85 =15'b0;

   // m194_86 = W*in
   wire signed [14:0] m194_86;
   assign m194_86 =15'b0;

   // m194_87 = W*in
   wire signed [14:0] m194_87;
   assign m194_87 =15'b0;

   // m194_88 = W*in
   wire signed [14:0] m194_88;
   assign m194_88 =15'b0;

   // m194_89 = W*in
   wire signed [14:0] m194_89;
   assign m194_89 =15'b0;

   // m194_90 = W*in
   wire signed [14:0] m194_90;
   assign m194_90 =15'b0;

   // m194_91 = W*in
   wire signed [14:0] m194_91;
   assign m194_91 =15'b0;

   // m194_92 = W*in
   wire signed [14:0] m194_92;
   assign m194_92 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_93 = W*in
   wire signed [14:0] m194_93;
   assign m194_93 =15'b0;

   // m194_94 = W*in
   wire signed [14:0] m194_94;
   assign m194_94 =15'b0;

   // m194_95 = W*in
   wire signed [14:0] m194_95;
   assign m194_95 =15'b0;

   // m194_96 = W*in
   wire signed [14:0] m194_96;
   assign m194_96 ={ {3{in194[14]}} , in194[14:3] };

   // m194_97 = W*in
   wire signed [14:0] m194_97;
   assign m194_97 ={ {3{neg194[14]}} , neg194[14:3] };

   // m194_98 = W*in
   wire signed [14:0] m194_98;
   assign m194_98 =15'b0;

   // m194_99 = W*in
   wire signed [14:0] m194_99;
   assign m194_99 ={ {3{in194[14]}} , in194[14:3] };

   // m194_100 = W*in
   wire signed [14:0] m194_100;
   assign m194_100 =15'b0;

   // m195_1 = W*in
   wire signed [14:0] m195_1;
   assign m195_1 =15'b0;

   // m195_2 = W*in
   wire signed [14:0] m195_2;
   assign m195_2 =15'b0;

   // m195_3 = W*in
   wire signed [14:0] m195_3;
   assign m195_3 =15'b0;

   // m195_4 = W*in
   wire signed [14:0] m195_4;
   assign m195_4 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_5 = W*in
   wire signed [14:0] m195_5;
   assign m195_5 =15'b0;

   // m195_6 = W*in
   wire signed [14:0] m195_6;
   assign m195_6 =15'b0;

   // m195_7 = W*in
   wire signed [14:0] m195_7;
   assign m195_7 =15'b0;

   // m195_8 = W*in
   wire signed [14:0] m195_8;
   assign m195_8 =15'b0;

   // m195_9 = W*in
   wire signed [14:0] m195_9;
   assign m195_9 =15'b0;

   // m195_10 = W*in
   wire signed [14:0] m195_10;
   assign m195_10 =15'b0;

   // m195_11 = W*in
   wire signed [14:0] m195_11;
   assign m195_11 =15'b0;

   // m195_12 = W*in
   wire signed [14:0] m195_12;
   assign m195_12 =15'b0;

   // m195_13 = W*in
   wire signed [14:0] m195_13;
   assign m195_13 =15'b0;

   // m195_14 = W*in
   wire signed [14:0] m195_14;
   assign m195_14 =15'b0;

   // m195_15 = W*in
   wire signed [14:0] m195_15;
   assign m195_15 =15'b0;

   // m195_16 = W*in
   wire signed [14:0] m195_16;
   assign m195_16 =15'b0;

   // m195_17 = W*in
   wire signed [14:0] m195_17;
   assign m195_17 =15'b0;

   // m195_18 = W*in
   wire signed [14:0] m195_18;
   assign m195_18 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_19 = W*in
   wire signed [14:0] m195_19;
   assign m195_19 ={ {4{in195[14]}} , in195[14:4] };

   // m195_20 = W*in
   wire signed [14:0] m195_20;
   assign m195_20 =15'b0;

   // m195_21 = W*in
   wire signed [14:0] m195_21;
   assign m195_21 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_22 = W*in
   wire signed [14:0] m195_22;
   assign m195_22 =15'b0;

   // m195_23 = W*in
   wire signed [14:0] m195_23;
   assign m195_23 =15'b0;

   // m195_24 = W*in
   wire signed [14:0] m195_24;
   assign m195_24 =15'b0;

   // m195_25 = W*in
   wire signed [14:0] m195_25;
   assign m195_25 =15'b0;

   // m195_26 = W*in
   wire signed [14:0] m195_26;
   assign m195_26 =15'b0;

   // m195_27 = W*in
   wire signed [14:0] m195_27;
   assign m195_27 =15'b0;

   // m195_28 = W*in
   wire signed [14:0] m195_28;
   assign m195_28 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_29 = W*in
   wire signed [14:0] m195_29;
   assign m195_29 =15'b0;

   // m195_30 = W*in
   wire signed [14:0] m195_30;
   assign m195_30 =15'b0;

   // m195_31 = W*in
   wire signed [14:0] m195_31;
   assign m195_31 =15'b0;

   // m195_32 = W*in
   wire signed [14:0] m195_32;
   assign m195_32 =15'b0;

   // m195_33 = W*in
   wire signed [14:0] m195_33;
   assign m195_33 ={ {4{in195[14]}} , in195[14:4] };

   // m195_34 = W*in
   wire signed [14:0] m195_34;
   assign m195_34 =15'b0;

   // m195_35 = W*in
   wire signed [14:0] m195_35;
   assign m195_35 =15'b0;

   // m195_36 = W*in
   wire signed [14:0] m195_36;
   assign m195_36 =15'b0;

   // m195_37 = W*in
   wire signed [14:0] m195_37;
   assign m195_37 =15'b0;

   // m195_38 = W*in
   wire signed [14:0] m195_38;
   assign m195_38 =15'b0;

   // m195_39 = W*in
   wire signed [14:0] m195_39;
   assign m195_39 =15'b0;

   // m195_40 = W*in
   wire signed [14:0] m195_40;
   assign m195_40 =15'b0;

   // m195_41 = W*in
   wire signed [14:0] m195_41;
   assign m195_41 ={ {3{neg195[14]}} , neg195[14:3] };

   // m195_42 = W*in
   wire signed [14:0] m195_42;
   assign m195_42 =15'b0;

   // m195_43 = W*in
   wire signed [14:0] m195_43;
   assign m195_43 =15'b0;

   // m195_44 = W*in
   wire signed [14:0] m195_44;
   assign m195_44 =15'b0;

   // m195_45 = W*in
   wire signed [14:0] m195_45;
   assign m195_45 =15'b0;

   // m195_46 = W*in
   wire signed [14:0] m195_46;
   assign m195_46 =15'b0;

   // m195_47 = W*in
   wire signed [14:0] m195_47;
   assign m195_47 =15'b0;

   // m195_48 = W*in
   wire signed [14:0] m195_48;
   assign m195_48 =15'b0;

   // m195_49 = W*in
   wire signed [14:0] m195_49;
   assign m195_49 =15'b0;

   // m195_50 = W*in
   wire signed [14:0] m195_50;
   assign m195_50 =15'b0;

   // m195_51 = W*in
   wire signed [14:0] m195_51;
   assign m195_51 =15'b0;

   // m195_52 = W*in
   wire signed [14:0] m195_52;
   assign m195_52 =15'b0;

   // m195_53 = W*in
   wire signed [14:0] m195_53;
   assign m195_53 =15'b0;

   // m195_54 = W*in
   wire signed [14:0] m195_54;
   assign m195_54 =15'b0;

   // m195_55 = W*in
   wire signed [14:0] m195_55;
   assign m195_55 =15'b0;

   // m195_56 = W*in
   wire signed [14:0] m195_56;
   assign m195_56 =15'b0;

   // m195_57 = W*in
   wire signed [14:0] m195_57;
   assign m195_57 =15'b0;

   // m195_58 = W*in
   wire signed [14:0] m195_58;
   assign m195_58 =15'b0;

   // m195_59 = W*in
   wire signed [14:0] m195_59;
   assign m195_59 ={ {4{in195[14]}} , in195[14:4] };

   // m195_60 = W*in
   wire signed [14:0] m195_60;
   assign m195_60 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_61 = W*in
   wire signed [14:0] m195_61;
   assign m195_61 =15'b0;

   // m195_62 = W*in
   wire signed [14:0] m195_62;
   assign m195_62 =15'b0;

   // m195_63 = W*in
   wire signed [14:0] m195_63;
   assign m195_63 ={ {3{in195[14]}} , in195[14:3] };

   // m195_64 = W*in
   wire signed [14:0] m195_64;
   assign m195_64 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_65 = W*in
   wire signed [14:0] m195_65;
   assign m195_65 =15'b0;

   // m195_66 = W*in
   wire signed [14:0] m195_66;
   assign m195_66 ={ {4{in195[14]}} , in195[14:4] };

   // m195_67 = W*in
   wire signed [14:0] m195_67;
   assign m195_67 =15'b0;

   // m195_68 = W*in
   wire signed [14:0] m195_68;
   assign m195_68 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_69 = W*in
   wire signed [14:0] m195_69;
   assign m195_69 =15'b0;

   // m195_70 = W*in
   wire signed [14:0] m195_70;
   assign m195_70 =15'b0;

   // m195_71 = W*in
   wire signed [14:0] m195_71;
   assign m195_71 =15'b0;

   // m195_72 = W*in
   wire signed [14:0] m195_72;
   assign m195_72 =15'b0;

   // m195_73 = W*in
   wire signed [14:0] m195_73;
   assign m195_73 =15'b0;

   // m195_74 = W*in
   wire signed [14:0] m195_74;
   assign m195_74 =15'b0;

   // m195_75 = W*in
   wire signed [14:0] m195_75;
   assign m195_75 =15'b0;

   // m195_76 = W*in
   wire signed [14:0] m195_76;
   assign m195_76 =15'b0;

   // m195_77 = W*in
   wire signed [14:0] m195_77;
   assign m195_77 =15'b0;

   // m195_78 = W*in
   wire signed [14:0] m195_78;
   assign m195_78 ={ {3{neg195[14]}} , neg195[14:3] };

   // m195_79 = W*in
   wire signed [14:0] m195_79;
   assign m195_79 =15'b0;

   // m195_80 = W*in
   wire signed [14:0] m195_80;
   assign m195_80 =15'b0;

   // m195_81 = W*in
   wire signed [14:0] m195_81;
   assign m195_81 =15'b0;

   // m195_82 = W*in
   wire signed [14:0] m195_82;
   assign m195_82 =15'b0;

   // m195_83 = W*in
   wire signed [14:0] m195_83;
   assign m195_83 =15'b0;

   // m195_84 = W*in
   wire signed [14:0] m195_84;
   assign m195_84 =15'b0;

   // m195_85 = W*in
   wire signed [14:0] m195_85;
   assign m195_85 =15'b0;

   // m195_86 = W*in
   wire signed [14:0] m195_86;
   assign m195_86 =15'b0;

   // m195_87 = W*in
   wire signed [14:0] m195_87;
   assign m195_87 =15'b0;

   // m195_88 = W*in
   wire signed [14:0] m195_88;
   assign m195_88 =15'b0;

   // m195_89 = W*in
   wire signed [14:0] m195_89;
   assign m195_89 =15'b0;

   // m195_90 = W*in
   wire signed [14:0] m195_90;
   assign m195_90 =15'b0;

   // m195_91 = W*in
   wire signed [14:0] m195_91;
   assign m195_91 =15'b0;

   // m195_92 = W*in
   wire signed [14:0] m195_92;
   assign m195_92 =15'b0;

   // m195_93 = W*in
   wire signed [14:0] m195_93;
   assign m195_93 =15'b0;

   // m195_94 = W*in
   wire signed [14:0] m195_94;
   assign m195_94 =15'b0;

   // m195_95 = W*in
   wire signed [14:0] m195_95;
   assign m195_95 =15'b0;

   // m195_96 = W*in
   wire signed [14:0] m195_96;
   assign m195_96 ={ {4{neg195[14]}} , neg195[14:4] };

   // m195_97 = W*in
   wire signed [14:0] m195_97;
   assign m195_97 =15'b0;

   // m195_98 = W*in
   wire signed [14:0] m195_98;
   assign m195_98 =15'b0;

   // m195_99 = W*in
   wire signed [14:0] m195_99;
   assign m195_99 =15'b0;

   // m195_100 = W*in
   wire signed [14:0] m195_100;
   assign m195_100 =15'b0;

   // m196_1 = W*in
   wire signed [14:0] m196_1;
   assign m196_1 =15'b0;

   // m196_2 = W*in
   wire signed [14:0] m196_2;
   assign m196_2 =15'b0;

   // m196_3 = W*in
   wire signed [14:0] m196_3;
   assign m196_3 =15'b0;

   // m196_4 = W*in
   wire signed [14:0] m196_4;
   assign m196_4 ={ {4{in196[14]}} , in196[14:4] };

   // m196_5 = W*in
   wire signed [14:0] m196_5;
   assign m196_5 =15'b0;

   // m196_6 = W*in
   wire signed [14:0] m196_6;
   assign m196_6 =15'b0;

   // m196_7 = W*in
   wire signed [14:0] m196_7;
   assign m196_7 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_8 = W*in
   wire signed [14:0] m196_8;
   assign m196_8 =15'b0;

   // m196_9 = W*in
   wire signed [14:0] m196_9;
   assign m196_9 =15'b0;

   // m196_10 = W*in
   wire signed [14:0] m196_10;
   assign m196_10 =15'b0;

   // m196_11 = W*in
   wire signed [14:0] m196_11;
   assign m196_11 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_12 = W*in
   wire signed [14:0] m196_12;
   assign m196_12 =15'b0;

   // m196_13 = W*in
   wire signed [14:0] m196_13;
   assign m196_13 =15'b0;

   // m196_14 = W*in
   wire signed [14:0] m196_14;
   assign m196_14 =15'b0;

   // m196_15 = W*in
   wire signed [14:0] m196_15;
   assign m196_15 =15'b0;

   // m196_16 = W*in
   wire signed [14:0] m196_16;
   assign m196_16 =15'b0;

   // m196_17 = W*in
   wire signed [14:0] m196_17;
   assign m196_17 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_18 = W*in
   wire signed [14:0] m196_18;
   assign m196_18 =15'b0;

   // m196_19 = W*in
   wire signed [14:0] m196_19;
   assign m196_19 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_20 = W*in
   wire signed [14:0] m196_20;
   assign m196_20 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_21 = W*in
   wire signed [14:0] m196_21;
   assign m196_21 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_22 = W*in
   wire signed [14:0] m196_22;
   assign m196_22 ={ {3{in196[14]}} , in196[14:3] };

   // m196_23 = W*in
   wire signed [14:0] m196_23;
   assign m196_23 =15'b0;

   // m196_24 = W*in
   wire signed [14:0] m196_24;
   assign m196_24 =15'b0;

   // m196_25 = W*in
   wire signed [14:0] m196_25;
   assign m196_25 =15'b0;

   // m196_26 = W*in
   wire signed [14:0] m196_26;
   assign m196_26 ={ {3{in196[14]}} , in196[14:3] };

   // m196_27 = W*in
   wire signed [14:0] m196_27;
   assign m196_27 =15'b0;

   // m196_28 = W*in
   wire signed [14:0] m196_28;
   assign m196_28 =15'b0;

   // m196_29 = W*in
   wire signed [14:0] m196_29;
   assign m196_29 =15'b0;

   // m196_30 = W*in
   wire signed [14:0] m196_30;
   assign m196_30 =15'b0;

   // m196_31 = W*in
   wire signed [14:0] m196_31;
   assign m196_31 =15'b0;

   // m196_32 = W*in
   wire signed [14:0] m196_32;
   assign m196_32 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_33 = W*in
   wire signed [14:0] m196_33;
   assign m196_33 =15'b0;

   // m196_34 = W*in
   wire signed [14:0] m196_34;
   assign m196_34 =15'b0;

   // m196_35 = W*in
   wire signed [14:0] m196_35;
   assign m196_35 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_36 = W*in
   wire signed [14:0] m196_36;
   assign m196_36 =15'b0;

   // m196_37 = W*in
   wire signed [14:0] m196_37;
   assign m196_37 =15'b0;

   // m196_38 = W*in
   wire signed [14:0] m196_38;
   assign m196_38 =15'b0;

   // m196_39 = W*in
   wire signed [14:0] m196_39;
   assign m196_39 =15'b0;

   // m196_40 = W*in
   wire signed [14:0] m196_40;
   assign m196_40 =15'b0;

   // m196_41 = W*in
   wire signed [14:0] m196_41;
   assign m196_41 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_42 = W*in
   wire signed [14:0] m196_42;
   assign m196_42 =15'b0;

   // m196_43 = W*in
   wire signed [14:0] m196_43;
   assign m196_43 =15'b0;

   // m196_44 = W*in
   wire signed [14:0] m196_44;
   assign m196_44 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_45 = W*in
   wire signed [14:0] m196_45;
   assign m196_45 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_46 = W*in
   wire signed [14:0] m196_46;
   assign m196_46 =15'b0;

   // m196_47 = W*in
   wire signed [14:0] m196_47;
   assign m196_47 =15'b0;

   // m196_48 = W*in
   wire signed [14:0] m196_48;
   assign m196_48 =15'b0;

   // m196_49 = W*in
   wire signed [14:0] m196_49;
   assign m196_49 =15'b0;

   // m196_50 = W*in
   wire signed [14:0] m196_50;
   assign m196_50 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_51 = W*in
   wire signed [14:0] m196_51;
   assign m196_51 =15'b0;

   // m196_52 = W*in
   wire signed [14:0] m196_52;
   assign m196_52 =15'b0;

   // m196_53 = W*in
   wire signed [14:0] m196_53;
   assign m196_53 =15'b0;

   // m196_54 = W*in
   wire signed [14:0] m196_54;
   assign m196_54 =15'b0;

   // m196_55 = W*in
   wire signed [14:0] m196_55;
   assign m196_55 =15'b0;

   // m196_56 = W*in
   wire signed [14:0] m196_56;
   assign m196_56 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_57 = W*in
   wire signed [14:0] m196_57;
   assign m196_57 ={ {3{in196[14]}} , in196[14:3] };

   // m196_58 = W*in
   wire signed [14:0] m196_58;
   assign m196_58 =15'b0;

   // m196_59 = W*in
   wire signed [14:0] m196_59;
   assign m196_59 =15'b0;

   // m196_60 = W*in
   wire signed [14:0] m196_60;
   assign m196_60 =15'b0;

   // m196_61 = W*in
   wire signed [14:0] m196_61;
   assign m196_61 ={ {4{in196[14]}} , in196[14:4] };

   // m196_62 = W*in
   wire signed [14:0] m196_62;
   assign m196_62 ={ {3{in196[14]}} , in196[14:3] };

   // m196_63 = W*in
   wire signed [14:0] m196_63;
   assign m196_63 ={ {3{in196[14]}} , in196[14:3] };

   // m196_64 = W*in
   wire signed [14:0] m196_64;
   assign m196_64 =15'b0;

   // m196_65 = W*in
   wire signed [14:0] m196_65;
   assign m196_65 =15'b0;

   // m196_66 = W*in
   wire signed [14:0] m196_66;
   assign m196_66 =15'b0;

   // m196_67 = W*in
   wire signed [14:0] m196_67;
   assign m196_67 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_68 = W*in
   wire signed [14:0] m196_68;
   assign m196_68 =15'b0;

   // m196_69 = W*in
   wire signed [14:0] m196_69;
   assign m196_69 ={ {4{neg196[14]}} , neg196[14:4] };

   // m196_70 = W*in
   wire signed [14:0] m196_70;
   assign m196_70 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_71 = W*in
   wire signed [14:0] m196_71;
   assign m196_71 =15'b0;

   // m196_72 = W*in
   wire signed [14:0] m196_72;
   assign m196_72 =15'b0;

   // m196_73 = W*in
   wire signed [14:0] m196_73;
   assign m196_73 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_74 = W*in
   wire signed [14:0] m196_74;
   assign m196_74 ={ {4{neg196[14]}} , neg196[14:4] };

   // m196_75 = W*in
   wire signed [14:0] m196_75;
   assign m196_75 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_76 = W*in
   wire signed [14:0] m196_76;
   assign m196_76 =15'b0;

   // m196_77 = W*in
   wire signed [14:0] m196_77;
   assign m196_77 =15'b0;

   // m196_78 = W*in
   wire signed [14:0] m196_78;
   assign m196_78 =15'b0;

   // m196_79 = W*in
   wire signed [14:0] m196_79;
   assign m196_79 =15'b0;

   // m196_80 = W*in
   wire signed [14:0] m196_80;
   assign m196_80 ={ {4{in196[14]}} , in196[14:4] };

   // m196_81 = W*in
   wire signed [14:0] m196_81;
   assign m196_81 =15'b0;

   // m196_82 = W*in
   wire signed [14:0] m196_82;
   assign m196_82 =15'b0;

   // m196_83 = W*in
   wire signed [14:0] m196_83;
   assign m196_83 =15'b0;

   // m196_84 = W*in
   wire signed [14:0] m196_84;
   assign m196_84 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_85 = W*in
   wire signed [14:0] m196_85;
   assign m196_85 =15'b0;

   // m196_86 = W*in
   wire signed [14:0] m196_86;
   assign m196_86 =15'b0;

   // m196_87 = W*in
   wire signed [14:0] m196_87;
   assign m196_87 =15'b0;

   // m196_88 = W*in
   wire signed [14:0] m196_88;
   assign m196_88 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_89 = W*in
   wire signed [14:0] m196_89;
   assign m196_89 =15'b0;

   // m196_90 = W*in
   wire signed [14:0] m196_90;
   assign m196_90 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_91 = W*in
   wire signed [14:0] m196_91;
   assign m196_91 ={ {3{in196[14]}} , in196[14:3] };

   // m196_92 = W*in
   wire signed [14:0] m196_92;
   assign m196_92 ={ {3{in196[14]}} , in196[14:3] };

   // m196_93 = W*in
   wire signed [14:0] m196_93;
   assign m196_93 ={ {3{in196[14]}} , in196[14:3] };

   // m196_94 = W*in
   wire signed [14:0] m196_94;
   assign m196_94 =15'b0;

   // m196_95 = W*in
   wire signed [14:0] m196_95;
   assign m196_95 ={ {3{neg196[14]}} , neg196[14:3] };

   // m196_96 = W*in
   wire signed [14:0] m196_96;
   assign m196_96 =15'b0;

   // m196_97 = W*in
   wire signed [14:0] m196_97;
   assign m196_97 =15'b0;

   // m196_98 = W*in
   wire signed [14:0] m196_98;
   assign m196_98 ={ {2{neg196[14]}} , neg196[14:2] };

   // m196_99 = W*in
   wire signed [14:0] m196_99;
   assign m196_99 =15'b0;

   // m196_100 = W*in
   wire signed [14:0] m196_100;
   assign m196_100 ={ {3{in196[14]}} , in196[14:3] };

   // m197_1 = W*in
   wire signed [14:0] m197_1;
   assign m197_1 =15'b0;

   // m197_2 = W*in
   wire signed [14:0] m197_2;
   assign m197_2 =15'b0;

   // m197_3 = W*in
   wire signed [14:0] m197_3;
   assign m197_3 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_4 = W*in
   wire signed [14:0] m197_4;
   assign m197_4 =15'b0;

   // m197_5 = W*in
   wire signed [14:0] m197_5;
   assign m197_5 ={ {4{in197[14]}} , in197[14:4] };

   // m197_6 = W*in
   wire signed [14:0] m197_6;
   assign m197_6 =15'b0;

   // m197_7 = W*in
   wire signed [14:0] m197_7;
   assign m197_7 =15'b0;

   // m197_8 = W*in
   wire signed [14:0] m197_8;
   assign m197_8 =15'b0;

   // m197_9 = W*in
   wire signed [14:0] m197_9;
   assign m197_9 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_10 = W*in
   wire signed [14:0] m197_10;
   assign m197_10 ={ {3{in197[14]}} , in197[14:3] };

   // m197_11 = W*in
   wire signed [14:0] m197_11;
   assign m197_11 =15'b0;

   // m197_12 = W*in
   wire signed [14:0] m197_12;
   assign m197_12 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_13 = W*in
   wire signed [14:0] m197_13;
   assign m197_13 =15'b0;

   // m197_14 = W*in
   wire signed [14:0] m197_14;
   assign m197_14 =15'b0;

   // m197_15 = W*in
   wire signed [14:0] m197_15;
   assign m197_15 ={ {3{in197[14]}} , in197[14:3] };

   // m197_16 = W*in
   wire signed [14:0] m197_16;
   assign m197_16 ={ {3{in197[14]}} , in197[14:3] };

   // m197_17 = W*in
   wire signed [14:0] m197_17;
   assign m197_17 =15'b0;

   // m197_18 = W*in
   wire signed [14:0] m197_18;
   assign m197_18 ={ {3{in197[14]}} , in197[14:3] };

   // m197_19 = W*in
   wire signed [14:0] m197_19;
   assign m197_19 =15'b0;

   // m197_20 = W*in
   wire signed [14:0] m197_20;
   assign m197_20 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_21 = W*in
   wire signed [14:0] m197_21;
   assign m197_21 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_22 = W*in
   wire signed [14:0] m197_22;
   assign m197_22 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_23 = W*in
   wire signed [14:0] m197_23;
   assign m197_23 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_24 = W*in
   wire signed [14:0] m197_24;
   assign m197_24 =15'b0;

   // m197_25 = W*in
   wire signed [14:0] m197_25;
   assign m197_25 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_26 = W*in
   wire signed [14:0] m197_26;
   assign m197_26 =15'b0;

   // m197_27 = W*in
   wire signed [14:0] m197_27;
   assign m197_27 =15'b0;

   // m197_28 = W*in
   wire signed [14:0] m197_28;
   assign m197_28 =15'b0;

   // m197_29 = W*in
   wire signed [14:0] m197_29;
   assign m197_29 =15'b0;

   // m197_30 = W*in
   wire signed [14:0] m197_30;
   assign m197_30 ={ {3{in197[14]}} , in197[14:3] };

   // m197_31 = W*in
   wire signed [14:0] m197_31;
   assign m197_31 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_32 = W*in
   wire signed [14:0] m197_32;
   assign m197_32 ={ {4{in197[14]}} , in197[14:4] };

   // m197_33 = W*in
   wire signed [14:0] m197_33;
   assign m197_33 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_34 = W*in
   wire signed [14:0] m197_34;
   assign m197_34 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_35 = W*in
   wire signed [14:0] m197_35;
   assign m197_35 =15'b0;

   // m197_36 = W*in
   wire signed [14:0] m197_36;
   assign m197_36 =15'b0;

   // m197_37 = W*in
   wire signed [14:0] m197_37;
   assign m197_37 =15'b0;

   // m197_38 = W*in
   wire signed [14:0] m197_38;
   assign m197_38 =15'b0;

   // m197_39 = W*in
   wire signed [14:0] m197_39;
   assign m197_39 =15'b0;

   // m197_40 = W*in
   wire signed [14:0] m197_40;
   assign m197_40 =15'b0;

   // m197_41 = W*in
   wire signed [14:0] m197_41;
   assign m197_41 =15'b0;

   // m197_42 = W*in
   wire signed [14:0] m197_42;
   assign m197_42 ={ {3{in197[14]}} , in197[14:3] };

   // m197_43 = W*in
   wire signed [14:0] m197_43;
   assign m197_43 ={ {3{in197[14]}} , in197[14:3] };

   // m197_44 = W*in
   wire signed [14:0] m197_44;
   assign m197_44 =15'b0;

   // m197_45 = W*in
   wire signed [14:0] m197_45;
   assign m197_45 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_46 = W*in
   wire signed [14:0] m197_46;
   assign m197_46 =15'b0;

   // m197_47 = W*in
   wire signed [14:0] m197_47;
   assign m197_47 =15'b0;

   // m197_48 = W*in
   wire signed [14:0] m197_48;
   assign m197_48 ={ {3{in197[14]}} , in197[14:3] };

   // m197_49 = W*in
   wire signed [14:0] m197_49;
   assign m197_49 =15'b0;

   // m197_50 = W*in
   wire signed [14:0] m197_50;
   assign m197_50 =15'b0;

   // m197_51 = W*in
   wire signed [14:0] m197_51;
   assign m197_51 =15'b0;

   // m197_52 = W*in
   wire signed [14:0] m197_52;
   assign m197_52 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_53 = W*in
   wire signed [14:0] m197_53;
   assign m197_53 =15'b0;

   // m197_54 = W*in
   wire signed [14:0] m197_54;
   assign m197_54 =15'b0;

   // m197_55 = W*in
   wire signed [14:0] m197_55;
   assign m197_55 =15'b0;

   // m197_56 = W*in
   wire signed [14:0] m197_56;
   assign m197_56 =15'b0;

   // m197_57 = W*in
   wire signed [14:0] m197_57;
   assign m197_57 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_58 = W*in
   wire signed [14:0] m197_58;
   assign m197_58 =15'b0;

   // m197_59 = W*in
   wire signed [14:0] m197_59;
   assign m197_59 ={ {4{neg197[14]}} , neg197[14:4] };

   // m197_60 = W*in
   wire signed [14:0] m197_60;
   assign m197_60 =15'b0;

   // m197_61 = W*in
   wire signed [14:0] m197_61;
   assign m197_61 ={ {3{in197[14]}} , in197[14:3] };

   // m197_62 = W*in
   wire signed [14:0] m197_62;
   assign m197_62 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_63 = W*in
   wire signed [14:0] m197_63;
   assign m197_63 ={ {3{in197[14]}} , in197[14:3] };

   // m197_64 = W*in
   wire signed [14:0] m197_64;
   assign m197_64 =15'b0;

   // m197_65 = W*in
   wire signed [14:0] m197_65;
   assign m197_65 ={ {3{in197[14]}} , in197[14:3] };

   // m197_66 = W*in
   wire signed [14:0] m197_66;
   assign m197_66 =15'b0;

   // m197_67 = W*in
   wire signed [14:0] m197_67;
   assign m197_67 ={ {3{in197[14]}} , in197[14:3] };

   // m197_68 = W*in
   wire signed [14:0] m197_68;
   assign m197_68 =15'b0;

   // m197_69 = W*in
   wire signed [14:0] m197_69;
   assign m197_69 ={ {4{in197[14]}} , in197[14:4] };

   // m197_70 = W*in
   wire signed [14:0] m197_70;
   assign m197_70 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_71 = W*in
   wire signed [14:0] m197_71;
   assign m197_71 =15'b0;

   // m197_72 = W*in
   wire signed [14:0] m197_72;
   assign m197_72 =15'b0;

   // m197_73 = W*in
   wire signed [14:0] m197_73;
   assign m197_73 =15'b0;

   // m197_74 = W*in
   wire signed [14:0] m197_74;
   assign m197_74 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_75 = W*in
   wire signed [14:0] m197_75;
   assign m197_75 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_76 = W*in
   wire signed [14:0] m197_76;
   assign m197_76 =15'b0;

   // m197_77 = W*in
   wire signed [14:0] m197_77;
   assign m197_77 =15'b0;

   // m197_78 = W*in
   wire signed [14:0] m197_78;
   assign m197_78 ={ {3{in197[14]}} , in197[14:3] };

   // m197_79 = W*in
   wire signed [14:0] m197_79;
   assign m197_79 =15'b0;

   // m197_80 = W*in
   wire signed [14:0] m197_80;
   assign m197_80 =15'b0;

   // m197_81 = W*in
   wire signed [14:0] m197_81;
   assign m197_81 =15'b0;

   // m197_82 = W*in
   wire signed [14:0] m197_82;
   assign m197_82 ={ {3{in197[14]}} , in197[14:3] };

   // m197_83 = W*in
   wire signed [14:0] m197_83;
   assign m197_83 =15'b0;

   // m197_84 = W*in
   wire signed [14:0] m197_84;
   assign m197_84 =15'b0;

   // m197_85 = W*in
   wire signed [14:0] m197_85;
   assign m197_85 =15'b0;

   // m197_86 = W*in
   wire signed [14:0] m197_86;
   assign m197_86 =15'b0;

   // m197_87 = W*in
   wire signed [14:0] m197_87;
   assign m197_87 =15'b0;

   // m197_88 = W*in
   wire signed [14:0] m197_88;
   assign m197_88 ={ {3{neg197[14]}} , neg197[14:3] };

   // m197_89 = W*in
   wire signed [14:0] m197_89;
   assign m197_89 =15'b0;

   // m197_90 = W*in
   wire signed [14:0] m197_90;
   assign m197_90 =15'b0;

   // m197_91 = W*in
   wire signed [14:0] m197_91;
   assign m197_91 =15'b0;

   // m197_92 = W*in
   wire signed [14:0] m197_92;
   assign m197_92 =15'b0;

   // m197_93 = W*in
   wire signed [14:0] m197_93;
   assign m197_93 =15'b0;

   // m197_94 = W*in
   wire signed [14:0] m197_94;
   assign m197_94 =15'b0;

   // m197_95 = W*in
   wire signed [14:0] m197_95;
   assign m197_95 =15'b0;

   // m197_96 = W*in
   wire signed [14:0] m197_96;
   assign m197_96 =15'b0;

   // m197_97 = W*in
   wire signed [14:0] m197_97;
   assign m197_97 =15'b0;

   // m197_98 = W*in
   wire signed [14:0] m197_98;
   assign m197_98 =15'b0;

   // m197_99 = W*in
   wire signed [14:0] m197_99;
   assign m197_99 =15'b0;

   // m197_100 = W*in
   wire signed [14:0] m197_100;
   assign m197_100 =15'b0;

   // m198_1 = W*in
   wire signed [14:0] m198_1;
   assign m198_1 =15'b0;

   // m198_2 = W*in
   wire signed [14:0] m198_2;
   assign m198_2 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_3 = W*in
   wire signed [14:0] m198_3;
   assign m198_3 =15'b0;

   // m198_4 = W*in
   wire signed [14:0] m198_4;
   assign m198_4 =15'b0;

   // m198_5 = W*in
   wire signed [14:0] m198_5;
   assign m198_5 =15'b0;

   // m198_6 = W*in
   wire signed [14:0] m198_6;
   assign m198_6 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_7 = W*in
   wire signed [14:0] m198_7;
   assign m198_7 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_8 = W*in
   wire signed [14:0] m198_8;
   assign m198_8 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_9 = W*in
   wire signed [14:0] m198_9;
   assign m198_9 =15'b0;

   // m198_10 = W*in
   wire signed [14:0] m198_10;
   assign m198_10 =15'b0;

   // m198_11 = W*in
   wire signed [14:0] m198_11;
   assign m198_11 =15'b0;

   // m198_12 = W*in
   wire signed [14:0] m198_12;
   assign m198_12 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_13 = W*in
   wire signed [14:0] m198_13;
   assign m198_13 =15'b0;

   // m198_14 = W*in
   wire signed [14:0] m198_14;
   assign m198_14 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_15 = W*in
   wire signed [14:0] m198_15;
   assign m198_15 =15'b0;

   // m198_16 = W*in
   wire signed [14:0] m198_16;
   assign m198_16 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_17 = W*in
   wire signed [14:0] m198_17;
   assign m198_17 =15'b0;

   // m198_18 = W*in
   wire signed [14:0] m198_18;
   assign m198_18 =15'b0;

   // m198_19 = W*in
   wire signed [14:0] m198_19;
   assign m198_19 ={ {4{in198[14]}} , in198[14:4] };

   // m198_20 = W*in
   wire signed [14:0] m198_20;
   assign m198_20 =15'b0;

   // m198_21 = W*in
   wire signed [14:0] m198_21;
   assign m198_21 ={ {3{in198[14]}} , in198[14:3] };

   // m198_22 = W*in
   wire signed [14:0] m198_22;
   assign m198_22 ={ {4{neg198[14]}} , neg198[14:4] };

   // m198_23 = W*in
   wire signed [14:0] m198_23;
   assign m198_23 =15'b0;

   // m198_24 = W*in
   wire signed [14:0] m198_24;
   assign m198_24 =15'b0;

   // m198_25 = W*in
   wire signed [14:0] m198_25;
   assign m198_25 ={ {4{neg198[14]}} , neg198[14:4] };

   // m198_26 = W*in
   wire signed [14:0] m198_26;
   assign m198_26 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_27 = W*in
   wire signed [14:0] m198_27;
   assign m198_27 ={ {4{neg198[14]}} , neg198[14:4] };

   // m198_28 = W*in
   wire signed [14:0] m198_28;
   assign m198_28 =15'b0;

   // m198_29 = W*in
   wire signed [14:0] m198_29;
   assign m198_29 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_30 = W*in
   wire signed [14:0] m198_30;
   assign m198_30 =15'b0;

   // m198_31 = W*in
   wire signed [14:0] m198_31;
   assign m198_31 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_32 = W*in
   wire signed [14:0] m198_32;
   assign m198_32 =15'b0;

   // m198_33 = W*in
   wire signed [14:0] m198_33;
   assign m198_33 ={ {4{neg198[14]}} , neg198[14:4] };

   // m198_34 = W*in
   wire signed [14:0] m198_34;
   assign m198_34 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_35 = W*in
   wire signed [14:0] m198_35;
   assign m198_35 =15'b0;

   // m198_36 = W*in
   wire signed [14:0] m198_36;
   assign m198_36 =15'b0;

   // m198_37 = W*in
   wire signed [14:0] m198_37;
   assign m198_37 =15'b0;

   // m198_38 = W*in
   wire signed [14:0] m198_38;
   assign m198_38 =15'b0;

   // m198_39 = W*in
   wire signed [14:0] m198_39;
   assign m198_39 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_40 = W*in
   wire signed [14:0] m198_40;
   assign m198_40 =15'b0;

   // m198_41 = W*in
   wire signed [14:0] m198_41;
   assign m198_41 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_42 = W*in
   wire signed [14:0] m198_42;
   assign m198_42 =15'b0;

   // m198_43 = W*in
   wire signed [14:0] m198_43;
   assign m198_43 =15'b0;

   // m198_44 = W*in
   wire signed [14:0] m198_44;
   assign m198_44 =15'b0;

   // m198_45 = W*in
   wire signed [14:0] m198_45;
   assign m198_45 =15'b0;

   // m198_46 = W*in
   wire signed [14:0] m198_46;
   assign m198_46 =15'b0;

   // m198_47 = W*in
   wire signed [14:0] m198_47;
   assign m198_47 =15'b0;

   // m198_48 = W*in
   wire signed [14:0] m198_48;
   assign m198_48 =15'b0;

   // m198_49 = W*in
   wire signed [14:0] m198_49;
   assign m198_49 =15'b0;

   // m198_50 = W*in
   wire signed [14:0] m198_50;
   assign m198_50 =15'b0;

   // m198_51 = W*in
   wire signed [14:0] m198_51;
   assign m198_51 =15'b0;

   // m198_52 = W*in
   wire signed [14:0] m198_52;
   assign m198_52 =15'b0;

   // m198_53 = W*in
   wire signed [14:0] m198_53;
   assign m198_53 =15'b0;

   // m198_54 = W*in
   wire signed [14:0] m198_54;
   assign m198_54 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_55 = W*in
   wire signed [14:0] m198_55;
   assign m198_55 =15'b0;

   // m198_56 = W*in
   wire signed [14:0] m198_56;
   assign m198_56 ={ {3{in198[14]}} , in198[14:3] };

   // m198_57 = W*in
   wire signed [14:0] m198_57;
   assign m198_57 ={ {3{in198[14]}} , in198[14:3] };

   // m198_58 = W*in
   wire signed [14:0] m198_58;
   assign m198_58 =15'b0;

   // m198_59 = W*in
   wire signed [14:0] m198_59;
   assign m198_59 ={ {3{in198[14]}} , in198[14:3] };

   // m198_60 = W*in
   wire signed [14:0] m198_60;
   assign m198_60 ={ {4{neg198[14]}} , neg198[14:4] };

   // m198_61 = W*in
   wire signed [14:0] m198_61;
   assign m198_61 ={ {3{in198[14]}} , in198[14:3] };

   // m198_62 = W*in
   wire signed [14:0] m198_62;
   assign m198_62 ={ {3{in198[14]}} , in198[14:3] };

   // m198_63 = W*in
   wire signed [14:0] m198_63;
   assign m198_63 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_64 = W*in
   wire signed [14:0] m198_64;
   assign m198_64 ={ {2{in198[14]}} , in198[14:2] };

   // m198_65 = W*in
   wire signed [14:0] m198_65;
   assign m198_65 =15'b0;

   // m198_66 = W*in
   wire signed [14:0] m198_66;
   assign m198_66 ={ {4{neg198[14]}} , neg198[14:4] };

   // m198_67 = W*in
   wire signed [14:0] m198_67;
   assign m198_67 =15'b0;

   // m198_68 = W*in
   wire signed [14:0] m198_68;
   assign m198_68 =15'b0;

   // m198_69 = W*in
   wire signed [14:0] m198_69;
   assign m198_69 =15'b0;

   // m198_70 = W*in
   wire signed [14:0] m198_70;
   assign m198_70 =15'b0;

   // m198_71 = W*in
   wire signed [14:0] m198_71;
   assign m198_71 =15'b0;

   // m198_72 = W*in
   wire signed [14:0] m198_72;
   assign m198_72 =15'b0;

   // m198_73 = W*in
   wire signed [14:0] m198_73;
   assign m198_73 =15'b0;

   // m198_74 = W*in
   wire signed [14:0] m198_74;
   assign m198_74 =15'b0;

   // m198_75 = W*in
   wire signed [14:0] m198_75;
   assign m198_75 ={ {3{in198[14]}} , in198[14:3] };

   // m198_76 = W*in
   wire signed [14:0] m198_76;
   assign m198_76 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_77 = W*in
   wire signed [14:0] m198_77;
   assign m198_77 =15'b0;

   // m198_78 = W*in
   wire signed [14:0] m198_78;
   assign m198_78 =15'b0;

   // m198_79 = W*in
   wire signed [14:0] m198_79;
   assign m198_79 =15'b0;

   // m198_80 = W*in
   wire signed [14:0] m198_80;
   assign m198_80 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_81 = W*in
   wire signed [14:0] m198_81;
   assign m198_81 =15'b0;

   // m198_82 = W*in
   wire signed [14:0] m198_82;
   assign m198_82 =15'b0;

   // m198_83 = W*in
   wire signed [14:0] m198_83;
   assign m198_83 =15'b0;

   // m198_84 = W*in
   wire signed [14:0] m198_84;
   assign m198_84 =15'b0;

   // m198_85 = W*in
   wire signed [14:0] m198_85;
   assign m198_85 =15'b0;

   // m198_86 = W*in
   wire signed [14:0] m198_86;
   assign m198_86 =15'b0;

   // m198_87 = W*in
   wire signed [14:0] m198_87;
   assign m198_87 ={ {3{in198[14]}} , in198[14:3] };

   // m198_88 = W*in
   wire signed [14:0] m198_88;
   assign m198_88 =15'b0;

   // m198_89 = W*in
   wire signed [14:0] m198_89;
   assign m198_89 =15'b0;

   // m198_90 = W*in
   wire signed [14:0] m198_90;
   assign m198_90 =15'b0;

   // m198_91 = W*in
   wire signed [14:0] m198_91;
   assign m198_91 =15'b0;

   // m198_92 = W*in
   wire signed [14:0] m198_92;
   assign m198_92 ={ {2{in198[14]}} , in198[14:2] };

   // m198_93 = W*in
   wire signed [14:0] m198_93;
   assign m198_93 =15'b0;

   // m198_94 = W*in
   wire signed [14:0] m198_94;
   assign m198_94 =15'b0;

   // m198_95 = W*in
   wire signed [14:0] m198_95;
   assign m198_95 =15'b0;

   // m198_96 = W*in
   wire signed [14:0] m198_96;
   assign m198_96 ={ {3{neg198[14]}} , neg198[14:3] };

   // m198_97 = W*in
   wire signed [14:0] m198_97;
   assign m198_97 =15'b0;

   // m198_98 = W*in
   wire signed [14:0] m198_98;
   assign m198_98 =15'b0;

   // m198_99 = W*in
   wire signed [14:0] m198_99;
   assign m198_99 ={ {3{in198[14]}} , in198[14:3] };

   // m198_100 = W*in
   wire signed [14:0] m198_100;
   assign m198_100 =15'b0;

   // m199_1 = W*in
   wire signed [14:0] m199_1;
   assign m199_1 ={ {4{neg199[14]}} , neg199[14:4] };

   // m199_2 = W*in
   wire signed [14:0] m199_2;
   assign m199_2 =15'b0;

   // m199_3 = W*in
   wire signed [14:0] m199_3;
   assign m199_3 =15'b0;

   // m199_4 = W*in
   wire signed [14:0] m199_4;
   assign m199_4 =15'b0;

   // m199_5 = W*in
   wire signed [14:0] m199_5;
   assign m199_5 =15'b0;

   // m199_6 = W*in
   wire signed [14:0] m199_6;
   assign m199_6 =15'b0;

   // m199_7 = W*in
   wire signed [14:0] m199_7;
   assign m199_7 =15'b0;

   // m199_8 = W*in
   wire signed [14:0] m199_8;
   assign m199_8 =15'b0;

   // m199_9 = W*in
   wire signed [14:0] m199_9;
   assign m199_9 =15'b0;

   // m199_10 = W*in
   wire signed [14:0] m199_10;
   assign m199_10 =15'b0;

   // m199_11 = W*in
   wire signed [14:0] m199_11;
   assign m199_11 =15'b0;

   // m199_12 = W*in
   wire signed [14:0] m199_12;
   assign m199_12 =15'b0;

   // m199_13 = W*in
   wire signed [14:0] m199_13;
   assign m199_13 =15'b0;

   // m199_14 = W*in
   wire signed [14:0] m199_14;
   assign m199_14 =15'b0;

   // m199_15 = W*in
   wire signed [14:0] m199_15;
   assign m199_15 =15'b0;

   // m199_16 = W*in
   wire signed [14:0] m199_16;
   assign m199_16 =15'b0;

   // m199_17 = W*in
   wire signed [14:0] m199_17;
   assign m199_17 =15'b0;

   // m199_18 = W*in
   wire signed [14:0] m199_18;
   assign m199_18 =15'b0;

   // m199_19 = W*in
   wire signed [14:0] m199_19;
   assign m199_19 =15'b0;

   // m199_20 = W*in
   wire signed [14:0] m199_20;
   assign m199_20 ={ {4{in199[14]}} , in199[14:4] };

   // m199_21 = W*in
   wire signed [14:0] m199_21;
   assign m199_21 =15'b0;

   // m199_22 = W*in
   wire signed [14:0] m199_22;
   assign m199_22 =15'b0;

   // m199_23 = W*in
   wire signed [14:0] m199_23;
   assign m199_23 =15'b0;

   // m199_24 = W*in
   wire signed [14:0] m199_24;
   assign m199_24 =15'b0;

   // m199_25 = W*in
   wire signed [14:0] m199_25;
   assign m199_25 =15'b0;

   // m199_26 = W*in
   wire signed [14:0] m199_26;
   assign m199_26 =15'b0;

   // m199_27 = W*in
   wire signed [14:0] m199_27;
   assign m199_27 =15'b0;

   // m199_28 = W*in
   wire signed [14:0] m199_28;
   assign m199_28 =15'b0;

   // m199_29 = W*in
   wire signed [14:0] m199_29;
   assign m199_29 =15'b0;

   // m199_30 = W*in
   wire signed [14:0] m199_30;
   assign m199_30 =15'b0;

   // m199_31 = W*in
   wire signed [14:0] m199_31;
   assign m199_31 =15'b0;

   // m199_32 = W*in
   wire signed [14:0] m199_32;
   assign m199_32 =15'b0;

   // m199_33 = W*in
   wire signed [14:0] m199_33;
   assign m199_33 =15'b0;

   // m199_34 = W*in
   wire signed [14:0] m199_34;
   assign m199_34 =15'b0;

   // m199_35 = W*in
   wire signed [14:0] m199_35;
   assign m199_35 =15'b0;

   // m199_36 = W*in
   wire signed [14:0] m199_36;
   assign m199_36 =15'b0;

   // m199_37 = W*in
   wire signed [14:0] m199_37;
   assign m199_37 =15'b0;

   // m199_38 = W*in
   wire signed [14:0] m199_38;
   assign m199_38 =15'b0;

   // m199_39 = W*in
   wire signed [14:0] m199_39;
   assign m199_39 =15'b0;

   // m199_40 = W*in
   wire signed [14:0] m199_40;
   assign m199_40 =15'b0;

   // m199_41 = W*in
   wire signed [14:0] m199_41;
   assign m199_41 =15'b0;

   // m199_42 = W*in
   wire signed [14:0] m199_42;
   assign m199_42 =15'b0;

   // m199_43 = W*in
   wire signed [14:0] m199_43;
   assign m199_43 =15'b0;

   // m199_44 = W*in
   wire signed [14:0] m199_44;
   assign m199_44 =15'b0;

   // m199_45 = W*in
   wire signed [14:0] m199_45;
   assign m199_45 =15'b0;

   // m199_46 = W*in
   wire signed [14:0] m199_46;
   assign m199_46 =15'b0;

   // m199_47 = W*in
   wire signed [14:0] m199_47;
   assign m199_47 =15'b0;

   // m199_48 = W*in
   wire signed [14:0] m199_48;
   assign m199_48 =15'b0;

   // m199_49 = W*in
   wire signed [14:0] m199_49;
   assign m199_49 =15'b0;

   // m199_50 = W*in
   wire signed [14:0] m199_50;
   assign m199_50 =15'b0;

   // m199_51 = W*in
   wire signed [14:0] m199_51;
   assign m199_51 =15'b0;

   // m199_52 = W*in
   wire signed [14:0] m199_52;
   assign m199_52 =15'b0;

   // m199_53 = W*in
   wire signed [14:0] m199_53;
   assign m199_53 =15'b0;

   // m199_54 = W*in
   wire signed [14:0] m199_54;
   assign m199_54 =15'b0;

   // m199_55 = W*in
   wire signed [14:0] m199_55;
   assign m199_55 =15'b0;

   // m199_56 = W*in
   wire signed [14:0] m199_56;
   assign m199_56 =15'b0;

   // m199_57 = W*in
   wire signed [14:0] m199_57;
   assign m199_57 =15'b0;

   // m199_58 = W*in
   wire signed [14:0] m199_58;
   assign m199_58 =15'b0;

   // m199_59 = W*in
   wire signed [14:0] m199_59;
   assign m199_59 =15'b0;

   // m199_60 = W*in
   wire signed [14:0] m199_60;
   assign m199_60 ={ {4{in199[14]}} , in199[14:4] };

   // m199_61 = W*in
   wire signed [14:0] m199_61;
   assign m199_61 =15'b0;

   // m199_62 = W*in
   wire signed [14:0] m199_62;
   assign m199_62 =15'b0;

   // m199_63 = W*in
   wire signed [14:0] m199_63;
   assign m199_63 =15'b0;

   // m199_64 = W*in
   wire signed [14:0] m199_64;
   assign m199_64 =15'b0;

   // m199_65 = W*in
   wire signed [14:0] m199_65;
   assign m199_65 =15'b0;

   // m199_66 = W*in
   wire signed [14:0] m199_66;
   assign m199_66 =15'b0;

   // m199_67 = W*in
   wire signed [14:0] m199_67;
   assign m199_67 =15'b0;

   // m199_68 = W*in
   wire signed [14:0] m199_68;
   assign m199_68 =15'b0;

   // m199_69 = W*in
   wire signed [14:0] m199_69;
   assign m199_69 =15'b0;

   // m199_70 = W*in
   wire signed [14:0] m199_70;
   assign m199_70 =15'b0;

   // m199_71 = W*in
   wire signed [14:0] m199_71;
   assign m199_71 =15'b0;

   // m199_72 = W*in
   wire signed [14:0] m199_72;
   assign m199_72 =15'b0;

   // m199_73 = W*in
   wire signed [14:0] m199_73;
   assign m199_73 =15'b0;

   // m199_74 = W*in
   wire signed [14:0] m199_74;
   assign m199_74 ={ {3{in199[14]}} , in199[14:3] };

   // m199_75 = W*in
   wire signed [14:0] m199_75;
   assign m199_75 =15'b0;

   // m199_76 = W*in
   wire signed [14:0] m199_76;
   assign m199_76 ={ {4{neg199[14]}} , neg199[14:4] };

   // m199_77 = W*in
   wire signed [14:0] m199_77;
   assign m199_77 =15'b0;

   // m199_78 = W*in
   wire signed [14:0] m199_78;
   assign m199_78 ={ {3{in199[14]}} , in199[14:3] };

   // m199_79 = W*in
   wire signed [14:0] m199_79;
   assign m199_79 =15'b0;

   // m199_80 = W*in
   wire signed [14:0] m199_80;
   assign m199_80 =15'b0;

   // m199_81 = W*in
   wire signed [14:0] m199_81;
   assign m199_81 =15'b0;

   // m199_82 = W*in
   wire signed [14:0] m199_82;
   assign m199_82 =15'b0;

   // m199_83 = W*in
   wire signed [14:0] m199_83;
   assign m199_83 =15'b0;

   // m199_84 = W*in
   wire signed [14:0] m199_84;
   assign m199_84 =15'b0;

   // m199_85 = W*in
   wire signed [14:0] m199_85;
   assign m199_85 =15'b0;

   // m199_86 = W*in
   wire signed [14:0] m199_86;
   assign m199_86 =15'b0;

   // m199_87 = W*in
   wire signed [14:0] m199_87;
   assign m199_87 =15'b0;

   // m199_88 = W*in
   wire signed [14:0] m199_88;
   assign m199_88 =15'b0;

   // m199_89 = W*in
   wire signed [14:0] m199_89;
   assign m199_89 =15'b0;

   // m199_90 = W*in
   wire signed [14:0] m199_90;
   assign m199_90 =15'b0;

   // m199_91 = W*in
   wire signed [14:0] m199_91;
   assign m199_91 =15'b0;

   // m199_92 = W*in
   wire signed [14:0] m199_92;
   assign m199_92 =15'b0;

   // m199_93 = W*in
   wire signed [14:0] m199_93;
   assign m199_93 =15'b0;

   // m199_94 = W*in
   wire signed [14:0] m199_94;
   assign m199_94 =15'b0;

   // m199_95 = W*in
   wire signed [14:0] m199_95;
   assign m199_95 =15'b0;

   // m199_96 = W*in
   wire signed [14:0] m199_96;
   assign m199_96 =15'b0;

   // m199_97 = W*in
   wire signed [14:0] m199_97;
   assign m199_97 =15'b0;

   // m199_98 = W*in
   wire signed [14:0] m199_98;
   assign m199_98 =15'b0;

   // m199_99 = W*in
   wire signed [14:0] m199_99;
   assign m199_99 =15'b0;

   // m199_100 = W*in
   wire signed [14:0] m199_100;
   assign m199_100 =15'b0;

   // m200_1 = W*in
   wire signed [14:0] m200_1;
   assign m200_1 =15'b0;

   // m200_2 = W*in
   wire signed [14:0] m200_2;
   assign m200_2 =15'b0;

   // m200_3 = W*in
   wire signed [14:0] m200_3;
   assign m200_3 =15'b0;

   // m200_4 = W*in
   wire signed [14:0] m200_4;
   assign m200_4 =15'b0;

   // m200_5 = W*in
   wire signed [14:0] m200_5;
   assign m200_5 =15'b0;

   // m200_6 = W*in
   wire signed [14:0] m200_6;
   assign m200_6 =15'b0;

   // m200_7 = W*in
   wire signed [14:0] m200_7;
   assign m200_7 =15'b0;

   // m200_8 = W*in
   wire signed [14:0] m200_8;
   assign m200_8 =15'b0;

   // m200_9 = W*in
   wire signed [14:0] m200_9;
   assign m200_9 =15'b0;

   // m200_10 = W*in
   wire signed [14:0] m200_10;
   assign m200_10 ={ {3{in200[14]}} , in200[14:3] };

   // m200_11 = W*in
   wire signed [14:0] m200_11;
   assign m200_11 =15'b0;

   // m200_12 = W*in
   wire signed [14:0] m200_12;
   assign m200_12 =15'b0;

   // m200_13 = W*in
   wire signed [14:0] m200_13;
   assign m200_13 =15'b0;

   // m200_14 = W*in
   wire signed [14:0] m200_14;
   assign m200_14 =15'b0;

   // m200_15 = W*in
   wire signed [14:0] m200_15;
   assign m200_15 =15'b0;

   // m200_16 = W*in
   wire signed [14:0] m200_16;
   assign m200_16 ={ {3{neg200[14]}} , neg200[14:3] };

   // m200_17 = W*in
   wire signed [14:0] m200_17;
   assign m200_17 =15'b0;

   // m200_18 = W*in
   wire signed [14:0] m200_18;
   assign m200_18 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_19 = W*in
   wire signed [14:0] m200_19;
   assign m200_19 ={ {4{in200[14]}} , in200[14:4] };

   // m200_20 = W*in
   wire signed [14:0] m200_20;
   assign m200_20 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_21 = W*in
   wire signed [14:0] m200_21;
   assign m200_21 =15'b0;

   // m200_22 = W*in
   wire signed [14:0] m200_22;
   assign m200_22 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_23 = W*in
   wire signed [14:0] m200_23;
   assign m200_23 =15'b0;

   // m200_24 = W*in
   wire signed [14:0] m200_24;
   assign m200_24 =15'b0;

   // m200_25 = W*in
   wire signed [14:0] m200_25;
   assign m200_25 ={ {3{in200[14]}} , in200[14:3] };

   // m200_26 = W*in
   wire signed [14:0] m200_26;
   assign m200_26 ={ {3{neg200[14]}} , neg200[14:3] };

   // m200_27 = W*in
   wire signed [14:0] m200_27;
   assign m200_27 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_28 = W*in
   wire signed [14:0] m200_28;
   assign m200_28 =15'b0;

   // m200_29 = W*in
   wire signed [14:0] m200_29;
   assign m200_29 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_30 = W*in
   wire signed [14:0] m200_30;
   assign m200_30 =15'b0;

   // m200_31 = W*in
   wire signed [14:0] m200_31;
   assign m200_31 ={ {4{in200[14]}} , in200[14:4] };

   // m200_32 = W*in
   wire signed [14:0] m200_32;
   assign m200_32 =15'b0;

   // m200_33 = W*in
   wire signed [14:0] m200_33;
   assign m200_33 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_34 = W*in
   wire signed [14:0] m200_34;
   assign m200_34 =15'b0;

   // m200_35 = W*in
   wire signed [14:0] m200_35;
   assign m200_35 =15'b0;

   // m200_36 = W*in
   wire signed [14:0] m200_36;
   assign m200_36 =15'b0;

   // m200_37 = W*in
   wire signed [14:0] m200_37;
   assign m200_37 =15'b0;

   // m200_38 = W*in
   wire signed [14:0] m200_38;
   assign m200_38 =15'b0;

   // m200_39 = W*in
   wire signed [14:0] m200_39;
   assign m200_39 ={ {3{in200[14]}} , in200[14:3] };

   // m200_40 = W*in
   wire signed [14:0] m200_40;
   assign m200_40 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_41 = W*in
   wire signed [14:0] m200_41;
   assign m200_41 =15'b0;

   // m200_42 = W*in
   wire signed [14:0] m200_42;
   assign m200_42 =15'b0;

   // m200_43 = W*in
   wire signed [14:0] m200_43;
   assign m200_43 =15'b0;

   // m200_44 = W*in
   wire signed [14:0] m200_44;
   assign m200_44 ={ {3{in200[14]}} , in200[14:3] };

   // m200_45 = W*in
   wire signed [14:0] m200_45;
   assign m200_45 =15'b0;

   // m200_46 = W*in
   wire signed [14:0] m200_46;
   assign m200_46 =15'b0;

   // m200_47 = W*in
   wire signed [14:0] m200_47;
   assign m200_47 ={ {3{in200[14]}} , in200[14:3] };

   // m200_48 = W*in
   wire signed [14:0] m200_48;
   assign m200_48 =15'b0;

   // m200_49 = W*in
   wire signed [14:0] m200_49;
   assign m200_49 =15'b0;

   // m200_50 = W*in
   wire signed [14:0] m200_50;
   assign m200_50 =15'b0;

   // m200_51 = W*in
   wire signed [14:0] m200_51;
   assign m200_51 =15'b0;

   // m200_52 = W*in
   wire signed [14:0] m200_52;
   assign m200_52 =15'b0;

   // m200_53 = W*in
   wire signed [14:0] m200_53;
   assign m200_53 =15'b0;

   // m200_54 = W*in
   wire signed [14:0] m200_54;
   assign m200_54 =15'b0;

   // m200_55 = W*in
   wire signed [14:0] m200_55;
   assign m200_55 =15'b0;

   // m200_56 = W*in
   wire signed [14:0] m200_56;
   assign m200_56 =15'b0;

   // m200_57 = W*in
   wire signed [14:0] m200_57;
   assign m200_57 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_58 = W*in
   wire signed [14:0] m200_58;
   assign m200_58 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_59 = W*in
   wire signed [14:0] m200_59;
   assign m200_59 =15'b0;

   // m200_60 = W*in
   wire signed [14:0] m200_60;
   assign m200_60 ={ {4{neg200[14]}} , neg200[14:4] };

   // m200_61 = W*in
   wire signed [14:0] m200_61;
   assign m200_61 =15'b0;

   // m200_62 = W*in
   wire signed [14:0] m200_62;
   assign m200_62 =15'b0;

   // m200_63 = W*in
   wire signed [14:0] m200_63;
   assign m200_63 =15'b0;

   // m200_64 = W*in
   wire signed [14:0] m200_64;
   assign m200_64 =15'b0;

   // m200_65 = W*in
   wire signed [14:0] m200_65;
   assign m200_65 ={ {3{neg200[14]}} , neg200[14:3] };

   // m200_66 = W*in
   wire signed [14:0] m200_66;
   assign m200_66 =15'b0;

   // m200_67 = W*in
   wire signed [14:0] m200_67;
   assign m200_67 =15'b0;

   // m200_68 = W*in
   wire signed [14:0] m200_68;
   assign m200_68 =15'b0;

   // m200_69 = W*in
   wire signed [14:0] m200_69;
   assign m200_69 =15'b0;

   // m200_70 = W*in
   wire signed [14:0] m200_70;
   assign m200_70 =15'b0;

   // m200_71 = W*in
   wire signed [14:0] m200_71;
   assign m200_71 ={ {3{in200[14]}} , in200[14:3] };

   // m200_72 = W*in
   wire signed [14:0] m200_72;
   assign m200_72 =15'b0;

   // m200_73 = W*in
   wire signed [14:0] m200_73;
   assign m200_73 =15'b0;

   // m200_74 = W*in
   wire signed [14:0] m200_74;
   assign m200_74 =15'b0;

   // m200_75 = W*in
   wire signed [14:0] m200_75;
   assign m200_75 =15'b0;

   // m200_76 = W*in
   wire signed [14:0] m200_76;
   assign m200_76 =15'b0;

   // m200_77 = W*in
   wire signed [14:0] m200_77;
   assign m200_77 =15'b0;

   // m200_78 = W*in
   wire signed [14:0] m200_78;
   assign m200_78 =15'b0;

   // m200_79 = W*in
   wire signed [14:0] m200_79;
   assign m200_79 ={ {3{in200[14]}} , in200[14:3] };

   // m200_80 = W*in
   wire signed [14:0] m200_80;
   assign m200_80 =15'b0;

   // m200_81 = W*in
   wire signed [14:0] m200_81;
   assign m200_81 =15'b0;

   // m200_82 = W*in
   wire signed [14:0] m200_82;
   assign m200_82 =15'b0;

   // m200_83 = W*in
   wire signed [14:0] m200_83;
   assign m200_83 =15'b0;

   // m200_84 = W*in
   wire signed [14:0] m200_84;
   assign m200_84 ={ {3{neg200[14]}} , neg200[14:3] };

   // m200_85 = W*in
   wire signed [14:0] m200_85;
   assign m200_85 =15'b0;

   // m200_86 = W*in
   wire signed [14:0] m200_86;
   assign m200_86 =15'b0;

   // m200_87 = W*in
   wire signed [14:0] m200_87;
   assign m200_87 =15'b0;

   // m200_88 = W*in
   wire signed [14:0] m200_88;
   assign m200_88 =15'b0;

   // m200_89 = W*in
   wire signed [14:0] m200_89;
   assign m200_89 =15'b0;

   // m200_90 = W*in
   wire signed [14:0] m200_90;
   assign m200_90 =15'b0;

   // m200_91 = W*in
   wire signed [14:0] m200_91;
   assign m200_91 =15'b0;

   // m200_92 = W*in
   wire signed [14:0] m200_92;
   assign m200_92 =15'b0;

   // m200_93 = W*in
   wire signed [14:0] m200_93;
   assign m200_93 =15'b0;

   // m200_94 = W*in
   wire signed [14:0] m200_94;
   assign m200_94 =15'b0;

   // m200_95 = W*in
   wire signed [14:0] m200_95;
   assign m200_95 =15'b0;

   // m200_96 = W*in
   wire signed [14:0] m200_96;
   assign m200_96 =15'b0;

   // m200_97 = W*in
   wire signed [14:0] m200_97;
   assign m200_97 =15'b0;

   // m200_98 = W*in
   wire signed [14:0] m200_98;
   assign m200_98 =15'b0;

   // m200_99 = W*in
   wire signed [14:0] m200_99;
   assign m200_99 =15'b0;

   // m200_100 = W*in
   wire signed [14:0] m200_100;
   assign m200_100 =15'b0;

   // m201_1 = W*in
   wire signed [14:0] m201_1;
   assign m201_1 ={ {4{in201[14]}} , in201[14:4] };

   // m201_2 = W*in
   wire signed [14:0] m201_2;
   assign m201_2 =15'b0;

   // m201_3 = W*in
   wire signed [14:0] m201_3;
   assign m201_3 =15'b0;

   // m201_4 = W*in
   wire signed [14:0] m201_4;
   assign m201_4 ={ {4{neg201[14]}} , neg201[14:4] };

   // m201_5 = W*in
   wire signed [14:0] m201_5;
   assign m201_5 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_6 = W*in
   wire signed [14:0] m201_6;
   assign m201_6 =15'b0;

   // m201_7 = W*in
   wire signed [14:0] m201_7;
   assign m201_7 =15'b0;

   // m201_8 = W*in
   wire signed [14:0] m201_8;
   assign m201_8 =15'b0;

   // m201_9 = W*in
   wire signed [14:0] m201_9;
   assign m201_9 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_10 = W*in
   wire signed [14:0] m201_10;
   assign m201_10 =15'b0;

   // m201_11 = W*in
   wire signed [14:0] m201_11;
   assign m201_11 ={ {3{in201[14]}} , in201[14:3] };

   // m201_12 = W*in
   wire signed [14:0] m201_12;
   assign m201_12 =15'b0;

   // m201_13 = W*in
   wire signed [14:0] m201_13;
   assign m201_13 =15'b0;

   // m201_14 = W*in
   wire signed [14:0] m201_14;
   assign m201_14 =15'b0;

   // m201_15 = W*in
   wire signed [14:0] m201_15;
   assign m201_15 =15'b0;

   // m201_16 = W*in
   wire signed [14:0] m201_16;
   assign m201_16 =15'b0;

   // m201_17 = W*in
   wire signed [14:0] m201_17;
   assign m201_17 =15'b0;

   // m201_18 = W*in
   wire signed [14:0] m201_18;
   assign m201_18 ={ {3{in201[14]}} , in201[14:3] };

   // m201_19 = W*in
   wire signed [14:0] m201_19;
   assign m201_19 =15'b0;

   // m201_20 = W*in
   wire signed [14:0] m201_20;
   assign m201_20 =15'b0;

   // m201_21 = W*in
   wire signed [14:0] m201_21;
   assign m201_21 ={ {3{in201[14]}} , in201[14:3] };

   // m201_22 = W*in
   wire signed [14:0] m201_22;
   assign m201_22 =15'b0;

   // m201_23 = W*in
   wire signed [14:0] m201_23;
   assign m201_23 =15'b0;

   // m201_24 = W*in
   wire signed [14:0] m201_24;
   assign m201_24 =15'b0;

   // m201_25 = W*in
   wire signed [14:0] m201_25;
   assign m201_25 =15'b0;

   // m201_26 = W*in
   wire signed [14:0] m201_26;
   assign m201_26 =15'b0;

   // m201_27 = W*in
   wire signed [14:0] m201_27;
   assign m201_27 =15'b0;

   // m201_28 = W*in
   wire signed [14:0] m201_28;
   assign m201_28 =15'b0;

   // m201_29 = W*in
   wire signed [14:0] m201_29;
   assign m201_29 =15'b0;

   // m201_30 = W*in
   wire signed [14:0] m201_30;
   assign m201_30 =15'b0;

   // m201_31 = W*in
   wire signed [14:0] m201_31;
   assign m201_31 =15'b0;

   // m201_32 = W*in
   wire signed [14:0] m201_32;
   assign m201_32 =15'b0;

   // m201_33 = W*in
   wire signed [14:0] m201_33;
   assign m201_33 =15'b0;

   // m201_34 = W*in
   wire signed [14:0] m201_34;
   assign m201_34 =15'b0;

   // m201_35 = W*in
   wire signed [14:0] m201_35;
   assign m201_35 =15'b0;

   // m201_36 = W*in
   wire signed [14:0] m201_36;
   assign m201_36 =15'b0;

   // m201_37 = W*in
   wire signed [14:0] m201_37;
   assign m201_37 =15'b0;

   // m201_38 = W*in
   wire signed [14:0] m201_38;
   assign m201_38 =15'b0;

   // m201_39 = W*in
   wire signed [14:0] m201_39;
   assign m201_39 =15'b0;

   // m201_40 = W*in
   wire signed [14:0] m201_40;
   assign m201_40 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_41 = W*in
   wire signed [14:0] m201_41;
   assign m201_41 =15'b0;

   // m201_42 = W*in
   wire signed [14:0] m201_42;
   assign m201_42 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_43 = W*in
   wire signed [14:0] m201_43;
   assign m201_43 =15'b0;

   // m201_44 = W*in
   wire signed [14:0] m201_44;
   assign m201_44 =15'b0;

   // m201_45 = W*in
   wire signed [14:0] m201_45;
   assign m201_45 =15'b0;

   // m201_46 = W*in
   wire signed [14:0] m201_46;
   assign m201_46 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_47 = W*in
   wire signed [14:0] m201_47;
   assign m201_47 =15'b0;

   // m201_48 = W*in
   wire signed [14:0] m201_48;
   assign m201_48 =15'b0;

   // m201_49 = W*in
   wire signed [14:0] m201_49;
   assign m201_49 =15'b0;

   // m201_50 = W*in
   wire signed [14:0] m201_50;
   assign m201_50 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_51 = W*in
   wire signed [14:0] m201_51;
   assign m201_51 =15'b0;

   // m201_52 = W*in
   wire signed [14:0] m201_52;
   assign m201_52 =15'b0;

   // m201_53 = W*in
   wire signed [14:0] m201_53;
   assign m201_53 =15'b0;

   // m201_54 = W*in
   wire signed [14:0] m201_54;
   assign m201_54 =15'b0;

   // m201_55 = W*in
   wire signed [14:0] m201_55;
   assign m201_55 =15'b0;

   // m201_56 = W*in
   wire signed [14:0] m201_56;
   assign m201_56 =15'b0;

   // m201_57 = W*in
   wire signed [14:0] m201_57;
   assign m201_57 =15'b0;

   // m201_58 = W*in
   wire signed [14:0] m201_58;
   assign m201_58 =15'b0;

   // m201_59 = W*in
   wire signed [14:0] m201_59;
   assign m201_59 ={ {4{in201[14]}} , in201[14:4] };

   // m201_60 = W*in
   wire signed [14:0] m201_60;
   assign m201_60 ={ {3{in201[14]}} , in201[14:3] };

   // m201_61 = W*in
   wire signed [14:0] m201_61;
   assign m201_61 =15'b0;

   // m201_62 = W*in
   wire signed [14:0] m201_62;
   assign m201_62 =15'b0;

   // m201_63 = W*in
   wire signed [14:0] m201_63;
   assign m201_63 ={ {4{neg201[14]}} , neg201[14:4] };

   // m201_64 = W*in
   wire signed [14:0] m201_64;
   assign m201_64 =15'b0;

   // m201_65 = W*in
   wire signed [14:0] m201_65;
   assign m201_65 =15'b0;

   // m201_66 = W*in
   wire signed [14:0] m201_66;
   assign m201_66 =15'b0;

   // m201_67 = W*in
   wire signed [14:0] m201_67;
   assign m201_67 =15'b0;

   // m201_68 = W*in
   wire signed [14:0] m201_68;
   assign m201_68 =15'b0;

   // m201_69 = W*in
   wire signed [14:0] m201_69;
   assign m201_69 =15'b0;

   // m201_70 = W*in
   wire signed [14:0] m201_70;
   assign m201_70 =15'b0;

   // m201_71 = W*in
   wire signed [14:0] m201_71;
   assign m201_71 =15'b0;

   // m201_72 = W*in
   wire signed [14:0] m201_72;
   assign m201_72 =15'b0;

   // m201_73 = W*in
   wire signed [14:0] m201_73;
   assign m201_73 =15'b0;

   // m201_74 = W*in
   wire signed [14:0] m201_74;
   assign m201_74 =15'b0;

   // m201_75 = W*in
   wire signed [14:0] m201_75;
   assign m201_75 =15'b0;

   // m201_76 = W*in
   wire signed [14:0] m201_76;
   assign m201_76 ={ {3{neg201[14]}} , neg201[14:3] };

   // m201_77 = W*in
   wire signed [14:0] m201_77;
   assign m201_77 ={ {4{in201[14]}} , in201[14:4] };

   // m201_78 = W*in
   wire signed [14:0] m201_78;
   assign m201_78 ={ {3{in201[14]}} , in201[14:3] };

   // m201_79 = W*in
   wire signed [14:0] m201_79;
   assign m201_79 =15'b0;

   // m201_80 = W*in
   wire signed [14:0] m201_80;
   assign m201_80 =15'b0;

   // m201_81 = W*in
   wire signed [14:0] m201_81;
   assign m201_81 =15'b0;

   // m201_82 = W*in
   wire signed [14:0] m201_82;
   assign m201_82 =15'b0;

   // m201_83 = W*in
   wire signed [14:0] m201_83;
   assign m201_83 =15'b0;

   // m201_84 = W*in
   wire signed [14:0] m201_84;
   assign m201_84 =15'b0;

   // m201_85 = W*in
   wire signed [14:0] m201_85;
   assign m201_85 =15'b0;

   // m201_86 = W*in
   wire signed [14:0] m201_86;
   assign m201_86 =15'b0;

   // m201_87 = W*in
   wire signed [14:0] m201_87;
   assign m201_87 =15'b0;

   // m201_88 = W*in
   wire signed [14:0] m201_88;
   assign m201_88 ={ {3{in201[14]}} , in201[14:3] };

   // m201_89 = W*in
   wire signed [14:0] m201_89;
   assign m201_89 =15'b0;

   // m201_90 = W*in
   wire signed [14:0] m201_90;
   assign m201_90 =15'b0;

   // m201_91 = W*in
   wire signed [14:0] m201_91;
   assign m201_91 =15'b0;

   // m201_92 = W*in
   wire signed [14:0] m201_92;
   assign m201_92 ={ {3{in201[14]}} , in201[14:3] };

   // m201_93 = W*in
   wire signed [14:0] m201_93;
   assign m201_93 =15'b0;

   // m201_94 = W*in
   wire signed [14:0] m201_94;
   assign m201_94 =15'b0;

   // m201_95 = W*in
   wire signed [14:0] m201_95;
   assign m201_95 ={ {4{neg201[14]}} , neg201[14:4] };

   // m201_96 = W*in
   wire signed [14:0] m201_96;
   assign m201_96 =15'b0;

   // m201_97 = W*in
   wire signed [14:0] m201_97;
   assign m201_97 =15'b0;

   // m201_98 = W*in
   wire signed [14:0] m201_98;
   assign m201_98 =15'b0;

   // m201_99 = W*in
   wire signed [14:0] m201_99;
   assign m201_99 =15'b0;

   // m201_100 = W*in
   wire signed [14:0] m201_100;
   assign m201_100 =15'b0;

   // m202_1 = W*in
   wire signed [14:0] m202_1;
   assign m202_1 =15'b0;

   // m202_2 = W*in
   wire signed [14:0] m202_2;
   assign m202_2 =15'b0;

   // m202_3 = W*in
   wire signed [14:0] m202_3;
   assign m202_3 ={ {3{in202[14]}} , in202[14:3] };

   // m202_4 = W*in
   wire signed [14:0] m202_4;
   assign m202_4 =15'b0;

   // m202_5 = W*in
   wire signed [14:0] m202_5;
   assign m202_5 =15'b0;

   // m202_6 = W*in
   wire signed [14:0] m202_6;
   assign m202_6 =15'b0;

   // m202_7 = W*in
   wire signed [14:0] m202_7;
   assign m202_7 =15'b0;

   // m202_8 = W*in
   wire signed [14:0] m202_8;
   assign m202_8 =15'b0;

   // m202_9 = W*in
   wire signed [14:0] m202_9;
   assign m202_9 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_10 = W*in
   wire signed [14:0] m202_10;
   assign m202_10 =15'b0;

   // m202_11 = W*in
   wire signed [14:0] m202_11;
   assign m202_11 =15'b0;

   // m202_12 = W*in
   wire signed [14:0] m202_12;
   assign m202_12 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_13 = W*in
   wire signed [14:0] m202_13;
   assign m202_13 =15'b0;

   // m202_14 = W*in
   wire signed [14:0] m202_14;
   assign m202_14 =15'b0;

   // m202_15 = W*in
   wire signed [14:0] m202_15;
   assign m202_15 =15'b0;

   // m202_16 = W*in
   wire signed [14:0] m202_16;
   assign m202_16 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_17 = W*in
   wire signed [14:0] m202_17;
   assign m202_17 ={ {3{in202[14]}} , in202[14:3] };

   // m202_18 = W*in
   wire signed [14:0] m202_18;
   assign m202_18 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_19 = W*in
   wire signed [14:0] m202_19;
   assign m202_19 =15'b0;

   // m202_20 = W*in
   wire signed [14:0] m202_20;
   assign m202_20 =15'b0;

   // m202_21 = W*in
   wire signed [14:0] m202_21;
   assign m202_21 =15'b0;

   // m202_22 = W*in
   wire signed [14:0] m202_22;
   assign m202_22 ={ {4{neg202[14]}} , neg202[14:4] };

   // m202_23 = W*in
   wire signed [14:0] m202_23;
   assign m202_23 =15'b0;

   // m202_24 = W*in
   wire signed [14:0] m202_24;
   assign m202_24 =15'b0;

   // m202_25 = W*in
   wire signed [14:0] m202_25;
   assign m202_25 =15'b0;

   // m202_26 = W*in
   wire signed [14:0] m202_26;
   assign m202_26 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_27 = W*in
   wire signed [14:0] m202_27;
   assign m202_27 =15'b0;

   // m202_28 = W*in
   wire signed [14:0] m202_28;
   assign m202_28 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_29 = W*in
   wire signed [14:0] m202_29;
   assign m202_29 =15'b0;

   // m202_30 = W*in
   wire signed [14:0] m202_30;
   assign m202_30 =15'b0;

   // m202_31 = W*in
   wire signed [14:0] m202_31;
   assign m202_31 =15'b0;

   // m202_32 = W*in
   wire signed [14:0] m202_32;
   assign m202_32 =15'b0;

   // m202_33 = W*in
   wire signed [14:0] m202_33;
   assign m202_33 ={ {4{neg202[14]}} , neg202[14:4] };

   // m202_34 = W*in
   wire signed [14:0] m202_34;
   assign m202_34 =15'b0;

   // m202_35 = W*in
   wire signed [14:0] m202_35;
   assign m202_35 =15'b0;

   // m202_36 = W*in
   wire signed [14:0] m202_36;
   assign m202_36 =15'b0;

   // m202_37 = W*in
   wire signed [14:0] m202_37;
   assign m202_37 =15'b0;

   // m202_38 = W*in
   wire signed [14:0] m202_38;
   assign m202_38 =15'b0;

   // m202_39 = W*in
   wire signed [14:0] m202_39;
   assign m202_39 ={ {3{in202[14]}} , in202[14:3] };

   // m202_40 = W*in
   wire signed [14:0] m202_40;
   assign m202_40 =15'b0;

   // m202_41 = W*in
   wire signed [14:0] m202_41;
   assign m202_41 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_42 = W*in
   wire signed [14:0] m202_42;
   assign m202_42 =15'b0;

   // m202_43 = W*in
   wire signed [14:0] m202_43;
   assign m202_43 =15'b0;

   // m202_44 = W*in
   wire signed [14:0] m202_44;
   assign m202_44 ={ {3{in202[14]}} , in202[14:3] };

   // m202_45 = W*in
   wire signed [14:0] m202_45;
   assign m202_45 =15'b0;

   // m202_46 = W*in
   wire signed [14:0] m202_46;
   assign m202_46 =15'b0;

   // m202_47 = W*in
   wire signed [14:0] m202_47;
   assign m202_47 =15'b0;

   // m202_48 = W*in
   wire signed [14:0] m202_48;
   assign m202_48 ={ {4{neg202[14]}} , neg202[14:4] };

   // m202_49 = W*in
   wire signed [14:0] m202_49;
   assign m202_49 =15'b0;

   // m202_50 = W*in
   wire signed [14:0] m202_50;
   assign m202_50 =15'b0;

   // m202_51 = W*in
   wire signed [14:0] m202_51;
   assign m202_51 =15'b0;

   // m202_52 = W*in
   wire signed [14:0] m202_52;
   assign m202_52 =15'b0;

   // m202_53 = W*in
   wire signed [14:0] m202_53;
   assign m202_53 =15'b0;

   // m202_54 = W*in
   wire signed [14:0] m202_54;
   assign m202_54 ={ {3{in202[14]}} , in202[14:3] };

   // m202_55 = W*in
   wire signed [14:0] m202_55;
   assign m202_55 =15'b0;

   // m202_56 = W*in
   wire signed [14:0] m202_56;
   assign m202_56 =15'b0;

   // m202_57 = W*in
   wire signed [14:0] m202_57;
   assign m202_57 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_58 = W*in
   wire signed [14:0] m202_58;
   assign m202_58 =15'b0;

   // m202_59 = W*in
   wire signed [14:0] m202_59;
   assign m202_59 =15'b0;

   // m202_60 = W*in
   wire signed [14:0] m202_60;
   assign m202_60 =15'b0;

   // m202_61 = W*in
   wire signed [14:0] m202_61;
   assign m202_61 ={ {4{neg202[14]}} , neg202[14:4] };

   // m202_62 = W*in
   wire signed [14:0] m202_62;
   assign m202_62 =15'b0;

   // m202_63 = W*in
   wire signed [14:0] m202_63;
   assign m202_63 =15'b0;

   // m202_64 = W*in
   wire signed [14:0] m202_64;
   assign m202_64 =15'b0;

   // m202_65 = W*in
   wire signed [14:0] m202_65;
   assign m202_65 =15'b0;

   // m202_66 = W*in
   wire signed [14:0] m202_66;
   assign m202_66 ={ {3{in202[14]}} , in202[14:3] };

   // m202_67 = W*in
   wire signed [14:0] m202_67;
   assign m202_67 =15'b0;

   // m202_68 = W*in
   wire signed [14:0] m202_68;
   assign m202_68 ={ {4{neg202[14]}} , neg202[14:4] };

   // m202_69 = W*in
   wire signed [14:0] m202_69;
   assign m202_69 =15'b0;

   // m202_70 = W*in
   wire signed [14:0] m202_70;
   assign m202_70 ={ {3{in202[14]}} , in202[14:3] };

   // m202_71 = W*in
   wire signed [14:0] m202_71;
   assign m202_71 =15'b0;

   // m202_72 = W*in
   wire signed [14:0] m202_72;
   assign m202_72 =15'b0;

   // m202_73 = W*in
   wire signed [14:0] m202_73;
   assign m202_73 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_74 = W*in
   wire signed [14:0] m202_74;
   assign m202_74 =15'b0;

   // m202_75 = W*in
   wire signed [14:0] m202_75;
   assign m202_75 =15'b0;

   // m202_76 = W*in
   wire signed [14:0] m202_76;
   assign m202_76 =15'b0;

   // m202_77 = W*in
   wire signed [14:0] m202_77;
   assign m202_77 =15'b0;

   // m202_78 = W*in
   wire signed [14:0] m202_78;
   assign m202_78 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_79 = W*in
   wire signed [14:0] m202_79;
   assign m202_79 =15'b0;

   // m202_80 = W*in
   wire signed [14:0] m202_80;
   assign m202_80 =15'b0;

   // m202_81 = W*in
   wire signed [14:0] m202_81;
   assign m202_81 =15'b0;

   // m202_82 = W*in
   wire signed [14:0] m202_82;
   assign m202_82 =15'b0;

   // m202_83 = W*in
   wire signed [14:0] m202_83;
   assign m202_83 =15'b0;

   // m202_84 = W*in
   wire signed [14:0] m202_84;
   assign m202_84 =15'b0;

   // m202_85 = W*in
   wire signed [14:0] m202_85;
   assign m202_85 =15'b0;

   // m202_86 = W*in
   wire signed [14:0] m202_86;
   assign m202_86 ={ {3{in202[14]}} , in202[14:3] };

   // m202_87 = W*in
   wire signed [14:0] m202_87;
   assign m202_87 =15'b0;

   // m202_88 = W*in
   wire signed [14:0] m202_88;
   assign m202_88 =15'b0;

   // m202_89 = W*in
   wire signed [14:0] m202_89;
   assign m202_89 =15'b0;

   // m202_90 = W*in
   wire signed [14:0] m202_90;
   assign m202_90 =15'b0;

   // m202_91 = W*in
   wire signed [14:0] m202_91;
   assign m202_91 =15'b0;

   // m202_92 = W*in
   wire signed [14:0] m202_92;
   assign m202_92 =15'b0;

   // m202_93 = W*in
   wire signed [14:0] m202_93;
   assign m202_93 =15'b0;

   // m202_94 = W*in
   wire signed [14:0] m202_94;
   assign m202_94 ={ {3{in202[14]}} , in202[14:3] };

   // m202_95 = W*in
   wire signed [14:0] m202_95;
   assign m202_95 ={ {3{in202[14]}} , in202[14:3] };

   // m202_96 = W*in
   wire signed [14:0] m202_96;
   assign m202_96 =15'b0;

   // m202_97 = W*in
   wire signed [14:0] m202_97;
   assign m202_97 ={ {3{neg202[14]}} , neg202[14:3] };

   // m202_98 = W*in
   wire signed [14:0] m202_98;
   assign m202_98 =15'b0;

   // m202_99 = W*in
   wire signed [14:0] m202_99;
   assign m202_99 =15'b0;

   // m202_100 = W*in
   wire signed [14:0] m202_100;
   assign m202_100 =15'b0;

   // m203_1 = W*in
   wire signed [14:0] m203_1;
   assign m203_1 =15'b0;

   // m203_2 = W*in
   wire signed [14:0] m203_2;
   assign m203_2 =15'b0;

   // m203_3 = W*in
   wire signed [14:0] m203_3;
   assign m203_3 =15'b0;

   // m203_4 = W*in
   wire signed [14:0] m203_4;
   assign m203_4 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_5 = W*in
   wire signed [14:0] m203_5;
   assign m203_5 ={ {4{in203[14]}} , in203[14:4] };

   // m203_6 = W*in
   wire signed [14:0] m203_6;
   assign m203_6 =15'b0;

   // m203_7 = W*in
   wire signed [14:0] m203_7;
   assign m203_7 =15'b0;

   // m203_8 = W*in
   wire signed [14:0] m203_8;
   assign m203_8 =15'b0;

   // m203_9 = W*in
   wire signed [14:0] m203_9;
   assign m203_9 =15'b0;

   // m203_10 = W*in
   wire signed [14:0] m203_10;
   assign m203_10 =15'b0;

   // m203_11 = W*in
   wire signed [14:0] m203_11;
   assign m203_11 =15'b0;

   // m203_12 = W*in
   wire signed [14:0] m203_12;
   assign m203_12 =15'b0;

   // m203_13 = W*in
   wire signed [14:0] m203_13;
   assign m203_13 =15'b0;

   // m203_14 = W*in
   wire signed [14:0] m203_14;
   assign m203_14 =15'b0;

   // m203_15 = W*in
   wire signed [14:0] m203_15;
   assign m203_15 =15'b0;

   // m203_16 = W*in
   wire signed [14:0] m203_16;
   assign m203_16 =15'b0;

   // m203_17 = W*in
   wire signed [14:0] m203_17;
   assign m203_17 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_18 = W*in
   wire signed [14:0] m203_18;
   assign m203_18 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_19 = W*in
   wire signed [14:0] m203_19;
   assign m203_19 ={ {4{in203[14]}} , in203[14:4] };

   // m203_20 = W*in
   wire signed [14:0] m203_20;
   assign m203_20 =15'b0;

   // m203_21 = W*in
   wire signed [14:0] m203_21;
   assign m203_21 ={ {4{in203[14]}} , in203[14:4] };

   // m203_22 = W*in
   wire signed [14:0] m203_22;
   assign m203_22 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_23 = W*in
   wire signed [14:0] m203_23;
   assign m203_23 =15'b0;

   // m203_24 = W*in
   wire signed [14:0] m203_24;
   assign m203_24 =15'b0;

   // m203_25 = W*in
   wire signed [14:0] m203_25;
   assign m203_25 ={ {3{in203[14]}} , in203[14:3] };

   // m203_26 = W*in
   wire signed [14:0] m203_26;
   assign m203_26 ={ {3{in203[14]}} , in203[14:3] };

   // m203_27 = W*in
   wire signed [14:0] m203_27;
   assign m203_27 ={ {4{in203[14]}} , in203[14:4] };

   // m203_28 = W*in
   wire signed [14:0] m203_28;
   assign m203_28 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_29 = W*in
   wire signed [14:0] m203_29;
   assign m203_29 ={ {4{in203[14]}} , in203[14:4] };

   // m203_30 = W*in
   wire signed [14:0] m203_30;
   assign m203_30 ={ {3{in203[14]}} , in203[14:3] };

   // m203_31 = W*in
   wire signed [14:0] m203_31;
   assign m203_31 =15'b0;

   // m203_32 = W*in
   wire signed [14:0] m203_32;
   assign m203_32 ={ {3{in203[14]}} , in203[14:3] };

   // m203_33 = W*in
   wire signed [14:0] m203_33;
   assign m203_33 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_34 = W*in
   wire signed [14:0] m203_34;
   assign m203_34 =15'b0;

   // m203_35 = W*in
   wire signed [14:0] m203_35;
   assign m203_35 =15'b0;

   // m203_36 = W*in
   wire signed [14:0] m203_36;
   assign m203_36 =15'b0;

   // m203_37 = W*in
   wire signed [14:0] m203_37;
   assign m203_37 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_38 = W*in
   wire signed [14:0] m203_38;
   assign m203_38 =15'b0;

   // m203_39 = W*in
   wire signed [14:0] m203_39;
   assign m203_39 =15'b0;

   // m203_40 = W*in
   wire signed [14:0] m203_40;
   assign m203_40 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_41 = W*in
   wire signed [14:0] m203_41;
   assign m203_41 =15'b0;

   // m203_42 = W*in
   wire signed [14:0] m203_42;
   assign m203_42 =15'b0;

   // m203_43 = W*in
   wire signed [14:0] m203_43;
   assign m203_43 ={ {3{in203[14]}} , in203[14:3] };

   // m203_44 = W*in
   wire signed [14:0] m203_44;
   assign m203_44 =15'b0;

   // m203_45 = W*in
   wire signed [14:0] m203_45;
   assign m203_45 =15'b0;

   // m203_46 = W*in
   wire signed [14:0] m203_46;
   assign m203_46 =15'b0;

   // m203_47 = W*in
   wire signed [14:0] m203_47;
   assign m203_47 =15'b0;

   // m203_48 = W*in
   wire signed [14:0] m203_48;
   assign m203_48 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_49 = W*in
   wire signed [14:0] m203_49;
   assign m203_49 =15'b0;

   // m203_50 = W*in
   wire signed [14:0] m203_50;
   assign m203_50 =15'b0;

   // m203_51 = W*in
   wire signed [14:0] m203_51;
   assign m203_51 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_52 = W*in
   wire signed [14:0] m203_52;
   assign m203_52 =15'b0;

   // m203_53 = W*in
   wire signed [14:0] m203_53;
   assign m203_53 =15'b0;

   // m203_54 = W*in
   wire signed [14:0] m203_54;
   assign m203_54 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_55 = W*in
   wire signed [14:0] m203_55;
   assign m203_55 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_56 = W*in
   wire signed [14:0] m203_56;
   assign m203_56 =15'b0;

   // m203_57 = W*in
   wire signed [14:0] m203_57;
   assign m203_57 =15'b0;

   // m203_58 = W*in
   wire signed [14:0] m203_58;
   assign m203_58 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_59 = W*in
   wire signed [14:0] m203_59;
   assign m203_59 =15'b0;

   // m203_60 = W*in
   wire signed [14:0] m203_60;
   assign m203_60 =15'b0;

   // m203_61 = W*in
   wire signed [14:0] m203_61;
   assign m203_61 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_62 = W*in
   wire signed [14:0] m203_62;
   assign m203_62 =15'b0;

   // m203_63 = W*in
   wire signed [14:0] m203_63;
   assign m203_63 =15'b0;

   // m203_64 = W*in
   wire signed [14:0] m203_64;
   assign m203_64 =15'b0;

   // m203_65 = W*in
   wire signed [14:0] m203_65;
   assign m203_65 ={ {3{in203[14]}} , in203[14:3] };

   // m203_66 = W*in
   wire signed [14:0] m203_66;
   assign m203_66 =15'b0;

   // m203_67 = W*in
   wire signed [14:0] m203_67;
   assign m203_67 ={ {4{in203[14]}} , in203[14:4] };

   // m203_68 = W*in
   wire signed [14:0] m203_68;
   assign m203_68 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_69 = W*in
   wire signed [14:0] m203_69;
   assign m203_69 ={ {3{in203[14]}} , in203[14:3] };

   // m203_70 = W*in
   wire signed [14:0] m203_70;
   assign m203_70 ={ {4{neg203[14]}} , neg203[14:4] };

   // m203_71 = W*in
   wire signed [14:0] m203_71;
   assign m203_71 =15'b0;

   // m203_72 = W*in
   wire signed [14:0] m203_72;
   assign m203_72 =15'b0;

   // m203_73 = W*in
   wire signed [14:0] m203_73;
   assign m203_73 =15'b0;

   // m203_74 = W*in
   wire signed [14:0] m203_74;
   assign m203_74 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_75 = W*in
   wire signed [14:0] m203_75;
   assign m203_75 =15'b0;

   // m203_76 = W*in
   wire signed [14:0] m203_76;
   assign m203_76 =15'b0;

   // m203_77 = W*in
   wire signed [14:0] m203_77;
   assign m203_77 ={ {3{in203[14]}} , in203[14:3] };

   // m203_78 = W*in
   wire signed [14:0] m203_78;
   assign m203_78 =15'b0;

   // m203_79 = W*in
   wire signed [14:0] m203_79;
   assign m203_79 =15'b0;

   // m203_80 = W*in
   wire signed [14:0] m203_80;
   assign m203_80 =15'b0;

   // m203_81 = W*in
   wire signed [14:0] m203_81;
   assign m203_81 =15'b0;

   // m203_82 = W*in
   wire signed [14:0] m203_82;
   assign m203_82 =15'b0;

   // m203_83 = W*in
   wire signed [14:0] m203_83;
   assign m203_83 =15'b0;

   // m203_84 = W*in
   wire signed [14:0] m203_84;
   assign m203_84 =15'b0;

   // m203_85 = W*in
   wire signed [14:0] m203_85;
   assign m203_85 =15'b0;

   // m203_86 = W*in
   wire signed [14:0] m203_86;
   assign m203_86 =15'b0;

   // m203_87 = W*in
   wire signed [14:0] m203_87;
   assign m203_87 =15'b0;

   // m203_88 = W*in
   wire signed [14:0] m203_88;
   assign m203_88 =15'b0;

   // m203_89 = W*in
   wire signed [14:0] m203_89;
   assign m203_89 ={ {3{neg203[14]}} , neg203[14:3] };

   // m203_90 = W*in
   wire signed [14:0] m203_90;
   assign m203_90 ={ {3{in203[14]}} , in203[14:3] };

   // m203_91 = W*in
   wire signed [14:0] m203_91;
   assign m203_91 =15'b0;

   // m203_92 = W*in
   wire signed [14:0] m203_92;
   assign m203_92 =15'b0;

   // m203_93 = W*in
   wire signed [14:0] m203_93;
   assign m203_93 =15'b0;

   // m203_94 = W*in
   wire signed [14:0] m203_94;
   assign m203_94 =15'b0;

   // m203_95 = W*in
   wire signed [14:0] m203_95;
   assign m203_95 =15'b0;

   // m203_96 = W*in
   wire signed [14:0] m203_96;
   assign m203_96 =15'b0;

   // m203_97 = W*in
   wire signed [14:0] m203_97;
   assign m203_97 =15'b0;

   // m203_98 = W*in
   wire signed [14:0] m203_98;
   assign m203_98 =15'b0;

   // m203_99 = W*in
   wire signed [14:0] m203_99;
   assign m203_99 =15'b0;

   // m203_100 = W*in
   wire signed [14:0] m203_100;
   assign m203_100 =15'b0;

   // m204_1 = W*in
   wire signed [14:0] m204_1;
   assign m204_1 =15'b0;

   // m204_2 = W*in
   wire signed [14:0] m204_2;
   assign m204_2 =15'b0;

   // m204_3 = W*in
   wire signed [14:0] m204_3;
   assign m204_3 =15'b0;

   // m204_4 = W*in
   wire signed [14:0] m204_4;
   assign m204_4 =15'b0;

   // m204_5 = W*in
   wire signed [14:0] m204_5;
   assign m204_5 =15'b0;

   // m204_6 = W*in
   wire signed [14:0] m204_6;
   assign m204_6 =15'b0;

   // m204_7 = W*in
   wire signed [14:0] m204_7;
   assign m204_7 =15'b0;

   // m204_8 = W*in
   wire signed [14:0] m204_8;
   assign m204_8 =15'b0;

   // m204_9 = W*in
   wire signed [14:0] m204_9;
   assign m204_9 =15'b0;

   // m204_10 = W*in
   wire signed [14:0] m204_10;
   assign m204_10 =15'b0;

   // m204_11 = W*in
   wire signed [14:0] m204_11;
   assign m204_11 =15'b0;

   // m204_12 = W*in
   wire signed [14:0] m204_12;
   assign m204_12 =15'b0;

   // m204_13 = W*in
   wire signed [14:0] m204_13;
   assign m204_13 =15'b0;

   // m204_14 = W*in
   wire signed [14:0] m204_14;
   assign m204_14 =15'b0;

   // m204_15 = W*in
   wire signed [14:0] m204_15;
   assign m204_15 =15'b0;

   // m204_16 = W*in
   wire signed [14:0] m204_16;
   assign m204_16 =15'b0;

   // m204_17 = W*in
   wire signed [14:0] m204_17;
   assign m204_17 =15'b0;

   // m204_18 = W*in
   wire signed [14:0] m204_18;
   assign m204_18 =15'b0;

   // m204_19 = W*in
   wire signed [14:0] m204_19;
   assign m204_19 ={ {4{in204[14]}} , in204[14:4] };

   // m204_20 = W*in
   wire signed [14:0] m204_20;
   assign m204_20 =15'b0;

   // m204_21 = W*in
   wire signed [14:0] m204_21;
   assign m204_21 =15'b0;

   // m204_22 = W*in
   wire signed [14:0] m204_22;
   assign m204_22 =15'b0;

   // m204_23 = W*in
   wire signed [14:0] m204_23;
   assign m204_23 =15'b0;

   // m204_24 = W*in
   wire signed [14:0] m204_24;
   assign m204_24 =15'b0;

   // m204_25 = W*in
   wire signed [14:0] m204_25;
   assign m204_25 =15'b0;

   // m204_26 = W*in
   wire signed [14:0] m204_26;
   assign m204_26 ={ {4{neg204[14]}} , neg204[14:4] };

   // m204_27 = W*in
   wire signed [14:0] m204_27;
   assign m204_27 =15'b0;

   // m204_28 = W*in
   wire signed [14:0] m204_28;
   assign m204_28 =15'b0;

   // m204_29 = W*in
   wire signed [14:0] m204_29;
   assign m204_29 ={ {4{neg204[14]}} , neg204[14:4] };

   // m204_30 = W*in
   wire signed [14:0] m204_30;
   assign m204_30 =15'b0;

   // m204_31 = W*in
   wire signed [14:0] m204_31;
   assign m204_31 ={ {4{neg204[14]}} , neg204[14:4] };

   // m204_32 = W*in
   wire signed [14:0] m204_32;
   assign m204_32 =15'b0;

   // m204_33 = W*in
   wire signed [14:0] m204_33;
   assign m204_33 =15'b0;

   // m204_34 = W*in
   wire signed [14:0] m204_34;
   assign m204_34 =15'b0;

   // m204_35 = W*in
   wire signed [14:0] m204_35;
   assign m204_35 =15'b0;

   // m204_36 = W*in
   wire signed [14:0] m204_36;
   assign m204_36 =15'b0;

   // m204_37 = W*in
   wire signed [14:0] m204_37;
   assign m204_37 =15'b0;

   // m204_38 = W*in
   wire signed [14:0] m204_38;
   assign m204_38 =15'b0;

   // m204_39 = W*in
   wire signed [14:0] m204_39;
   assign m204_39 =15'b0;

   // m204_40 = W*in
   wire signed [14:0] m204_40;
   assign m204_40 =15'b0;

   // m204_41 = W*in
   wire signed [14:0] m204_41;
   assign m204_41 =15'b0;

   // m204_42 = W*in
   wire signed [14:0] m204_42;
   assign m204_42 =15'b0;

   // m204_43 = W*in
   wire signed [14:0] m204_43;
   assign m204_43 =15'b0;

   // m204_44 = W*in
   wire signed [14:0] m204_44;
   assign m204_44 =15'b0;

   // m204_45 = W*in
   wire signed [14:0] m204_45;
   assign m204_45 =15'b0;

   // m204_46 = W*in
   wire signed [14:0] m204_46;
   assign m204_46 =15'b0;

   // m204_47 = W*in
   wire signed [14:0] m204_47;
   assign m204_47 =15'b0;

   // m204_48 = W*in
   wire signed [14:0] m204_48;
   assign m204_48 =15'b0;

   // m204_49 = W*in
   wire signed [14:0] m204_49;
   assign m204_49 =15'b0;

   // m204_50 = W*in
   wire signed [14:0] m204_50;
   assign m204_50 =15'b0;

   // m204_51 = W*in
   wire signed [14:0] m204_51;
   assign m204_51 =15'b0;

   // m204_52 = W*in
   wire signed [14:0] m204_52;
   assign m204_52 =15'b0;

   // m204_53 = W*in
   wire signed [14:0] m204_53;
   assign m204_53 =15'b0;

   // m204_54 = W*in
   wire signed [14:0] m204_54;
   assign m204_54 =15'b0;

   // m204_55 = W*in
   wire signed [14:0] m204_55;
   assign m204_55 =15'b0;

   // m204_56 = W*in
   wire signed [14:0] m204_56;
   assign m204_56 =15'b0;

   // m204_57 = W*in
   wire signed [14:0] m204_57;
   assign m204_57 =15'b0;

   // m204_58 = W*in
   wire signed [14:0] m204_58;
   assign m204_58 =15'b0;

   // m204_59 = W*in
   wire signed [14:0] m204_59;
   assign m204_59 ={ {4{in204[14]}} , in204[14:4] };

   // m204_60 = W*in
   wire signed [14:0] m204_60;
   assign m204_60 =15'b0;

   // m204_61 = W*in
   wire signed [14:0] m204_61;
   assign m204_61 ={ {4{in204[14]}} , in204[14:4] };

   // m204_62 = W*in
   wire signed [14:0] m204_62;
   assign m204_62 =15'b0;

   // m204_63 = W*in
   wire signed [14:0] m204_63;
   assign m204_63 =15'b0;

   // m204_64 = W*in
   wire signed [14:0] m204_64;
   assign m204_64 ={ {4{in204[14]}} , in204[14:4] };

   // m204_65 = W*in
   wire signed [14:0] m204_65;
   assign m204_65 =15'b0;

   // m204_66 = W*in
   wire signed [14:0] m204_66;
   assign m204_66 =15'b0;

   // m204_67 = W*in
   wire signed [14:0] m204_67;
   assign m204_67 ={ {4{in204[14]}} , in204[14:4] };

   // m204_68 = W*in
   wire signed [14:0] m204_68;
   assign m204_68 =15'b0;

   // m204_69 = W*in
   wire signed [14:0] m204_69;
   assign m204_69 =15'b0;

   // m204_70 = W*in
   wire signed [14:0] m204_70;
   assign m204_70 =15'b0;

   // m204_71 = W*in
   wire signed [14:0] m204_71;
   assign m204_71 =15'b0;

   // m204_72 = W*in
   wire signed [14:0] m204_72;
   assign m204_72 =15'b0;

   // m204_73 = W*in
   wire signed [14:0] m204_73;
   assign m204_73 =15'b0;

   // m204_74 = W*in
   wire signed [14:0] m204_74;
   assign m204_74 =15'b0;

   // m204_75 = W*in
   wire signed [14:0] m204_75;
   assign m204_75 =15'b0;

   // m204_76 = W*in
   wire signed [14:0] m204_76;
   assign m204_76 =15'b0;

   // m204_77 = W*in
   wire signed [14:0] m204_77;
   assign m204_77 =15'b0;

   // m204_78 = W*in
   wire signed [14:0] m204_78;
   assign m204_78 =15'b0;

   // m204_79 = W*in
   wire signed [14:0] m204_79;
   assign m204_79 =15'b0;

   // m204_80 = W*in
   wire signed [14:0] m204_80;
   assign m204_80 =15'b0;

   // m204_81 = W*in
   wire signed [14:0] m204_81;
   assign m204_81 =15'b0;

   // m204_82 = W*in
   wire signed [14:0] m204_82;
   assign m204_82 =15'b0;

   // m204_83 = W*in
   wire signed [14:0] m204_83;
   assign m204_83 =15'b0;

   // m204_84 = W*in
   wire signed [14:0] m204_84;
   assign m204_84 =15'b0;

   // m204_85 = W*in
   wire signed [14:0] m204_85;
   assign m204_85 =15'b0;

   // m204_86 = W*in
   wire signed [14:0] m204_86;
   assign m204_86 =15'b0;

   // m204_87 = W*in
   wire signed [14:0] m204_87;
   assign m204_87 =15'b0;

   // m204_88 = W*in
   wire signed [14:0] m204_88;
   assign m204_88 =15'b0;

   // m204_89 = W*in
   wire signed [14:0] m204_89;
   assign m204_89 =15'b0;

   // m204_90 = W*in
   wire signed [14:0] m204_90;
   assign m204_90 =15'b0;

   // m204_91 = W*in
   wire signed [14:0] m204_91;
   assign m204_91 =15'b0;

   // m204_92 = W*in
   wire signed [14:0] m204_92;
   assign m204_92 =15'b0;

   // m204_93 = W*in
   wire signed [14:0] m204_93;
   assign m204_93 =15'b0;

   // m204_94 = W*in
   wire signed [14:0] m204_94;
   assign m204_94 =15'b0;

   // m204_95 = W*in
   wire signed [14:0] m204_95;
   assign m204_95 =15'b0;

   // m204_96 = W*in
   wire signed [14:0] m204_96;
   assign m204_96 =15'b0;

   // m204_97 = W*in
   wire signed [14:0] m204_97;
   assign m204_97 =15'b0;

   // m204_98 = W*in
   wire signed [14:0] m204_98;
   assign m204_98 =15'b0;

   // m204_99 = W*in
   wire signed [14:0] m204_99;
   assign m204_99 =15'b0;

   // m204_100 = W*in
   wire signed [14:0] m204_100;
   assign m204_100 =15'b0;

   // m205_1 = W*in
   wire signed [14:0] m205_1;
   assign m205_1 =15'b0;

   // m205_2 = W*in
   wire signed [14:0] m205_2;
   assign m205_2 =15'b0;

   // m205_3 = W*in
   wire signed [14:0] m205_3;
   assign m205_3 =15'b0;

   // m205_4 = W*in
   wire signed [14:0] m205_4;
   assign m205_4 =15'b0;

   // m205_5 = W*in
   wire signed [14:0] m205_5;
   assign m205_5 =15'b0;

   // m205_6 = W*in
   wire signed [14:0] m205_6;
   assign m205_6 =15'b0;

   // m205_7 = W*in
   wire signed [14:0] m205_7;
   assign m205_7 =15'b0;

   // m205_8 = W*in
   wire signed [14:0] m205_8;
   assign m205_8 =15'b0;

   // m205_9 = W*in
   wire signed [14:0] m205_9;
   assign m205_9 =15'b0;

   // m205_10 = W*in
   wire signed [14:0] m205_10;
   assign m205_10 =15'b0;

   // m205_11 = W*in
   wire signed [14:0] m205_11;
   assign m205_11 =15'b0;

   // m205_12 = W*in
   wire signed [14:0] m205_12;
   assign m205_12 =15'b0;

   // m205_13 = W*in
   wire signed [14:0] m205_13;
   assign m205_13 =15'b0;

   // m205_14 = W*in
   wire signed [14:0] m205_14;
   assign m205_14 =15'b0;

   // m205_15 = W*in
   wire signed [14:0] m205_15;
   assign m205_15 =15'b0;

   // m205_16 = W*in
   wire signed [14:0] m205_16;
   assign m205_16 =15'b0;

   // m205_17 = W*in
   wire signed [14:0] m205_17;
   assign m205_17 ={ {4{neg205[14]}} , neg205[14:4] };

   // m205_18 = W*in
   wire signed [14:0] m205_18;
   assign m205_18 =15'b0;

   // m205_19 = W*in
   wire signed [14:0] m205_19;
   assign m205_19 ={ {4{neg205[14]}} , neg205[14:4] };

   // m205_20 = W*in
   wire signed [14:0] m205_20;
   assign m205_20 =15'b0;

   // m205_21 = W*in
   wire signed [14:0] m205_21;
   assign m205_21 =15'b0;

   // m205_22 = W*in
   wire signed [14:0] m205_22;
   assign m205_22 =15'b0;

   // m205_23 = W*in
   wire signed [14:0] m205_23;
   assign m205_23 =15'b0;

   // m205_24 = W*in
   wire signed [14:0] m205_24;
   assign m205_24 =15'b0;

   // m205_25 = W*in
   wire signed [14:0] m205_25;
   assign m205_25 =15'b0;

   // m205_26 = W*in
   wire signed [14:0] m205_26;
   assign m205_26 =15'b0;

   // m205_27 = W*in
   wire signed [14:0] m205_27;
   assign m205_27 ={ {4{in205[14]}} , in205[14:4] };

   // m205_28 = W*in
   wire signed [14:0] m205_28;
   assign m205_28 =15'b0;

   // m205_29 = W*in
   wire signed [14:0] m205_29;
   assign m205_29 =15'b0;

   // m205_30 = W*in
   wire signed [14:0] m205_30;
   assign m205_30 =15'b0;

   // m205_31 = W*in
   wire signed [14:0] m205_31;
   assign m205_31 =15'b0;

   // m205_32 = W*in
   wire signed [14:0] m205_32;
   assign m205_32 =15'b0;

   // m205_33 = W*in
   wire signed [14:0] m205_33;
   assign m205_33 =15'b0;

   // m205_34 = W*in
   wire signed [14:0] m205_34;
   assign m205_34 =15'b0;

   // m205_35 = W*in
   wire signed [14:0] m205_35;
   assign m205_35 =15'b0;

   // m205_36 = W*in
   wire signed [14:0] m205_36;
   assign m205_36 ={ {3{in205[14]}} , in205[14:3] };

   // m205_37 = W*in
   wire signed [14:0] m205_37;
   assign m205_37 =15'b0;

   // m205_38 = W*in
   wire signed [14:0] m205_38;
   assign m205_38 =15'b0;

   // m205_39 = W*in
   wire signed [14:0] m205_39;
   assign m205_39 =15'b0;

   // m205_40 = W*in
   wire signed [14:0] m205_40;
   assign m205_40 =15'b0;

   // m205_41 = W*in
   wire signed [14:0] m205_41;
   assign m205_41 =15'b0;

   // m205_42 = W*in
   wire signed [14:0] m205_42;
   assign m205_42 =15'b0;

   // m205_43 = W*in
   wire signed [14:0] m205_43;
   assign m205_43 ={ {3{neg205[14]}} , neg205[14:3] };

   // m205_44 = W*in
   wire signed [14:0] m205_44;
   assign m205_44 =15'b0;

   // m205_45 = W*in
   wire signed [14:0] m205_45;
   assign m205_45 =15'b0;

   // m205_46 = W*in
   wire signed [14:0] m205_46;
   assign m205_46 =15'b0;

   // m205_47 = W*in
   wire signed [14:0] m205_47;
   assign m205_47 =15'b0;

   // m205_48 = W*in
   wire signed [14:0] m205_48;
   assign m205_48 =15'b0;

   // m205_49 = W*in
   wire signed [14:0] m205_49;
   assign m205_49 =15'b0;

   // m205_50 = W*in
   wire signed [14:0] m205_50;
   assign m205_50 =15'b0;

   // m205_51 = W*in
   wire signed [14:0] m205_51;
   assign m205_51 =15'b0;

   // m205_52 = W*in
   wire signed [14:0] m205_52;
   assign m205_52 =15'b0;

   // m205_53 = W*in
   wire signed [14:0] m205_53;
   assign m205_53 =15'b0;

   // m205_54 = W*in
   wire signed [14:0] m205_54;
   assign m205_54 =15'b0;

   // m205_55 = W*in
   wire signed [14:0] m205_55;
   assign m205_55 =15'b0;

   // m205_56 = W*in
   wire signed [14:0] m205_56;
   assign m205_56 =15'b0;

   // m205_57 = W*in
   wire signed [14:0] m205_57;
   assign m205_57 =15'b0;

   // m205_58 = W*in
   wire signed [14:0] m205_58;
   assign m205_58 =15'b0;

   // m205_59 = W*in
   wire signed [14:0] m205_59;
   assign m205_59 =15'b0;

   // m205_60 = W*in
   wire signed [14:0] m205_60;
   assign m205_60 =15'b0;

   // m205_61 = W*in
   wire signed [14:0] m205_61;
   assign m205_61 =15'b0;

   // m205_62 = W*in
   wire signed [14:0] m205_62;
   assign m205_62 ={ {4{in205[14]}} , in205[14:4] };

   // m205_63 = W*in
   wire signed [14:0] m205_63;
   assign m205_63 =15'b0;

   // m205_64 = W*in
   wire signed [14:0] m205_64;
   assign m205_64 ={ {4{in205[14]}} , in205[14:4] };

   // m205_65 = W*in
   wire signed [14:0] m205_65;
   assign m205_65 =15'b0;

   // m205_66 = W*in
   wire signed [14:0] m205_66;
   assign m205_66 =15'b0;

   // m205_67 = W*in
   wire signed [14:0] m205_67;
   assign m205_67 =15'b0;

   // m205_68 = W*in
   wire signed [14:0] m205_68;
   assign m205_68 =15'b0;

   // m205_69 = W*in
   wire signed [14:0] m205_69;
   assign m205_69 =15'b0;

   // m205_70 = W*in
   wire signed [14:0] m205_70;
   assign m205_70 =15'b0;

   // m205_71 = W*in
   wire signed [14:0] m205_71;
   assign m205_71 =15'b0;

   // m205_72 = W*in
   wire signed [14:0] m205_72;
   assign m205_72 =15'b0;

   // m205_73 = W*in
   wire signed [14:0] m205_73;
   assign m205_73 ={ {3{in205[14]}} , in205[14:3] };

   // m205_74 = W*in
   wire signed [14:0] m205_74;
   assign m205_74 ={ {3{neg205[14]}} , neg205[14:3] };

   // m205_75 = W*in
   wire signed [14:0] m205_75;
   assign m205_75 =15'b0;

   // m205_76 = W*in
   wire signed [14:0] m205_76;
   assign m205_76 =15'b0;

   // m205_77 = W*in
   wire signed [14:0] m205_77;
   assign m205_77 =15'b0;

   // m205_78 = W*in
   wire signed [14:0] m205_78;
   assign m205_78 =15'b0;

   // m205_79 = W*in
   wire signed [14:0] m205_79;
   assign m205_79 =15'b0;

   // m205_80 = W*in
   wire signed [14:0] m205_80;
   assign m205_80 =15'b0;

   // m205_81 = W*in
   wire signed [14:0] m205_81;
   assign m205_81 =15'b0;

   // m205_82 = W*in
   wire signed [14:0] m205_82;
   assign m205_82 =15'b0;

   // m205_83 = W*in
   wire signed [14:0] m205_83;
   assign m205_83 =15'b0;

   // m205_84 = W*in
   wire signed [14:0] m205_84;
   assign m205_84 ={ {3{neg205[14]}} , neg205[14:3] };

   // m205_85 = W*in
   wire signed [14:0] m205_85;
   assign m205_85 =15'b0;

   // m205_86 = W*in
   wire signed [14:0] m205_86;
   assign m205_86 =15'b0;

   // m205_87 = W*in
   wire signed [14:0] m205_87;
   assign m205_87 =15'b0;

   // m205_88 = W*in
   wire signed [14:0] m205_88;
   assign m205_88 =15'b0;

   // m205_89 = W*in
   wire signed [14:0] m205_89;
   assign m205_89 =15'b0;

   // m205_90 = W*in
   wire signed [14:0] m205_90;
   assign m205_90 =15'b0;

   // m205_91 = W*in
   wire signed [14:0] m205_91;
   assign m205_91 =15'b0;

   // m205_92 = W*in
   wire signed [14:0] m205_92;
   assign m205_92 =15'b0;

   // m205_93 = W*in
   wire signed [14:0] m205_93;
   assign m205_93 =15'b0;

   // m205_94 = W*in
   wire signed [14:0] m205_94;
   assign m205_94 =15'b0;

   // m205_95 = W*in
   wire signed [14:0] m205_95;
   assign m205_95 =15'b0;

   // m205_96 = W*in
   wire signed [14:0] m205_96;
   assign m205_96 =15'b0;

   // m205_97 = W*in
   wire signed [14:0] m205_97;
   assign m205_97 ={ {4{in205[14]}} , in205[14:4] };

   // m205_98 = W*in
   wire signed [14:0] m205_98;
   assign m205_98 =15'b0;

   // m205_99 = W*in
   wire signed [14:0] m205_99;
   assign m205_99 =15'b0;

   // m205_100 = W*in
   wire signed [14:0] m205_100;
   assign m205_100 =15'b0;

   // m206_1 = W*in
   wire signed [14:0] m206_1;
   assign m206_1 =15'b0;

   // m206_2 = W*in
   wire signed [14:0] m206_2;
   assign m206_2 =15'b0;

   // m206_3 = W*in
   wire signed [14:0] m206_3;
   assign m206_3 =15'b0;

   // m206_4 = W*in
   wire signed [14:0] m206_4;
   assign m206_4 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_5 = W*in
   wire signed [14:0] m206_5;
   assign m206_5 ={ {2{in206[14]}} , in206[14:2] };

   // m206_6 = W*in
   wire signed [14:0] m206_6;
   assign m206_6 =15'b0;

   // m206_7 = W*in
   wire signed [14:0] m206_7;
   assign m206_7 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_8 = W*in
   wire signed [14:0] m206_8;
   assign m206_8 =15'b0;

   // m206_9 = W*in
   wire signed [14:0] m206_9;
   assign m206_9 =15'b0;

   // m206_10 = W*in
   wire signed [14:0] m206_10;
   assign m206_10 =15'b0;

   // m206_11 = W*in
   wire signed [14:0] m206_11;
   assign m206_11 =15'b0;

   // m206_12 = W*in
   wire signed [14:0] m206_12;
   assign m206_12 ={ {4{in206[14]}} , in206[14:4] };

   // m206_13 = W*in
   wire signed [14:0] m206_13;
   assign m206_13 =15'b0;

   // m206_14 = W*in
   wire signed [14:0] m206_14;
   assign m206_14 =15'b0;

   // m206_15 = W*in
   wire signed [14:0] m206_15;
   assign m206_15 =15'b0;

   // m206_16 = W*in
   wire signed [14:0] m206_16;
   assign m206_16 =15'b0;

   // m206_17 = W*in
   wire signed [14:0] m206_17;
   assign m206_17 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_18 = W*in
   wire signed [14:0] m206_18;
   assign m206_18 =15'b0;

   // m206_19 = W*in
   wire signed [14:0] m206_19;
   assign m206_19 ={ {3{in206[14]}} , in206[14:3] };

   // m206_20 = W*in
   wire signed [14:0] m206_20;
   assign m206_20 =15'b0;

   // m206_21 = W*in
   wire signed [14:0] m206_21;
   assign m206_21 =15'b0;

   // m206_22 = W*in
   wire signed [14:0] m206_22;
   assign m206_22 =15'b0;

   // m206_23 = W*in
   wire signed [14:0] m206_23;
   assign m206_23 =15'b0;

   // m206_24 = W*in
   wire signed [14:0] m206_24;
   assign m206_24 =15'b0;

   // m206_25 = W*in
   wire signed [14:0] m206_25;
   assign m206_25 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_26 = W*in
   wire signed [14:0] m206_26;
   assign m206_26 =15'b0;

   // m206_27 = W*in
   wire signed [14:0] m206_27;
   assign m206_27 =15'b0;

   // m206_28 = W*in
   wire signed [14:0] m206_28;
   assign m206_28 =15'b0;

   // m206_29 = W*in
   wire signed [14:0] m206_29;
   assign m206_29 =15'b0;

   // m206_30 = W*in
   wire signed [14:0] m206_30;
   assign m206_30 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_31 = W*in
   wire signed [14:0] m206_31;
   assign m206_31 =15'b0;

   // m206_32 = W*in
   wire signed [14:0] m206_32;
   assign m206_32 =15'b0;

   // m206_33 = W*in
   wire signed [14:0] m206_33;
   assign m206_33 =15'b0;

   // m206_34 = W*in
   wire signed [14:0] m206_34;
   assign m206_34 =15'b0;

   // m206_35 = W*in
   wire signed [14:0] m206_35;
   assign m206_35 =15'b0;

   // m206_36 = W*in
   wire signed [14:0] m206_36;
   assign m206_36 =15'b0;

   // m206_37 = W*in
   wire signed [14:0] m206_37;
   assign m206_37 =15'b0;

   // m206_38 = W*in
   wire signed [14:0] m206_38;
   assign m206_38 =15'b0;

   // m206_39 = W*in
   wire signed [14:0] m206_39;
   assign m206_39 =15'b0;

   // m206_40 = W*in
   wire signed [14:0] m206_40;
   assign m206_40 =15'b0;

   // m206_41 = W*in
   wire signed [14:0] m206_41;
   assign m206_41 =15'b0;

   // m206_42 = W*in
   wire signed [14:0] m206_42;
   assign m206_42 =15'b0;

   // m206_43 = W*in
   wire signed [14:0] m206_43;
   assign m206_43 ={ {3{neg206[14]}} , neg206[14:3] };

   // m206_44 = W*in
   wire signed [14:0] m206_44;
   assign m206_44 =15'b0;

   // m206_45 = W*in
   wire signed [14:0] m206_45;
   assign m206_45 =15'b0;

   // m206_46 = W*in
   wire signed [14:0] m206_46;
   assign m206_46 =15'b0;

   // m206_47 = W*in
   wire signed [14:0] m206_47;
   assign m206_47 =15'b0;

   // m206_48 = W*in
   wire signed [14:0] m206_48;
   assign m206_48 =15'b0;

   // m206_49 = W*in
   wire signed [14:0] m206_49;
   assign m206_49 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_50 = W*in
   wire signed [14:0] m206_50;
   assign m206_50 =15'b0;

   // m206_51 = W*in
   wire signed [14:0] m206_51;
   assign m206_51 =15'b0;

   // m206_52 = W*in
   wire signed [14:0] m206_52;
   assign m206_52 =15'b0;

   // m206_53 = W*in
   wire signed [14:0] m206_53;
   assign m206_53 =15'b0;

   // m206_54 = W*in
   wire signed [14:0] m206_54;
   assign m206_54 =15'b0;

   // m206_55 = W*in
   wire signed [14:0] m206_55;
   assign m206_55 =15'b0;

   // m206_56 = W*in
   wire signed [14:0] m206_56;
   assign m206_56 =15'b0;

   // m206_57 = W*in
   wire signed [14:0] m206_57;
   assign m206_57 =15'b0;

   // m206_58 = W*in
   wire signed [14:0] m206_58;
   assign m206_58 =15'b0;

   // m206_59 = W*in
   wire signed [14:0] m206_59;
   assign m206_59 =15'b0;

   // m206_60 = W*in
   wire signed [14:0] m206_60;
   assign m206_60 =15'b0;

   // m206_61 = W*in
   wire signed [14:0] m206_61;
   assign m206_61 =15'b0;

   // m206_62 = W*in
   wire signed [14:0] m206_62;
   assign m206_62 ={ {4{in206[14]}} , in206[14:4] };

   // m206_63 = W*in
   wire signed [14:0] m206_63;
   assign m206_63 =15'b0;

   // m206_64 = W*in
   wire signed [14:0] m206_64;
   assign m206_64 =15'b0;

   // m206_65 = W*in
   wire signed [14:0] m206_65;
   assign m206_65 ={ {3{neg206[14]}} , neg206[14:3] };

   // m206_66 = W*in
   wire signed [14:0] m206_66;
   assign m206_66 ={ {3{neg206[14]}} , neg206[14:3] };

   // m206_67 = W*in
   wire signed [14:0] m206_67;
   assign m206_67 =15'b0;

   // m206_68 = W*in
   wire signed [14:0] m206_68;
   assign m206_68 ={ {4{neg206[14]}} , neg206[14:4] };

   // m206_69 = W*in
   wire signed [14:0] m206_69;
   assign m206_69 =15'b0;

   // m206_70 = W*in
   wire signed [14:0] m206_70;
   assign m206_70 =15'b0;

   // m206_71 = W*in
   wire signed [14:0] m206_71;
   assign m206_71 =15'b0;

   // m206_72 = W*in
   wire signed [14:0] m206_72;
   assign m206_72 =15'b0;

   // m206_73 = W*in
   wire signed [14:0] m206_73;
   assign m206_73 =15'b0;

   // m206_74 = W*in
   wire signed [14:0] m206_74;
   assign m206_74 =15'b0;

   // m206_75 = W*in
   wire signed [14:0] m206_75;
   assign m206_75 ={ {4{in206[14]}} , in206[14:4] };

   // m206_76 = W*in
   wire signed [14:0] m206_76;
   assign m206_76 =15'b0;

   // m206_77 = W*in
   wire signed [14:0] m206_77;
   assign m206_77 =15'b0;

   // m206_78 = W*in
   wire signed [14:0] m206_78;
   assign m206_78 =15'b0;

   // m206_79 = W*in
   wire signed [14:0] m206_79;
   assign m206_79 =15'b0;

   // m206_80 = W*in
   wire signed [14:0] m206_80;
   assign m206_80 =15'b0;

   // m206_81 = W*in
   wire signed [14:0] m206_81;
   assign m206_81 =15'b0;

   // m206_82 = W*in
   wire signed [14:0] m206_82;
   assign m206_82 =15'b0;

   // m206_83 = W*in
   wire signed [14:0] m206_83;
   assign m206_83 ={ {3{in206[14]}} , in206[14:3] };

   // m206_84 = W*in
   wire signed [14:0] m206_84;
   assign m206_84 =15'b0;

   // m206_85 = W*in
   wire signed [14:0] m206_85;
   assign m206_85 =15'b0;

   // m206_86 = W*in
   wire signed [14:0] m206_86;
   assign m206_86 =15'b0;

   // m206_87 = W*in
   wire signed [14:0] m206_87;
   assign m206_87 =15'b0;

   // m206_88 = W*in
   wire signed [14:0] m206_88;
   assign m206_88 =15'b0;

   // m206_89 = W*in
   wire signed [14:0] m206_89;
   assign m206_89 =15'b0;

   // m206_90 = W*in
   wire signed [14:0] m206_90;
   assign m206_90 =15'b0;

   // m206_91 = W*in
   wire signed [14:0] m206_91;
   assign m206_91 =15'b0;

   // m206_92 = W*in
   wire signed [14:0] m206_92;
   assign m206_92 =15'b0;

   // m206_93 = W*in
   wire signed [14:0] m206_93;
   assign m206_93 =15'b0;

   // m206_94 = W*in
   wire signed [14:0] m206_94;
   assign m206_94 =15'b0;

   // m206_95 = W*in
   wire signed [14:0] m206_95;
   assign m206_95 =15'b0;

   // m206_96 = W*in
   wire signed [14:0] m206_96;
   assign m206_96 =15'b0;

   // m206_97 = W*in
   wire signed [14:0] m206_97;
   assign m206_97 =15'b0;

   // m206_98 = W*in
   wire signed [14:0] m206_98;
   assign m206_98 =15'b0;

   // m206_99 = W*in
   wire signed [14:0] m206_99;
   assign m206_99 =15'b0;

   // m206_100 = W*in
   wire signed [14:0] m206_100;
   assign m206_100 =15'b0;

   // m207_1 = W*in
   wire signed [14:0] m207_1;
   assign m207_1 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_2 = W*in
   wire signed [14:0] m207_2;
   assign m207_2 =15'b0;

   // m207_3 = W*in
   wire signed [14:0] m207_3;
   assign m207_3 =15'b0;

   // m207_4 = W*in
   wire signed [14:0] m207_4;
   assign m207_4 =15'b0;

   // m207_5 = W*in
   wire signed [14:0] m207_5;
   assign m207_5 =15'b0;

   // m207_6 = W*in
   wire signed [14:0] m207_6;
   assign m207_6 =15'b0;

   // m207_7 = W*in
   wire signed [14:0] m207_7;
   assign m207_7 =15'b0;

   // m207_8 = W*in
   wire signed [14:0] m207_8;
   assign m207_8 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_9 = W*in
   wire signed [14:0] m207_9;
   assign m207_9 =15'b0;

   // m207_10 = W*in
   wire signed [14:0] m207_10;
   assign m207_10 =15'b0;

   // m207_11 = W*in
   wire signed [14:0] m207_11;
   assign m207_11 =15'b0;

   // m207_12 = W*in
   wire signed [14:0] m207_12;
   assign m207_12 ={ {3{in207[14]}} , in207[14:3] };

   // m207_13 = W*in
   wire signed [14:0] m207_13;
   assign m207_13 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_14 = W*in
   wire signed [14:0] m207_14;
   assign m207_14 =15'b0;

   // m207_15 = W*in
   wire signed [14:0] m207_15;
   assign m207_15 =15'b0;

   // m207_16 = W*in
   wire signed [14:0] m207_16;
   assign m207_16 ={ {3{in207[14]}} , in207[14:3] };

   // m207_17 = W*in
   wire signed [14:0] m207_17;
   assign m207_17 =15'b0;

   // m207_18 = W*in
   wire signed [14:0] m207_18;
   assign m207_18 =15'b0;

   // m207_19 = W*in
   wire signed [14:0] m207_19;
   assign m207_19 =15'b0;

   // m207_20 = W*in
   wire signed [14:0] m207_20;
   assign m207_20 ={ {4{neg207[14]}} , neg207[14:4] };

   // m207_21 = W*in
   wire signed [14:0] m207_21;
   assign m207_21 =15'b0;

   // m207_22 = W*in
   wire signed [14:0] m207_22;
   assign m207_22 =15'b0;

   // m207_23 = W*in
   wire signed [14:0] m207_23;
   assign m207_23 =15'b0;

   // m207_24 = W*in
   wire signed [14:0] m207_24;
   assign m207_24 =15'b0;

   // m207_25 = W*in
   wire signed [14:0] m207_25;
   assign m207_25 ={ {3{in207[14]}} , in207[14:3] };

   // m207_26 = W*in
   wire signed [14:0] m207_26;
   assign m207_26 ={ {3{in207[14]}} , in207[14:3] };

   // m207_27 = W*in
   wire signed [14:0] m207_27;
   assign m207_27 =15'b0;

   // m207_28 = W*in
   wire signed [14:0] m207_28;
   assign m207_28 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_29 = W*in
   wire signed [14:0] m207_29;
   assign m207_29 =15'b0;

   // m207_30 = W*in
   wire signed [14:0] m207_30;
   assign m207_30 ={ {3{in207[14]}} , in207[14:3] };

   // m207_31 = W*in
   wire signed [14:0] m207_31;
   assign m207_31 =15'b0;

   // m207_32 = W*in
   wire signed [14:0] m207_32;
   assign m207_32 =15'b0;

   // m207_33 = W*in
   wire signed [14:0] m207_33;
   assign m207_33 =15'b0;

   // m207_34 = W*in
   wire signed [14:0] m207_34;
   assign m207_34 =15'b0;

   // m207_35 = W*in
   wire signed [14:0] m207_35;
   assign m207_35 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_36 = W*in
   wire signed [14:0] m207_36;
   assign m207_36 ={ {3{in207[14]}} , in207[14:3] };

   // m207_37 = W*in
   wire signed [14:0] m207_37;
   assign m207_37 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_38 = W*in
   wire signed [14:0] m207_38;
   assign m207_38 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_39 = W*in
   wire signed [14:0] m207_39;
   assign m207_39 =15'b0;

   // m207_40 = W*in
   wire signed [14:0] m207_40;
   assign m207_40 =15'b0;

   // m207_41 = W*in
   wire signed [14:0] m207_41;
   assign m207_41 =15'b0;

   // m207_42 = W*in
   wire signed [14:0] m207_42;
   assign m207_42 =15'b0;

   // m207_43 = W*in
   wire signed [14:0] m207_43;
   assign m207_43 ={ {3{in207[14]}} , in207[14:3] };

   // m207_44 = W*in
   wire signed [14:0] m207_44;
   assign m207_44 =15'b0;

   // m207_45 = W*in
   wire signed [14:0] m207_45;
   assign m207_45 =15'b0;

   // m207_46 = W*in
   wire signed [14:0] m207_46;
   assign m207_46 =15'b0;

   // m207_47 = W*in
   wire signed [14:0] m207_47;
   assign m207_47 =15'b0;

   // m207_48 = W*in
   wire signed [14:0] m207_48;
   assign m207_48 =15'b0;

   // m207_49 = W*in
   wire signed [14:0] m207_49;
   assign m207_49 ={ {3{in207[14]}} , in207[14:3] };

   // m207_50 = W*in
   wire signed [14:0] m207_50;
   assign m207_50 =15'b0;

   // m207_51 = W*in
   wire signed [14:0] m207_51;
   assign m207_51 =15'b0;

   // m207_52 = W*in
   wire signed [14:0] m207_52;
   assign m207_52 =15'b0;

   // m207_53 = W*in
   wire signed [14:0] m207_53;
   assign m207_53 =15'b0;

   // m207_54 = W*in
   wire signed [14:0] m207_54;
   assign m207_54 =15'b0;

   // m207_55 = W*in
   wire signed [14:0] m207_55;
   assign m207_55 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_56 = W*in
   wire signed [14:0] m207_56;
   assign m207_56 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_57 = W*in
   wire signed [14:0] m207_57;
   assign m207_57 =15'b0;

   // m207_58 = W*in
   wire signed [14:0] m207_58;
   assign m207_58 =15'b0;

   // m207_59 = W*in
   wire signed [14:0] m207_59;
   assign m207_59 =15'b0;

   // m207_60 = W*in
   wire signed [14:0] m207_60;
   assign m207_60 =15'b0;

   // m207_61 = W*in
   wire signed [14:0] m207_61;
   assign m207_61 =15'b0;

   // m207_62 = W*in
   wire signed [14:0] m207_62;
   assign m207_62 =15'b0;

   // m207_63 = W*in
   wire signed [14:0] m207_63;
   assign m207_63 =15'b0;

   // m207_64 = W*in
   wire signed [14:0] m207_64;
   assign m207_64 =15'b0;

   // m207_65 = W*in
   wire signed [14:0] m207_65;
   assign m207_65 =15'b0;

   // m207_66 = W*in
   wire signed [14:0] m207_66;
   assign m207_66 =15'b0;

   // m207_67 = W*in
   wire signed [14:0] m207_67;
   assign m207_67 =15'b0;

   // m207_68 = W*in
   wire signed [14:0] m207_68;
   assign m207_68 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_69 = W*in
   wire signed [14:0] m207_69;
   assign m207_69 ={ {3{in207[14]}} , in207[14:3] };

   // m207_70 = W*in
   wire signed [14:0] m207_70;
   assign m207_70 =15'b0;

   // m207_71 = W*in
   wire signed [14:0] m207_71;
   assign m207_71 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_72 = W*in
   wire signed [14:0] m207_72;
   assign m207_72 =15'b0;

   // m207_73 = W*in
   wire signed [14:0] m207_73;
   assign m207_73 =15'b0;

   // m207_74 = W*in
   wire signed [14:0] m207_74;
   assign m207_74 ={ {4{neg207[14]}} , neg207[14:4] };

   // m207_75 = W*in
   wire signed [14:0] m207_75;
   assign m207_75 =15'b0;

   // m207_76 = W*in
   wire signed [14:0] m207_76;
   assign m207_76 =15'b0;

   // m207_77 = W*in
   wire signed [14:0] m207_77;
   assign m207_77 =15'b0;

   // m207_78 = W*in
   wire signed [14:0] m207_78;
   assign m207_78 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_79 = W*in
   wire signed [14:0] m207_79;
   assign m207_79 ={ {3{in207[14]}} , in207[14:3] };

   // m207_80 = W*in
   wire signed [14:0] m207_80;
   assign m207_80 =15'b0;

   // m207_81 = W*in
   wire signed [14:0] m207_81;
   assign m207_81 =15'b0;

   // m207_82 = W*in
   wire signed [14:0] m207_82;
   assign m207_82 =15'b0;

   // m207_83 = W*in
   wire signed [14:0] m207_83;
   assign m207_83 ={ {3{neg207[14]}} , neg207[14:3] };

   // m207_84 = W*in
   wire signed [14:0] m207_84;
   assign m207_84 =15'b0;

   // m207_85 = W*in
   wire signed [14:0] m207_85;
   assign m207_85 =15'b0;

   // m207_86 = W*in
   wire signed [14:0] m207_86;
   assign m207_86 =15'b0;

   // m207_87 = W*in
   wire signed [14:0] m207_87;
   assign m207_87 =15'b0;

   // m207_88 = W*in
   wire signed [14:0] m207_88;
   assign m207_88 =15'b0;

   // m207_89 = W*in
   wire signed [14:0] m207_89;
   assign m207_89 ={ {4{neg207[14]}} , neg207[14:4] };

   // m207_90 = W*in
   wire signed [14:0] m207_90;
   assign m207_90 =15'b0;

   // m207_91 = W*in
   wire signed [14:0] m207_91;
   assign m207_91 ={ {4{in207[14]}} , in207[14:4] };

   // m207_92 = W*in
   wire signed [14:0] m207_92;
   assign m207_92 ={ {3{in207[14]}} , in207[14:3] };

   // m207_93 = W*in
   wire signed [14:0] m207_93;
   assign m207_93 =15'b0;

   // m207_94 = W*in
   wire signed [14:0] m207_94;
   assign m207_94 =15'b0;

   // m207_95 = W*in
   wire signed [14:0] m207_95;
   assign m207_95 =15'b0;

   // m207_96 = W*in
   wire signed [14:0] m207_96;
   assign m207_96 =15'b0;

   // m207_97 = W*in
   wire signed [14:0] m207_97;
   assign m207_97 =15'b0;

   // m207_98 = W*in
   wire signed [14:0] m207_98;
   assign m207_98 =15'b0;

   // m207_99 = W*in
   wire signed [14:0] m207_99;
   assign m207_99 =15'b0;

   // m207_100 = W*in
   wire signed [14:0] m207_100;
   assign m207_100 =15'b0;

   // m208_1 = W*in
   wire signed [14:0] m208_1;
   assign m208_1 =15'b0;

   // m208_2 = W*in
   wire signed [14:0] m208_2;
   assign m208_2 =15'b0;

   // m208_3 = W*in
   wire signed [14:0] m208_3;
   assign m208_3 =15'b0;

   // m208_4 = W*in
   wire signed [14:0] m208_4;
   assign m208_4 =15'b0;

   // m208_5 = W*in
   wire signed [14:0] m208_5;
   assign m208_5 =15'b0;

   // m208_6 = W*in
   wire signed [14:0] m208_6;
   assign m208_6 =15'b0;

   // m208_7 = W*in
   wire signed [14:0] m208_7;
   assign m208_7 =15'b0;

   // m208_8 = W*in
   wire signed [14:0] m208_8;
   assign m208_8 =15'b0;

   // m208_9 = W*in
   wire signed [14:0] m208_9;
   assign m208_9 =15'b0;

   // m208_10 = W*in
   wire signed [14:0] m208_10;
   assign m208_10 =15'b0;

   // m208_11 = W*in
   wire signed [14:0] m208_11;
   assign m208_11 =15'b0;

   // m208_12 = W*in
   wire signed [14:0] m208_12;
   assign m208_12 =15'b0;

   // m208_13 = W*in
   wire signed [14:0] m208_13;
   assign m208_13 =15'b0;

   // m208_14 = W*in
   wire signed [14:0] m208_14;
   assign m208_14 =15'b0;

   // m208_15 = W*in
   wire signed [14:0] m208_15;
   assign m208_15 =15'b0;

   // m208_16 = W*in
   wire signed [14:0] m208_16;
   assign m208_16 =15'b0;

   // m208_17 = W*in
   wire signed [14:0] m208_17;
   assign m208_17 =15'b0;

   // m208_18 = W*in
   wire signed [14:0] m208_18;
   assign m208_18 =15'b0;

   // m208_19 = W*in
   wire signed [14:0] m208_19;
   assign m208_19 =15'b0;

   // m208_20 = W*in
   wire signed [14:0] m208_20;
   assign m208_20 =15'b0;

   // m208_21 = W*in
   wire signed [14:0] m208_21;
   assign m208_21 =15'b0;

   // m208_22 = W*in
   wire signed [14:0] m208_22;
   assign m208_22 =15'b0;

   // m208_23 = W*in
   wire signed [14:0] m208_23;
   assign m208_23 =15'b0;

   // m208_24 = W*in
   wire signed [14:0] m208_24;
   assign m208_24 =15'b0;

   // m208_25 = W*in
   wire signed [14:0] m208_25;
   assign m208_25 =15'b0;

   // m208_26 = W*in
   wire signed [14:0] m208_26;
   assign m208_26 =15'b0;

   // m208_27 = W*in
   wire signed [14:0] m208_27;
   assign m208_27 =15'b0;

   // m208_28 = W*in
   wire signed [14:0] m208_28;
   assign m208_28 =15'b0;

   // m208_29 = W*in
   wire signed [14:0] m208_29;
   assign m208_29 ={ {4{neg208[14]}} , neg208[14:4] };

   // m208_30 = W*in
   wire signed [14:0] m208_30;
   assign m208_30 ={ {3{neg208[14]}} , neg208[14:3] };

   // m208_31 = W*in
   wire signed [14:0] m208_31;
   assign m208_31 =15'b0;

   // m208_32 = W*in
   wire signed [14:0] m208_32;
   assign m208_32 ={ {3{in208[14]}} , in208[14:3] };

   // m208_33 = W*in
   wire signed [14:0] m208_33;
   assign m208_33 =15'b0;

   // m208_34 = W*in
   wire signed [14:0] m208_34;
   assign m208_34 =15'b0;

   // m208_35 = W*in
   wire signed [14:0] m208_35;
   assign m208_35 =15'b0;

   // m208_36 = W*in
   wire signed [14:0] m208_36;
   assign m208_36 =15'b0;

   // m208_37 = W*in
   wire signed [14:0] m208_37;
   assign m208_37 =15'b0;

   // m208_38 = W*in
   wire signed [14:0] m208_38;
   assign m208_38 =15'b0;

   // m208_39 = W*in
   wire signed [14:0] m208_39;
   assign m208_39 =15'b0;

   // m208_40 = W*in
   wire signed [14:0] m208_40;
   assign m208_40 =15'b0;

   // m208_41 = W*in
   wire signed [14:0] m208_41;
   assign m208_41 ={ {4{neg208[14]}} , neg208[14:4] };

   // m208_42 = W*in
   wire signed [14:0] m208_42;
   assign m208_42 =15'b0;

   // m208_43 = W*in
   wire signed [14:0] m208_43;
   assign m208_43 =15'b0;

   // m208_44 = W*in
   wire signed [14:0] m208_44;
   assign m208_44 =15'b0;

   // m208_45 = W*in
   wire signed [14:0] m208_45;
   assign m208_45 =15'b0;

   // m208_46 = W*in
   wire signed [14:0] m208_46;
   assign m208_46 ={ {4{in208[14]}} , in208[14:4] };

   // m208_47 = W*in
   wire signed [14:0] m208_47;
   assign m208_47 =15'b0;

   // m208_48 = W*in
   wire signed [14:0] m208_48;
   assign m208_48 =15'b0;

   // m208_49 = W*in
   wire signed [14:0] m208_49;
   assign m208_49 =15'b0;

   // m208_50 = W*in
   wire signed [14:0] m208_50;
   assign m208_50 =15'b0;

   // m208_51 = W*in
   wire signed [14:0] m208_51;
   assign m208_51 =15'b0;

   // m208_52 = W*in
   wire signed [14:0] m208_52;
   assign m208_52 =15'b0;

   // m208_53 = W*in
   wire signed [14:0] m208_53;
   assign m208_53 =15'b0;

   // m208_54 = W*in
   wire signed [14:0] m208_54;
   assign m208_54 =15'b0;

   // m208_55 = W*in
   wire signed [14:0] m208_55;
   assign m208_55 =15'b0;

   // m208_56 = W*in
   wire signed [14:0] m208_56;
   assign m208_56 ={ {3{in208[14]}} , in208[14:3] };

   // m208_57 = W*in
   wire signed [14:0] m208_57;
   assign m208_57 =15'b0;

   // m208_58 = W*in
   wire signed [14:0] m208_58;
   assign m208_58 =15'b0;

   // m208_59 = W*in
   wire signed [14:0] m208_59;
   assign m208_59 =15'b0;

   // m208_60 = W*in
   wire signed [14:0] m208_60;
   assign m208_60 =15'b0;

   // m208_61 = W*in
   wire signed [14:0] m208_61;
   assign m208_61 =15'b0;

   // m208_62 = W*in
   wire signed [14:0] m208_62;
   assign m208_62 =15'b0;

   // m208_63 = W*in
   wire signed [14:0] m208_63;
   assign m208_63 =15'b0;

   // m208_64 = W*in
   wire signed [14:0] m208_64;
   assign m208_64 =15'b0;

   // m208_65 = W*in
   wire signed [14:0] m208_65;
   assign m208_65 =15'b0;

   // m208_66 = W*in
   wire signed [14:0] m208_66;
   assign m208_66 =15'b0;

   // m208_67 = W*in
   wire signed [14:0] m208_67;
   assign m208_67 =15'b0;

   // m208_68 = W*in
   wire signed [14:0] m208_68;
   assign m208_68 =15'b0;

   // m208_69 = W*in
   wire signed [14:0] m208_69;
   assign m208_69 =15'b0;

   // m208_70 = W*in
   wire signed [14:0] m208_70;
   assign m208_70 =15'b0;

   // m208_71 = W*in
   wire signed [14:0] m208_71;
   assign m208_71 =15'b0;

   // m208_72 = W*in
   wire signed [14:0] m208_72;
   assign m208_72 =15'b0;

   // m208_73 = W*in
   wire signed [14:0] m208_73;
   assign m208_73 =15'b0;

   // m208_74 = W*in
   wire signed [14:0] m208_74;
   assign m208_74 =15'b0;

   // m208_75 = W*in
   wire signed [14:0] m208_75;
   assign m208_75 =15'b0;

   // m208_76 = W*in
   wire signed [14:0] m208_76;
   assign m208_76 ={ {3{neg208[14]}} , neg208[14:3] };

   // m208_77 = W*in
   wire signed [14:0] m208_77;
   assign m208_77 =15'b0;

   // m208_78 = W*in
   wire signed [14:0] m208_78;
   assign m208_78 ={ {4{neg208[14]}} , neg208[14:4] };

   // m208_79 = W*in
   wire signed [14:0] m208_79;
   assign m208_79 =15'b0;

   // m208_80 = W*in
   wire signed [14:0] m208_80;
   assign m208_80 =15'b0;

   // m208_81 = W*in
   wire signed [14:0] m208_81;
   assign m208_81 =15'b0;

   // m208_82 = W*in
   wire signed [14:0] m208_82;
   assign m208_82 =15'b0;

   // m208_83 = W*in
   wire signed [14:0] m208_83;
   assign m208_83 ={ {4{in208[14]}} , in208[14:4] };

   // m208_84 = W*in
   wire signed [14:0] m208_84;
   assign m208_84 =15'b0;

   // m208_85 = W*in
   wire signed [14:0] m208_85;
   assign m208_85 =15'b0;

   // m208_86 = W*in
   wire signed [14:0] m208_86;
   assign m208_86 =15'b0;

   // m208_87 = W*in
   wire signed [14:0] m208_87;
   assign m208_87 =15'b0;

   // m208_88 = W*in
   wire signed [14:0] m208_88;
   assign m208_88 =15'b0;

   // m208_89 = W*in
   wire signed [14:0] m208_89;
   assign m208_89 =15'b0;

   // m208_90 = W*in
   wire signed [14:0] m208_90;
   assign m208_90 =15'b0;

   // m208_91 = W*in
   wire signed [14:0] m208_91;
   assign m208_91 =15'b0;

   // m208_92 = W*in
   wire signed [14:0] m208_92;
   assign m208_92 ={ {3{in208[14]}} , in208[14:3] };

   // m208_93 = W*in
   wire signed [14:0] m208_93;
   assign m208_93 =15'b0;

   // m208_94 = W*in
   wire signed [14:0] m208_94;
   assign m208_94 ={ {3{in208[14]}} , in208[14:3] };

   // m208_95 = W*in
   wire signed [14:0] m208_95;
   assign m208_95 =15'b0;

   // m208_96 = W*in
   wire signed [14:0] m208_96;
   assign m208_96 =15'b0;

   // m208_97 = W*in
   wire signed [14:0] m208_97;
   assign m208_97 =15'b0;

   // m208_98 = W*in
   wire signed [14:0] m208_98;
   assign m208_98 =15'b0;

   // m208_99 = W*in
   wire signed [14:0] m208_99;
   assign m208_99 =15'b0;

   // m208_100 = W*in
   wire signed [14:0] m208_100;
   assign m208_100 =15'b0;

   // m209_1 = W*in
   wire signed [14:0] m209_1;
   assign m209_1 =15'b0;

   // m209_2 = W*in
   wire signed [14:0] m209_2;
   assign m209_2 ={ {3{in209[14]}} , in209[14:3] };

   // m209_3 = W*in
   wire signed [14:0] m209_3;
   assign m209_3 =15'b0;

   // m209_4 = W*in
   wire signed [14:0] m209_4;
   assign m209_4 ={ {3{in209[14]}} , in209[14:3] };

   // m209_5 = W*in
   wire signed [14:0] m209_5;
   assign m209_5 =15'b0;

   // m209_6 = W*in
   wire signed [14:0] m209_6;
   assign m209_6 =15'b0;

   // m209_7 = W*in
   wire signed [14:0] m209_7;
   assign m209_7 =15'b0;

   // m209_8 = W*in
   wire signed [14:0] m209_8;
   assign m209_8 =15'b0;

   // m209_9 = W*in
   wire signed [14:0] m209_9;
   assign m209_9 =15'b0;

   // m209_10 = W*in
   wire signed [14:0] m209_10;
   assign m209_10 =15'b0;

   // m209_11 = W*in
   wire signed [14:0] m209_11;
   assign m209_11 =15'b0;

   // m209_12 = W*in
   wire signed [14:0] m209_12;
   assign m209_12 =15'b0;

   // m209_13 = W*in
   wire signed [14:0] m209_13;
   assign m209_13 ={ {2{in209[14]}} , in209[14:2] };

   // m209_14 = W*in
   wire signed [14:0] m209_14;
   assign m209_14 =15'b0;

   // m209_15 = W*in
   wire signed [14:0] m209_15;
   assign m209_15 =15'b0;

   // m209_16 = W*in
   wire signed [14:0] m209_16;
   assign m209_16 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_17 = W*in
   wire signed [14:0] m209_17;
   assign m209_17 ={ {4{in209[14]}} , in209[14:4] };

   // m209_18 = W*in
   wire signed [14:0] m209_18;
   assign m209_18 ={ {3{in209[14]}} , in209[14:3] };

   // m209_19 = W*in
   wire signed [14:0] m209_19;
   assign m209_19 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_20 = W*in
   wire signed [14:0] m209_20;
   assign m209_20 ={ {4{in209[14]}} , in209[14:4] };

   // m209_21 = W*in
   wire signed [14:0] m209_21;
   assign m209_21 ={ {3{in209[14]}} , in209[14:3] };

   // m209_22 = W*in
   wire signed [14:0] m209_22;
   assign m209_22 ={ {3{in209[14]}} , in209[14:3] };

   // m209_23 = W*in
   wire signed [14:0] m209_23;
   assign m209_23 =15'b0;

   // m209_24 = W*in
   wire signed [14:0] m209_24;
   assign m209_24 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_25 = W*in
   wire signed [14:0] m209_25;
   assign m209_25 ={ {3{in209[14]}} , in209[14:3] };

   // m209_26 = W*in
   wire signed [14:0] m209_26;
   assign m209_26 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_27 = W*in
   wire signed [14:0] m209_27;
   assign m209_27 =15'b0;

   // m209_28 = W*in
   wire signed [14:0] m209_28;
   assign m209_28 ={ {3{in209[14]}} , in209[14:3] };

   // m209_29 = W*in
   wire signed [14:0] m209_29;
   assign m209_29 =15'b0;

   // m209_30 = W*in
   wire signed [14:0] m209_30;
   assign m209_30 =15'b0;

   // m209_31 = W*in
   wire signed [14:0] m209_31;
   assign m209_31 =15'b0;

   // m209_32 = W*in
   wire signed [14:0] m209_32;
   assign m209_32 ={ {4{neg209[14]}} , neg209[14:4] };

   // m209_33 = W*in
   wire signed [14:0] m209_33;
   assign m209_33 =15'b0;

   // m209_34 = W*in
   wire signed [14:0] m209_34;
   assign m209_34 ={ {3{in209[14]}} , in209[14:3] };

   // m209_35 = W*in
   wire signed [14:0] m209_35;
   assign m209_35 =15'b0;

   // m209_36 = W*in
   wire signed [14:0] m209_36;
   assign m209_36 =15'b0;

   // m209_37 = W*in
   wire signed [14:0] m209_37;
   assign m209_37 =15'b0;

   // m209_38 = W*in
   wire signed [14:0] m209_38;
   assign m209_38 ={ {3{in209[14]}} , in209[14:3] };

   // m209_39 = W*in
   wire signed [14:0] m209_39;
   assign m209_39 =15'b0;

   // m209_40 = W*in
   wire signed [14:0] m209_40;
   assign m209_40 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_41 = W*in
   wire signed [14:0] m209_41;
   assign m209_41 =15'b0;

   // m209_42 = W*in
   wire signed [14:0] m209_42;
   assign m209_42 =15'b0;

   // m209_43 = W*in
   wire signed [14:0] m209_43;
   assign m209_43 =15'b0;

   // m209_44 = W*in
   wire signed [14:0] m209_44;
   assign m209_44 =15'b0;

   // m209_45 = W*in
   wire signed [14:0] m209_45;
   assign m209_45 =15'b0;

   // m209_46 = W*in
   wire signed [14:0] m209_46;
   assign m209_46 ={ {4{neg209[14]}} , neg209[14:4] };

   // m209_47 = W*in
   wire signed [14:0] m209_47;
   assign m209_47 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_48 = W*in
   wire signed [14:0] m209_48;
   assign m209_48 ={ {4{neg209[14]}} , neg209[14:4] };

   // m209_49 = W*in
   wire signed [14:0] m209_49;
   assign m209_49 =15'b0;

   // m209_50 = W*in
   wire signed [14:0] m209_50;
   assign m209_50 =15'b0;

   // m209_51 = W*in
   wire signed [14:0] m209_51;
   assign m209_51 =15'b0;

   // m209_52 = W*in
   wire signed [14:0] m209_52;
   assign m209_52 =15'b0;

   // m209_53 = W*in
   wire signed [14:0] m209_53;
   assign m209_53 =15'b0;

   // m209_54 = W*in
   wire signed [14:0] m209_54;
   assign m209_54 =15'b0;

   // m209_55 = W*in
   wire signed [14:0] m209_55;
   assign m209_55 =15'b0;

   // m209_56 = W*in
   wire signed [14:0] m209_56;
   assign m209_56 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_57 = W*in
   wire signed [14:0] m209_57;
   assign m209_57 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_58 = W*in
   wire signed [14:0] m209_58;
   assign m209_58 =15'b0;

   // m209_59 = W*in
   wire signed [14:0] m209_59;
   assign m209_59 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_60 = W*in
   wire signed [14:0] m209_60;
   assign m209_60 ={ {4{in209[14]}} , in209[14:4] };

   // m209_61 = W*in
   wire signed [14:0] m209_61;
   assign m209_61 =15'b0;

   // m209_62 = W*in
   wire signed [14:0] m209_62;
   assign m209_62 =15'b0;

   // m209_63 = W*in
   wire signed [14:0] m209_63;
   assign m209_63 =15'b0;

   // m209_64 = W*in
   wire signed [14:0] m209_64;
   assign m209_64 =15'b0;

   // m209_65 = W*in
   wire signed [14:0] m209_65;
   assign m209_65 =15'b0;

   // m209_66 = W*in
   wire signed [14:0] m209_66;
   assign m209_66 =15'b0;

   // m209_67 = W*in
   wire signed [14:0] m209_67;
   assign m209_67 =15'b0;

   // m209_68 = W*in
   wire signed [14:0] m209_68;
   assign m209_68 =15'b0;

   // m209_69 = W*in
   wire signed [14:0] m209_69;
   assign m209_69 =15'b0;

   // m209_70 = W*in
   wire signed [14:0] m209_70;
   assign m209_70 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_71 = W*in
   wire signed [14:0] m209_71;
   assign m209_71 =15'b0;

   // m209_72 = W*in
   wire signed [14:0] m209_72;
   assign m209_72 ={ {3{in209[14]}} , in209[14:3] };

   // m209_73 = W*in
   wire signed [14:0] m209_73;
   assign m209_73 =15'b0;

   // m209_74 = W*in
   wire signed [14:0] m209_74;
   assign m209_74 ={ {4{neg209[14]}} , neg209[14:4] };

   // m209_75 = W*in
   wire signed [14:0] m209_75;
   assign m209_75 =15'b0;

   // m209_76 = W*in
   wire signed [14:0] m209_76;
   assign m209_76 =15'b0;

   // m209_77 = W*in
   wire signed [14:0] m209_77;
   assign m209_77 =15'b0;

   // m209_78 = W*in
   wire signed [14:0] m209_78;
   assign m209_78 ={ {3{in209[14]}} , in209[14:3] };

   // m209_79 = W*in
   wire signed [14:0] m209_79;
   assign m209_79 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_80 = W*in
   wire signed [14:0] m209_80;
   assign m209_80 =15'b0;

   // m209_81 = W*in
   wire signed [14:0] m209_81;
   assign m209_81 =15'b0;

   // m209_82 = W*in
   wire signed [14:0] m209_82;
   assign m209_82 ={ {3{in209[14]}} , in209[14:3] };

   // m209_83 = W*in
   wire signed [14:0] m209_83;
   assign m209_83 =15'b0;

   // m209_84 = W*in
   wire signed [14:0] m209_84;
   assign m209_84 =15'b0;

   // m209_85 = W*in
   wire signed [14:0] m209_85;
   assign m209_85 =15'b0;

   // m209_86 = W*in
   wire signed [14:0] m209_86;
   assign m209_86 =15'b0;

   // m209_87 = W*in
   wire signed [14:0] m209_87;
   assign m209_87 =15'b0;

   // m209_88 = W*in
   wire signed [14:0] m209_88;
   assign m209_88 =15'b0;

   // m209_89 = W*in
   wire signed [14:0] m209_89;
   assign m209_89 =15'b0;

   // m209_90 = W*in
   wire signed [14:0] m209_90;
   assign m209_90 =15'b0;

   // m209_91 = W*in
   wire signed [14:0] m209_91;
   assign m209_91 =15'b0;

   // m209_92 = W*in
   wire signed [14:0] m209_92;
   assign m209_92 =15'b0;

   // m209_93 = W*in
   wire signed [14:0] m209_93;
   assign m209_93 =15'b0;

   // m209_94 = W*in
   wire signed [14:0] m209_94;
   assign m209_94 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_95 = W*in
   wire signed [14:0] m209_95;
   assign m209_95 =15'b0;

   // m209_96 = W*in
   wire signed [14:0] m209_96;
   assign m209_96 ={ {3{in209[14]}} , in209[14:3] };

   // m209_97 = W*in
   wire signed [14:0] m209_97;
   assign m209_97 =15'b0;

   // m209_98 = W*in
   wire signed [14:0] m209_98;
   assign m209_98 ={ {3{neg209[14]}} , neg209[14:3] };

   // m209_99 = W*in
   wire signed [14:0] m209_99;
   assign m209_99 =15'b0;

   // m209_100 = W*in
   wire signed [14:0] m209_100;
   assign m209_100 =15'b0;

   // m210_1 = W*in
   wire signed [14:0] m210_1;
   assign m210_1 =15'b0;

   // m210_2 = W*in
   wire signed [14:0] m210_2;
   assign m210_2 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_3 = W*in
   wire signed [14:0] m210_3;
   assign m210_3 ={ {4{neg210[14]}} , neg210[14:4] };

   // m210_4 = W*in
   wire signed [14:0] m210_4;
   assign m210_4 ={ {3{in210[14]}} , in210[14:3] };

   // m210_5 = W*in
   wire signed [14:0] m210_5;
   assign m210_5 =15'b0;

   // m210_6 = W*in
   wire signed [14:0] m210_6;
   assign m210_6 ={ {3{in210[14]}} , in210[14:3] };

   // m210_7 = W*in
   wire signed [14:0] m210_7;
   assign m210_7 =15'b0;

   // m210_8 = W*in
   wire signed [14:0] m210_8;
   assign m210_8 ={ {3{in210[14]}} , in210[14:3] };

   // m210_9 = W*in
   wire signed [14:0] m210_9;
   assign m210_9 ={ {3{in210[14]}} , in210[14:3] };

   // m210_10 = W*in
   wire signed [14:0] m210_10;
   assign m210_10 =15'b0;

   // m210_11 = W*in
   wire signed [14:0] m210_11;
   assign m210_11 =15'b0;

   // m210_12 = W*in
   wire signed [14:0] m210_12;
   assign m210_12 =15'b0;

   // m210_13 = W*in
   wire signed [14:0] m210_13;
   assign m210_13 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_14 = W*in
   wire signed [14:0] m210_14;
   assign m210_14 =15'b0;

   // m210_15 = W*in
   wire signed [14:0] m210_15;
   assign m210_15 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_16 = W*in
   wire signed [14:0] m210_16;
   assign m210_16 =15'b0;

   // m210_17 = W*in
   wire signed [14:0] m210_17;
   assign m210_17 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_18 = W*in
   wire signed [14:0] m210_18;
   assign m210_18 =15'b0;

   // m210_19 = W*in
   wire signed [14:0] m210_19;
   assign m210_19 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_20 = W*in
   wire signed [14:0] m210_20;
   assign m210_20 =15'b0;

   // m210_21 = W*in
   wire signed [14:0] m210_21;
   assign m210_21 =15'b0;

   // m210_22 = W*in
   wire signed [14:0] m210_22;
   assign m210_22 =15'b0;

   // m210_23 = W*in
   wire signed [14:0] m210_23;
   assign m210_23 =15'b0;

   // m210_24 = W*in
   wire signed [14:0] m210_24;
   assign m210_24 ={ {3{in210[14]}} , in210[14:3] };

   // m210_25 = W*in
   wire signed [14:0] m210_25;
   assign m210_25 ={ {3{in210[14]}} , in210[14:3] };

   // m210_26 = W*in
   wire signed [14:0] m210_26;
   assign m210_26 =15'b0;

   // m210_27 = W*in
   wire signed [14:0] m210_27;
   assign m210_27 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_28 = W*in
   wire signed [14:0] m210_28;
   assign m210_28 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_29 = W*in
   wire signed [14:0] m210_29;
   assign m210_29 ={ {3{in210[14]}} , in210[14:3] };

   // m210_30 = W*in
   wire signed [14:0] m210_30;
   assign m210_30 =15'b0;

   // m210_31 = W*in
   wire signed [14:0] m210_31;
   assign m210_31 ={ {3{in210[14]}} , in210[14:3] };

   // m210_32 = W*in
   wire signed [14:0] m210_32;
   assign m210_32 =15'b0;

   // m210_33 = W*in
   wire signed [14:0] m210_33;
   assign m210_33 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_34 = W*in
   wire signed [14:0] m210_34;
   assign m210_34 ={ {3{in210[14]}} , in210[14:3] };

   // m210_35 = W*in
   wire signed [14:0] m210_35;
   assign m210_35 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_36 = W*in
   wire signed [14:0] m210_36;
   assign m210_36 =15'b0;

   // m210_37 = W*in
   wire signed [14:0] m210_37;
   assign m210_37 =15'b0;

   // m210_38 = W*in
   wire signed [14:0] m210_38;
   assign m210_38 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_39 = W*in
   wire signed [14:0] m210_39;
   assign m210_39 =15'b0;

   // m210_40 = W*in
   wire signed [14:0] m210_40;
   assign m210_40 =15'b0;

   // m210_41 = W*in
   wire signed [14:0] m210_41;
   assign m210_41 ={ {3{in210[14]}} , in210[14:3] };

   // m210_42 = W*in
   wire signed [14:0] m210_42;
   assign m210_42 =15'b0;

   // m210_43 = W*in
   wire signed [14:0] m210_43;
   assign m210_43 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_44 = W*in
   wire signed [14:0] m210_44;
   assign m210_44 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_45 = W*in
   wire signed [14:0] m210_45;
   assign m210_45 =15'b0;

   // m210_46 = W*in
   wire signed [14:0] m210_46;
   assign m210_46 =15'b0;

   // m210_47 = W*in
   wire signed [14:0] m210_47;
   assign m210_47 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_48 = W*in
   wire signed [14:0] m210_48;
   assign m210_48 =15'b0;

   // m210_49 = W*in
   wire signed [14:0] m210_49;
   assign m210_49 =15'b0;

   // m210_50 = W*in
   wire signed [14:0] m210_50;
   assign m210_50 =15'b0;

   // m210_51 = W*in
   wire signed [14:0] m210_51;
   assign m210_51 =15'b0;

   // m210_52 = W*in
   wire signed [14:0] m210_52;
   assign m210_52 =15'b0;

   // m210_53 = W*in
   wire signed [14:0] m210_53;
   assign m210_53 =15'b0;

   // m210_54 = W*in
   wire signed [14:0] m210_54;
   assign m210_54 =15'b0;

   // m210_55 = W*in
   wire signed [14:0] m210_55;
   assign m210_55 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_56 = W*in
   wire signed [14:0] m210_56;
   assign m210_56 =15'b0;

   // m210_57 = W*in
   wire signed [14:0] m210_57;
   assign m210_57 =15'b0;

   // m210_58 = W*in
   wire signed [14:0] m210_58;
   assign m210_58 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_59 = W*in
   wire signed [14:0] m210_59;
   assign m210_59 =15'b0;

   // m210_60 = W*in
   wire signed [14:0] m210_60;
   assign m210_60 ={ {3{in210[14]}} , in210[14:3] };

   // m210_61 = W*in
   wire signed [14:0] m210_61;
   assign m210_61 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_62 = W*in
   wire signed [14:0] m210_62;
   assign m210_62 =15'b0;

   // m210_63 = W*in
   wire signed [14:0] m210_63;
   assign m210_63 =15'b0;

   // m210_64 = W*in
   wire signed [14:0] m210_64;
   assign m210_64 =15'b0;

   // m210_65 = W*in
   wire signed [14:0] m210_65;
   assign m210_65 =15'b0;

   // m210_66 = W*in
   wire signed [14:0] m210_66;
   assign m210_66 =15'b0;

   // m210_67 = W*in
   wire signed [14:0] m210_67;
   assign m210_67 =15'b0;

   // m210_68 = W*in
   wire signed [14:0] m210_68;
   assign m210_68 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_69 = W*in
   wire signed [14:0] m210_69;
   assign m210_69 =15'b0;

   // m210_70 = W*in
   wire signed [14:0] m210_70;
   assign m210_70 =15'b0;

   // m210_71 = W*in
   wire signed [14:0] m210_71;
   assign m210_71 =15'b0;

   // m210_72 = W*in
   wire signed [14:0] m210_72;
   assign m210_72 =15'b0;

   // m210_73 = W*in
   wire signed [14:0] m210_73;
   assign m210_73 =15'b0;

   // m210_74 = W*in
   wire signed [14:0] m210_74;
   assign m210_74 =15'b0;

   // m210_75 = W*in
   wire signed [14:0] m210_75;
   assign m210_75 =15'b0;

   // m210_76 = W*in
   wire signed [14:0] m210_76;
   assign m210_76 =15'b0;

   // m210_77 = W*in
   wire signed [14:0] m210_77;
   assign m210_77 =15'b0;

   // m210_78 = W*in
   wire signed [14:0] m210_78;
   assign m210_78 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_79 = W*in
   wire signed [14:0] m210_79;
   assign m210_79 ={ {3{in210[14]}} , in210[14:3] };

   // m210_80 = W*in
   wire signed [14:0] m210_80;
   assign m210_80 ={ {3{in210[14]}} , in210[14:3] };

   // m210_81 = W*in
   wire signed [14:0] m210_81;
   assign m210_81 =15'b0;

   // m210_82 = W*in
   wire signed [14:0] m210_82;
   assign m210_82 =15'b0;

   // m210_83 = W*in
   wire signed [14:0] m210_83;
   assign m210_83 =15'b0;

   // m210_84 = W*in
   wire signed [14:0] m210_84;
   assign m210_84 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_85 = W*in
   wire signed [14:0] m210_85;
   assign m210_85 =15'b0;

   // m210_86 = W*in
   wire signed [14:0] m210_86;
   assign m210_86 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_87 = W*in
   wire signed [14:0] m210_87;
   assign m210_87 =15'b0;

   // m210_88 = W*in
   wire signed [14:0] m210_88;
   assign m210_88 =15'b0;

   // m210_89 = W*in
   wire signed [14:0] m210_89;
   assign m210_89 =15'b0;

   // m210_90 = W*in
   wire signed [14:0] m210_90;
   assign m210_90 =15'b0;

   // m210_91 = W*in
   wire signed [14:0] m210_91;
   assign m210_91 =15'b0;

   // m210_92 = W*in
   wire signed [14:0] m210_92;
   assign m210_92 =15'b0;

   // m210_93 = W*in
   wire signed [14:0] m210_93;
   assign m210_93 =15'b0;

   // m210_94 = W*in
   wire signed [14:0] m210_94;
   assign m210_94 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_95 = W*in
   wire signed [14:0] m210_95;
   assign m210_95 =15'b0;

   // m210_96 = W*in
   wire signed [14:0] m210_96;
   assign m210_96 ={ {3{in210[14]}} , in210[14:3] };

   // m210_97 = W*in
   wire signed [14:0] m210_97;
   assign m210_97 ={ {3{neg210[14]}} , neg210[14:3] };

   // m210_98 = W*in
   wire signed [14:0] m210_98;
   assign m210_98 =15'b0;

   // m210_99 = W*in
   wire signed [14:0] m210_99;
   assign m210_99 =15'b0;

   // m210_100 = W*in
   wire signed [14:0] m210_100;
   assign m210_100 =15'b0;

   // m211_1 = W*in
   wire signed [14:0] m211_1;
   assign m211_1 =15'b0;

   // m211_2 = W*in
   wire signed [14:0] m211_2;
   assign m211_2 =15'b0;

   // m211_3 = W*in
   wire signed [14:0] m211_3;
   assign m211_3 =15'b0;

   // m211_4 = W*in
   wire signed [14:0] m211_4;
   assign m211_4 =15'b0;

   // m211_5 = W*in
   wire signed [14:0] m211_5;
   assign m211_5 =15'b0;

   // m211_6 = W*in
   wire signed [14:0] m211_6;
   assign m211_6 =15'b0;

   // m211_7 = W*in
   wire signed [14:0] m211_7;
   assign m211_7 =15'b0;

   // m211_8 = W*in
   wire signed [14:0] m211_8;
   assign m211_8 =15'b0;

   // m211_9 = W*in
   wire signed [14:0] m211_9;
   assign m211_9 =15'b0;

   // m211_10 = W*in
   wire signed [14:0] m211_10;
   assign m211_10 =15'b0;

   // m211_11 = W*in
   wire signed [14:0] m211_11;
   assign m211_11 =15'b0;

   // m211_12 = W*in
   wire signed [14:0] m211_12;
   assign m211_12 =15'b0;

   // m211_13 = W*in
   wire signed [14:0] m211_13;
   assign m211_13 =15'b0;

   // m211_14 = W*in
   wire signed [14:0] m211_14;
   assign m211_14 ={ {4{neg211[14]}} , neg211[14:4] };

   // m211_15 = W*in
   wire signed [14:0] m211_15;
   assign m211_15 =15'b0;

   // m211_16 = W*in
   wire signed [14:0] m211_16;
   assign m211_16 =15'b0;

   // m211_17 = W*in
   wire signed [14:0] m211_17;
   assign m211_17 =15'b0;

   // m211_18 = W*in
   wire signed [14:0] m211_18;
   assign m211_18 =15'b0;

   // m211_19 = W*in
   wire signed [14:0] m211_19;
   assign m211_19 =15'b0;

   // m211_20 = W*in
   wire signed [14:0] m211_20;
   assign m211_20 =15'b0;

   // m211_21 = W*in
   wire signed [14:0] m211_21;
   assign m211_21 =15'b0;

   // m211_22 = W*in
   wire signed [14:0] m211_22;
   assign m211_22 =15'b0;

   // m211_23 = W*in
   wire signed [14:0] m211_23;
   assign m211_23 =15'b0;

   // m211_24 = W*in
   wire signed [14:0] m211_24;
   assign m211_24 =15'b0;

   // m211_25 = W*in
   wire signed [14:0] m211_25;
   assign m211_25 =15'b0;

   // m211_26 = W*in
   wire signed [14:0] m211_26;
   assign m211_26 =15'b0;

   // m211_27 = W*in
   wire signed [14:0] m211_27;
   assign m211_27 =15'b0;

   // m211_28 = W*in
   wire signed [14:0] m211_28;
   assign m211_28 =15'b0;

   // m211_29 = W*in
   wire signed [14:0] m211_29;
   assign m211_29 =15'b0;

   // m211_30 = W*in
   wire signed [14:0] m211_30;
   assign m211_30 ={ {3{neg211[14]}} , neg211[14:3] };

   // m211_31 = W*in
   wire signed [14:0] m211_31;
   assign m211_31 =15'b0;

   // m211_32 = W*in
   wire signed [14:0] m211_32;
   assign m211_32 =15'b0;

   // m211_33 = W*in
   wire signed [14:0] m211_33;
   assign m211_33 =15'b0;

   // m211_34 = W*in
   wire signed [14:0] m211_34;
   assign m211_34 =15'b0;

   // m211_35 = W*in
   wire signed [14:0] m211_35;
   assign m211_35 =15'b0;

   // m211_36 = W*in
   wire signed [14:0] m211_36;
   assign m211_36 =15'b0;

   // m211_37 = W*in
   wire signed [14:0] m211_37;
   assign m211_37 =15'b0;

   // m211_38 = W*in
   wire signed [14:0] m211_38;
   assign m211_38 =15'b0;

   // m211_39 = W*in
   wire signed [14:0] m211_39;
   assign m211_39 =15'b0;

   // m211_40 = W*in
   wire signed [14:0] m211_40;
   assign m211_40 =15'b0;

   // m211_41 = W*in
   wire signed [14:0] m211_41;
   assign m211_41 =15'b0;

   // m211_42 = W*in
   wire signed [14:0] m211_42;
   assign m211_42 =15'b0;

   // m211_43 = W*in
   wire signed [14:0] m211_43;
   assign m211_43 =15'b0;

   // m211_44 = W*in
   wire signed [14:0] m211_44;
   assign m211_44 =15'b0;

   // m211_45 = W*in
   wire signed [14:0] m211_45;
   assign m211_45 =15'b0;

   // m211_46 = W*in
   wire signed [14:0] m211_46;
   assign m211_46 =15'b0;

   // m211_47 = W*in
   wire signed [14:0] m211_47;
   assign m211_47 =15'b0;

   // m211_48 = W*in
   wire signed [14:0] m211_48;
   assign m211_48 =15'b0;

   // m211_49 = W*in
   wire signed [14:0] m211_49;
   assign m211_49 =15'b0;

   // m211_50 = W*in
   wire signed [14:0] m211_50;
   assign m211_50 =15'b0;

   // m211_51 = W*in
   wire signed [14:0] m211_51;
   assign m211_51 =15'b0;

   // m211_52 = W*in
   wire signed [14:0] m211_52;
   assign m211_52 =15'b0;

   // m211_53 = W*in
   wire signed [14:0] m211_53;
   assign m211_53 =15'b0;

   // m211_54 = W*in
   wire signed [14:0] m211_54;
   assign m211_54 =15'b0;

   // m211_55 = W*in
   wire signed [14:0] m211_55;
   assign m211_55 =15'b0;

   // m211_56 = W*in
   wire signed [14:0] m211_56;
   assign m211_56 =15'b0;

   // m211_57 = W*in
   wire signed [14:0] m211_57;
   assign m211_57 =15'b0;

   // m211_58 = W*in
   wire signed [14:0] m211_58;
   assign m211_58 ={ {4{in211[14]}} , in211[14:4] };

   // m211_59 = W*in
   wire signed [14:0] m211_59;
   assign m211_59 =15'b0;

   // m211_60 = W*in
   wire signed [14:0] m211_60;
   assign m211_60 =15'b0;

   // m211_61 = W*in
   wire signed [14:0] m211_61;
   assign m211_61 =15'b0;

   // m211_62 = W*in
   wire signed [14:0] m211_62;
   assign m211_62 =15'b0;

   // m211_63 = W*in
   wire signed [14:0] m211_63;
   assign m211_63 ={ {4{in211[14]}} , in211[14:4] };

   // m211_64 = W*in
   wire signed [14:0] m211_64;
   assign m211_64 =15'b0;

   // m211_65 = W*in
   wire signed [14:0] m211_65;
   assign m211_65 =15'b0;

   // m211_66 = W*in
   wire signed [14:0] m211_66;
   assign m211_66 =15'b0;

   // m211_67 = W*in
   wire signed [14:0] m211_67;
   assign m211_67 ={ {3{neg211[14]}} , neg211[14:3] };

   // m211_68 = W*in
   wire signed [14:0] m211_68;
   assign m211_68 =15'b0;

   // m211_69 = W*in
   wire signed [14:0] m211_69;
   assign m211_69 =15'b0;

   // m211_70 = W*in
   wire signed [14:0] m211_70;
   assign m211_70 =15'b0;

   // m211_71 = W*in
   wire signed [14:0] m211_71;
   assign m211_71 =15'b0;

   // m211_72 = W*in
   wire signed [14:0] m211_72;
   assign m211_72 =15'b0;

   // m211_73 = W*in
   wire signed [14:0] m211_73;
   assign m211_73 =15'b0;

   // m211_74 = W*in
   wire signed [14:0] m211_74;
   assign m211_74 =15'b0;

   // m211_75 = W*in
   wire signed [14:0] m211_75;
   assign m211_75 =15'b0;

   // m211_76 = W*in
   wire signed [14:0] m211_76;
   assign m211_76 =15'b0;

   // m211_77 = W*in
   wire signed [14:0] m211_77;
   assign m211_77 =15'b0;

   // m211_78 = W*in
   wire signed [14:0] m211_78;
   assign m211_78 =15'b0;

   // m211_79 = W*in
   wire signed [14:0] m211_79;
   assign m211_79 =15'b0;

   // m211_80 = W*in
   wire signed [14:0] m211_80;
   assign m211_80 =15'b0;

   // m211_81 = W*in
   wire signed [14:0] m211_81;
   assign m211_81 =15'b0;

   // m211_82 = W*in
   wire signed [14:0] m211_82;
   assign m211_82 ={ {3{in211[14]}} , in211[14:3] };

   // m211_83 = W*in
   wire signed [14:0] m211_83;
   assign m211_83 =15'b0;

   // m211_84 = W*in
   wire signed [14:0] m211_84;
   assign m211_84 =15'b0;

   // m211_85 = W*in
   wire signed [14:0] m211_85;
   assign m211_85 =15'b0;

   // m211_86 = W*in
   wire signed [14:0] m211_86;
   assign m211_86 ={ {3{neg211[14]}} , neg211[14:3] };

   // m211_87 = W*in
   wire signed [14:0] m211_87;
   assign m211_87 =15'b0;

   // m211_88 = W*in
   wire signed [14:0] m211_88;
   assign m211_88 =15'b0;

   // m211_89 = W*in
   wire signed [14:0] m211_89;
   assign m211_89 =15'b0;

   // m211_90 = W*in
   wire signed [14:0] m211_90;
   assign m211_90 =15'b0;

   // m211_91 = W*in
   wire signed [14:0] m211_91;
   assign m211_91 =15'b0;

   // m211_92 = W*in
   wire signed [14:0] m211_92;
   assign m211_92 =15'b0;

   // m211_93 = W*in
   wire signed [14:0] m211_93;
   assign m211_93 ={ {3{in211[14]}} , in211[14:3] };

   // m211_94 = W*in
   wire signed [14:0] m211_94;
   assign m211_94 =15'b0;

   // m211_95 = W*in
   wire signed [14:0] m211_95;
   assign m211_95 ={ {3{neg211[14]}} , neg211[14:3] };

   // m211_96 = W*in
   wire signed [14:0] m211_96;
   assign m211_96 =15'b0;

   // m211_97 = W*in
   wire signed [14:0] m211_97;
   assign m211_97 =15'b0;

   // m211_98 = W*in
   wire signed [14:0] m211_98;
   assign m211_98 =15'b0;

   // m211_99 = W*in
   wire signed [14:0] m211_99;
   assign m211_99 =15'b0;

   // m211_100 = W*in
   wire signed [14:0] m211_100;
   assign m211_100 ={ {2{in211[14]}} , in211[14:2] };

   // m212_1 = W*in
   wire signed [14:0] m212_1;
   assign m212_1 =15'b0;

   // m212_2 = W*in
   wire signed [14:0] m212_2;
   assign m212_2 =15'b0;

   // m212_3 = W*in
   wire signed [14:0] m212_3;
   assign m212_3 =15'b0;

   // m212_4 = W*in
   wire signed [14:0] m212_4;
   assign m212_4 ={ {3{in212[14]}} , in212[14:3] };

   // m212_5 = W*in
   wire signed [14:0] m212_5;
   assign m212_5 =15'b0;

   // m212_6 = W*in
   wire signed [14:0] m212_6;
   assign m212_6 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_7 = W*in
   wire signed [14:0] m212_7;
   assign m212_7 =15'b0;

   // m212_8 = W*in
   wire signed [14:0] m212_8;
   assign m212_8 =15'b0;

   // m212_9 = W*in
   wire signed [14:0] m212_9;
   assign m212_9 =15'b0;

   // m212_10 = W*in
   wire signed [14:0] m212_10;
   assign m212_10 =15'b0;

   // m212_11 = W*in
   wire signed [14:0] m212_11;
   assign m212_11 =15'b0;

   // m212_12 = W*in
   wire signed [14:0] m212_12;
   assign m212_12 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_13 = W*in
   wire signed [14:0] m212_13;
   assign m212_13 =15'b0;

   // m212_14 = W*in
   wire signed [14:0] m212_14;
   assign m212_14 =15'b0;

   // m212_15 = W*in
   wire signed [14:0] m212_15;
   assign m212_15 =15'b0;

   // m212_16 = W*in
   wire signed [14:0] m212_16;
   assign m212_16 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_17 = W*in
   wire signed [14:0] m212_17;
   assign m212_17 =15'b0;

   // m212_18 = W*in
   wire signed [14:0] m212_18;
   assign m212_18 =15'b0;

   // m212_19 = W*in
   wire signed [14:0] m212_19;
   assign m212_19 ={ {4{neg212[14]}} , neg212[14:4] };

   // m212_20 = W*in
   wire signed [14:0] m212_20;
   assign m212_20 =15'b0;

   // m212_21 = W*in
   wire signed [14:0] m212_21;
   assign m212_21 ={ {3{in212[14]}} , in212[14:3] };

   // m212_22 = W*in
   wire signed [14:0] m212_22;
   assign m212_22 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_23 = W*in
   wire signed [14:0] m212_23;
   assign m212_23 =15'b0;

   // m212_24 = W*in
   wire signed [14:0] m212_24;
   assign m212_24 =15'b0;

   // m212_25 = W*in
   wire signed [14:0] m212_25;
   assign m212_25 =15'b0;

   // m212_26 = W*in
   wire signed [14:0] m212_26;
   assign m212_26 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_27 = W*in
   wire signed [14:0] m212_27;
   assign m212_27 =15'b0;

   // m212_28 = W*in
   wire signed [14:0] m212_28;
   assign m212_28 =15'b0;

   // m212_29 = W*in
   wire signed [14:0] m212_29;
   assign m212_29 =15'b0;

   // m212_30 = W*in
   wire signed [14:0] m212_30;
   assign m212_30 =15'b0;

   // m212_31 = W*in
   wire signed [14:0] m212_31;
   assign m212_31 =15'b0;

   // m212_32 = W*in
   wire signed [14:0] m212_32;
   assign m212_32 =15'b0;

   // m212_33 = W*in
   wire signed [14:0] m212_33;
   assign m212_33 =15'b0;

   // m212_34 = W*in
   wire signed [14:0] m212_34;
   assign m212_34 =15'b0;

   // m212_35 = W*in
   wire signed [14:0] m212_35;
   assign m212_35 =15'b0;

   // m212_36 = W*in
   wire signed [14:0] m212_36;
   assign m212_36 =15'b0;

   // m212_37 = W*in
   wire signed [14:0] m212_37;
   assign m212_37 =15'b0;

   // m212_38 = W*in
   wire signed [14:0] m212_38;
   assign m212_38 =15'b0;

   // m212_39 = W*in
   wire signed [14:0] m212_39;
   assign m212_39 =15'b0;

   // m212_40 = W*in
   wire signed [14:0] m212_40;
   assign m212_40 =15'b0;

   // m212_41 = W*in
   wire signed [14:0] m212_41;
   assign m212_41 =15'b0;

   // m212_42 = W*in
   wire signed [14:0] m212_42;
   assign m212_42 =15'b0;

   // m212_43 = W*in
   wire signed [14:0] m212_43;
   assign m212_43 =15'b0;

   // m212_44 = W*in
   wire signed [14:0] m212_44;
   assign m212_44 =15'b0;

   // m212_45 = W*in
   wire signed [14:0] m212_45;
   assign m212_45 =15'b0;

   // m212_46 = W*in
   wire signed [14:0] m212_46;
   assign m212_46 =15'b0;

   // m212_47 = W*in
   wire signed [14:0] m212_47;
   assign m212_47 =15'b0;

   // m212_48 = W*in
   wire signed [14:0] m212_48;
   assign m212_48 =15'b0;

   // m212_49 = W*in
   wire signed [14:0] m212_49;
   assign m212_49 ={ {4{in212[14]}} , in212[14:4] };

   // m212_50 = W*in
   wire signed [14:0] m212_50;
   assign m212_50 =15'b0;

   // m212_51 = W*in
   wire signed [14:0] m212_51;
   assign m212_51 =15'b0;

   // m212_52 = W*in
   wire signed [14:0] m212_52;
   assign m212_52 =15'b0;

   // m212_53 = W*in
   wire signed [14:0] m212_53;
   assign m212_53 =15'b0;

   // m212_54 = W*in
   wire signed [14:0] m212_54;
   assign m212_54 =15'b0;

   // m212_55 = W*in
   wire signed [14:0] m212_55;
   assign m212_55 =15'b0;

   // m212_56 = W*in
   wire signed [14:0] m212_56;
   assign m212_56 =15'b0;

   // m212_57 = W*in
   wire signed [14:0] m212_57;
   assign m212_57 =15'b0;

   // m212_58 = W*in
   wire signed [14:0] m212_58;
   assign m212_58 =15'b0;

   // m212_59 = W*in
   wire signed [14:0] m212_59;
   assign m212_59 =15'b0;

   // m212_60 = W*in
   wire signed [14:0] m212_60;
   assign m212_60 ={ {3{in212[14]}} , in212[14:3] };

   // m212_61 = W*in
   wire signed [14:0] m212_61;
   assign m212_61 =15'b0;

   // m212_62 = W*in
   wire signed [14:0] m212_62;
   assign m212_62 =15'b0;

   // m212_63 = W*in
   wire signed [14:0] m212_63;
   assign m212_63 =15'b0;

   // m212_64 = W*in
   wire signed [14:0] m212_64;
   assign m212_64 =15'b0;

   // m212_65 = W*in
   wire signed [14:0] m212_65;
   assign m212_65 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_66 = W*in
   wire signed [14:0] m212_66;
   assign m212_66 =15'b0;

   // m212_67 = W*in
   wire signed [14:0] m212_67;
   assign m212_67 =15'b0;

   // m212_68 = W*in
   wire signed [14:0] m212_68;
   assign m212_68 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_69 = W*in
   wire signed [14:0] m212_69;
   assign m212_69 =15'b0;

   // m212_70 = W*in
   wire signed [14:0] m212_70;
   assign m212_70 =15'b0;

   // m212_71 = W*in
   wire signed [14:0] m212_71;
   assign m212_71 =15'b0;

   // m212_72 = W*in
   wire signed [14:0] m212_72;
   assign m212_72 ={ {3{in212[14]}} , in212[14:3] };

   // m212_73 = W*in
   wire signed [14:0] m212_73;
   assign m212_73 =15'b0;

   // m212_74 = W*in
   wire signed [14:0] m212_74;
   assign m212_74 =15'b0;

   // m212_75 = W*in
   wire signed [14:0] m212_75;
   assign m212_75 =15'b0;

   // m212_76 = W*in
   wire signed [14:0] m212_76;
   assign m212_76 =15'b0;

   // m212_77 = W*in
   wire signed [14:0] m212_77;
   assign m212_77 ={ {3{in212[14]}} , in212[14:3] };

   // m212_78 = W*in
   wire signed [14:0] m212_78;
   assign m212_78 =15'b0;

   // m212_79 = W*in
   wire signed [14:0] m212_79;
   assign m212_79 =15'b0;

   // m212_80 = W*in
   wire signed [14:0] m212_80;
   assign m212_80 =15'b0;

   // m212_81 = W*in
   wire signed [14:0] m212_81;
   assign m212_81 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_82 = W*in
   wire signed [14:0] m212_82;
   assign m212_82 =15'b0;

   // m212_83 = W*in
   wire signed [14:0] m212_83;
   assign m212_83 =15'b0;

   // m212_84 = W*in
   wire signed [14:0] m212_84;
   assign m212_84 =15'b0;

   // m212_85 = W*in
   wire signed [14:0] m212_85;
   assign m212_85 =15'b0;

   // m212_86 = W*in
   wire signed [14:0] m212_86;
   assign m212_86 =15'b0;

   // m212_87 = W*in
   wire signed [14:0] m212_87;
   assign m212_87 =15'b0;

   // m212_88 = W*in
   wire signed [14:0] m212_88;
   assign m212_88 =15'b0;

   // m212_89 = W*in
   wire signed [14:0] m212_89;
   assign m212_89 =15'b0;

   // m212_90 = W*in
   wire signed [14:0] m212_90;
   assign m212_90 =15'b0;

   // m212_91 = W*in
   wire signed [14:0] m212_91;
   assign m212_91 =15'b0;

   // m212_92 = W*in
   wire signed [14:0] m212_92;
   assign m212_92 =15'b0;

   // m212_93 = W*in
   wire signed [14:0] m212_93;
   assign m212_93 =15'b0;

   // m212_94 = W*in
   wire signed [14:0] m212_94;
   assign m212_94 =15'b0;

   // m212_95 = W*in
   wire signed [14:0] m212_95;
   assign m212_95 ={ {3{neg212[14]}} , neg212[14:3] };

   // m212_96 = W*in
   wire signed [14:0] m212_96;
   assign m212_96 ={ {3{in212[14]}} , in212[14:3] };

   // m212_97 = W*in
   wire signed [14:0] m212_97;
   assign m212_97 ={ {4{in212[14]}} , in212[14:4] };

   // m212_98 = W*in
   wire signed [14:0] m212_98;
   assign m212_98 =15'b0;

   // m212_99 = W*in
   wire signed [14:0] m212_99;
   assign m212_99 =15'b0;

   // m212_100 = W*in
   wire signed [14:0] m212_100;
   assign m212_100 ={ {4{neg212[14]}} , neg212[14:4] };

   // m213_1 = W*in
   wire signed [14:0] m213_1;
   assign m213_1 =15'b0;

   // m213_2 = W*in
   wire signed [14:0] m213_2;
   assign m213_2 =15'b0;

   // m213_3 = W*in
   wire signed [14:0] m213_3;
   assign m213_3 =15'b0;

   // m213_4 = W*in
   wire signed [14:0] m213_4;
   assign m213_4 ={ {4{in213[14]}} , in213[14:4] };

   // m213_5 = W*in
   wire signed [14:0] m213_5;
   assign m213_5 =15'b0;

   // m213_6 = W*in
   wire signed [14:0] m213_6;
   assign m213_6 =15'b0;

   // m213_7 = W*in
   wire signed [14:0] m213_7;
   assign m213_7 =15'b0;

   // m213_8 = W*in
   wire signed [14:0] m213_8;
   assign m213_8 ={ {3{in213[14]}} , in213[14:3] };

   // m213_9 = W*in
   wire signed [14:0] m213_9;
   assign m213_9 =15'b0;

   // m213_10 = W*in
   wire signed [14:0] m213_10;
   assign m213_10 =15'b0;

   // m213_11 = W*in
   wire signed [14:0] m213_11;
   assign m213_11 =15'b0;

   // m213_12 = W*in
   wire signed [14:0] m213_12;
   assign m213_12 =15'b0;

   // m213_13 = W*in
   wire signed [14:0] m213_13;
   assign m213_13 =15'b0;

   // m213_14 = W*in
   wire signed [14:0] m213_14;
   assign m213_14 =15'b0;

   // m213_15 = W*in
   wire signed [14:0] m213_15;
   assign m213_15 =15'b0;

   // m213_16 = W*in
   wire signed [14:0] m213_16;
   assign m213_16 =15'b0;

   // m213_17 = W*in
   wire signed [14:0] m213_17;
   assign m213_17 =15'b0;

   // m213_18 = W*in
   wire signed [14:0] m213_18;
   assign m213_18 =15'b0;

   // m213_19 = W*in
   wire signed [14:0] m213_19;
   assign m213_19 =15'b0;

   // m213_20 = W*in
   wire signed [14:0] m213_20;
   assign m213_20 =15'b0;

   // m213_21 = W*in
   wire signed [14:0] m213_21;
   assign m213_21 =15'b0;

   // m213_22 = W*in
   wire signed [14:0] m213_22;
   assign m213_22 =15'b0;

   // m213_23 = W*in
   wire signed [14:0] m213_23;
   assign m213_23 =15'b0;

   // m213_24 = W*in
   wire signed [14:0] m213_24;
   assign m213_24 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_25 = W*in
   wire signed [14:0] m213_25;
   assign m213_25 =15'b0;

   // m213_26 = W*in
   wire signed [14:0] m213_26;
   assign m213_26 =15'b0;

   // m213_27 = W*in
   wire signed [14:0] m213_27;
   assign m213_27 =15'b0;

   // m213_28 = W*in
   wire signed [14:0] m213_28;
   assign m213_28 ={ {3{in213[14]}} , in213[14:3] };

   // m213_29 = W*in
   wire signed [14:0] m213_29;
   assign m213_29 =15'b0;

   // m213_30 = W*in
   wire signed [14:0] m213_30;
   assign m213_30 =15'b0;

   // m213_31 = W*in
   wire signed [14:0] m213_31;
   assign m213_31 ={ {3{in213[14]}} , in213[14:3] };

   // m213_32 = W*in
   wire signed [14:0] m213_32;
   assign m213_32 =15'b0;

   // m213_33 = W*in
   wire signed [14:0] m213_33;
   assign m213_33 =15'b0;

   // m213_34 = W*in
   wire signed [14:0] m213_34;
   assign m213_34 =15'b0;

   // m213_35 = W*in
   wire signed [14:0] m213_35;
   assign m213_35 =15'b0;

   // m213_36 = W*in
   wire signed [14:0] m213_36;
   assign m213_36 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_37 = W*in
   wire signed [14:0] m213_37;
   assign m213_37 =15'b0;

   // m213_38 = W*in
   wire signed [14:0] m213_38;
   assign m213_38 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_39 = W*in
   wire signed [14:0] m213_39;
   assign m213_39 =15'b0;

   // m213_40 = W*in
   wire signed [14:0] m213_40;
   assign m213_40 =15'b0;

   // m213_41 = W*in
   wire signed [14:0] m213_41;
   assign m213_41 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_42 = W*in
   wire signed [14:0] m213_42;
   assign m213_42 =15'b0;

   // m213_43 = W*in
   wire signed [14:0] m213_43;
   assign m213_43 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_44 = W*in
   wire signed [14:0] m213_44;
   assign m213_44 =15'b0;

   // m213_45 = W*in
   wire signed [14:0] m213_45;
   assign m213_45 =15'b0;

   // m213_46 = W*in
   wire signed [14:0] m213_46;
   assign m213_46 =15'b0;

   // m213_47 = W*in
   wire signed [14:0] m213_47;
   assign m213_47 =15'b0;

   // m213_48 = W*in
   wire signed [14:0] m213_48;
   assign m213_48 =15'b0;

   // m213_49 = W*in
   wire signed [14:0] m213_49;
   assign m213_49 =15'b0;

   // m213_50 = W*in
   wire signed [14:0] m213_50;
   assign m213_50 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_51 = W*in
   wire signed [14:0] m213_51;
   assign m213_51 =15'b0;

   // m213_52 = W*in
   wire signed [14:0] m213_52;
   assign m213_52 =15'b0;

   // m213_53 = W*in
   wire signed [14:0] m213_53;
   assign m213_53 ={ {3{in213[14]}} , in213[14:3] };

   // m213_54 = W*in
   wire signed [14:0] m213_54;
   assign m213_54 =15'b0;

   // m213_55 = W*in
   wire signed [14:0] m213_55;
   assign m213_55 =15'b0;

   // m213_56 = W*in
   wire signed [14:0] m213_56;
   assign m213_56 =15'b0;

   // m213_57 = W*in
   wire signed [14:0] m213_57;
   assign m213_57 =15'b0;

   // m213_58 = W*in
   wire signed [14:0] m213_58;
   assign m213_58 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_59 = W*in
   wire signed [14:0] m213_59;
   assign m213_59 =15'b0;

   // m213_60 = W*in
   wire signed [14:0] m213_60;
   assign m213_60 =15'b0;

   // m213_61 = W*in
   wire signed [14:0] m213_61;
   assign m213_61 =15'b0;

   // m213_62 = W*in
   wire signed [14:0] m213_62;
   assign m213_62 =15'b0;

   // m213_63 = W*in
   wire signed [14:0] m213_63;
   assign m213_63 =15'b0;

   // m213_64 = W*in
   wire signed [14:0] m213_64;
   assign m213_64 =15'b0;

   // m213_65 = W*in
   wire signed [14:0] m213_65;
   assign m213_65 =15'b0;

   // m213_66 = W*in
   wire signed [14:0] m213_66;
   assign m213_66 =15'b0;

   // m213_67 = W*in
   wire signed [14:0] m213_67;
   assign m213_67 =15'b0;

   // m213_68 = W*in
   wire signed [14:0] m213_68;
   assign m213_68 ={ {4{in213[14]}} , in213[14:4] };

   // m213_69 = W*in
   wire signed [14:0] m213_69;
   assign m213_69 ={ {4{in213[14]}} , in213[14:4] };

   // m213_70 = W*in
   wire signed [14:0] m213_70;
   assign m213_70 =15'b0;

   // m213_71 = W*in
   wire signed [14:0] m213_71;
   assign m213_71 =15'b0;

   // m213_72 = W*in
   wire signed [14:0] m213_72;
   assign m213_72 =15'b0;

   // m213_73 = W*in
   wire signed [14:0] m213_73;
   assign m213_73 ={ {3{in213[14]}} , in213[14:3] };

   // m213_74 = W*in
   wire signed [14:0] m213_74;
   assign m213_74 ={ {4{in213[14]}} , in213[14:4] };

   // m213_75 = W*in
   wire signed [14:0] m213_75;
   assign m213_75 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_76 = W*in
   wire signed [14:0] m213_76;
   assign m213_76 ={ {4{neg213[14]}} , neg213[14:4] };

   // m213_77 = W*in
   wire signed [14:0] m213_77;
   assign m213_77 =15'b0;

   // m213_78 = W*in
   wire signed [14:0] m213_78;
   assign m213_78 ={ {3{in213[14]}} , in213[14:3] };

   // m213_79 = W*in
   wire signed [14:0] m213_79;
   assign m213_79 =15'b0;

   // m213_80 = W*in
   wire signed [14:0] m213_80;
   assign m213_80 =15'b0;

   // m213_81 = W*in
   wire signed [14:0] m213_81;
   assign m213_81 =15'b0;

   // m213_82 = W*in
   wire signed [14:0] m213_82;
   assign m213_82 =15'b0;

   // m213_83 = W*in
   wire signed [14:0] m213_83;
   assign m213_83 =15'b0;

   // m213_84 = W*in
   wire signed [14:0] m213_84;
   assign m213_84 =15'b0;

   // m213_85 = W*in
   wire signed [14:0] m213_85;
   assign m213_85 =15'b0;

   // m213_86 = W*in
   wire signed [14:0] m213_86;
   assign m213_86 =15'b0;

   // m213_87 = W*in
   wire signed [14:0] m213_87;
   assign m213_87 =15'b0;

   // m213_88 = W*in
   wire signed [14:0] m213_88;
   assign m213_88 =15'b0;

   // m213_89 = W*in
   wire signed [14:0] m213_89;
   assign m213_89 =15'b0;

   // m213_90 = W*in
   wire signed [14:0] m213_90;
   assign m213_90 =15'b0;

   // m213_91 = W*in
   wire signed [14:0] m213_91;
   assign m213_91 =15'b0;

   // m213_92 = W*in
   wire signed [14:0] m213_92;
   assign m213_92 =15'b0;

   // m213_93 = W*in
   wire signed [14:0] m213_93;
   assign m213_93 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_94 = W*in
   wire signed [14:0] m213_94;
   assign m213_94 =15'b0;

   // m213_95 = W*in
   wire signed [14:0] m213_95;
   assign m213_95 =15'b0;

   // m213_96 = W*in
   wire signed [14:0] m213_96;
   assign m213_96 ={ {3{neg213[14]}} , neg213[14:3] };

   // m213_97 = W*in
   wire signed [14:0] m213_97;
   assign m213_97 =15'b0;

   // m213_98 = W*in
   wire signed [14:0] m213_98;
   assign m213_98 =15'b0;

   // m213_99 = W*in
   wire signed [14:0] m213_99;
   assign m213_99 =15'b0;

   // m213_100 = W*in
   wire signed [14:0] m213_100;
   assign m213_100 ={ {3{neg213[14]}} , neg213[14:3] };

   // m214_1 = W*in
   wire signed [14:0] m214_1;
   assign m214_1 =15'b0;

   // m214_2 = W*in
   wire signed [14:0] m214_2;
   assign m214_2 =15'b0;

   // m214_3 = W*in
   wire signed [14:0] m214_3;
   assign m214_3 =15'b0;

   // m214_4 = W*in
   wire signed [14:0] m214_4;
   assign m214_4 =15'b0;

   // m214_5 = W*in
   wire signed [14:0] m214_5;
   assign m214_5 =15'b0;

   // m214_6 = W*in
   wire signed [14:0] m214_6;
   assign m214_6 =15'b0;

   // m214_7 = W*in
   wire signed [14:0] m214_7;
   assign m214_7 =15'b0;

   // m214_8 = W*in
   wire signed [14:0] m214_8;
   assign m214_8 =15'b0;

   // m214_9 = W*in
   wire signed [14:0] m214_9;
   assign m214_9 =15'b0;

   // m214_10 = W*in
   wire signed [14:0] m214_10;
   assign m214_10 =15'b0;

   // m214_11 = W*in
   wire signed [14:0] m214_11;
   assign m214_11 =15'b0;

   // m214_12 = W*in
   wire signed [14:0] m214_12;
   assign m214_12 =15'b0;

   // m214_13 = W*in
   wire signed [14:0] m214_13;
   assign m214_13 =15'b0;

   // m214_14 = W*in
   wire signed [14:0] m214_14;
   assign m214_14 =15'b0;

   // m214_15 = W*in
   wire signed [14:0] m214_15;
   assign m214_15 =15'b0;

   // m214_16 = W*in
   wire signed [14:0] m214_16;
   assign m214_16 =15'b0;

   // m214_17 = W*in
   wire signed [14:0] m214_17;
   assign m214_17 =15'b0;

   // m214_18 = W*in
   wire signed [14:0] m214_18;
   assign m214_18 =15'b0;

   // m214_19 = W*in
   wire signed [14:0] m214_19;
   assign m214_19 =15'b0;

   // m214_20 = W*in
   wire signed [14:0] m214_20;
   assign m214_20 =15'b0;

   // m214_21 = W*in
   wire signed [14:0] m214_21;
   assign m214_21 =15'b0;

   // m214_22 = W*in
   wire signed [14:0] m214_22;
   assign m214_22 =15'b0;

   // m214_23 = W*in
   wire signed [14:0] m214_23;
   assign m214_23 =15'b0;

   // m214_24 = W*in
   wire signed [14:0] m214_24;
   assign m214_24 =15'b0;

   // m214_25 = W*in
   wire signed [14:0] m214_25;
   assign m214_25 ={ {4{neg214[14]}} , neg214[14:4] };

   // m214_26 = W*in
   wire signed [14:0] m214_26;
   assign m214_26 =15'b0;

   // m214_27 = W*in
   wire signed [14:0] m214_27;
   assign m214_27 ={ {4{in214[14]}} , in214[14:4] };

   // m214_28 = W*in
   wire signed [14:0] m214_28;
   assign m214_28 =15'b0;

   // m214_29 = W*in
   wire signed [14:0] m214_29;
   assign m214_29 =15'b0;

   // m214_30 = W*in
   wire signed [14:0] m214_30;
   assign m214_30 =15'b0;

   // m214_31 = W*in
   wire signed [14:0] m214_31;
   assign m214_31 =15'b0;

   // m214_32 = W*in
   wire signed [14:0] m214_32;
   assign m214_32 =15'b0;

   // m214_33 = W*in
   wire signed [14:0] m214_33;
   assign m214_33 ={ {3{in214[14]}} , in214[14:3] };

   // m214_34 = W*in
   wire signed [14:0] m214_34;
   assign m214_34 =15'b0;

   // m214_35 = W*in
   wire signed [14:0] m214_35;
   assign m214_35 =15'b0;

   // m214_36 = W*in
   wire signed [14:0] m214_36;
   assign m214_36 =15'b0;

   // m214_37 = W*in
   wire signed [14:0] m214_37;
   assign m214_37 =15'b0;

   // m214_38 = W*in
   wire signed [14:0] m214_38;
   assign m214_38 ={ {3{in214[14]}} , in214[14:3] };

   // m214_39 = W*in
   wire signed [14:0] m214_39;
   assign m214_39 =15'b0;

   // m214_40 = W*in
   wire signed [14:0] m214_40;
   assign m214_40 =15'b0;

   // m214_41 = W*in
   wire signed [14:0] m214_41;
   assign m214_41 =15'b0;

   // m214_42 = W*in
   wire signed [14:0] m214_42;
   assign m214_42 =15'b0;

   // m214_43 = W*in
   wire signed [14:0] m214_43;
   assign m214_43 ={ {3{neg214[14]}} , neg214[14:3] };

   // m214_44 = W*in
   wire signed [14:0] m214_44;
   assign m214_44 =15'b0;

   // m214_45 = W*in
   wire signed [14:0] m214_45;
   assign m214_45 =15'b0;

   // m214_46 = W*in
   wire signed [14:0] m214_46;
   assign m214_46 =15'b0;

   // m214_47 = W*in
   wire signed [14:0] m214_47;
   assign m214_47 =15'b0;

   // m214_48 = W*in
   wire signed [14:0] m214_48;
   assign m214_48 =15'b0;

   // m214_49 = W*in
   wire signed [14:0] m214_49;
   assign m214_49 =15'b0;

   // m214_50 = W*in
   wire signed [14:0] m214_50;
   assign m214_50 =15'b0;

   // m214_51 = W*in
   wire signed [14:0] m214_51;
   assign m214_51 =15'b0;

   // m214_52 = W*in
   wire signed [14:0] m214_52;
   assign m214_52 ={ {3{neg214[14]}} , neg214[14:3] };

   // m214_53 = W*in
   wire signed [14:0] m214_53;
   assign m214_53 =15'b0;

   // m214_54 = W*in
   wire signed [14:0] m214_54;
   assign m214_54 =15'b0;

   // m214_55 = W*in
   wire signed [14:0] m214_55;
   assign m214_55 =15'b0;

   // m214_56 = W*in
   wire signed [14:0] m214_56;
   assign m214_56 ={ {3{in214[14]}} , in214[14:3] };

   // m214_57 = W*in
   wire signed [14:0] m214_57;
   assign m214_57 =15'b0;

   // m214_58 = W*in
   wire signed [14:0] m214_58;
   assign m214_58 =15'b0;

   // m214_59 = W*in
   wire signed [14:0] m214_59;
   assign m214_59 =15'b0;

   // m214_60 = W*in
   wire signed [14:0] m214_60;
   assign m214_60 =15'b0;

   // m214_61 = W*in
   wire signed [14:0] m214_61;
   assign m214_61 =15'b0;

   // m214_62 = W*in
   wire signed [14:0] m214_62;
   assign m214_62 =15'b0;

   // m214_63 = W*in
   wire signed [14:0] m214_63;
   assign m214_63 =15'b0;

   // m214_64 = W*in
   wire signed [14:0] m214_64;
   assign m214_64 =15'b0;

   // m214_65 = W*in
   wire signed [14:0] m214_65;
   assign m214_65 ={ {4{neg214[14]}} , neg214[14:4] };

   // m214_66 = W*in
   wire signed [14:0] m214_66;
   assign m214_66 =15'b0;

   // m214_67 = W*in
   wire signed [14:0] m214_67;
   assign m214_67 =15'b0;

   // m214_68 = W*in
   wire signed [14:0] m214_68;
   assign m214_68 =15'b0;

   // m214_69 = W*in
   wire signed [14:0] m214_69;
   assign m214_69 =15'b0;

   // m214_70 = W*in
   wire signed [14:0] m214_70;
   assign m214_70 =15'b0;

   // m214_71 = W*in
   wire signed [14:0] m214_71;
   assign m214_71 =15'b0;

   // m214_72 = W*in
   wire signed [14:0] m214_72;
   assign m214_72 ={ {3{neg214[14]}} , neg214[14:3] };

   // m214_73 = W*in
   wire signed [14:0] m214_73;
   assign m214_73 =15'b0;

   // m214_74 = W*in
   wire signed [14:0] m214_74;
   assign m214_74 =15'b0;

   // m214_75 = W*in
   wire signed [14:0] m214_75;
   assign m214_75 =15'b0;

   // m214_76 = W*in
   wire signed [14:0] m214_76;
   assign m214_76 =15'b0;

   // m214_77 = W*in
   wire signed [14:0] m214_77;
   assign m214_77 =15'b0;

   // m214_78 = W*in
   wire signed [14:0] m214_78;
   assign m214_78 ={ {3{in214[14]}} , in214[14:3] };

   // m214_79 = W*in
   wire signed [14:0] m214_79;
   assign m214_79 =15'b0;

   // m214_80 = W*in
   wire signed [14:0] m214_80;
   assign m214_80 ={ {3{neg214[14]}} , neg214[14:3] };

   // m214_81 = W*in
   wire signed [14:0] m214_81;
   assign m214_81 =15'b0;

   // m214_82 = W*in
   wire signed [14:0] m214_82;
   assign m214_82 =15'b0;

   // m214_83 = W*in
   wire signed [14:0] m214_83;
   assign m214_83 =15'b0;

   // m214_84 = W*in
   wire signed [14:0] m214_84;
   assign m214_84 =15'b0;

   // m214_85 = W*in
   wire signed [14:0] m214_85;
   assign m214_85 =15'b0;

   // m214_86 = W*in
   wire signed [14:0] m214_86;
   assign m214_86 =15'b0;

   // m214_87 = W*in
   wire signed [14:0] m214_87;
   assign m214_87 =15'b0;

   // m214_88 = W*in
   wire signed [14:0] m214_88;
   assign m214_88 =15'b0;

   // m214_89 = W*in
   wire signed [14:0] m214_89;
   assign m214_89 =15'b0;

   // m214_90 = W*in
   wire signed [14:0] m214_90;
   assign m214_90 =15'b0;

   // m214_91 = W*in
   wire signed [14:0] m214_91;
   assign m214_91 =15'b0;

   // m214_92 = W*in
   wire signed [14:0] m214_92;
   assign m214_92 =15'b0;

   // m214_93 = W*in
   wire signed [14:0] m214_93;
   assign m214_93 =15'b0;

   // m214_94 = W*in
   wire signed [14:0] m214_94;
   assign m214_94 =15'b0;

   // m214_95 = W*in
   wire signed [14:0] m214_95;
   assign m214_95 =15'b0;

   // m214_96 = W*in
   wire signed [14:0] m214_96;
   assign m214_96 =15'b0;

   // m214_97 = W*in
   wire signed [14:0] m214_97;
   assign m214_97 =15'b0;

   // m214_98 = W*in
   wire signed [14:0] m214_98;
   assign m214_98 =15'b0;

   // m214_99 = W*in
   wire signed [14:0] m214_99;
   assign m214_99 =15'b0;

   // m214_100 = W*in
   wire signed [14:0] m214_100;
   assign m214_100 =15'b0;

   // m215_1 = W*in
   wire signed [14:0] m215_1;
   assign m215_1 =15'b0;

   // m215_2 = W*in
   wire signed [14:0] m215_2;
   assign m215_2 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_3 = W*in
   wire signed [14:0] m215_3;
   assign m215_3 =15'b0;

   // m215_4 = W*in
   wire signed [14:0] m215_4;
   assign m215_4 =15'b0;

   // m215_5 = W*in
   wire signed [14:0] m215_5;
   assign m215_5 ={ {4{neg215[14]}} , neg215[14:4] };

   // m215_6 = W*in
   wire signed [14:0] m215_6;
   assign m215_6 =15'b0;

   // m215_7 = W*in
   wire signed [14:0] m215_7;
   assign m215_7 =15'b0;

   // m215_8 = W*in
   wire signed [14:0] m215_8;
   assign m215_8 ={ {3{in215[14]}} , in215[14:3] };

   // m215_9 = W*in
   wire signed [14:0] m215_9;
   assign m215_9 =15'b0;

   // m215_10 = W*in
   wire signed [14:0] m215_10;
   assign m215_10 =15'b0;

   // m215_11 = W*in
   wire signed [14:0] m215_11;
   assign m215_11 =15'b0;

   // m215_12 = W*in
   wire signed [14:0] m215_12;
   assign m215_12 =15'b0;

   // m215_13 = W*in
   wire signed [14:0] m215_13;
   assign m215_13 =15'b0;

   // m215_14 = W*in
   wire signed [14:0] m215_14;
   assign m215_14 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_15 = W*in
   wire signed [14:0] m215_15;
   assign m215_15 =15'b0;

   // m215_16 = W*in
   wire signed [14:0] m215_16;
   assign m215_16 =15'b0;

   // m215_17 = W*in
   wire signed [14:0] m215_17;
   assign m215_17 =15'b0;

   // m215_18 = W*in
   wire signed [14:0] m215_18;
   assign m215_18 =15'b0;

   // m215_19 = W*in
   wire signed [14:0] m215_19;
   assign m215_19 ={ {4{neg215[14]}} , neg215[14:4] };

   // m215_20 = W*in
   wire signed [14:0] m215_20;
   assign m215_20 =15'b0;

   // m215_21 = W*in
   wire signed [14:0] m215_21;
   assign m215_21 =15'b0;

   // m215_22 = W*in
   wire signed [14:0] m215_22;
   assign m215_22 =15'b0;

   // m215_23 = W*in
   wire signed [14:0] m215_23;
   assign m215_23 =15'b0;

   // m215_24 = W*in
   wire signed [14:0] m215_24;
   assign m215_24 =15'b0;

   // m215_25 = W*in
   wire signed [14:0] m215_25;
   assign m215_25 ={ {3{in215[14]}} , in215[14:3] };

   // m215_26 = W*in
   wire signed [14:0] m215_26;
   assign m215_26 =15'b0;

   // m215_27 = W*in
   wire signed [14:0] m215_27;
   assign m215_27 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_28 = W*in
   wire signed [14:0] m215_28;
   assign m215_28 ={ {4{neg215[14]}} , neg215[14:4] };

   // m215_29 = W*in
   wire signed [14:0] m215_29;
   assign m215_29 =15'b0;

   // m215_30 = W*in
   wire signed [14:0] m215_30;
   assign m215_30 =15'b0;

   // m215_31 = W*in
   wire signed [14:0] m215_31;
   assign m215_31 ={ {4{in215[14]}} , in215[14:4] };

   // m215_32 = W*in
   wire signed [14:0] m215_32;
   assign m215_32 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_33 = W*in
   wire signed [14:0] m215_33;
   assign m215_33 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_34 = W*in
   wire signed [14:0] m215_34;
   assign m215_34 =15'b0;

   // m215_35 = W*in
   wire signed [14:0] m215_35;
   assign m215_35 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_36 = W*in
   wire signed [14:0] m215_36;
   assign m215_36 =15'b0;

   // m215_37 = W*in
   wire signed [14:0] m215_37;
   assign m215_37 =15'b0;

   // m215_38 = W*in
   wire signed [14:0] m215_38;
   assign m215_38 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_39 = W*in
   wire signed [14:0] m215_39;
   assign m215_39 =15'b0;

   // m215_40 = W*in
   wire signed [14:0] m215_40;
   assign m215_40 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_41 = W*in
   wire signed [14:0] m215_41;
   assign m215_41 =15'b0;

   // m215_42 = W*in
   wire signed [14:0] m215_42;
   assign m215_42 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_43 = W*in
   wire signed [14:0] m215_43;
   assign m215_43 =15'b0;

   // m215_44 = W*in
   wire signed [14:0] m215_44;
   assign m215_44 =15'b0;

   // m215_45 = W*in
   wire signed [14:0] m215_45;
   assign m215_45 =15'b0;

   // m215_46 = W*in
   wire signed [14:0] m215_46;
   assign m215_46 =15'b0;

   // m215_47 = W*in
   wire signed [14:0] m215_47;
   assign m215_47 =15'b0;

   // m215_48 = W*in
   wire signed [14:0] m215_48;
   assign m215_48 =15'b0;

   // m215_49 = W*in
   wire signed [14:0] m215_49;
   assign m215_49 ={ {3{in215[14]}} , in215[14:3] };

   // m215_50 = W*in
   wire signed [14:0] m215_50;
   assign m215_50 =15'b0;

   // m215_51 = W*in
   wire signed [14:0] m215_51;
   assign m215_51 =15'b0;

   // m215_52 = W*in
   wire signed [14:0] m215_52;
   assign m215_52 =15'b0;

   // m215_53 = W*in
   wire signed [14:0] m215_53;
   assign m215_53 =15'b0;

   // m215_54 = W*in
   wire signed [14:0] m215_54;
   assign m215_54 =15'b0;

   // m215_55 = W*in
   wire signed [14:0] m215_55;
   assign m215_55 =15'b0;

   // m215_56 = W*in
   wire signed [14:0] m215_56;
   assign m215_56 =15'b0;

   // m215_57 = W*in
   wire signed [14:0] m215_57;
   assign m215_57 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_58 = W*in
   wire signed [14:0] m215_58;
   assign m215_58 =15'b0;

   // m215_59 = W*in
   wire signed [14:0] m215_59;
   assign m215_59 =15'b0;

   // m215_60 = W*in
   wire signed [14:0] m215_60;
   assign m215_60 ={ {4{in215[14]}} , in215[14:4] };

   // m215_61 = W*in
   wire signed [14:0] m215_61;
   assign m215_61 =15'b0;

   // m215_62 = W*in
   wire signed [14:0] m215_62;
   assign m215_62 =15'b0;

   // m215_63 = W*in
   wire signed [14:0] m215_63;
   assign m215_63 =15'b0;

   // m215_64 = W*in
   wire signed [14:0] m215_64;
   assign m215_64 =15'b0;

   // m215_65 = W*in
   wire signed [14:0] m215_65;
   assign m215_65 ={ {3{in215[14]}} , in215[14:3] };

   // m215_66 = W*in
   wire signed [14:0] m215_66;
   assign m215_66 =15'b0;

   // m215_67 = W*in
   wire signed [14:0] m215_67;
   assign m215_67 =15'b0;

   // m215_68 = W*in
   wire signed [14:0] m215_68;
   assign m215_68 ={ {3{in215[14]}} , in215[14:3] };

   // m215_69 = W*in
   wire signed [14:0] m215_69;
   assign m215_69 ={ {3{in215[14]}} , in215[14:3] };

   // m215_70 = W*in
   wire signed [14:0] m215_70;
   assign m215_70 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_71 = W*in
   wire signed [14:0] m215_71;
   assign m215_71 =15'b0;

   // m215_72 = W*in
   wire signed [14:0] m215_72;
   assign m215_72 ={ {3{in215[14]}} , in215[14:3] };

   // m215_73 = W*in
   wire signed [14:0] m215_73;
   assign m215_73 ={ {3{in215[14]}} , in215[14:3] };

   // m215_74 = W*in
   wire signed [14:0] m215_74;
   assign m215_74 =15'b0;

   // m215_75 = W*in
   wire signed [14:0] m215_75;
   assign m215_75 =15'b0;

   // m215_76 = W*in
   wire signed [14:0] m215_76;
   assign m215_76 =15'b0;

   // m215_77 = W*in
   wire signed [14:0] m215_77;
   assign m215_77 ={ {3{in215[14]}} , in215[14:3] };

   // m215_78 = W*in
   wire signed [14:0] m215_78;
   assign m215_78 =15'b0;

   // m215_79 = W*in
   wire signed [14:0] m215_79;
   assign m215_79 =15'b0;

   // m215_80 = W*in
   wire signed [14:0] m215_80;
   assign m215_80 =15'b0;

   // m215_81 = W*in
   wire signed [14:0] m215_81;
   assign m215_81 =15'b0;

   // m215_82 = W*in
   wire signed [14:0] m215_82;
   assign m215_82 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_83 = W*in
   wire signed [14:0] m215_83;
   assign m215_83 =15'b0;

   // m215_84 = W*in
   wire signed [14:0] m215_84;
   assign m215_84 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_85 = W*in
   wire signed [14:0] m215_85;
   assign m215_85 =15'b0;

   // m215_86 = W*in
   wire signed [14:0] m215_86;
   assign m215_86 =15'b0;

   // m215_87 = W*in
   wire signed [14:0] m215_87;
   assign m215_87 =15'b0;

   // m215_88 = W*in
   wire signed [14:0] m215_88;
   assign m215_88 =15'b0;

   // m215_89 = W*in
   wire signed [14:0] m215_89;
   assign m215_89 =15'b0;

   // m215_90 = W*in
   wire signed [14:0] m215_90;
   assign m215_90 =15'b0;

   // m215_91 = W*in
   wire signed [14:0] m215_91;
   assign m215_91 =15'b0;

   // m215_92 = W*in
   wire signed [14:0] m215_92;
   assign m215_92 =15'b0;

   // m215_93 = W*in
   wire signed [14:0] m215_93;
   assign m215_93 =15'b0;

   // m215_94 = W*in
   wire signed [14:0] m215_94;
   assign m215_94 ={ {3{neg215[14]}} , neg215[14:3] };

   // m215_95 = W*in
   wire signed [14:0] m215_95;
   assign m215_95 =15'b0;

   // m215_96 = W*in
   wire signed [14:0] m215_96;
   assign m215_96 =15'b0;

   // m215_97 = W*in
   wire signed [14:0] m215_97;
   assign m215_97 =15'b0;

   // m215_98 = W*in
   wire signed [14:0] m215_98;
   assign m215_98 =15'b0;

   // m215_99 = W*in
   wire signed [14:0] m215_99;
   assign m215_99 =15'b0;

   // m215_100 = W*in
   wire signed [14:0] m215_100;
   assign m215_100 =15'b0;

   // m216_1 = W*in
   wire signed [14:0] m216_1;
   assign m216_1 =15'b0;

   // m216_2 = W*in
   wire signed [14:0] m216_2;
   assign m216_2 =15'b0;

   // m216_3 = W*in
   wire signed [14:0] m216_3;
   assign m216_3 =15'b0;

   // m216_4 = W*in
   wire signed [14:0] m216_4;
   assign m216_4 =15'b0;

   // m216_5 = W*in
   wire signed [14:0] m216_5;
   assign m216_5 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_6 = W*in
   wire signed [14:0] m216_6;
   assign m216_6 =15'b0;

   // m216_7 = W*in
   wire signed [14:0] m216_7;
   assign m216_7 =15'b0;

   // m216_8 = W*in
   wire signed [14:0] m216_8;
   assign m216_8 =15'b0;

   // m216_9 = W*in
   wire signed [14:0] m216_9;
   assign m216_9 =15'b0;

   // m216_10 = W*in
   wire signed [14:0] m216_10;
   assign m216_10 =15'b0;

   // m216_11 = W*in
   wire signed [14:0] m216_11;
   assign m216_11 =15'b0;

   // m216_12 = W*in
   wire signed [14:0] m216_12;
   assign m216_12 =15'b0;

   // m216_13 = W*in
   wire signed [14:0] m216_13;
   assign m216_13 =15'b0;

   // m216_14 = W*in
   wire signed [14:0] m216_14;
   assign m216_14 =15'b0;

   // m216_15 = W*in
   wire signed [14:0] m216_15;
   assign m216_15 =15'b0;

   // m216_16 = W*in
   wire signed [14:0] m216_16;
   assign m216_16 =15'b0;

   // m216_17 = W*in
   wire signed [14:0] m216_17;
   assign m216_17 ={ {3{in216[14]}} , in216[14:3] };

   // m216_18 = W*in
   wire signed [14:0] m216_18;
   assign m216_18 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_19 = W*in
   wire signed [14:0] m216_19;
   assign m216_19 =15'b0;

   // m216_20 = W*in
   wire signed [14:0] m216_20;
   assign m216_20 =15'b0;

   // m216_21 = W*in
   wire signed [14:0] m216_21;
   assign m216_21 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_22 = W*in
   wire signed [14:0] m216_22;
   assign m216_22 =15'b0;

   // m216_23 = W*in
   wire signed [14:0] m216_23;
   assign m216_23 =15'b0;

   // m216_24 = W*in
   wire signed [14:0] m216_24;
   assign m216_24 =15'b0;

   // m216_25 = W*in
   wire signed [14:0] m216_25;
   assign m216_25 =15'b0;

   // m216_26 = W*in
   wire signed [14:0] m216_26;
   assign m216_26 =15'b0;

   // m216_27 = W*in
   wire signed [14:0] m216_27;
   assign m216_27 =15'b0;

   // m216_28 = W*in
   wire signed [14:0] m216_28;
   assign m216_28 =15'b0;

   // m216_29 = W*in
   wire signed [14:0] m216_29;
   assign m216_29 =15'b0;

   // m216_30 = W*in
   wire signed [14:0] m216_30;
   assign m216_30 =15'b0;

   // m216_31 = W*in
   wire signed [14:0] m216_31;
   assign m216_31 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_32 = W*in
   wire signed [14:0] m216_32;
   assign m216_32 =15'b0;

   // m216_33 = W*in
   wire signed [14:0] m216_33;
   assign m216_33 =15'b0;

   // m216_34 = W*in
   wire signed [14:0] m216_34;
   assign m216_34 =15'b0;

   // m216_35 = W*in
   wire signed [14:0] m216_35;
   assign m216_35 =15'b0;

   // m216_36 = W*in
   wire signed [14:0] m216_36;
   assign m216_36 =15'b0;

   // m216_37 = W*in
   wire signed [14:0] m216_37;
   assign m216_37 =15'b0;

   // m216_38 = W*in
   wire signed [14:0] m216_38;
   assign m216_38 =15'b0;

   // m216_39 = W*in
   wire signed [14:0] m216_39;
   assign m216_39 ={ {3{in216[14]}} , in216[14:3] };

   // m216_40 = W*in
   wire signed [14:0] m216_40;
   assign m216_40 =15'b0;

   // m216_41 = W*in
   wire signed [14:0] m216_41;
   assign m216_41 =15'b0;

   // m216_42 = W*in
   wire signed [14:0] m216_42;
   assign m216_42 =15'b0;

   // m216_43 = W*in
   wire signed [14:0] m216_43;
   assign m216_43 =15'b0;

   // m216_44 = W*in
   wire signed [14:0] m216_44;
   assign m216_44 =15'b0;

   // m216_45 = W*in
   wire signed [14:0] m216_45;
   assign m216_45 =15'b0;

   // m216_46 = W*in
   wire signed [14:0] m216_46;
   assign m216_46 =15'b0;

   // m216_47 = W*in
   wire signed [14:0] m216_47;
   assign m216_47 =15'b0;

   // m216_48 = W*in
   wire signed [14:0] m216_48;
   assign m216_48 =15'b0;

   // m216_49 = W*in
   wire signed [14:0] m216_49;
   assign m216_49 =15'b0;

   // m216_50 = W*in
   wire signed [14:0] m216_50;
   assign m216_50 =15'b0;

   // m216_51 = W*in
   wire signed [14:0] m216_51;
   assign m216_51 =15'b0;

   // m216_52 = W*in
   wire signed [14:0] m216_52;
   assign m216_52 =15'b0;

   // m216_53 = W*in
   wire signed [14:0] m216_53;
   assign m216_53 =15'b0;

   // m216_54 = W*in
   wire signed [14:0] m216_54;
   assign m216_54 =15'b0;

   // m216_55 = W*in
   wire signed [14:0] m216_55;
   assign m216_55 =15'b0;

   // m216_56 = W*in
   wire signed [14:0] m216_56;
   assign m216_56 =15'b0;

   // m216_57 = W*in
   wire signed [14:0] m216_57;
   assign m216_57 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_58 = W*in
   wire signed [14:0] m216_58;
   assign m216_58 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_59 = W*in
   wire signed [14:0] m216_59;
   assign m216_59 =15'b0;

   // m216_60 = W*in
   wire signed [14:0] m216_60;
   assign m216_60 =15'b0;

   // m216_61 = W*in
   wire signed [14:0] m216_61;
   assign m216_61 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_62 = W*in
   wire signed [14:0] m216_62;
   assign m216_62 =15'b0;

   // m216_63 = W*in
   wire signed [14:0] m216_63;
   assign m216_63 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_64 = W*in
   wire signed [14:0] m216_64;
   assign m216_64 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_65 = W*in
   wire signed [14:0] m216_65;
   assign m216_65 =15'b0;

   // m216_66 = W*in
   wire signed [14:0] m216_66;
   assign m216_66 =15'b0;

   // m216_67 = W*in
   wire signed [14:0] m216_67;
   assign m216_67 =15'b0;

   // m216_68 = W*in
   wire signed [14:0] m216_68;
   assign m216_68 ={ {4{neg216[14]}} , neg216[14:4] };

   // m216_69 = W*in
   wire signed [14:0] m216_69;
   assign m216_69 =15'b0;

   // m216_70 = W*in
   wire signed [14:0] m216_70;
   assign m216_70 ={ {4{in216[14]}} , in216[14:4] };

   // m216_71 = W*in
   wire signed [14:0] m216_71;
   assign m216_71 =15'b0;

   // m216_72 = W*in
   wire signed [14:0] m216_72;
   assign m216_72 =15'b0;

   // m216_73 = W*in
   wire signed [14:0] m216_73;
   assign m216_73 =15'b0;

   // m216_74 = W*in
   wire signed [14:0] m216_74;
   assign m216_74 =15'b0;

   // m216_75 = W*in
   wire signed [14:0] m216_75;
   assign m216_75 =15'b0;

   // m216_76 = W*in
   wire signed [14:0] m216_76;
   assign m216_76 =15'b0;

   // m216_77 = W*in
   wire signed [14:0] m216_77;
   assign m216_77 =15'b0;

   // m216_78 = W*in
   wire signed [14:0] m216_78;
   assign m216_78 =15'b0;

   // m216_79 = W*in
   wire signed [14:0] m216_79;
   assign m216_79 =15'b0;

   // m216_80 = W*in
   wire signed [14:0] m216_80;
   assign m216_80 =15'b0;

   // m216_81 = W*in
   wire signed [14:0] m216_81;
   assign m216_81 =15'b0;

   // m216_82 = W*in
   wire signed [14:0] m216_82;
   assign m216_82 =15'b0;

   // m216_83 = W*in
   wire signed [14:0] m216_83;
   assign m216_83 =15'b0;

   // m216_84 = W*in
   wire signed [14:0] m216_84;
   assign m216_84 =15'b0;

   // m216_85 = W*in
   wire signed [14:0] m216_85;
   assign m216_85 =15'b0;

   // m216_86 = W*in
   wire signed [14:0] m216_86;
   assign m216_86 =15'b0;

   // m216_87 = W*in
   wire signed [14:0] m216_87;
   assign m216_87 =15'b0;

   // m216_88 = W*in
   wire signed [14:0] m216_88;
   assign m216_88 =15'b0;

   // m216_89 = W*in
   wire signed [14:0] m216_89;
   assign m216_89 =15'b0;

   // m216_90 = W*in
   wire signed [14:0] m216_90;
   assign m216_90 =15'b0;

   // m216_91 = W*in
   wire signed [14:0] m216_91;
   assign m216_91 =15'b0;

   // m216_92 = W*in
   wire signed [14:0] m216_92;
   assign m216_92 =15'b0;

   // m216_93 = W*in
   wire signed [14:0] m216_93;
   assign m216_93 =15'b0;

   // m216_94 = W*in
   wire signed [14:0] m216_94;
   assign m216_94 ={ {3{in216[14]}} , in216[14:3] };

   // m216_95 = W*in
   wire signed [14:0] m216_95;
   assign m216_95 =15'b0;

   // m216_96 = W*in
   wire signed [14:0] m216_96;
   assign m216_96 =15'b0;

   // m216_97 = W*in
   wire signed [14:0] m216_97;
   assign m216_97 =15'b0;

   // m216_98 = W*in
   wire signed [14:0] m216_98;
   assign m216_98 =15'b0;

   // m216_99 = W*in
   wire signed [14:0] m216_99;
   assign m216_99 =15'b0;

   // m216_100 = W*in
   wire signed [14:0] m216_100;
   assign m216_100 =15'b0;

   // m217_1 = W*in
   wire signed [14:0] m217_1;
   assign m217_1 =15'b0;

   // m217_2 = W*in
   wire signed [14:0] m217_2;
   assign m217_2 =15'b0;

   // m217_3 = W*in
   wire signed [14:0] m217_3;
   assign m217_3 =15'b0;

   // m217_4 = W*in
   wire signed [14:0] m217_4;
   assign m217_4 =15'b0;

   // m217_5 = W*in
   wire signed [14:0] m217_5;
   assign m217_5 =15'b0;

   // m217_6 = W*in
   wire signed [14:0] m217_6;
   assign m217_6 =15'b0;

   // m217_7 = W*in
   wire signed [14:0] m217_7;
   assign m217_7 =15'b0;

   // m217_8 = W*in
   wire signed [14:0] m217_8;
   assign m217_8 =15'b0;

   // m217_9 = W*in
   wire signed [14:0] m217_9;
   assign m217_9 =15'b0;

   // m217_10 = W*in
   wire signed [14:0] m217_10;
   assign m217_10 =15'b0;

   // m217_11 = W*in
   wire signed [14:0] m217_11;
   assign m217_11 =15'b0;

   // m217_12 = W*in
   wire signed [14:0] m217_12;
   assign m217_12 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_13 = W*in
   wire signed [14:0] m217_13;
   assign m217_13 =15'b0;

   // m217_14 = W*in
   wire signed [14:0] m217_14;
   assign m217_14 =15'b0;

   // m217_15 = W*in
   wire signed [14:0] m217_15;
   assign m217_15 =15'b0;

   // m217_16 = W*in
   wire signed [14:0] m217_16;
   assign m217_16 =15'b0;

   // m217_17 = W*in
   wire signed [14:0] m217_17;
   assign m217_17 =15'b0;

   // m217_18 = W*in
   wire signed [14:0] m217_18;
   assign m217_18 =15'b0;

   // m217_19 = W*in
   wire signed [14:0] m217_19;
   assign m217_19 =15'b0;

   // m217_20 = W*in
   wire signed [14:0] m217_20;
   assign m217_20 =15'b0;

   // m217_21 = W*in
   wire signed [14:0] m217_21;
   assign m217_21 =15'b0;

   // m217_22 = W*in
   wire signed [14:0] m217_22;
   assign m217_22 =15'b0;

   // m217_23 = W*in
   wire signed [14:0] m217_23;
   assign m217_23 =15'b0;

   // m217_24 = W*in
   wire signed [14:0] m217_24;
   assign m217_24 =15'b0;

   // m217_25 = W*in
   wire signed [14:0] m217_25;
   assign m217_25 =15'b0;

   // m217_26 = W*in
   wire signed [14:0] m217_26;
   assign m217_26 =15'b0;

   // m217_27 = W*in
   wire signed [14:0] m217_27;
   assign m217_27 =15'b0;

   // m217_28 = W*in
   wire signed [14:0] m217_28;
   assign m217_28 =15'b0;

   // m217_29 = W*in
   wire signed [14:0] m217_29;
   assign m217_29 ={ {4{neg217[14]}} , neg217[14:4] };

   // m217_30 = W*in
   wire signed [14:0] m217_30;
   assign m217_30 =15'b0;

   // m217_31 = W*in
   wire signed [14:0] m217_31;
   assign m217_31 =15'b0;

   // m217_32 = W*in
   wire signed [14:0] m217_32;
   assign m217_32 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_33 = W*in
   wire signed [14:0] m217_33;
   assign m217_33 =15'b0;

   // m217_34 = W*in
   wire signed [14:0] m217_34;
   assign m217_34 =15'b0;

   // m217_35 = W*in
   wire signed [14:0] m217_35;
   assign m217_35 =15'b0;

   // m217_36 = W*in
   wire signed [14:0] m217_36;
   assign m217_36 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_37 = W*in
   wire signed [14:0] m217_37;
   assign m217_37 =15'b0;

   // m217_38 = W*in
   wire signed [14:0] m217_38;
   assign m217_38 ={ {3{in217[14]}} , in217[14:3] };

   // m217_39 = W*in
   wire signed [14:0] m217_39;
   assign m217_39 =15'b0;

   // m217_40 = W*in
   wire signed [14:0] m217_40;
   assign m217_40 =15'b0;

   // m217_41 = W*in
   wire signed [14:0] m217_41;
   assign m217_41 =15'b0;

   // m217_42 = W*in
   wire signed [14:0] m217_42;
   assign m217_42 =15'b0;

   // m217_43 = W*in
   wire signed [14:0] m217_43;
   assign m217_43 =15'b0;

   // m217_44 = W*in
   wire signed [14:0] m217_44;
   assign m217_44 =15'b0;

   // m217_45 = W*in
   wire signed [14:0] m217_45;
   assign m217_45 ={ {2{in217[14]}} , in217[14:2] };

   // m217_46 = W*in
   wire signed [14:0] m217_46;
   assign m217_46 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_47 = W*in
   wire signed [14:0] m217_47;
   assign m217_47 =15'b0;

   // m217_48 = W*in
   wire signed [14:0] m217_48;
   assign m217_48 =15'b0;

   // m217_49 = W*in
   wire signed [14:0] m217_49;
   assign m217_49 =15'b0;

   // m217_50 = W*in
   wire signed [14:0] m217_50;
   assign m217_50 =15'b0;

   // m217_51 = W*in
   wire signed [14:0] m217_51;
   assign m217_51 =15'b0;

   // m217_52 = W*in
   wire signed [14:0] m217_52;
   assign m217_52 =15'b0;

   // m217_53 = W*in
   wire signed [14:0] m217_53;
   assign m217_53 =15'b0;

   // m217_54 = W*in
   wire signed [14:0] m217_54;
   assign m217_54 =15'b0;

   // m217_55 = W*in
   wire signed [14:0] m217_55;
   assign m217_55 =15'b0;

   // m217_56 = W*in
   wire signed [14:0] m217_56;
   assign m217_56 =15'b0;

   // m217_57 = W*in
   wire signed [14:0] m217_57;
   assign m217_57 =15'b0;

   // m217_58 = W*in
   wire signed [14:0] m217_58;
   assign m217_58 ={ {3{in217[14]}} , in217[14:3] };

   // m217_59 = W*in
   wire signed [14:0] m217_59;
   assign m217_59 =15'b0;

   // m217_60 = W*in
   wire signed [14:0] m217_60;
   assign m217_60 =15'b0;

   // m217_61 = W*in
   wire signed [14:0] m217_61;
   assign m217_61 =15'b0;

   // m217_62 = W*in
   wire signed [14:0] m217_62;
   assign m217_62 =15'b0;

   // m217_63 = W*in
   wire signed [14:0] m217_63;
   assign m217_63 =15'b0;

   // m217_64 = W*in
   wire signed [14:0] m217_64;
   assign m217_64 ={ {3{in217[14]}} , in217[14:3] };

   // m217_65 = W*in
   wire signed [14:0] m217_65;
   assign m217_65 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_66 = W*in
   wire signed [14:0] m217_66;
   assign m217_66 =15'b0;

   // m217_67 = W*in
   wire signed [14:0] m217_67;
   assign m217_67 =15'b0;

   // m217_68 = W*in
   wire signed [14:0] m217_68;
   assign m217_68 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_69 = W*in
   wire signed [14:0] m217_69;
   assign m217_69 =15'b0;

   // m217_70 = W*in
   wire signed [14:0] m217_70;
   assign m217_70 =15'b0;

   // m217_71 = W*in
   wire signed [14:0] m217_71;
   assign m217_71 =15'b0;

   // m217_72 = W*in
   wire signed [14:0] m217_72;
   assign m217_72 =15'b0;

   // m217_73 = W*in
   wire signed [14:0] m217_73;
   assign m217_73 =15'b0;

   // m217_74 = W*in
   wire signed [14:0] m217_74;
   assign m217_74 ={ {3{in217[14]}} , in217[14:3] };

   // m217_75 = W*in
   wire signed [14:0] m217_75;
   assign m217_75 =15'b0;

   // m217_76 = W*in
   wire signed [14:0] m217_76;
   assign m217_76 =15'b0;

   // m217_77 = W*in
   wire signed [14:0] m217_77;
   assign m217_77 =15'b0;

   // m217_78 = W*in
   wire signed [14:0] m217_78;
   assign m217_78 =15'b0;

   // m217_79 = W*in
   wire signed [14:0] m217_79;
   assign m217_79 =15'b0;

   // m217_80 = W*in
   wire signed [14:0] m217_80;
   assign m217_80 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_81 = W*in
   wire signed [14:0] m217_81;
   assign m217_81 =15'b0;

   // m217_82 = W*in
   wire signed [14:0] m217_82;
   assign m217_82 =15'b0;

   // m217_83 = W*in
   wire signed [14:0] m217_83;
   assign m217_83 =15'b0;

   // m217_84 = W*in
   wire signed [14:0] m217_84;
   assign m217_84 =15'b0;

   // m217_85 = W*in
   wire signed [14:0] m217_85;
   assign m217_85 =15'b0;

   // m217_86 = W*in
   wire signed [14:0] m217_86;
   assign m217_86 =15'b0;

   // m217_87 = W*in
   wire signed [14:0] m217_87;
   assign m217_87 =15'b0;

   // m217_88 = W*in
   wire signed [14:0] m217_88;
   assign m217_88 =15'b0;

   // m217_89 = W*in
   wire signed [14:0] m217_89;
   assign m217_89 =15'b0;

   // m217_90 = W*in
   wire signed [14:0] m217_90;
   assign m217_90 =15'b0;

   // m217_91 = W*in
   wire signed [14:0] m217_91;
   assign m217_91 =15'b0;

   // m217_92 = W*in
   wire signed [14:0] m217_92;
   assign m217_92 ={ {3{in217[14]}} , in217[14:3] };

   // m217_93 = W*in
   wire signed [14:0] m217_93;
   assign m217_93 ={ {3{neg217[14]}} , neg217[14:3] };

   // m217_94 = W*in
   wire signed [14:0] m217_94;
   assign m217_94 =15'b0;

   // m217_95 = W*in
   wire signed [14:0] m217_95;
   assign m217_95 =15'b0;

   // m217_96 = W*in
   wire signed [14:0] m217_96;
   assign m217_96 =15'b0;

   // m217_97 = W*in
   wire signed [14:0] m217_97;
   assign m217_97 =15'b0;

   // m217_98 = W*in
   wire signed [14:0] m217_98;
   assign m217_98 =15'b0;

   // m217_99 = W*in
   wire signed [14:0] m217_99;
   assign m217_99 ={ {3{in217[14]}} , in217[14:3] };

   // m217_100 = W*in
   wire signed [14:0] m217_100;
   assign m217_100 =15'b0;

   // m218_1 = W*in
   wire signed [14:0] m218_1;
   assign m218_1 =15'b0;

   // m218_2 = W*in
   wire signed [14:0] m218_2;
   assign m218_2 =15'b0;

   // m218_3 = W*in
   wire signed [14:0] m218_3;
   assign m218_3 =15'b0;

   // m218_4 = W*in
   wire signed [14:0] m218_4;
   assign m218_4 =15'b0;

   // m218_5 = W*in
   wire signed [14:0] m218_5;
   assign m218_5 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_6 = W*in
   wire signed [14:0] m218_6;
   assign m218_6 =15'b0;

   // m218_7 = W*in
   wire signed [14:0] m218_7;
   assign m218_7 =15'b0;

   // m218_8 = W*in
   wire signed [14:0] m218_8;
   assign m218_8 =15'b0;

   // m218_9 = W*in
   wire signed [14:0] m218_9;
   assign m218_9 =15'b0;

   // m218_10 = W*in
   wire signed [14:0] m218_10;
   assign m218_10 =15'b0;

   // m218_11 = W*in
   wire signed [14:0] m218_11;
   assign m218_11 ={ {3{in218[14]}} , in218[14:3] };

   // m218_12 = W*in
   wire signed [14:0] m218_12;
   assign m218_12 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_13 = W*in
   wire signed [14:0] m218_13;
   assign m218_13 ={ {4{neg218[14]}} , neg218[14:4] };

   // m218_14 = W*in
   wire signed [14:0] m218_14;
   assign m218_14 =15'b0;

   // m218_15 = W*in
   wire signed [14:0] m218_15;
   assign m218_15 =15'b0;

   // m218_16 = W*in
   wire signed [14:0] m218_16;
   assign m218_16 =15'b0;

   // m218_17 = W*in
   wire signed [14:0] m218_17;
   assign m218_17 =15'b0;

   // m218_18 = W*in
   wire signed [14:0] m218_18;
   assign m218_18 =15'b0;

   // m218_19 = W*in
   wire signed [14:0] m218_19;
   assign m218_19 =15'b0;

   // m218_20 = W*in
   wire signed [14:0] m218_20;
   assign m218_20 =15'b0;

   // m218_21 = W*in
   wire signed [14:0] m218_21;
   assign m218_21 ={ {3{in218[14]}} , in218[14:3] };

   // m218_22 = W*in
   wire signed [14:0] m218_22;
   assign m218_22 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_23 = W*in
   wire signed [14:0] m218_23;
   assign m218_23 ={ {3{in218[14]}} , in218[14:3] };

   // m218_24 = W*in
   wire signed [14:0] m218_24;
   assign m218_24 =15'b0;

   // m218_25 = W*in
   wire signed [14:0] m218_25;
   assign m218_25 =15'b0;

   // m218_26 = W*in
   wire signed [14:0] m218_26;
   assign m218_26 =15'b0;

   // m218_27 = W*in
   wire signed [14:0] m218_27;
   assign m218_27 ={ {2{neg218[14]}} , neg218[14:2] };

   // m218_28 = W*in
   wire signed [14:0] m218_28;
   assign m218_28 =15'b0;

   // m218_29 = W*in
   wire signed [14:0] m218_29;
   assign m218_29 =15'b0;

   // m218_30 = W*in
   wire signed [14:0] m218_30;
   assign m218_30 =15'b0;

   // m218_31 = W*in
   wire signed [14:0] m218_31;
   assign m218_31 ={ {4{neg218[14]}} , neg218[14:4] };

   // m218_32 = W*in
   wire signed [14:0] m218_32;
   assign m218_32 =15'b0;

   // m218_33 = W*in
   wire signed [14:0] m218_33;
   assign m218_33 =15'b0;

   // m218_34 = W*in
   wire signed [14:0] m218_34;
   assign m218_34 =15'b0;

   // m218_35 = W*in
   wire signed [14:0] m218_35;
   assign m218_35 =15'b0;

   // m218_36 = W*in
   wire signed [14:0] m218_36;
   assign m218_36 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_37 = W*in
   wire signed [14:0] m218_37;
   assign m218_37 ={ {4{in218[14]}} , in218[14:4] };

   // m218_38 = W*in
   wire signed [14:0] m218_38;
   assign m218_38 =15'b0;

   // m218_39 = W*in
   wire signed [14:0] m218_39;
   assign m218_39 =15'b0;

   // m218_40 = W*in
   wire signed [14:0] m218_40;
   assign m218_40 =15'b0;

   // m218_41 = W*in
   wire signed [14:0] m218_41;
   assign m218_41 =15'b0;

   // m218_42 = W*in
   wire signed [14:0] m218_42;
   assign m218_42 =15'b0;

   // m218_43 = W*in
   wire signed [14:0] m218_43;
   assign m218_43 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_44 = W*in
   wire signed [14:0] m218_44;
   assign m218_44 =15'b0;

   // m218_45 = W*in
   wire signed [14:0] m218_45;
   assign m218_45 ={ {3{in218[14]}} , in218[14:3] };

   // m218_46 = W*in
   wire signed [14:0] m218_46;
   assign m218_46 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_47 = W*in
   wire signed [14:0] m218_47;
   assign m218_47 =15'b0;

   // m218_48 = W*in
   wire signed [14:0] m218_48;
   assign m218_48 =15'b0;

   // m218_49 = W*in
   wire signed [14:0] m218_49;
   assign m218_49 =15'b0;

   // m218_50 = W*in
   wire signed [14:0] m218_50;
   assign m218_50 =15'b0;

   // m218_51 = W*in
   wire signed [14:0] m218_51;
   assign m218_51 =15'b0;

   // m218_52 = W*in
   wire signed [14:0] m218_52;
   assign m218_52 =15'b0;

   // m218_53 = W*in
   wire signed [14:0] m218_53;
   assign m218_53 =15'b0;

   // m218_54 = W*in
   wire signed [14:0] m218_54;
   assign m218_54 =15'b0;

   // m218_55 = W*in
   wire signed [14:0] m218_55;
   assign m218_55 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_56 = W*in
   wire signed [14:0] m218_56;
   assign m218_56 ={ {3{in218[14]}} , in218[14:3] };

   // m218_57 = W*in
   wire signed [14:0] m218_57;
   assign m218_57 =15'b0;

   // m218_58 = W*in
   wire signed [14:0] m218_58;
   assign m218_58 =15'b0;

   // m218_59 = W*in
   wire signed [14:0] m218_59;
   assign m218_59 =15'b0;

   // m218_60 = W*in
   wire signed [14:0] m218_60;
   assign m218_60 ={ {4{neg218[14]}} , neg218[14:4] };

   // m218_61 = W*in
   wire signed [14:0] m218_61;
   assign m218_61 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_62 = W*in
   wire signed [14:0] m218_62;
   assign m218_62 =15'b0;

   // m218_63 = W*in
   wire signed [14:0] m218_63;
   assign m218_63 =15'b0;

   // m218_64 = W*in
   wire signed [14:0] m218_64;
   assign m218_64 =15'b0;

   // m218_65 = W*in
   wire signed [14:0] m218_65;
   assign m218_65 =15'b0;

   // m218_66 = W*in
   wire signed [14:0] m218_66;
   assign m218_66 =15'b0;

   // m218_67 = W*in
   wire signed [14:0] m218_67;
   assign m218_67 =15'b0;

   // m218_68 = W*in
   wire signed [14:0] m218_68;
   assign m218_68 =15'b0;

   // m218_69 = W*in
   wire signed [14:0] m218_69;
   assign m218_69 =15'b0;

   // m218_70 = W*in
   wire signed [14:0] m218_70;
   assign m218_70 =15'b0;

   // m218_71 = W*in
   wire signed [14:0] m218_71;
   assign m218_71 =15'b0;

   // m218_72 = W*in
   wire signed [14:0] m218_72;
   assign m218_72 =15'b0;

   // m218_73 = W*in
   wire signed [14:0] m218_73;
   assign m218_73 =15'b0;

   // m218_74 = W*in
   wire signed [14:0] m218_74;
   assign m218_74 ={ {4{in218[14]}} , in218[14:4] };

   // m218_75 = W*in
   wire signed [14:0] m218_75;
   assign m218_75 =15'b0;

   // m218_76 = W*in
   wire signed [14:0] m218_76;
   assign m218_76 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_77 = W*in
   wire signed [14:0] m218_77;
   assign m218_77 =15'b0;

   // m218_78 = W*in
   wire signed [14:0] m218_78;
   assign m218_78 =15'b0;

   // m218_79 = W*in
   wire signed [14:0] m218_79;
   assign m218_79 =15'b0;

   // m218_80 = W*in
   wire signed [14:0] m218_80;
   assign m218_80 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_81 = W*in
   wire signed [14:0] m218_81;
   assign m218_81 =15'b0;

   // m218_82 = W*in
   wire signed [14:0] m218_82;
   assign m218_82 ={ {3{neg218[14]}} , neg218[14:3] };

   // m218_83 = W*in
   wire signed [14:0] m218_83;
   assign m218_83 =15'b0;

   // m218_84 = W*in
   wire signed [14:0] m218_84;
   assign m218_84 =15'b0;

   // m218_85 = W*in
   wire signed [14:0] m218_85;
   assign m218_85 =15'b0;

   // m218_86 = W*in
   wire signed [14:0] m218_86;
   assign m218_86 ={ {3{in218[14]}} , in218[14:3] };

   // m218_87 = W*in
   wire signed [14:0] m218_87;
   assign m218_87 =15'b0;

   // m218_88 = W*in
   wire signed [14:0] m218_88;
   assign m218_88 =15'b0;

   // m218_89 = W*in
   wire signed [14:0] m218_89;
   assign m218_89 ={ {3{in218[14]}} , in218[14:3] };

   // m218_90 = W*in
   wire signed [14:0] m218_90;
   assign m218_90 =15'b0;

   // m218_91 = W*in
   wire signed [14:0] m218_91;
   assign m218_91 =15'b0;

   // m218_92 = W*in
   wire signed [14:0] m218_92;
   assign m218_92 =15'b0;

   // m218_93 = W*in
   wire signed [14:0] m218_93;
   assign m218_93 =15'b0;

   // m218_94 = W*in
   wire signed [14:0] m218_94;
   assign m218_94 =15'b0;

   // m218_95 = W*in
   wire signed [14:0] m218_95;
   assign m218_95 =15'b0;

   // m218_96 = W*in
   wire signed [14:0] m218_96;
   assign m218_96 =15'b0;

   // m218_97 = W*in
   wire signed [14:0] m218_97;
   assign m218_97 =15'b0;

   // m218_98 = W*in
   wire signed [14:0] m218_98;
   assign m218_98 =15'b0;

   // m218_99 = W*in
   wire signed [14:0] m218_99;
   assign m218_99 =15'b0;

   // m218_100 = W*in
   wire signed [14:0] m218_100;
   assign m218_100 =15'b0;

   // m219_1 = W*in
   wire signed [14:0] m219_1;
   assign m219_1 =15'b0;

   // m219_2 = W*in
   wire signed [14:0] m219_2;
   assign m219_2 =15'b0;

   // m219_3 = W*in
   wire signed [14:0] m219_3;
   assign m219_3 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_4 = W*in
   wire signed [14:0] m219_4;
   assign m219_4 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_5 = W*in
   wire signed [14:0] m219_5;
   assign m219_5 =15'b0;

   // m219_6 = W*in
   wire signed [14:0] m219_6;
   assign m219_6 =15'b0;

   // m219_7 = W*in
   wire signed [14:0] m219_7;
   assign m219_7 =15'b0;

   // m219_8 = W*in
   wire signed [14:0] m219_8;
   assign m219_8 ={ {3{in219[14]}} , in219[14:3] };

   // m219_9 = W*in
   wire signed [14:0] m219_9;
   assign m219_9 =15'b0;

   // m219_10 = W*in
   wire signed [14:0] m219_10;
   assign m219_10 ={ {3{in219[14]}} , in219[14:3] };

   // m219_11 = W*in
   wire signed [14:0] m219_11;
   assign m219_11 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_12 = W*in
   wire signed [14:0] m219_12;
   assign m219_12 =15'b0;

   // m219_13 = W*in
   wire signed [14:0] m219_13;
   assign m219_13 =15'b0;

   // m219_14 = W*in
   wire signed [14:0] m219_14;
   assign m219_14 =15'b0;

   // m219_15 = W*in
   wire signed [14:0] m219_15;
   assign m219_15 =15'b0;

   // m219_16 = W*in
   wire signed [14:0] m219_16;
   assign m219_16 =15'b0;

   // m219_17 = W*in
   wire signed [14:0] m219_17;
   assign m219_17 =15'b0;

   // m219_18 = W*in
   wire signed [14:0] m219_18;
   assign m219_18 =15'b0;

   // m219_19 = W*in
   wire signed [14:0] m219_19;
   assign m219_19 =15'b0;

   // m219_20 = W*in
   wire signed [14:0] m219_20;
   assign m219_20 =15'b0;

   // m219_21 = W*in
   wire signed [14:0] m219_21;
   assign m219_21 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_22 = W*in
   wire signed [14:0] m219_22;
   assign m219_22 =15'b0;

   // m219_23 = W*in
   wire signed [14:0] m219_23;
   assign m219_23 =15'b0;

   // m219_24 = W*in
   wire signed [14:0] m219_24;
   assign m219_24 =15'b0;

   // m219_25 = W*in
   wire signed [14:0] m219_25;
   assign m219_25 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_26 = W*in
   wire signed [14:0] m219_26;
   assign m219_26 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_27 = W*in
   wire signed [14:0] m219_27;
   assign m219_27 =15'b0;

   // m219_28 = W*in
   wire signed [14:0] m219_28;
   assign m219_28 =15'b0;

   // m219_29 = W*in
   wire signed [14:0] m219_29;
   assign m219_29 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_30 = W*in
   wire signed [14:0] m219_30;
   assign m219_30 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_31 = W*in
   wire signed [14:0] m219_31;
   assign m219_31 ={ {3{in219[14]}} , in219[14:3] };

   // m219_32 = W*in
   wire signed [14:0] m219_32;
   assign m219_32 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_33 = W*in
   wire signed [14:0] m219_33;
   assign m219_33 =15'b0;

   // m219_34 = W*in
   wire signed [14:0] m219_34;
   assign m219_34 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_35 = W*in
   wire signed [14:0] m219_35;
   assign m219_35 =15'b0;

   // m219_36 = W*in
   wire signed [14:0] m219_36;
   assign m219_36 =15'b0;

   // m219_37 = W*in
   wire signed [14:0] m219_37;
   assign m219_37 =15'b0;

   // m219_38 = W*in
   wire signed [14:0] m219_38;
   assign m219_38 =15'b0;

   // m219_39 = W*in
   wire signed [14:0] m219_39;
   assign m219_39 ={ {3{in219[14]}} , in219[14:3] };

   // m219_40 = W*in
   wire signed [14:0] m219_40;
   assign m219_40 =15'b0;

   // m219_41 = W*in
   wire signed [14:0] m219_41;
   assign m219_41 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_42 = W*in
   wire signed [14:0] m219_42;
   assign m219_42 =15'b0;

   // m219_43 = W*in
   wire signed [14:0] m219_43;
   assign m219_43 =15'b0;

   // m219_44 = W*in
   wire signed [14:0] m219_44;
   assign m219_44 =15'b0;

   // m219_45 = W*in
   wire signed [14:0] m219_45;
   assign m219_45 =15'b0;

   // m219_46 = W*in
   wire signed [14:0] m219_46;
   assign m219_46 =15'b0;

   // m219_47 = W*in
   wire signed [14:0] m219_47;
   assign m219_47 =15'b0;

   // m219_48 = W*in
   wire signed [14:0] m219_48;
   assign m219_48 ={ {4{in219[14]}} , in219[14:4] };

   // m219_49 = W*in
   wire signed [14:0] m219_49;
   assign m219_49 =15'b0;

   // m219_50 = W*in
   wire signed [14:0] m219_50;
   assign m219_50 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_51 = W*in
   wire signed [14:0] m219_51;
   assign m219_51 ={ {3{in219[14]}} , in219[14:3] };

   // m219_52 = W*in
   wire signed [14:0] m219_52;
   assign m219_52 =15'b0;

   // m219_53 = W*in
   wire signed [14:0] m219_53;
   assign m219_53 =15'b0;

   // m219_54 = W*in
   wire signed [14:0] m219_54;
   assign m219_54 =15'b0;

   // m219_55 = W*in
   wire signed [14:0] m219_55;
   assign m219_55 =15'b0;

   // m219_56 = W*in
   wire signed [14:0] m219_56;
   assign m219_56 =15'b0;

   // m219_57 = W*in
   wire signed [14:0] m219_57;
   assign m219_57 =15'b0;

   // m219_58 = W*in
   wire signed [14:0] m219_58;
   assign m219_58 =15'b0;

   // m219_59 = W*in
   wire signed [14:0] m219_59;
   assign m219_59 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_60 = W*in
   wire signed [14:0] m219_60;
   assign m219_60 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_61 = W*in
   wire signed [14:0] m219_61;
   assign m219_61 =15'b0;

   // m219_62 = W*in
   wire signed [14:0] m219_62;
   assign m219_62 =15'b0;

   // m219_63 = W*in
   wire signed [14:0] m219_63;
   assign m219_63 ={ {4{in219[14]}} , in219[14:4] };

   // m219_64 = W*in
   wire signed [14:0] m219_64;
   assign m219_64 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_65 = W*in
   wire signed [14:0] m219_65;
   assign m219_65 =15'b0;

   // m219_66 = W*in
   wire signed [14:0] m219_66;
   assign m219_66 ={ {4{in219[14]}} , in219[14:4] };

   // m219_67 = W*in
   wire signed [14:0] m219_67;
   assign m219_67 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_68 = W*in
   wire signed [14:0] m219_68;
   assign m219_68 =15'b0;

   // m219_69 = W*in
   wire signed [14:0] m219_69;
   assign m219_69 =15'b0;

   // m219_70 = W*in
   wire signed [14:0] m219_70;
   assign m219_70 =15'b0;

   // m219_71 = W*in
   wire signed [14:0] m219_71;
   assign m219_71 ={ {3{in219[14]}} , in219[14:3] };

   // m219_72 = W*in
   wire signed [14:0] m219_72;
   assign m219_72 =15'b0;

   // m219_73 = W*in
   wire signed [14:0] m219_73;
   assign m219_73 =15'b0;

   // m219_74 = W*in
   wire signed [14:0] m219_74;
   assign m219_74 =15'b0;

   // m219_75 = W*in
   wire signed [14:0] m219_75;
   assign m219_75 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_76 = W*in
   wire signed [14:0] m219_76;
   assign m219_76 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_77 = W*in
   wire signed [14:0] m219_77;
   assign m219_77 =15'b0;

   // m219_78 = W*in
   wire signed [14:0] m219_78;
   assign m219_78 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_79 = W*in
   wire signed [14:0] m219_79;
   assign m219_79 =15'b0;

   // m219_80 = W*in
   wire signed [14:0] m219_80;
   assign m219_80 ={ {4{neg219[14]}} , neg219[14:4] };

   // m219_81 = W*in
   wire signed [14:0] m219_81;
   assign m219_81 =15'b0;

   // m219_82 = W*in
   wire signed [14:0] m219_82;
   assign m219_82 =15'b0;

   // m219_83 = W*in
   wire signed [14:0] m219_83;
   assign m219_83 ={ {3{in219[14]}} , in219[14:3] };

   // m219_84 = W*in
   wire signed [14:0] m219_84;
   assign m219_84 =15'b0;

   // m219_85 = W*in
   wire signed [14:0] m219_85;
   assign m219_85 =15'b0;

   // m219_86 = W*in
   wire signed [14:0] m219_86;
   assign m219_86 =15'b0;

   // m219_87 = W*in
   wire signed [14:0] m219_87;
   assign m219_87 =15'b0;

   // m219_88 = W*in
   wire signed [14:0] m219_88;
   assign m219_88 =15'b0;

   // m219_89 = W*in
   wire signed [14:0] m219_89;
   assign m219_89 ={ {3{in219[14]}} , in219[14:3] };

   // m219_90 = W*in
   wire signed [14:0] m219_90;
   assign m219_90 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_91 = W*in
   wire signed [14:0] m219_91;
   assign m219_91 =15'b0;

   // m219_92 = W*in
   wire signed [14:0] m219_92;
   assign m219_92 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_93 = W*in
   wire signed [14:0] m219_93;
   assign m219_93 =15'b0;

   // m219_94 = W*in
   wire signed [14:0] m219_94;
   assign m219_94 =15'b0;

   // m219_95 = W*in
   wire signed [14:0] m219_95;
   assign m219_95 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_96 = W*in
   wire signed [14:0] m219_96;
   assign m219_96 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_97 = W*in
   wire signed [14:0] m219_97;
   assign m219_97 =15'b0;

   // m219_98 = W*in
   wire signed [14:0] m219_98;
   assign m219_98 ={ {3{neg219[14]}} , neg219[14:3] };

   // m219_99 = W*in
   wire signed [14:0] m219_99;
   assign m219_99 =15'b0;

   // m219_100 = W*in
   wire signed [14:0] m219_100;
   assign m219_100 =15'b0;

   // m220_1 = W*in
   wire signed [14:0] m220_1;
   assign m220_1 =15'b0;

   // m220_2 = W*in
   wire signed [14:0] m220_2;
   assign m220_2 =15'b0;

   // m220_3 = W*in
   wire signed [14:0] m220_3;
   assign m220_3 =15'b0;

   // m220_4 = W*in
   wire signed [14:0] m220_4;
   assign m220_4 ={ {4{in220[14]}} , in220[14:4] };

   // m220_5 = W*in
   wire signed [14:0] m220_5;
   assign m220_5 =15'b0;

   // m220_6 = W*in
   wire signed [14:0] m220_6;
   assign m220_6 =15'b0;

   // m220_7 = W*in
   wire signed [14:0] m220_7;
   assign m220_7 =15'b0;

   // m220_8 = W*in
   wire signed [14:0] m220_8;
   assign m220_8 =15'b0;

   // m220_9 = W*in
   wire signed [14:0] m220_9;
   assign m220_9 =15'b0;

   // m220_10 = W*in
   wire signed [14:0] m220_10;
   assign m220_10 =15'b0;

   // m220_11 = W*in
   wire signed [14:0] m220_11;
   assign m220_11 =15'b0;

   // m220_12 = W*in
   wire signed [14:0] m220_12;
   assign m220_12 =15'b0;

   // m220_13 = W*in
   wire signed [14:0] m220_13;
   assign m220_13 =15'b0;

   // m220_14 = W*in
   wire signed [14:0] m220_14;
   assign m220_14 =15'b0;

   // m220_15 = W*in
   wire signed [14:0] m220_15;
   assign m220_15 =15'b0;

   // m220_16 = W*in
   wire signed [14:0] m220_16;
   assign m220_16 =15'b0;

   // m220_17 = W*in
   wire signed [14:0] m220_17;
   assign m220_17 =15'b0;

   // m220_18 = W*in
   wire signed [14:0] m220_18;
   assign m220_18 ={ {4{in220[14]}} , in220[14:4] };

   // m220_19 = W*in
   wire signed [14:0] m220_19;
   assign m220_19 =15'b0;

   // m220_20 = W*in
   wire signed [14:0] m220_20;
   assign m220_20 =15'b0;

   // m220_21 = W*in
   wire signed [14:0] m220_21;
   assign m220_21 =15'b0;

   // m220_22 = W*in
   wire signed [14:0] m220_22;
   assign m220_22 =15'b0;

   // m220_23 = W*in
   wire signed [14:0] m220_23;
   assign m220_23 =15'b0;

   // m220_24 = W*in
   wire signed [14:0] m220_24;
   assign m220_24 =15'b0;

   // m220_25 = W*in
   wire signed [14:0] m220_25;
   assign m220_25 =15'b0;

   // m220_26 = W*in
   wire signed [14:0] m220_26;
   assign m220_26 ={ {4{in220[14]}} , in220[14:4] };

   // m220_27 = W*in
   wire signed [14:0] m220_27;
   assign m220_27 =15'b0;

   // m220_28 = W*in
   wire signed [14:0] m220_28;
   assign m220_28 =15'b0;

   // m220_29 = W*in
   wire signed [14:0] m220_29;
   assign m220_29 ={ {4{in220[14]}} , in220[14:4] };

   // m220_30 = W*in
   wire signed [14:0] m220_30;
   assign m220_30 =15'b0;

   // m220_31 = W*in
   wire signed [14:0] m220_31;
   assign m220_31 ={ {4{in220[14]}} , in220[14:4] };

   // m220_32 = W*in
   wire signed [14:0] m220_32;
   assign m220_32 =15'b0;

   // m220_33 = W*in
   wire signed [14:0] m220_33;
   assign m220_33 =15'b0;

   // m220_34 = W*in
   wire signed [14:0] m220_34;
   assign m220_34 =15'b0;

   // m220_35 = W*in
   wire signed [14:0] m220_35;
   assign m220_35 =15'b0;

   // m220_36 = W*in
   wire signed [14:0] m220_36;
   assign m220_36 =15'b0;

   // m220_37 = W*in
   wire signed [14:0] m220_37;
   assign m220_37 =15'b0;

   // m220_38 = W*in
   wire signed [14:0] m220_38;
   assign m220_38 =15'b0;

   // m220_39 = W*in
   wire signed [14:0] m220_39;
   assign m220_39 =15'b0;

   // m220_40 = W*in
   wire signed [14:0] m220_40;
   assign m220_40 =15'b0;

   // m220_41 = W*in
   wire signed [14:0] m220_41;
   assign m220_41 =15'b0;

   // m220_42 = W*in
   wire signed [14:0] m220_42;
   assign m220_42 =15'b0;

   // m220_43 = W*in
   wire signed [14:0] m220_43;
   assign m220_43 =15'b0;

   // m220_44 = W*in
   wire signed [14:0] m220_44;
   assign m220_44 =15'b0;

   // m220_45 = W*in
   wire signed [14:0] m220_45;
   assign m220_45 =15'b0;

   // m220_46 = W*in
   wire signed [14:0] m220_46;
   assign m220_46 =15'b0;

   // m220_47 = W*in
   wire signed [14:0] m220_47;
   assign m220_47 =15'b0;

   // m220_48 = W*in
   wire signed [14:0] m220_48;
   assign m220_48 =15'b0;

   // m220_49 = W*in
   wire signed [14:0] m220_49;
   assign m220_49 =15'b0;

   // m220_50 = W*in
   wire signed [14:0] m220_50;
   assign m220_50 =15'b0;

   // m220_51 = W*in
   wire signed [14:0] m220_51;
   assign m220_51 =15'b0;

   // m220_52 = W*in
   wire signed [14:0] m220_52;
   assign m220_52 =15'b0;

   // m220_53 = W*in
   wire signed [14:0] m220_53;
   assign m220_53 =15'b0;

   // m220_54 = W*in
   wire signed [14:0] m220_54;
   assign m220_54 =15'b0;

   // m220_55 = W*in
   wire signed [14:0] m220_55;
   assign m220_55 =15'b0;

   // m220_56 = W*in
   wire signed [14:0] m220_56;
   assign m220_56 =15'b0;

   // m220_57 = W*in
   wire signed [14:0] m220_57;
   assign m220_57 =15'b0;

   // m220_58 = W*in
   wire signed [14:0] m220_58;
   assign m220_58 =15'b0;

   // m220_59 = W*in
   wire signed [14:0] m220_59;
   assign m220_59 =15'b0;

   // m220_60 = W*in
   wire signed [14:0] m220_60;
   assign m220_60 =15'b0;

   // m220_61 = W*in
   wire signed [14:0] m220_61;
   assign m220_61 =15'b0;

   // m220_62 = W*in
   wire signed [14:0] m220_62;
   assign m220_62 =15'b0;

   // m220_63 = W*in
   wire signed [14:0] m220_63;
   assign m220_63 ={ {4{in220[14]}} , in220[14:4] };

   // m220_64 = W*in
   wire signed [14:0] m220_64;
   assign m220_64 ={ {4{neg220[14]}} , neg220[14:4] };

   // m220_65 = W*in
   wire signed [14:0] m220_65;
   assign m220_65 =15'b0;

   // m220_66 = W*in
   wire signed [14:0] m220_66;
   assign m220_66 ={ {3{in220[14]}} , in220[14:3] };

   // m220_67 = W*in
   wire signed [14:0] m220_67;
   assign m220_67 =15'b0;

   // m220_68 = W*in
   wire signed [14:0] m220_68;
   assign m220_68 =15'b0;

   // m220_69 = W*in
   wire signed [14:0] m220_69;
   assign m220_69 =15'b0;

   // m220_70 = W*in
   wire signed [14:0] m220_70;
   assign m220_70 =15'b0;

   // m220_71 = W*in
   wire signed [14:0] m220_71;
   assign m220_71 =15'b0;

   // m220_72 = W*in
   wire signed [14:0] m220_72;
   assign m220_72 =15'b0;

   // m220_73 = W*in
   wire signed [14:0] m220_73;
   assign m220_73 =15'b0;

   // m220_74 = W*in
   wire signed [14:0] m220_74;
   assign m220_74 =15'b0;

   // m220_75 = W*in
   wire signed [14:0] m220_75;
   assign m220_75 =15'b0;

   // m220_76 = W*in
   wire signed [14:0] m220_76;
   assign m220_76 =15'b0;

   // m220_77 = W*in
   wire signed [14:0] m220_77;
   assign m220_77 =15'b0;

   // m220_78 = W*in
   wire signed [14:0] m220_78;
   assign m220_78 =15'b0;

   // m220_79 = W*in
   wire signed [14:0] m220_79;
   assign m220_79 =15'b0;

   // m220_80 = W*in
   wire signed [14:0] m220_80;
   assign m220_80 =15'b0;

   // m220_81 = W*in
   wire signed [14:0] m220_81;
   assign m220_81 =15'b0;

   // m220_82 = W*in
   wire signed [14:0] m220_82;
   assign m220_82 =15'b0;

   // m220_83 = W*in
   wire signed [14:0] m220_83;
   assign m220_83 =15'b0;

   // m220_84 = W*in
   wire signed [14:0] m220_84;
   assign m220_84 =15'b0;

   // m220_85 = W*in
   wire signed [14:0] m220_85;
   assign m220_85 =15'b0;

   // m220_86 = W*in
   wire signed [14:0] m220_86;
   assign m220_86 =15'b0;

   // m220_87 = W*in
   wire signed [14:0] m220_87;
   assign m220_87 =15'b0;

   // m220_88 = W*in
   wire signed [14:0] m220_88;
   assign m220_88 =15'b0;

   // m220_89 = W*in
   wire signed [14:0] m220_89;
   assign m220_89 =15'b0;

   // m220_90 = W*in
   wire signed [14:0] m220_90;
   assign m220_90 =15'b0;

   // m220_91 = W*in
   wire signed [14:0] m220_91;
   assign m220_91 =15'b0;

   // m220_92 = W*in
   wire signed [14:0] m220_92;
   assign m220_92 =15'b0;

   // m220_93 = W*in
   wire signed [14:0] m220_93;
   assign m220_93 =15'b0;

   // m220_94 = W*in
   wire signed [14:0] m220_94;
   assign m220_94 =15'b0;

   // m220_95 = W*in
   wire signed [14:0] m220_95;
   assign m220_95 =15'b0;

   // m220_96 = W*in
   wire signed [14:0] m220_96;
   assign m220_96 =15'b0;

   // m220_97 = W*in
   wire signed [14:0] m220_97;
   assign m220_97 =15'b0;

   // m220_98 = W*in
   wire signed [14:0] m220_98;
   assign m220_98 =15'b0;

   // m220_99 = W*in
   wire signed [14:0] m220_99;
   assign m220_99 =15'b0;

   // m220_100 = W*in
   wire signed [14:0] m220_100;
   assign m220_100 =15'b0;

   // m221_1 = W*in
   wire signed [14:0] m221_1;
   assign m221_1 =15'b0;

   // m221_2 = W*in
   wire signed [14:0] m221_2;
   assign m221_2 =15'b0;

   // m221_3 = W*in
   wire signed [14:0] m221_3;
   assign m221_3 =15'b0;

   // m221_4 = W*in
   wire signed [14:0] m221_4;
   assign m221_4 ={ {4{neg221[14]}} , neg221[14:4] };

   // m221_5 = W*in
   wire signed [14:0] m221_5;
   assign m221_5 =15'b0;

   // m221_6 = W*in
   wire signed [14:0] m221_6;
   assign m221_6 =15'b0;

   // m221_7 = W*in
   wire signed [14:0] m221_7;
   assign m221_7 =15'b0;

   // m221_8 = W*in
   wire signed [14:0] m221_8;
   assign m221_8 =15'b0;

   // m221_9 = W*in
   wire signed [14:0] m221_9;
   assign m221_9 =15'b0;

   // m221_10 = W*in
   wire signed [14:0] m221_10;
   assign m221_10 =15'b0;

   // m221_11 = W*in
   wire signed [14:0] m221_11;
   assign m221_11 =15'b0;

   // m221_12 = W*in
   wire signed [14:0] m221_12;
   assign m221_12 =15'b0;

   // m221_13 = W*in
   wire signed [14:0] m221_13;
   assign m221_13 =15'b0;

   // m221_14 = W*in
   wire signed [14:0] m221_14;
   assign m221_14 =15'b0;

   // m221_15 = W*in
   wire signed [14:0] m221_15;
   assign m221_15 =15'b0;

   // m221_16 = W*in
   wire signed [14:0] m221_16;
   assign m221_16 =15'b0;

   // m221_17 = W*in
   wire signed [14:0] m221_17;
   assign m221_17 =15'b0;

   // m221_18 = W*in
   wire signed [14:0] m221_18;
   assign m221_18 =15'b0;

   // m221_19 = W*in
   wire signed [14:0] m221_19;
   assign m221_19 =15'b0;

   // m221_20 = W*in
   wire signed [14:0] m221_20;
   assign m221_20 =15'b0;

   // m221_21 = W*in
   wire signed [14:0] m221_21;
   assign m221_21 ={ {4{in221[14]}} , in221[14:4] };

   // m221_22 = W*in
   wire signed [14:0] m221_22;
   assign m221_22 =15'b0;

   // m221_23 = W*in
   wire signed [14:0] m221_23;
   assign m221_23 =15'b0;

   // m221_24 = W*in
   wire signed [14:0] m221_24;
   assign m221_24 =15'b0;

   // m221_25 = W*in
   wire signed [14:0] m221_25;
   assign m221_25 ={ {4{in221[14]}} , in221[14:4] };

   // m221_26 = W*in
   wire signed [14:0] m221_26;
   assign m221_26 =15'b0;

   // m221_27 = W*in
   wire signed [14:0] m221_27;
   assign m221_27 =15'b0;

   // m221_28 = W*in
   wire signed [14:0] m221_28;
   assign m221_28 ={ {4{neg221[14]}} , neg221[14:4] };

   // m221_29 = W*in
   wire signed [14:0] m221_29;
   assign m221_29 =15'b0;

   // m221_30 = W*in
   wire signed [14:0] m221_30;
   assign m221_30 =15'b0;

   // m221_31 = W*in
   wire signed [14:0] m221_31;
   assign m221_31 =15'b0;

   // m221_32 = W*in
   wire signed [14:0] m221_32;
   assign m221_32 ={ {4{neg221[14]}} , neg221[14:4] };

   // m221_33 = W*in
   wire signed [14:0] m221_33;
   assign m221_33 ={ {4{neg221[14]}} , neg221[14:4] };

   // m221_34 = W*in
   wire signed [14:0] m221_34;
   assign m221_34 =15'b0;

   // m221_35 = W*in
   wire signed [14:0] m221_35;
   assign m221_35 =15'b0;

   // m221_36 = W*in
   wire signed [14:0] m221_36;
   assign m221_36 =15'b0;

   // m221_37 = W*in
   wire signed [14:0] m221_37;
   assign m221_37 =15'b0;

   // m221_38 = W*in
   wire signed [14:0] m221_38;
   assign m221_38 =15'b0;

   // m221_39 = W*in
   wire signed [14:0] m221_39;
   assign m221_39 =15'b0;

   // m221_40 = W*in
   wire signed [14:0] m221_40;
   assign m221_40 ={ {4{neg221[14]}} , neg221[14:4] };

   // m221_41 = W*in
   wire signed [14:0] m221_41;
   assign m221_41 =15'b0;

   // m221_42 = W*in
   wire signed [14:0] m221_42;
   assign m221_42 =15'b0;

   // m221_43 = W*in
   wire signed [14:0] m221_43;
   assign m221_43 =15'b0;

   // m221_44 = W*in
   wire signed [14:0] m221_44;
   assign m221_44 =15'b0;

   // m221_45 = W*in
   wire signed [14:0] m221_45;
   assign m221_45 =15'b0;

   // m221_46 = W*in
   wire signed [14:0] m221_46;
   assign m221_46 =15'b0;

   // m221_47 = W*in
   wire signed [14:0] m221_47;
   assign m221_47 =15'b0;

   // m221_48 = W*in
   wire signed [14:0] m221_48;
   assign m221_48 =15'b0;

   // m221_49 = W*in
   wire signed [14:0] m221_49;
   assign m221_49 =15'b0;

   // m221_50 = W*in
   wire signed [14:0] m221_50;
   assign m221_50 =15'b0;

   // m221_51 = W*in
   wire signed [14:0] m221_51;
   assign m221_51 =15'b0;

   // m221_52 = W*in
   wire signed [14:0] m221_52;
   assign m221_52 =15'b0;

   // m221_53 = W*in
   wire signed [14:0] m221_53;
   assign m221_53 =15'b0;

   // m221_54 = W*in
   wire signed [14:0] m221_54;
   assign m221_54 =15'b0;

   // m221_55 = W*in
   wire signed [14:0] m221_55;
   assign m221_55 =15'b0;

   // m221_56 = W*in
   wire signed [14:0] m221_56;
   assign m221_56 =15'b0;

   // m221_57 = W*in
   wire signed [14:0] m221_57;
   assign m221_57 =15'b0;

   // m221_58 = W*in
   wire signed [14:0] m221_58;
   assign m221_58 ={ {4{in221[14]}} , in221[14:4] };

   // m221_59 = W*in
   wire signed [14:0] m221_59;
   assign m221_59 ={ {4{in221[14]}} , in221[14:4] };

   // m221_60 = W*in
   wire signed [14:0] m221_60;
   assign m221_60 =15'b0;

   // m221_61 = W*in
   wire signed [14:0] m221_61;
   assign m221_61 ={ {4{in221[14]}} , in221[14:4] };

   // m221_62 = W*in
   wire signed [14:0] m221_62;
   assign m221_62 =15'b0;

   // m221_63 = W*in
   wire signed [14:0] m221_63;
   assign m221_63 =15'b0;

   // m221_64 = W*in
   wire signed [14:0] m221_64;
   assign m221_64 ={ {4{in221[14]}} , in221[14:4] };

   // m221_65 = W*in
   wire signed [14:0] m221_65;
   assign m221_65 =15'b0;

   // m221_66 = W*in
   wire signed [14:0] m221_66;
   assign m221_66 =15'b0;

   // m221_67 = W*in
   wire signed [14:0] m221_67;
   assign m221_67 =15'b0;

   // m221_68 = W*in
   wire signed [14:0] m221_68;
   assign m221_68 =15'b0;

   // m221_69 = W*in
   wire signed [14:0] m221_69;
   assign m221_69 =15'b0;

   // m221_70 = W*in
   wire signed [14:0] m221_70;
   assign m221_70 =15'b0;

   // m221_71 = W*in
   wire signed [14:0] m221_71;
   assign m221_71 =15'b0;

   // m221_72 = W*in
   wire signed [14:0] m221_72;
   assign m221_72 =15'b0;

   // m221_73 = W*in
   wire signed [14:0] m221_73;
   assign m221_73 =15'b0;

   // m221_74 = W*in
   wire signed [14:0] m221_74;
   assign m221_74 =15'b0;

   // m221_75 = W*in
   wire signed [14:0] m221_75;
   assign m221_75 =15'b0;

   // m221_76 = W*in
   wire signed [14:0] m221_76;
   assign m221_76 ={ {4{neg221[14]}} , neg221[14:4] };

   // m221_77 = W*in
   wire signed [14:0] m221_77;
   assign m221_77 =15'b0;

   // m221_78 = W*in
   wire signed [14:0] m221_78;
   assign m221_78 =15'b0;

   // m221_79 = W*in
   wire signed [14:0] m221_79;
   assign m221_79 =15'b0;

   // m221_80 = W*in
   wire signed [14:0] m221_80;
   assign m221_80 =15'b0;

   // m221_81 = W*in
   wire signed [14:0] m221_81;
   assign m221_81 =15'b0;

   // m221_82 = W*in
   wire signed [14:0] m221_82;
   assign m221_82 =15'b0;

   // m221_83 = W*in
   wire signed [14:0] m221_83;
   assign m221_83 =15'b0;

   // m221_84 = W*in
   wire signed [14:0] m221_84;
   assign m221_84 =15'b0;

   // m221_85 = W*in
   wire signed [14:0] m221_85;
   assign m221_85 =15'b0;

   // m221_86 = W*in
   wire signed [14:0] m221_86;
   assign m221_86 =15'b0;

   // m221_87 = W*in
   wire signed [14:0] m221_87;
   assign m221_87 =15'b0;

   // m221_88 = W*in
   wire signed [14:0] m221_88;
   assign m221_88 =15'b0;

   // m221_89 = W*in
   wire signed [14:0] m221_89;
   assign m221_89 =15'b0;

   // m221_90 = W*in
   wire signed [14:0] m221_90;
   assign m221_90 =15'b0;

   // m221_91 = W*in
   wire signed [14:0] m221_91;
   assign m221_91 =15'b0;

   // m221_92 = W*in
   wire signed [14:0] m221_92;
   assign m221_92 =15'b0;

   // m221_93 = W*in
   wire signed [14:0] m221_93;
   assign m221_93 =15'b0;

   // m221_94 = W*in
   wire signed [14:0] m221_94;
   assign m221_94 =15'b0;

   // m221_95 = W*in
   wire signed [14:0] m221_95;
   assign m221_95 =15'b0;

   // m221_96 = W*in
   wire signed [14:0] m221_96;
   assign m221_96 =15'b0;

   // m221_97 = W*in
   wire signed [14:0] m221_97;
   assign m221_97 =15'b0;

   // m221_98 = W*in
   wire signed [14:0] m221_98;
   assign m221_98 =15'b0;

   // m221_99 = W*in
   wire signed [14:0] m221_99;
   assign m221_99 =15'b0;

   // m221_100 = W*in
   wire signed [14:0] m221_100;
   assign m221_100 =15'b0;

   // m222_1 = W*in
   wire signed [14:0] m222_1;
   assign m222_1 =15'b0;

   // m222_2 = W*in
   wire signed [14:0] m222_2;
   assign m222_2 =15'b0;

   // m222_3 = W*in
   wire signed [14:0] m222_3;
   assign m222_3 ={ {3{in222[14]}} , in222[14:3] };

   // m222_4 = W*in
   wire signed [14:0] m222_4;
   assign m222_4 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_5 = W*in
   wire signed [14:0] m222_5;
   assign m222_5 =15'b0;

   // m222_6 = W*in
   wire signed [14:0] m222_6;
   assign m222_6 ={ {3{in222[14]}} , in222[14:3] };

   // m222_7 = W*in
   wire signed [14:0] m222_7;
   assign m222_7 =15'b0;

   // m222_8 = W*in
   wire signed [14:0] m222_8;
   assign m222_8 =15'b0;

   // m222_9 = W*in
   wire signed [14:0] m222_9;
   assign m222_9 =15'b0;

   // m222_10 = W*in
   wire signed [14:0] m222_10;
   assign m222_10 =15'b0;

   // m222_11 = W*in
   wire signed [14:0] m222_11;
   assign m222_11 =15'b0;

   // m222_12 = W*in
   wire signed [14:0] m222_12;
   assign m222_12 =15'b0;

   // m222_13 = W*in
   wire signed [14:0] m222_13;
   assign m222_13 =15'b0;

   // m222_14 = W*in
   wire signed [14:0] m222_14;
   assign m222_14 =15'b0;

   // m222_15 = W*in
   wire signed [14:0] m222_15;
   assign m222_15 ={ {3{in222[14]}} , in222[14:3] };

   // m222_16 = W*in
   wire signed [14:0] m222_16;
   assign m222_16 ={ {3{in222[14]}} , in222[14:3] };

   // m222_17 = W*in
   wire signed [14:0] m222_17;
   assign m222_17 =15'b0;

   // m222_18 = W*in
   wire signed [14:0] m222_18;
   assign m222_18 =15'b0;

   // m222_19 = W*in
   wire signed [14:0] m222_19;
   assign m222_19 =15'b0;

   // m222_20 = W*in
   wire signed [14:0] m222_20;
   assign m222_20 =15'b0;

   // m222_21 = W*in
   wire signed [14:0] m222_21;
   assign m222_21 =15'b0;

   // m222_22 = W*in
   wire signed [14:0] m222_22;
   assign m222_22 =15'b0;

   // m222_23 = W*in
   wire signed [14:0] m222_23;
   assign m222_23 =15'b0;

   // m222_24 = W*in
   wire signed [14:0] m222_24;
   assign m222_24 ={ {3{in222[14]}} , in222[14:3] };

   // m222_25 = W*in
   wire signed [14:0] m222_25;
   assign m222_25 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_26 = W*in
   wire signed [14:0] m222_26;
   assign m222_26 ={ {3{in222[14]}} , in222[14:3] };

   // m222_27 = W*in
   wire signed [14:0] m222_27;
   assign m222_27 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_28 = W*in
   wire signed [14:0] m222_28;
   assign m222_28 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_29 = W*in
   wire signed [14:0] m222_29;
   assign m222_29 ={ {3{in222[14]}} , in222[14:3] };

   // m222_30 = W*in
   wire signed [14:0] m222_30;
   assign m222_30 =15'b0;

   // m222_31 = W*in
   wire signed [14:0] m222_31;
   assign m222_31 =15'b0;

   // m222_32 = W*in
   wire signed [14:0] m222_32;
   assign m222_32 =15'b0;

   // m222_33 = W*in
   wire signed [14:0] m222_33;
   assign m222_33 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_34 = W*in
   wire signed [14:0] m222_34;
   assign m222_34 ={ {3{in222[14]}} , in222[14:3] };

   // m222_35 = W*in
   wire signed [14:0] m222_35;
   assign m222_35 =15'b0;

   // m222_36 = W*in
   wire signed [14:0] m222_36;
   assign m222_36 =15'b0;

   // m222_37 = W*in
   wire signed [14:0] m222_37;
   assign m222_37 =15'b0;

   // m222_38 = W*in
   wire signed [14:0] m222_38;
   assign m222_38 =15'b0;

   // m222_39 = W*in
   wire signed [14:0] m222_39;
   assign m222_39 =15'b0;

   // m222_40 = W*in
   wire signed [14:0] m222_40;
   assign m222_40 =15'b0;

   // m222_41 = W*in
   wire signed [14:0] m222_41;
   assign m222_41 =15'b0;

   // m222_42 = W*in
   wire signed [14:0] m222_42;
   assign m222_42 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_43 = W*in
   wire signed [14:0] m222_43;
   assign m222_43 =15'b0;

   // m222_44 = W*in
   wire signed [14:0] m222_44;
   assign m222_44 =15'b0;

   // m222_45 = W*in
   wire signed [14:0] m222_45;
   assign m222_45 =15'b0;

   // m222_46 = W*in
   wire signed [14:0] m222_46;
   assign m222_46 ={ {4{in222[14]}} , in222[14:4] };

   // m222_47 = W*in
   wire signed [14:0] m222_47;
   assign m222_47 ={ {4{in222[14]}} , in222[14:4] };

   // m222_48 = W*in
   wire signed [14:0] m222_48;
   assign m222_48 =15'b0;

   // m222_49 = W*in
   wire signed [14:0] m222_49;
   assign m222_49 ={ {3{in222[14]}} , in222[14:3] };

   // m222_50 = W*in
   wire signed [14:0] m222_50;
   assign m222_50 =15'b0;

   // m222_51 = W*in
   wire signed [14:0] m222_51;
   assign m222_51 =15'b0;

   // m222_52 = W*in
   wire signed [14:0] m222_52;
   assign m222_52 =15'b0;

   // m222_53 = W*in
   wire signed [14:0] m222_53;
   assign m222_53 =15'b0;

   // m222_54 = W*in
   wire signed [14:0] m222_54;
   assign m222_54 =15'b0;

   // m222_55 = W*in
   wire signed [14:0] m222_55;
   assign m222_55 =15'b0;

   // m222_56 = W*in
   wire signed [14:0] m222_56;
   assign m222_56 =15'b0;

   // m222_57 = W*in
   wire signed [14:0] m222_57;
   assign m222_57 =15'b0;

   // m222_58 = W*in
   wire signed [14:0] m222_58;
   assign m222_58 =15'b0;

   // m222_59 = W*in
   wire signed [14:0] m222_59;
   assign m222_59 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_60 = W*in
   wire signed [14:0] m222_60;
   assign m222_60 ={ {4{in222[14]}} , in222[14:4] };

   // m222_61 = W*in
   wire signed [14:0] m222_61;
   assign m222_61 =15'b0;

   // m222_62 = W*in
   wire signed [14:0] m222_62;
   assign m222_62 =15'b0;

   // m222_63 = W*in
   wire signed [14:0] m222_63;
   assign m222_63 =15'b0;

   // m222_64 = W*in
   wire signed [14:0] m222_64;
   assign m222_64 ={ {4{in222[14]}} , in222[14:4] };

   // m222_65 = W*in
   wire signed [14:0] m222_65;
   assign m222_65 =15'b0;

   // m222_66 = W*in
   wire signed [14:0] m222_66;
   assign m222_66 =15'b0;

   // m222_67 = W*in
   wire signed [14:0] m222_67;
   assign m222_67 ={ {3{in222[14]}} , in222[14:3] };

   // m222_68 = W*in
   wire signed [14:0] m222_68;
   assign m222_68 =15'b0;

   // m222_69 = W*in
   wire signed [14:0] m222_69;
   assign m222_69 ={ {4{neg222[14]}} , neg222[14:4] };

   // m222_70 = W*in
   wire signed [14:0] m222_70;
   assign m222_70 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_71 = W*in
   wire signed [14:0] m222_71;
   assign m222_71 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_72 = W*in
   wire signed [14:0] m222_72;
   assign m222_72 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_73 = W*in
   wire signed [14:0] m222_73;
   assign m222_73 =15'b0;

   // m222_74 = W*in
   wire signed [14:0] m222_74;
   assign m222_74 ={ {4{neg222[14]}} , neg222[14:4] };

   // m222_75 = W*in
   wire signed [14:0] m222_75;
   assign m222_75 =15'b0;

   // m222_76 = W*in
   wire signed [14:0] m222_76;
   assign m222_76 ={ {4{neg222[14]}} , neg222[14:4] };

   // m222_77 = W*in
   wire signed [14:0] m222_77;
   assign m222_77 =15'b0;

   // m222_78 = W*in
   wire signed [14:0] m222_78;
   assign m222_78 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_79 = W*in
   wire signed [14:0] m222_79;
   assign m222_79 =15'b0;

   // m222_80 = W*in
   wire signed [14:0] m222_80;
   assign m222_80 =15'b0;

   // m222_81 = W*in
   wire signed [14:0] m222_81;
   assign m222_81 ={ {4{in222[14]}} , in222[14:4] };

   // m222_82 = W*in
   wire signed [14:0] m222_82;
   assign m222_82 =15'b0;

   // m222_83 = W*in
   wire signed [14:0] m222_83;
   assign m222_83 =15'b0;

   // m222_84 = W*in
   wire signed [14:0] m222_84;
   assign m222_84 =15'b0;

   // m222_85 = W*in
   wire signed [14:0] m222_85;
   assign m222_85 =15'b0;

   // m222_86 = W*in
   wire signed [14:0] m222_86;
   assign m222_86 =15'b0;

   // m222_87 = W*in
   wire signed [14:0] m222_87;
   assign m222_87 =15'b0;

   // m222_88 = W*in
   wire signed [14:0] m222_88;
   assign m222_88 =15'b0;

   // m222_89 = W*in
   wire signed [14:0] m222_89;
   assign m222_89 =15'b0;

   // m222_90 = W*in
   wire signed [14:0] m222_90;
   assign m222_90 =15'b0;

   // m222_91 = W*in
   wire signed [14:0] m222_91;
   assign m222_91 ={ {3{in222[14]}} , in222[14:3] };

   // m222_92 = W*in
   wire signed [14:0] m222_92;
   assign m222_92 =15'b0;

   // m222_93 = W*in
   wire signed [14:0] m222_93;
   assign m222_93 =15'b0;

   // m222_94 = W*in
   wire signed [14:0] m222_94;
   assign m222_94 =15'b0;

   // m222_95 = W*in
   wire signed [14:0] m222_95;
   assign m222_95 =15'b0;

   // m222_96 = W*in
   wire signed [14:0] m222_96;
   assign m222_96 =15'b0;

   // m222_97 = W*in
   wire signed [14:0] m222_97;
   assign m222_97 =15'b0;

   // m222_98 = W*in
   wire signed [14:0] m222_98;
   assign m222_98 =15'b0;

   // m222_99 = W*in
   wire signed [14:0] m222_99;
   assign m222_99 ={ {3{neg222[14]}} , neg222[14:3] };

   // m222_100 = W*in
   wire signed [14:0] m222_100;
   assign m222_100 =15'b0;

   // m223_1 = W*in
   wire signed [14:0] m223_1;
   assign m223_1 ={ {3{neg223[14]}} , neg223[14:3] };

   // m223_2 = W*in
   wire signed [14:0] m223_2;
   assign m223_2 =15'b0;

   // m223_3 = W*in
   wire signed [14:0] m223_3;
   assign m223_3 =15'b0;

   // m223_4 = W*in
   wire signed [14:0] m223_4;
   assign m223_4 =15'b0;

   // m223_5 = W*in
   wire signed [14:0] m223_5;
   assign m223_5 =15'b0;

   // m223_6 = W*in
   wire signed [14:0] m223_6;
   assign m223_6 =15'b0;

   // m223_7 = W*in
   wire signed [14:0] m223_7;
   assign m223_7 =15'b0;

   // m223_8 = W*in
   wire signed [14:0] m223_8;
   assign m223_8 =15'b0;

   // m223_9 = W*in
   wire signed [14:0] m223_9;
   assign m223_9 =15'b0;

   // m223_10 = W*in
   wire signed [14:0] m223_10;
   assign m223_10 =15'b0;

   // m223_11 = W*in
   wire signed [14:0] m223_11;
   assign m223_11 =15'b0;

   // m223_12 = W*in
   wire signed [14:0] m223_12;
   assign m223_12 =15'b0;

   // m223_13 = W*in
   wire signed [14:0] m223_13;
   assign m223_13 =15'b0;

   // m223_14 = W*in
   wire signed [14:0] m223_14;
   assign m223_14 =15'b0;

   // m223_15 = W*in
   wire signed [14:0] m223_15;
   assign m223_15 =15'b0;

   // m223_16 = W*in
   wire signed [14:0] m223_16;
   assign m223_16 =15'b0;

   // m223_17 = W*in
   wire signed [14:0] m223_17;
   assign m223_17 =15'b0;

   // m223_18 = W*in
   wire signed [14:0] m223_18;
   assign m223_18 =15'b0;

   // m223_19 = W*in
   wire signed [14:0] m223_19;
   assign m223_19 =15'b0;

   // m223_20 = W*in
   wire signed [14:0] m223_20;
   assign m223_20 =15'b0;

   // m223_21 = W*in
   wire signed [14:0] m223_21;
   assign m223_21 =15'b0;

   // m223_22 = W*in
   wire signed [14:0] m223_22;
   assign m223_22 =15'b0;

   // m223_23 = W*in
   wire signed [14:0] m223_23;
   assign m223_23 =15'b0;

   // m223_24 = W*in
   wire signed [14:0] m223_24;
   assign m223_24 =15'b0;

   // m223_25 = W*in
   wire signed [14:0] m223_25;
   assign m223_25 =15'b0;

   // m223_26 = W*in
   wire signed [14:0] m223_26;
   assign m223_26 =15'b0;

   // m223_27 = W*in
   wire signed [14:0] m223_27;
   assign m223_27 =15'b0;

   // m223_28 = W*in
   wire signed [14:0] m223_28;
   assign m223_28 =15'b0;

   // m223_29 = W*in
   wire signed [14:0] m223_29;
   assign m223_29 =15'b0;

   // m223_30 = W*in
   wire signed [14:0] m223_30;
   assign m223_30 =15'b0;

   // m223_31 = W*in
   wire signed [14:0] m223_31;
   assign m223_31 =15'b0;

   // m223_32 = W*in
   wire signed [14:0] m223_32;
   assign m223_32 =15'b0;

   // m223_33 = W*in
   wire signed [14:0] m223_33;
   assign m223_33 =15'b0;

   // m223_34 = W*in
   wire signed [14:0] m223_34;
   assign m223_34 =15'b0;

   // m223_35 = W*in
   wire signed [14:0] m223_35;
   assign m223_35 =15'b0;

   // m223_36 = W*in
   wire signed [14:0] m223_36;
   assign m223_36 =15'b0;

   // m223_37 = W*in
   wire signed [14:0] m223_37;
   assign m223_37 =15'b0;

   // m223_38 = W*in
   wire signed [14:0] m223_38;
   assign m223_38 =15'b0;

   // m223_39 = W*in
   wire signed [14:0] m223_39;
   assign m223_39 =15'b0;

   // m223_40 = W*in
   wire signed [14:0] m223_40;
   assign m223_40 =15'b0;

   // m223_41 = W*in
   wire signed [14:0] m223_41;
   assign m223_41 =15'b0;

   // m223_42 = W*in
   wire signed [14:0] m223_42;
   assign m223_42 =15'b0;

   // m223_43 = W*in
   wire signed [14:0] m223_43;
   assign m223_43 =15'b0;

   // m223_44 = W*in
   wire signed [14:0] m223_44;
   assign m223_44 ={ {4{neg223[14]}} , neg223[14:4] };

   // m223_45 = W*in
   wire signed [14:0] m223_45;
   assign m223_45 ={ {4{in223[14]}} , in223[14:4] };

   // m223_46 = W*in
   wire signed [14:0] m223_46;
   assign m223_46 =15'b0;

   // m223_47 = W*in
   wire signed [14:0] m223_47;
   assign m223_47 =15'b0;

   // m223_48 = W*in
   wire signed [14:0] m223_48;
   assign m223_48 =15'b0;

   // m223_49 = W*in
   wire signed [14:0] m223_49;
   assign m223_49 =15'b0;

   // m223_50 = W*in
   wire signed [14:0] m223_50;
   assign m223_50 =15'b0;

   // m223_51 = W*in
   wire signed [14:0] m223_51;
   assign m223_51 =15'b0;

   // m223_52 = W*in
   wire signed [14:0] m223_52;
   assign m223_52 =15'b0;

   // m223_53 = W*in
   wire signed [14:0] m223_53;
   assign m223_53 =15'b0;

   // m223_54 = W*in
   wire signed [14:0] m223_54;
   assign m223_54 =15'b0;

   // m223_55 = W*in
   wire signed [14:0] m223_55;
   assign m223_55 =15'b0;

   // m223_56 = W*in
   wire signed [14:0] m223_56;
   assign m223_56 =15'b0;

   // m223_57 = W*in
   wire signed [14:0] m223_57;
   assign m223_57 =15'b0;

   // m223_58 = W*in
   wire signed [14:0] m223_58;
   assign m223_58 ={ {2{neg223[14]}} , neg223[14:2] };

   // m223_59 = W*in
   wire signed [14:0] m223_59;
   assign m223_59 =15'b0;

   // m223_60 = W*in
   wire signed [14:0] m223_60;
   assign m223_60 =15'b0;

   // m223_61 = W*in
   wire signed [14:0] m223_61;
   assign m223_61 ={ {3{in223[14]}} , in223[14:3] };

   // m223_62 = W*in
   wire signed [14:0] m223_62;
   assign m223_62 =15'b0;

   // m223_63 = W*in
   wire signed [14:0] m223_63;
   assign m223_63 =15'b0;

   // m223_64 = W*in
   wire signed [14:0] m223_64;
   assign m223_64 ={ {4{in223[14]}} , in223[14:4] };

   // m223_65 = W*in
   wire signed [14:0] m223_65;
   assign m223_65 =15'b0;

   // m223_66 = W*in
   wire signed [14:0] m223_66;
   assign m223_66 =15'b0;

   // m223_67 = W*in
   wire signed [14:0] m223_67;
   assign m223_67 =15'b0;

   // m223_68 = W*in
   wire signed [14:0] m223_68;
   assign m223_68 =15'b0;

   // m223_69 = W*in
   wire signed [14:0] m223_69;
   assign m223_69 =15'b0;

   // m223_70 = W*in
   wire signed [14:0] m223_70;
   assign m223_70 =15'b0;

   // m223_71 = W*in
   wire signed [14:0] m223_71;
   assign m223_71 =15'b0;

   // m223_72 = W*in
   wire signed [14:0] m223_72;
   assign m223_72 =15'b0;

   // m223_73 = W*in
   wire signed [14:0] m223_73;
   assign m223_73 =15'b0;

   // m223_74 = W*in
   wire signed [14:0] m223_74;
   assign m223_74 =15'b0;

   // m223_75 = W*in
   wire signed [14:0] m223_75;
   assign m223_75 =15'b0;

   // m223_76 = W*in
   wire signed [14:0] m223_76;
   assign m223_76 ={ {4{neg223[14]}} , neg223[14:4] };

   // m223_77 = W*in
   wire signed [14:0] m223_77;
   assign m223_77 =15'b0;

   // m223_78 = W*in
   wire signed [14:0] m223_78;
   assign m223_78 =15'b0;

   // m223_79 = W*in
   wire signed [14:0] m223_79;
   assign m223_79 =15'b0;

   // m223_80 = W*in
   wire signed [14:0] m223_80;
   assign m223_80 =15'b0;

   // m223_81 = W*in
   wire signed [14:0] m223_81;
   assign m223_81 =15'b0;

   // m223_82 = W*in
   wire signed [14:0] m223_82;
   assign m223_82 =15'b0;

   // m223_83 = W*in
   wire signed [14:0] m223_83;
   assign m223_83 =15'b0;

   // m223_84 = W*in
   wire signed [14:0] m223_84;
   assign m223_84 =15'b0;

   // m223_85 = W*in
   wire signed [14:0] m223_85;
   assign m223_85 ={ {3{in223[14]}} , in223[14:3] };

   // m223_86 = W*in
   wire signed [14:0] m223_86;
   assign m223_86 =15'b0;

   // m223_87 = W*in
   wire signed [14:0] m223_87;
   assign m223_87 ={ {2{in223[14]}} , in223[14:2] };

   // m223_88 = W*in
   wire signed [14:0] m223_88;
   assign m223_88 ={ {3{neg223[14]}} , neg223[14:3] };

   // m223_89 = W*in
   wire signed [14:0] m223_89;
   assign m223_89 =15'b0;

   // m223_90 = W*in
   wire signed [14:0] m223_90;
   assign m223_90 =15'b0;

   // m223_91 = W*in
   wire signed [14:0] m223_91;
   assign m223_91 =15'b0;

   // m223_92 = W*in
   wire signed [14:0] m223_92;
   assign m223_92 ={ {4{neg223[14]}} , neg223[14:4] };

   // m223_93 = W*in
   wire signed [14:0] m223_93;
   assign m223_93 =15'b0;

   // m223_94 = W*in
   wire signed [14:0] m223_94;
   assign m223_94 =15'b0;

   // m223_95 = W*in
   wire signed [14:0] m223_95;
   assign m223_95 =15'b0;

   // m223_96 = W*in
   wire signed [14:0] m223_96;
   assign m223_96 =15'b0;

   // m223_97 = W*in
   wire signed [14:0] m223_97;
   assign m223_97 =15'b0;

   // m223_98 = W*in
   wire signed [14:0] m223_98;
   assign m223_98 =15'b0;

   // m223_99 = W*in
   wire signed [14:0] m223_99;
   assign m223_99 =15'b0;

   // m223_100 = W*in
   wire signed [14:0] m223_100;
   assign m223_100 =15'b0;

   // m224_1 = W*in
   wire signed [14:0] m224_1;
   assign m224_1 =15'b0;

   // m224_2 = W*in
   wire signed [14:0] m224_2;
   assign m224_2 =15'b0;

   // m224_3 = W*in
   wire signed [14:0] m224_3;
   assign m224_3 =15'b0;

   // m224_4 = W*in
   wire signed [14:0] m224_4;
   assign m224_4 =15'b0;

   // m224_5 = W*in
   wire signed [14:0] m224_5;
   assign m224_5 =15'b0;

   // m224_6 = W*in
   wire signed [14:0] m224_6;
   assign m224_6 =15'b0;

   // m224_7 = W*in
   wire signed [14:0] m224_7;
   assign m224_7 =15'b0;

   // m224_8 = W*in
   wire signed [14:0] m224_8;
   assign m224_8 =15'b0;

   // m224_9 = W*in
   wire signed [14:0] m224_9;
   assign m224_9 =15'b0;

   // m224_10 = W*in
   wire signed [14:0] m224_10;
   assign m224_10 =15'b0;

   // m224_11 = W*in
   wire signed [14:0] m224_11;
   assign m224_11 =15'b0;

   // m224_12 = W*in
   wire signed [14:0] m224_12;
   assign m224_12 =15'b0;

   // m224_13 = W*in
   wire signed [14:0] m224_13;
   assign m224_13 =15'b0;

   // m224_14 = W*in
   wire signed [14:0] m224_14;
   assign m224_14 =15'b0;

   // m224_15 = W*in
   wire signed [14:0] m224_15;
   assign m224_15 =15'b0;

   // m224_16 = W*in
   wire signed [14:0] m224_16;
   assign m224_16 =15'b0;

   // m224_17 = W*in
   wire signed [14:0] m224_17;
   assign m224_17 =15'b0;

   // m224_18 = W*in
   wire signed [14:0] m224_18;
   assign m224_18 =15'b0;

   // m224_19 = W*in
   wire signed [14:0] m224_19;
   assign m224_19 =15'b0;

   // m224_20 = W*in
   wire signed [14:0] m224_20;
   assign m224_20 =15'b0;

   // m224_21 = W*in
   wire signed [14:0] m224_21;
   assign m224_21 =15'b0;

   // m224_22 = W*in
   wire signed [14:0] m224_22;
   assign m224_22 =15'b0;

   // m224_23 = W*in
   wire signed [14:0] m224_23;
   assign m224_23 =15'b0;

   // m224_24 = W*in
   wire signed [14:0] m224_24;
   assign m224_24 =15'b0;

   // m224_25 = W*in
   wire signed [14:0] m224_25;
   assign m224_25 =15'b0;

   // m224_26 = W*in
   wire signed [14:0] m224_26;
   assign m224_26 =15'b0;

   // m224_27 = W*in
   wire signed [14:0] m224_27;
   assign m224_27 ={ {3{in224[14]}} , in224[14:3] };

   // m224_28 = W*in
   wire signed [14:0] m224_28;
   assign m224_28 =15'b0;

   // m224_29 = W*in
   wire signed [14:0] m224_29;
   assign m224_29 =15'b0;

   // m224_30 = W*in
   wire signed [14:0] m224_30;
   assign m224_30 =15'b0;

   // m224_31 = W*in
   wire signed [14:0] m224_31;
   assign m224_31 =15'b0;

   // m224_32 = W*in
   wire signed [14:0] m224_32;
   assign m224_32 =15'b0;

   // m224_33 = W*in
   wire signed [14:0] m224_33;
   assign m224_33 =15'b0;

   // m224_34 = W*in
   wire signed [14:0] m224_34;
   assign m224_34 =15'b0;

   // m224_35 = W*in
   wire signed [14:0] m224_35;
   assign m224_35 ={ {3{in224[14]}} , in224[14:3] };

   // m224_36 = W*in
   wire signed [14:0] m224_36;
   assign m224_36 =15'b0;

   // m224_37 = W*in
   wire signed [14:0] m224_37;
   assign m224_37 =15'b0;

   // m224_38 = W*in
   wire signed [14:0] m224_38;
   assign m224_38 =15'b0;

   // m224_39 = W*in
   wire signed [14:0] m224_39;
   assign m224_39 =15'b0;

   // m224_40 = W*in
   wire signed [14:0] m224_40;
   assign m224_40 ={ {3{in224[14]}} , in224[14:3] };

   // m224_41 = W*in
   wire signed [14:0] m224_41;
   assign m224_41 =15'b0;

   // m224_42 = W*in
   wire signed [14:0] m224_42;
   assign m224_42 =15'b0;

   // m224_43 = W*in
   wire signed [14:0] m224_43;
   assign m224_43 =15'b0;

   // m224_44 = W*in
   wire signed [14:0] m224_44;
   assign m224_44 =15'b0;

   // m224_45 = W*in
   wire signed [14:0] m224_45;
   assign m224_45 =15'b0;

   // m224_46 = W*in
   wire signed [14:0] m224_46;
   assign m224_46 =15'b0;

   // m224_47 = W*in
   wire signed [14:0] m224_47;
   assign m224_47 =15'b0;

   // m224_48 = W*in
   wire signed [14:0] m224_48;
   assign m224_48 =15'b0;

   // m224_49 = W*in
   wire signed [14:0] m224_49;
   assign m224_49 =15'b0;

   // m224_50 = W*in
   wire signed [14:0] m224_50;
   assign m224_50 =15'b0;

   // m224_51 = W*in
   wire signed [14:0] m224_51;
   assign m224_51 =15'b0;

   // m224_52 = W*in
   wire signed [14:0] m224_52;
   assign m224_52 =15'b0;

   // m224_53 = W*in
   wire signed [14:0] m224_53;
   assign m224_53 =15'b0;

   // m224_54 = W*in
   wire signed [14:0] m224_54;
   assign m224_54 =15'b0;

   // m224_55 = W*in
   wire signed [14:0] m224_55;
   assign m224_55 =15'b0;

   // m224_56 = W*in
   wire signed [14:0] m224_56;
   assign m224_56 =15'b0;

   // m224_57 = W*in
   wire signed [14:0] m224_57;
   assign m224_57 =15'b0;

   // m224_58 = W*in
   wire signed [14:0] m224_58;
   assign m224_58 ={ {3{neg224[14]}} , neg224[14:3] };

   // m224_59 = W*in
   wire signed [14:0] m224_59;
   assign m224_59 =15'b0;

   // m224_60 = W*in
   wire signed [14:0] m224_60;
   assign m224_60 =15'b0;

   // m224_61 = W*in
   wire signed [14:0] m224_61;
   assign m224_61 =15'b0;

   // m224_62 = W*in
   wire signed [14:0] m224_62;
   assign m224_62 =15'b0;

   // m224_63 = W*in
   wire signed [14:0] m224_63;
   assign m224_63 =15'b0;

   // m224_64 = W*in
   wire signed [14:0] m224_64;
   assign m224_64 =15'b0;

   // m224_65 = W*in
   wire signed [14:0] m224_65;
   assign m224_65 ={ {4{neg224[14]}} , neg224[14:4] };

   // m224_66 = W*in
   wire signed [14:0] m224_66;
   assign m224_66 =15'b0;

   // m224_67 = W*in
   wire signed [14:0] m224_67;
   assign m224_67 =15'b0;

   // m224_68 = W*in
   wire signed [14:0] m224_68;
   assign m224_68 =15'b0;

   // m224_69 = W*in
   wire signed [14:0] m224_69;
   assign m224_69 ={ {4{neg224[14]}} , neg224[14:4] };

   // m224_70 = W*in
   wire signed [14:0] m224_70;
   assign m224_70 =15'b0;

   // m224_71 = W*in
   wire signed [14:0] m224_71;
   assign m224_71 =15'b0;

   // m224_72 = W*in
   wire signed [14:0] m224_72;
   assign m224_72 =15'b0;

   // m224_73 = W*in
   wire signed [14:0] m224_73;
   assign m224_73 =15'b0;

   // m224_74 = W*in
   wire signed [14:0] m224_74;
   assign m224_74 =15'b0;

   // m224_75 = W*in
   wire signed [14:0] m224_75;
   assign m224_75 =15'b0;

   // m224_76 = W*in
   wire signed [14:0] m224_76;
   assign m224_76 =15'b0;

   // m224_77 = W*in
   wire signed [14:0] m224_77;
   assign m224_77 =15'b0;

   // m224_78 = W*in
   wire signed [14:0] m224_78;
   assign m224_78 =15'b0;

   // m224_79 = W*in
   wire signed [14:0] m224_79;
   assign m224_79 =15'b0;

   // m224_80 = W*in
   wire signed [14:0] m224_80;
   assign m224_80 =15'b0;

   // m224_81 = W*in
   wire signed [14:0] m224_81;
   assign m224_81 ={ {4{neg224[14]}} , neg224[14:4] };

   // m224_82 = W*in
   wire signed [14:0] m224_82;
   assign m224_82 =15'b0;

   // m224_83 = W*in
   wire signed [14:0] m224_83;
   assign m224_83 =15'b0;

   // m224_84 = W*in
   wire signed [14:0] m224_84;
   assign m224_84 =15'b0;

   // m224_85 = W*in
   wire signed [14:0] m224_85;
   assign m224_85 =15'b0;

   // m224_86 = W*in
   wire signed [14:0] m224_86;
   assign m224_86 =15'b0;

   // m224_87 = W*in
   wire signed [14:0] m224_87;
   assign m224_87 =15'b0;

   // m224_88 = W*in
   wire signed [14:0] m224_88;
   assign m224_88 =15'b0;

   // m224_89 = W*in
   wire signed [14:0] m224_89;
   assign m224_89 =15'b0;

   // m224_90 = W*in
   wire signed [14:0] m224_90;
   assign m224_90 =15'b0;

   // m224_91 = W*in
   wire signed [14:0] m224_91;
   assign m224_91 =15'b0;

   // m224_92 = W*in
   wire signed [14:0] m224_92;
   assign m224_92 =15'b0;

   // m224_93 = W*in
   wire signed [14:0] m224_93;
   assign m224_93 =15'b0;

   // m224_94 = W*in
   wire signed [14:0] m224_94;
   assign m224_94 ={ {3{in224[14]}} , in224[14:3] };

   // m224_95 = W*in
   wire signed [14:0] m224_95;
   assign m224_95 =15'b0;

   // m224_96 = W*in
   wire signed [14:0] m224_96;
   assign m224_96 =15'b0;

   // m224_97 = W*in
   wire signed [14:0] m224_97;
   assign m224_97 =15'b0;

   // m224_98 = W*in
   wire signed [14:0] m224_98;
   assign m224_98 =15'b0;

   // m224_99 = W*in
   wire signed [14:0] m224_99;
   assign m224_99 ={ {3{neg224[14]}} , neg224[14:3] };

   // m224_100 = W*in
   wire signed [14:0] m224_100;
   assign m224_100 =15'b0;

   // m225_1 = W*in
   wire signed [14:0] m225_1;
   assign m225_1 =15'b0;

   // m225_2 = W*in
   wire signed [14:0] m225_2;
   assign m225_2 =15'b0;

   // m225_3 = W*in
   wire signed [14:0] m225_3;
   assign m225_3 =15'b0;

   // m225_4 = W*in
   wire signed [14:0] m225_4;
   assign m225_4 =15'b0;

   // m225_5 = W*in
   wire signed [14:0] m225_5;
   assign m225_5 =15'b0;

   // m225_6 = W*in
   wire signed [14:0] m225_6;
   assign m225_6 =15'b0;

   // m225_7 = W*in
   wire signed [14:0] m225_7;
   assign m225_7 ={ {3{neg225[14]}} , neg225[14:3] };

   // m225_8 = W*in
   wire signed [14:0] m225_8;
   assign m225_8 =15'b0;

   // m225_9 = W*in
   wire signed [14:0] m225_9;
   assign m225_9 =15'b0;

   // m225_10 = W*in
   wire signed [14:0] m225_10;
   assign m225_10 =15'b0;

   // m225_11 = W*in
   wire signed [14:0] m225_11;
   assign m225_11 =15'b0;

   // m225_12 = W*in
   wire signed [14:0] m225_12;
   assign m225_12 =15'b0;

   // m225_13 = W*in
   wire signed [14:0] m225_13;
   assign m225_13 =15'b0;

   // m225_14 = W*in
   wire signed [14:0] m225_14;
   assign m225_14 =15'b0;

   // m225_15 = W*in
   wire signed [14:0] m225_15;
   assign m225_15 =15'b0;

   // m225_16 = W*in
   wire signed [14:0] m225_16;
   assign m225_16 =15'b0;

   // m225_17 = W*in
   wire signed [14:0] m225_17;
   assign m225_17 =15'b0;

   // m225_18 = W*in
   wire signed [14:0] m225_18;
   assign m225_18 =15'b0;

   // m225_19 = W*in
   wire signed [14:0] m225_19;
   assign m225_19 =15'b0;

   // m225_20 = W*in
   wire signed [14:0] m225_20;
   assign m225_20 =15'b0;

   // m225_21 = W*in
   wire signed [14:0] m225_21;
   assign m225_21 =15'b0;

   // m225_22 = W*in
   wire signed [14:0] m225_22;
   assign m225_22 =15'b0;

   // m225_23 = W*in
   wire signed [14:0] m225_23;
   assign m225_23 =15'b0;

   // m225_24 = W*in
   wire signed [14:0] m225_24;
   assign m225_24 =15'b0;

   // m225_25 = W*in
   wire signed [14:0] m225_25;
   assign m225_25 =15'b0;

   // m225_26 = W*in
   wire signed [14:0] m225_26;
   assign m225_26 =15'b0;

   // m225_27 = W*in
   wire signed [14:0] m225_27;
   assign m225_27 ={ {4{in225[14]}} , in225[14:4] };

   // m225_28 = W*in
   wire signed [14:0] m225_28;
   assign m225_28 =15'b0;

   // m225_29 = W*in
   wire signed [14:0] m225_29;
   assign m225_29 ={ {4{neg225[14]}} , neg225[14:4] };

   // m225_30 = W*in
   wire signed [14:0] m225_30;
   assign m225_30 =15'b0;

   // m225_31 = W*in
   wire signed [14:0] m225_31;
   assign m225_31 =15'b0;

   // m225_32 = W*in
   wire signed [14:0] m225_32;
   assign m225_32 ={ {4{neg225[14]}} , neg225[14:4] };

   // m225_33 = W*in
   wire signed [14:0] m225_33;
   assign m225_33 ={ {4{neg225[14]}} , neg225[14:4] };

   // m225_34 = W*in
   wire signed [14:0] m225_34;
   assign m225_34 =15'b0;

   // m225_35 = W*in
   wire signed [14:0] m225_35;
   assign m225_35 =15'b0;

   // m225_36 = W*in
   wire signed [14:0] m225_36;
   assign m225_36 =15'b0;

   // m225_37 = W*in
   wire signed [14:0] m225_37;
   assign m225_37 =15'b0;

   // m225_38 = W*in
   wire signed [14:0] m225_38;
   assign m225_38 =15'b0;

   // m225_39 = W*in
   wire signed [14:0] m225_39;
   assign m225_39 =15'b0;

   // m225_40 = W*in
   wire signed [14:0] m225_40;
   assign m225_40 =15'b0;

   // m225_41 = W*in
   wire signed [14:0] m225_41;
   assign m225_41 =15'b0;

   // m225_42 = W*in
   wire signed [14:0] m225_42;
   assign m225_42 =15'b0;

   // m225_43 = W*in
   wire signed [14:0] m225_43;
   assign m225_43 =15'b0;

   // m225_44 = W*in
   wire signed [14:0] m225_44;
   assign m225_44 =15'b0;

   // m225_45 = W*in
   wire signed [14:0] m225_45;
   assign m225_45 =15'b0;

   // m225_46 = W*in
   wire signed [14:0] m225_46;
   assign m225_46 =15'b0;

   // m225_47 = W*in
   wire signed [14:0] m225_47;
   assign m225_47 =15'b0;

   // m225_48 = W*in
   wire signed [14:0] m225_48;
   assign m225_48 =15'b0;

   // m225_49 = W*in
   wire signed [14:0] m225_49;
   assign m225_49 =15'b0;

   // m225_50 = W*in
   wire signed [14:0] m225_50;
   assign m225_50 =15'b0;

   // m225_51 = W*in
   wire signed [14:0] m225_51;
   assign m225_51 =15'b0;

   // m225_52 = W*in
   wire signed [14:0] m225_52;
   assign m225_52 =15'b0;

   // m225_53 = W*in
   wire signed [14:0] m225_53;
   assign m225_53 =15'b0;

   // m225_54 = W*in
   wire signed [14:0] m225_54;
   assign m225_54 =15'b0;

   // m225_55 = W*in
   wire signed [14:0] m225_55;
   assign m225_55 =15'b0;

   // m225_56 = W*in
   wire signed [14:0] m225_56;
   assign m225_56 =15'b0;

   // m225_57 = W*in
   wire signed [14:0] m225_57;
   assign m225_57 ={ {4{in225[14]}} , in225[14:4] };

   // m225_58 = W*in
   wire signed [14:0] m225_58;
   assign m225_58 ={ {4{in225[14]}} , in225[14:4] };

   // m225_59 = W*in
   wire signed [14:0] m225_59;
   assign m225_59 =15'b0;

   // m225_60 = W*in
   wire signed [14:0] m225_60;
   assign m225_60 =15'b0;

   // m225_61 = W*in
   wire signed [14:0] m225_61;
   assign m225_61 =15'b0;

   // m225_62 = W*in
   wire signed [14:0] m225_62;
   assign m225_62 ={ {3{in225[14]}} , in225[14:3] };

   // m225_63 = W*in
   wire signed [14:0] m225_63;
   assign m225_63 =15'b0;

   // m225_64 = W*in
   wire signed [14:0] m225_64;
   assign m225_64 ={ {3{in225[14]}} , in225[14:3] };

   // m225_65 = W*in
   wire signed [14:0] m225_65;
   assign m225_65 =15'b0;

   // m225_66 = W*in
   wire signed [14:0] m225_66;
   assign m225_66 ={ {4{neg225[14]}} , neg225[14:4] };

   // m225_67 = W*in
   wire signed [14:0] m225_67;
   assign m225_67 ={ {4{neg225[14]}} , neg225[14:4] };

   // m225_68 = W*in
   wire signed [14:0] m225_68;
   assign m225_68 =15'b0;

   // m225_69 = W*in
   wire signed [14:0] m225_69;
   assign m225_69 =15'b0;

   // m225_70 = W*in
   wire signed [14:0] m225_70;
   assign m225_70 =15'b0;

   // m225_71 = W*in
   wire signed [14:0] m225_71;
   assign m225_71 =15'b0;

   // m225_72 = W*in
   wire signed [14:0] m225_72;
   assign m225_72 =15'b0;

   // m225_73 = W*in
   wire signed [14:0] m225_73;
   assign m225_73 =15'b0;

   // m225_74 = W*in
   wire signed [14:0] m225_74;
   assign m225_74 =15'b0;

   // m225_75 = W*in
   wire signed [14:0] m225_75;
   assign m225_75 =15'b0;

   // m225_76 = W*in
   wire signed [14:0] m225_76;
   assign m225_76 =15'b0;

   // m225_77 = W*in
   wire signed [14:0] m225_77;
   assign m225_77 =15'b0;

   // m225_78 = W*in
   wire signed [14:0] m225_78;
   assign m225_78 =15'b0;

   // m225_79 = W*in
   wire signed [14:0] m225_79;
   assign m225_79 =15'b0;

   // m225_80 = W*in
   wire signed [14:0] m225_80;
   assign m225_80 =15'b0;

   // m225_81 = W*in
   wire signed [14:0] m225_81;
   assign m225_81 =15'b0;

   // m225_82 = W*in
   wire signed [14:0] m225_82;
   assign m225_82 =15'b0;

   // m225_83 = W*in
   wire signed [14:0] m225_83;
   assign m225_83 =15'b0;

   // m225_84 = W*in
   wire signed [14:0] m225_84;
   assign m225_84 =15'b0;

   // m225_85 = W*in
   wire signed [14:0] m225_85;
   assign m225_85 ={ {3{in225[14]}} , in225[14:3] };

   // m225_86 = W*in
   wire signed [14:0] m225_86;
   assign m225_86 =15'b0;

   // m225_87 = W*in
   wire signed [14:0] m225_87;
   assign m225_87 ={ {3{in225[14]}} , in225[14:3] };

   // m225_88 = W*in
   wire signed [14:0] m225_88;
   assign m225_88 =15'b0;

   // m225_89 = W*in
   wire signed [14:0] m225_89;
   assign m225_89 =15'b0;

   // m225_90 = W*in
   wire signed [14:0] m225_90;
   assign m225_90 =15'b0;

   // m225_91 = W*in
   wire signed [14:0] m225_91;
   assign m225_91 =15'b0;

   // m225_92 = W*in
   wire signed [14:0] m225_92;
   assign m225_92 =15'b0;

   // m225_93 = W*in
   wire signed [14:0] m225_93;
   assign m225_93 =15'b0;

   // m225_94 = W*in
   wire signed [14:0] m225_94;
   assign m225_94 =15'b0;

   // m225_95 = W*in
   wire signed [14:0] m225_95;
   assign m225_95 =15'b0;

   // m225_96 = W*in
   wire signed [14:0] m225_96;
   assign m225_96 =15'b0;

   // m225_97 = W*in
   wire signed [14:0] m225_97;
   assign m225_97 ={ {3{in225[14]}} , in225[14:3] };

   // m225_98 = W*in
   wire signed [14:0] m225_98;
   assign m225_98 =15'b0;

   // m225_99 = W*in
   wire signed [14:0] m225_99;
   assign m225_99 =15'b0;

   // m225_100 = W*in
   wire signed [14:0] m225_100;
   assign m225_100 =15'b0;

   // m226_1 = W*in
   wire signed [14:0] m226_1;
   assign m226_1 =15'b0;

   // m226_2 = W*in
   wire signed [14:0] m226_2;
   assign m226_2 ={ {3{in226[14]}} , in226[14:3] };

   // m226_3 = W*in
   wire signed [14:0] m226_3;
   assign m226_3 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_4 = W*in
   wire signed [14:0] m226_4;
   assign m226_4 =15'b0;

   // m226_5 = W*in
   wire signed [14:0] m226_5;
   assign m226_5 =15'b0;

   // m226_6 = W*in
   wire signed [14:0] m226_6;
   assign m226_6 =15'b0;

   // m226_7 = W*in
   wire signed [14:0] m226_7;
   assign m226_7 =15'b0;

   // m226_8 = W*in
   wire signed [14:0] m226_8;
   assign m226_8 =15'b0;

   // m226_9 = W*in
   wire signed [14:0] m226_9;
   assign m226_9 ={ {3{in226[14]}} , in226[14:3] };

   // m226_10 = W*in
   wire signed [14:0] m226_10;
   assign m226_10 =15'b0;

   // m226_11 = W*in
   wire signed [14:0] m226_11;
   assign m226_11 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_12 = W*in
   wire signed [14:0] m226_12;
   assign m226_12 =15'b0;

   // m226_13 = W*in
   wire signed [14:0] m226_13;
   assign m226_13 =15'b0;

   // m226_14 = W*in
   wire signed [14:0] m226_14;
   assign m226_14 =15'b0;

   // m226_15 = W*in
   wire signed [14:0] m226_15;
   assign m226_15 =15'b0;

   // m226_16 = W*in
   wire signed [14:0] m226_16;
   assign m226_16 =15'b0;

   // m226_17 = W*in
   wire signed [14:0] m226_17;
   assign m226_17 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_18 = W*in
   wire signed [14:0] m226_18;
   assign m226_18 =15'b0;

   // m226_19 = W*in
   wire signed [14:0] m226_19;
   assign m226_19 =15'b0;

   // m226_20 = W*in
   wire signed [14:0] m226_20;
   assign m226_20 =15'b0;

   // m226_21 = W*in
   wire signed [14:0] m226_21;
   assign m226_21 ={ {4{neg226[14]}} , neg226[14:4] };

   // m226_22 = W*in
   wire signed [14:0] m226_22;
   assign m226_22 =15'b0;

   // m226_23 = W*in
   wire signed [14:0] m226_23;
   assign m226_23 =15'b0;

   // m226_24 = W*in
   wire signed [14:0] m226_24;
   assign m226_24 ={ {3{in226[14]}} , in226[14:3] };

   // m226_25 = W*in
   wire signed [14:0] m226_25;
   assign m226_25 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_26 = W*in
   wire signed [14:0] m226_26;
   assign m226_26 =15'b0;

   // m226_27 = W*in
   wire signed [14:0] m226_27;
   assign m226_27 =15'b0;

   // m226_28 = W*in
   wire signed [14:0] m226_28;
   assign m226_28 =15'b0;

   // m226_29 = W*in
   wire signed [14:0] m226_29;
   assign m226_29 ={ {4{neg226[14]}} , neg226[14:4] };

   // m226_30 = W*in
   wire signed [14:0] m226_30;
   assign m226_30 =15'b0;

   // m226_31 = W*in
   wire signed [14:0] m226_31;
   assign m226_31 =15'b0;

   // m226_32 = W*in
   wire signed [14:0] m226_32;
   assign m226_32 =15'b0;

   // m226_33 = W*in
   wire signed [14:0] m226_33;
   assign m226_33 ={ {3{in226[14]}} , in226[14:3] };

   // m226_34 = W*in
   wire signed [14:0] m226_34;
   assign m226_34 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_35 = W*in
   wire signed [14:0] m226_35;
   assign m226_35 =15'b0;

   // m226_36 = W*in
   wire signed [14:0] m226_36;
   assign m226_36 =15'b0;

   // m226_37 = W*in
   wire signed [14:0] m226_37;
   assign m226_37 =15'b0;

   // m226_38 = W*in
   wire signed [14:0] m226_38;
   assign m226_38 =15'b0;

   // m226_39 = W*in
   wire signed [14:0] m226_39;
   assign m226_39 =15'b0;

   // m226_40 = W*in
   wire signed [14:0] m226_40;
   assign m226_40 ={ {3{in226[14]}} , in226[14:3] };

   // m226_41 = W*in
   wire signed [14:0] m226_41;
   assign m226_41 =15'b0;

   // m226_42 = W*in
   wire signed [14:0] m226_42;
   assign m226_42 =15'b0;

   // m226_43 = W*in
   wire signed [14:0] m226_43;
   assign m226_43 =15'b0;

   // m226_44 = W*in
   wire signed [14:0] m226_44;
   assign m226_44 =15'b0;

   // m226_45 = W*in
   wire signed [14:0] m226_45;
   assign m226_45 =15'b0;

   // m226_46 = W*in
   wire signed [14:0] m226_46;
   assign m226_46 =15'b0;

   // m226_47 = W*in
   wire signed [14:0] m226_47;
   assign m226_47 =15'b0;

   // m226_48 = W*in
   wire signed [14:0] m226_48;
   assign m226_48 =15'b0;

   // m226_49 = W*in
   wire signed [14:0] m226_49;
   assign m226_49 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_50 = W*in
   wire signed [14:0] m226_50;
   assign m226_50 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_51 = W*in
   wire signed [14:0] m226_51;
   assign m226_51 =15'b0;

   // m226_52 = W*in
   wire signed [14:0] m226_52;
   assign m226_52 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_53 = W*in
   wire signed [14:0] m226_53;
   assign m226_53 =15'b0;

   // m226_54 = W*in
   wire signed [14:0] m226_54;
   assign m226_54 =15'b0;

   // m226_55 = W*in
   wire signed [14:0] m226_55;
   assign m226_55 =15'b0;

   // m226_56 = W*in
   wire signed [14:0] m226_56;
   assign m226_56 =15'b0;

   // m226_57 = W*in
   wire signed [14:0] m226_57;
   assign m226_57 ={ {2{in226[14]}} , in226[14:2] };

   // m226_58 = W*in
   wire signed [14:0] m226_58;
   assign m226_58 =15'b0;

   // m226_59 = W*in
   wire signed [14:0] m226_59;
   assign m226_59 ={ {3{in226[14]}} , in226[14:3] };

   // m226_60 = W*in
   wire signed [14:0] m226_60;
   assign m226_60 ={ {4{neg226[14]}} , neg226[14:4] };

   // m226_61 = W*in
   wire signed [14:0] m226_61;
   assign m226_61 =15'b0;

   // m226_62 = W*in
   wire signed [14:0] m226_62;
   assign m226_62 =15'b0;

   // m226_63 = W*in
   wire signed [14:0] m226_63;
   assign m226_63 ={ {3{in226[14]}} , in226[14:3] };

   // m226_64 = W*in
   wire signed [14:0] m226_64;
   assign m226_64 =15'b0;

   // m226_65 = W*in
   wire signed [14:0] m226_65;
   assign m226_65 =15'b0;

   // m226_66 = W*in
   wire signed [14:0] m226_66;
   assign m226_66 =15'b0;

   // m226_67 = W*in
   wire signed [14:0] m226_67;
   assign m226_67 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_68 = W*in
   wire signed [14:0] m226_68;
   assign m226_68 =15'b0;

   // m226_69 = W*in
   wire signed [14:0] m226_69;
   assign m226_69 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_70 = W*in
   wire signed [14:0] m226_70;
   assign m226_70 ={ {4{in226[14]}} , in226[14:4] };

   // m226_71 = W*in
   wire signed [14:0] m226_71;
   assign m226_71 =15'b0;

   // m226_72 = W*in
   wire signed [14:0] m226_72;
   assign m226_72 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_73 = W*in
   wire signed [14:0] m226_73;
   assign m226_73 =15'b0;

   // m226_74 = W*in
   wire signed [14:0] m226_74;
   assign m226_74 ={ {4{in226[14]}} , in226[14:4] };

   // m226_75 = W*in
   wire signed [14:0] m226_75;
   assign m226_75 =15'b0;

   // m226_76 = W*in
   wire signed [14:0] m226_76;
   assign m226_76 ={ {4{in226[14]}} , in226[14:4] };

   // m226_77 = W*in
   wire signed [14:0] m226_77;
   assign m226_77 =15'b0;

   // m226_78 = W*in
   wire signed [14:0] m226_78;
   assign m226_78 =15'b0;

   // m226_79 = W*in
   wire signed [14:0] m226_79;
   assign m226_79 =15'b0;

   // m226_80 = W*in
   wire signed [14:0] m226_80;
   assign m226_80 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_81 = W*in
   wire signed [14:0] m226_81;
   assign m226_81 =15'b0;

   // m226_82 = W*in
   wire signed [14:0] m226_82;
   assign m226_82 ={ {3{in226[14]}} , in226[14:3] };

   // m226_83 = W*in
   wire signed [14:0] m226_83;
   assign m226_83 ={ {3{in226[14]}} , in226[14:3] };

   // m226_84 = W*in
   wire signed [14:0] m226_84;
   assign m226_84 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_85 = W*in
   wire signed [14:0] m226_85;
   assign m226_85 =15'b0;

   // m226_86 = W*in
   wire signed [14:0] m226_86;
   assign m226_86 =15'b0;

   // m226_87 = W*in
   wire signed [14:0] m226_87;
   assign m226_87 =15'b0;

   // m226_88 = W*in
   wire signed [14:0] m226_88;
   assign m226_88 =15'b0;

   // m226_89 = W*in
   wire signed [14:0] m226_89;
   assign m226_89 =15'b0;

   // m226_90 = W*in
   wire signed [14:0] m226_90;
   assign m226_90 =15'b0;

   // m226_91 = W*in
   wire signed [14:0] m226_91;
   assign m226_91 =15'b0;

   // m226_92 = W*in
   wire signed [14:0] m226_92;
   assign m226_92 ={ {3{in226[14]}} , in226[14:3] };

   // m226_93 = W*in
   wire signed [14:0] m226_93;
   assign m226_93 =15'b0;

   // m226_94 = W*in
   wire signed [14:0] m226_94;
   assign m226_94 =15'b0;

   // m226_95 = W*in
   wire signed [14:0] m226_95;
   assign m226_95 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_96 = W*in
   wire signed [14:0] m226_96;
   assign m226_96 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_97 = W*in
   wire signed [14:0] m226_97;
   assign m226_97 ={ {3{in226[14]}} , in226[14:3] };

   // m226_98 = W*in
   wire signed [14:0] m226_98;
   assign m226_98 ={ {3{neg226[14]}} , neg226[14:3] };

   // m226_99 = W*in
   wire signed [14:0] m226_99;
   assign m226_99 =15'b0;

   // m226_100 = W*in
   wire signed [14:0] m226_100;
   assign m226_100 ={ {3{in226[14]}} , in226[14:3] };

   // m227_1 = W*in
   wire signed [14:0] m227_1;
   assign m227_1 =15'b0;

   // m227_2 = W*in
   wire signed [14:0] m227_2;
   assign m227_2 ={ {3{in227[14]}} , in227[14:3] };

   // m227_3 = W*in
   wire signed [14:0] m227_3;
   assign m227_3 =15'b0;

   // m227_4 = W*in
   wire signed [14:0] m227_4;
   assign m227_4 ={ {4{neg227[14]}} , neg227[14:4] };

   // m227_5 = W*in
   wire signed [14:0] m227_5;
   assign m227_5 =15'b0;

   // m227_6 = W*in
   wire signed [14:0] m227_6;
   assign m227_6 =15'b0;

   // m227_7 = W*in
   wire signed [14:0] m227_7;
   assign m227_7 ={ {3{in227[14]}} , in227[14:3] };

   // m227_8 = W*in
   wire signed [14:0] m227_8;
   assign m227_8 ={ {3{neg227[14]}} , neg227[14:3] };

   // m227_9 = W*in
   wire signed [14:0] m227_9;
   assign m227_9 ={ {3{in227[14]}} , in227[14:3] };

   // m227_10 = W*in
   wire signed [14:0] m227_10;
   assign m227_10 =15'b0;

   // m227_11 = W*in
   wire signed [14:0] m227_11;
   assign m227_11 =15'b0;

   // m227_12 = W*in
   wire signed [14:0] m227_12;
   assign m227_12 ={ {3{in227[14]}} , in227[14:3] };

   // m227_13 = W*in
   wire signed [14:0] m227_13;
   assign m227_13 =15'b0;

   // m227_14 = W*in
   wire signed [14:0] m227_14;
   assign m227_14 =15'b0;

   // m227_15 = W*in
   wire signed [14:0] m227_15;
   assign m227_15 =15'b0;

   // m227_16 = W*in
   wire signed [14:0] m227_16;
   assign m227_16 =15'b0;

   // m227_17 = W*in
   wire signed [14:0] m227_17;
   assign m227_17 ={ {4{neg227[14]}} , neg227[14:4] };

   // m227_18 = W*in
   wire signed [14:0] m227_18;
   assign m227_18 =15'b0;

   // m227_19 = W*in
   wire signed [14:0] m227_19;
   assign m227_19 =15'b0;

   // m227_20 = W*in
   wire signed [14:0] m227_20;
   assign m227_20 =15'b0;

   // m227_21 = W*in
   wire signed [14:0] m227_21;
   assign m227_21 =15'b0;

   // m227_22 = W*in
   wire signed [14:0] m227_22;
   assign m227_22 =15'b0;

   // m227_23 = W*in
   wire signed [14:0] m227_23;
   assign m227_23 =15'b0;

   // m227_24 = W*in
   wire signed [14:0] m227_24;
   assign m227_24 =15'b0;

   // m227_25 = W*in
   wire signed [14:0] m227_25;
   assign m227_25 =15'b0;

   // m227_26 = W*in
   wire signed [14:0] m227_26;
   assign m227_26 =15'b0;

   // m227_27 = W*in
   wire signed [14:0] m227_27;
   assign m227_27 =15'b0;

   // m227_28 = W*in
   wire signed [14:0] m227_28;
   assign m227_28 =15'b0;

   // m227_29 = W*in
   wire signed [14:0] m227_29;
   assign m227_29 =15'b0;

   // m227_30 = W*in
   wire signed [14:0] m227_30;
   assign m227_30 =15'b0;

   // m227_31 = W*in
   wire signed [14:0] m227_31;
   assign m227_31 =15'b0;

   // m227_32 = W*in
   wire signed [14:0] m227_32;
   assign m227_32 =15'b0;

   // m227_33 = W*in
   wire signed [14:0] m227_33;
   assign m227_33 =15'b0;

   // m227_34 = W*in
   wire signed [14:0] m227_34;
   assign m227_34 =15'b0;

   // m227_35 = W*in
   wire signed [14:0] m227_35;
   assign m227_35 =15'b0;

   // m227_36 = W*in
   wire signed [14:0] m227_36;
   assign m227_36 =15'b0;

   // m227_37 = W*in
   wire signed [14:0] m227_37;
   assign m227_37 ={ {3{neg227[14]}} , neg227[14:3] };

   // m227_38 = W*in
   wire signed [14:0] m227_38;
   assign m227_38 =15'b0;

   // m227_39 = W*in
   wire signed [14:0] m227_39;
   assign m227_39 ={ {3{neg227[14]}} , neg227[14:3] };

   // m227_40 = W*in
   wire signed [14:0] m227_40;
   assign m227_40 =15'b0;

   // m227_41 = W*in
   wire signed [14:0] m227_41;
   assign m227_41 =15'b0;

   // m227_42 = W*in
   wire signed [14:0] m227_42;
   assign m227_42 =15'b0;

   // m227_43 = W*in
   wire signed [14:0] m227_43;
   assign m227_43 =15'b0;

   // m227_44 = W*in
   wire signed [14:0] m227_44;
   assign m227_44 =15'b0;

   // m227_45 = W*in
   wire signed [14:0] m227_45;
   assign m227_45 =15'b0;

   // m227_46 = W*in
   wire signed [14:0] m227_46;
   assign m227_46 =15'b0;

   // m227_47 = W*in
   wire signed [14:0] m227_47;
   assign m227_47 =15'b0;

   // m227_48 = W*in
   wire signed [14:0] m227_48;
   assign m227_48 =15'b0;

   // m227_49 = W*in
   wire signed [14:0] m227_49;
   assign m227_49 =15'b0;

   // m227_50 = W*in
   wire signed [14:0] m227_50;
   assign m227_50 =15'b0;

   // m227_51 = W*in
   wire signed [14:0] m227_51;
   assign m227_51 =15'b0;

   // m227_52 = W*in
   wire signed [14:0] m227_52;
   assign m227_52 =15'b0;

   // m227_53 = W*in
   wire signed [14:0] m227_53;
   assign m227_53 =15'b0;

   // m227_54 = W*in
   wire signed [14:0] m227_54;
   assign m227_54 =15'b0;

   // m227_55 = W*in
   wire signed [14:0] m227_55;
   assign m227_55 =15'b0;

   // m227_56 = W*in
   wire signed [14:0] m227_56;
   assign m227_56 =15'b0;

   // m227_57 = W*in
   wire signed [14:0] m227_57;
   assign m227_57 =15'b0;

   // m227_58 = W*in
   wire signed [14:0] m227_58;
   assign m227_58 =15'b0;

   // m227_59 = W*in
   wire signed [14:0] m227_59;
   assign m227_59 =15'b0;

   // m227_60 = W*in
   wire signed [14:0] m227_60;
   assign m227_60 =15'b0;

   // m227_61 = W*in
   wire signed [14:0] m227_61;
   assign m227_61 =15'b0;

   // m227_62 = W*in
   wire signed [14:0] m227_62;
   assign m227_62 =15'b0;

   // m227_63 = W*in
   wire signed [14:0] m227_63;
   assign m227_63 =15'b0;

   // m227_64 = W*in
   wire signed [14:0] m227_64;
   assign m227_64 =15'b0;

   // m227_65 = W*in
   wire signed [14:0] m227_65;
   assign m227_65 =15'b0;

   // m227_66 = W*in
   wire signed [14:0] m227_66;
   assign m227_66 =15'b0;

   // m227_67 = W*in
   wire signed [14:0] m227_67;
   assign m227_67 =15'b0;

   // m227_68 = W*in
   wire signed [14:0] m227_68;
   assign m227_68 ={ {4{neg227[14]}} , neg227[14:4] };

   // m227_69 = W*in
   wire signed [14:0] m227_69;
   assign m227_69 =15'b0;

   // m227_70 = W*in
   wire signed [14:0] m227_70;
   assign m227_70 =15'b0;

   // m227_71 = W*in
   wire signed [14:0] m227_71;
   assign m227_71 ={ {3{neg227[14]}} , neg227[14:3] };

   // m227_72 = W*in
   wire signed [14:0] m227_72;
   assign m227_72 =15'b0;

   // m227_73 = W*in
   wire signed [14:0] m227_73;
   assign m227_73 =15'b0;

   // m227_74 = W*in
   wire signed [14:0] m227_74;
   assign m227_74 =15'b0;

   // m227_75 = W*in
   wire signed [14:0] m227_75;
   assign m227_75 =15'b0;

   // m227_76 = W*in
   wire signed [14:0] m227_76;
   assign m227_76 =15'b0;

   // m227_77 = W*in
   wire signed [14:0] m227_77;
   assign m227_77 =15'b0;

   // m227_78 = W*in
   wire signed [14:0] m227_78;
   assign m227_78 =15'b0;

   // m227_79 = W*in
   wire signed [14:0] m227_79;
   assign m227_79 =15'b0;

   // m227_80 = W*in
   wire signed [14:0] m227_80;
   assign m227_80 =15'b0;

   // m227_81 = W*in
   wire signed [14:0] m227_81;
   assign m227_81 =15'b0;

   // m227_82 = W*in
   wire signed [14:0] m227_82;
   assign m227_82 =15'b0;

   // m227_83 = W*in
   wire signed [14:0] m227_83;
   assign m227_83 =15'b0;

   // m227_84 = W*in
   wire signed [14:0] m227_84;
   assign m227_84 =15'b0;

   // m227_85 = W*in
   wire signed [14:0] m227_85;
   assign m227_85 =15'b0;

   // m227_86 = W*in
   wire signed [14:0] m227_86;
   assign m227_86 =15'b0;

   // m227_87 = W*in
   wire signed [14:0] m227_87;
   assign m227_87 =15'b0;

   // m227_88 = W*in
   wire signed [14:0] m227_88;
   assign m227_88 =15'b0;

   // m227_89 = W*in
   wire signed [14:0] m227_89;
   assign m227_89 =15'b0;

   // m227_90 = W*in
   wire signed [14:0] m227_90;
   assign m227_90 =15'b0;

   // m227_91 = W*in
   wire signed [14:0] m227_91;
   assign m227_91 =15'b0;

   // m227_92 = W*in
   wire signed [14:0] m227_92;
   assign m227_92 =15'b0;

   // m227_93 = W*in
   wire signed [14:0] m227_93;
   assign m227_93 =15'b0;

   // m227_94 = W*in
   wire signed [14:0] m227_94;
   assign m227_94 =15'b0;

   // m227_95 = W*in
   wire signed [14:0] m227_95;
   assign m227_95 =15'b0;

   // m227_96 = W*in
   wire signed [14:0] m227_96;
   assign m227_96 =15'b0;

   // m227_97 = W*in
   wire signed [14:0] m227_97;
   assign m227_97 =15'b0;

   // m227_98 = W*in
   wire signed [14:0] m227_98;
   assign m227_98 =15'b0;

   // m227_99 = W*in
   wire signed [14:0] m227_99;
   assign m227_99 =15'b0;

   // m227_100 = W*in
   wire signed [14:0] m227_100;
   assign m227_100 =15'b0;

   // m228_1 = W*in
   wire signed [14:0] m228_1;
   assign m228_1 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_2 = W*in
   wire signed [14:0] m228_2;
   assign m228_2 =15'b0;

   // m228_3 = W*in
   wire signed [14:0] m228_3;
   assign m228_3 =15'b0;

   // m228_4 = W*in
   wire signed [14:0] m228_4;
   assign m228_4 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_5 = W*in
   wire signed [14:0] m228_5;
   assign m228_5 =15'b0;

   // m228_6 = W*in
   wire signed [14:0] m228_6;
   assign m228_6 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_7 = W*in
   wire signed [14:0] m228_7;
   assign m228_7 =15'b0;

   // m228_8 = W*in
   wire signed [14:0] m228_8;
   assign m228_8 =15'b0;

   // m228_9 = W*in
   wire signed [14:0] m228_9;
   assign m228_9 =15'b0;

   // m228_10 = W*in
   wire signed [14:0] m228_10;
   assign m228_10 =15'b0;

   // m228_11 = W*in
   wire signed [14:0] m228_11;
   assign m228_11 =15'b0;

   // m228_12 = W*in
   wire signed [14:0] m228_12;
   assign m228_12 =15'b0;

   // m228_13 = W*in
   wire signed [14:0] m228_13;
   assign m228_13 =15'b0;

   // m228_14 = W*in
   wire signed [14:0] m228_14;
   assign m228_14 =15'b0;

   // m228_15 = W*in
   wire signed [14:0] m228_15;
   assign m228_15 ={ {3{in228[14]}} , in228[14:3] };

   // m228_16 = W*in
   wire signed [14:0] m228_16;
   assign m228_16 =15'b0;

   // m228_17 = W*in
   wire signed [14:0] m228_17;
   assign m228_17 =15'b0;

   // m228_18 = W*in
   wire signed [14:0] m228_18;
   assign m228_18 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_19 = W*in
   wire signed [14:0] m228_19;
   assign m228_19 ={ {4{in228[14]}} , in228[14:4] };

   // m228_20 = W*in
   wire signed [14:0] m228_20;
   assign m228_20 =15'b0;

   // m228_21 = W*in
   wire signed [14:0] m228_21;
   assign m228_21 =15'b0;

   // m228_22 = W*in
   wire signed [14:0] m228_22;
   assign m228_22 =15'b0;

   // m228_23 = W*in
   wire signed [14:0] m228_23;
   assign m228_23 =15'b0;

   // m228_24 = W*in
   wire signed [14:0] m228_24;
   assign m228_24 =15'b0;

   // m228_25 = W*in
   wire signed [14:0] m228_25;
   assign m228_25 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_26 = W*in
   wire signed [14:0] m228_26;
   assign m228_26 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_27 = W*in
   wire signed [14:0] m228_27;
   assign m228_27 ={ {3{in228[14]}} , in228[14:3] };

   // m228_28 = W*in
   wire signed [14:0] m228_28;
   assign m228_28 =15'b0;

   // m228_29 = W*in
   wire signed [14:0] m228_29;
   assign m228_29 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_30 = W*in
   wire signed [14:0] m228_30;
   assign m228_30 =15'b0;

   // m228_31 = W*in
   wire signed [14:0] m228_31;
   assign m228_31 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_32 = W*in
   wire signed [14:0] m228_32;
   assign m228_32 =15'b0;

   // m228_33 = W*in
   wire signed [14:0] m228_33;
   assign m228_33 =15'b0;

   // m228_34 = W*in
   wire signed [14:0] m228_34;
   assign m228_34 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_35 = W*in
   wire signed [14:0] m228_35;
   assign m228_35 =15'b0;

   // m228_36 = W*in
   wire signed [14:0] m228_36;
   assign m228_36 =15'b0;

   // m228_37 = W*in
   wire signed [14:0] m228_37;
   assign m228_37 =15'b0;

   // m228_38 = W*in
   wire signed [14:0] m228_38;
   assign m228_38 =15'b0;

   // m228_39 = W*in
   wire signed [14:0] m228_39;
   assign m228_39 =15'b0;

   // m228_40 = W*in
   wire signed [14:0] m228_40;
   assign m228_40 =15'b0;

   // m228_41 = W*in
   wire signed [14:0] m228_41;
   assign m228_41 =15'b0;

   // m228_42 = W*in
   wire signed [14:0] m228_42;
   assign m228_42 =15'b0;

   // m228_43 = W*in
   wire signed [14:0] m228_43;
   assign m228_43 =15'b0;

   // m228_44 = W*in
   wire signed [14:0] m228_44;
   assign m228_44 =15'b0;

   // m228_45 = W*in
   wire signed [14:0] m228_45;
   assign m228_45 =15'b0;

   // m228_46 = W*in
   wire signed [14:0] m228_46;
   assign m228_46 ={ {4{in228[14]}} , in228[14:4] };

   // m228_47 = W*in
   wire signed [14:0] m228_47;
   assign m228_47 =15'b0;

   // m228_48 = W*in
   wire signed [14:0] m228_48;
   assign m228_48 ={ {4{in228[14]}} , in228[14:4] };

   // m228_49 = W*in
   wire signed [14:0] m228_49;
   assign m228_49 =15'b0;

   // m228_50 = W*in
   wire signed [14:0] m228_50;
   assign m228_50 =15'b0;

   // m228_51 = W*in
   wire signed [14:0] m228_51;
   assign m228_51 =15'b0;

   // m228_52 = W*in
   wire signed [14:0] m228_52;
   assign m228_52 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_53 = W*in
   wire signed [14:0] m228_53;
   assign m228_53 =15'b0;

   // m228_54 = W*in
   wire signed [14:0] m228_54;
   assign m228_54 =15'b0;

   // m228_55 = W*in
   wire signed [14:0] m228_55;
   assign m228_55 =15'b0;

   // m228_56 = W*in
   wire signed [14:0] m228_56;
   assign m228_56 ={ {3{in228[14]}} , in228[14:3] };

   // m228_57 = W*in
   wire signed [14:0] m228_57;
   assign m228_57 =15'b0;

   // m228_58 = W*in
   wire signed [14:0] m228_58;
   assign m228_58 =15'b0;

   // m228_59 = W*in
   wire signed [14:0] m228_59;
   assign m228_59 ={ {4{in228[14]}} , in228[14:4] };

   // m228_60 = W*in
   wire signed [14:0] m228_60;
   assign m228_60 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_61 = W*in
   wire signed [14:0] m228_61;
   assign m228_61 ={ {4{in228[14]}} , in228[14:4] };

   // m228_62 = W*in
   wire signed [14:0] m228_62;
   assign m228_62 =15'b0;

   // m228_63 = W*in
   wire signed [14:0] m228_63;
   assign m228_63 ={ {4{in228[14]}} , in228[14:4] };

   // m228_64 = W*in
   wire signed [14:0] m228_64;
   assign m228_64 =15'b0;

   // m228_65 = W*in
   wire signed [14:0] m228_65;
   assign m228_65 =15'b0;

   // m228_66 = W*in
   wire signed [14:0] m228_66;
   assign m228_66 =15'b0;

   // m228_67 = W*in
   wire signed [14:0] m228_67;
   assign m228_67 =15'b0;

   // m228_68 = W*in
   wire signed [14:0] m228_68;
   assign m228_68 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_69 = W*in
   wire signed [14:0] m228_69;
   assign m228_69 =15'b0;

   // m228_70 = W*in
   wire signed [14:0] m228_70;
   assign m228_70 ={ {4{in228[14]}} , in228[14:4] };

   // m228_71 = W*in
   wire signed [14:0] m228_71;
   assign m228_71 =15'b0;

   // m228_72 = W*in
   wire signed [14:0] m228_72;
   assign m228_72 =15'b0;

   // m228_73 = W*in
   wire signed [14:0] m228_73;
   assign m228_73 =15'b0;

   // m228_74 = W*in
   wire signed [14:0] m228_74;
   assign m228_74 =15'b0;

   // m228_75 = W*in
   wire signed [14:0] m228_75;
   assign m228_75 =15'b0;

   // m228_76 = W*in
   wire signed [14:0] m228_76;
   assign m228_76 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_77 = W*in
   wire signed [14:0] m228_77;
   assign m228_77 =15'b0;

   // m228_78 = W*in
   wire signed [14:0] m228_78;
   assign m228_78 ={ {4{neg228[14]}} , neg228[14:4] };

   // m228_79 = W*in
   wire signed [14:0] m228_79;
   assign m228_79 =15'b0;

   // m228_80 = W*in
   wire signed [14:0] m228_80;
   assign m228_80 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_81 = W*in
   wire signed [14:0] m228_81;
   assign m228_81 =15'b0;

   // m228_82 = W*in
   wire signed [14:0] m228_82;
   assign m228_82 =15'b0;

   // m228_83 = W*in
   wire signed [14:0] m228_83;
   assign m228_83 =15'b0;

   // m228_84 = W*in
   wire signed [14:0] m228_84;
   assign m228_84 =15'b0;

   // m228_85 = W*in
   wire signed [14:0] m228_85;
   assign m228_85 =15'b0;

   // m228_86 = W*in
   wire signed [14:0] m228_86;
   assign m228_86 =15'b0;

   // m228_87 = W*in
   wire signed [14:0] m228_87;
   assign m228_87 =15'b0;

   // m228_88 = W*in
   wire signed [14:0] m228_88;
   assign m228_88 =15'b0;

   // m228_89 = W*in
   wire signed [14:0] m228_89;
   assign m228_89 =15'b0;

   // m228_90 = W*in
   wire signed [14:0] m228_90;
   assign m228_90 =15'b0;

   // m228_91 = W*in
   wire signed [14:0] m228_91;
   assign m228_91 =15'b0;

   // m228_92 = W*in
   wire signed [14:0] m228_92;
   assign m228_92 =15'b0;

   // m228_93 = W*in
   wire signed [14:0] m228_93;
   assign m228_93 =15'b0;

   // m228_94 = W*in
   wire signed [14:0] m228_94;
   assign m228_94 =15'b0;

   // m228_95 = W*in
   wire signed [14:0] m228_95;
   assign m228_95 =15'b0;

   // m228_96 = W*in
   wire signed [14:0] m228_96;
   assign m228_96 ={ {3{neg228[14]}} , neg228[14:3] };

   // m228_97 = W*in
   wire signed [14:0] m228_97;
   assign m228_97 =15'b0;

   // m228_98 = W*in
   wire signed [14:0] m228_98;
   assign m228_98 =15'b0;

   // m228_99 = W*in
   wire signed [14:0] m228_99;
   assign m228_99 =15'b0;

   // m228_100 = W*in
   wire signed [14:0] m228_100;
   assign m228_100 =15'b0;

   // m229_1 = W*in
   wire signed [14:0] m229_1;
   assign m229_1 =15'b0;

   // m229_2 = W*in
   wire signed [14:0] m229_2;
   assign m229_2 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_3 = W*in
   wire signed [14:0] m229_3;
   assign m229_3 =15'b0;

   // m229_4 = W*in
   wire signed [14:0] m229_4;
   assign m229_4 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_5 = W*in
   wire signed [14:0] m229_5;
   assign m229_5 =15'b0;

   // m229_6 = W*in
   wire signed [14:0] m229_6;
   assign m229_6 =15'b0;

   // m229_7 = W*in
   wire signed [14:0] m229_7;
   assign m229_7 =15'b0;

   // m229_8 = W*in
   wire signed [14:0] m229_8;
   assign m229_8 =15'b0;

   // m229_9 = W*in
   wire signed [14:0] m229_9;
   assign m229_9 ={ {3{in229[14]}} , in229[14:3] };

   // m229_10 = W*in
   wire signed [14:0] m229_10;
   assign m229_10 =15'b0;

   // m229_11 = W*in
   wire signed [14:0] m229_11;
   assign m229_11 =15'b0;

   // m229_12 = W*in
   wire signed [14:0] m229_12;
   assign m229_12 =15'b0;

   // m229_13 = W*in
   wire signed [14:0] m229_13;
   assign m229_13 ={ {2{neg229[14]}} , neg229[14:2] };

   // m229_14 = W*in
   wire signed [14:0] m229_14;
   assign m229_14 =15'b0;

   // m229_15 = W*in
   wire signed [14:0] m229_15;
   assign m229_15 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_16 = W*in
   wire signed [14:0] m229_16;
   assign m229_16 =15'b0;

   // m229_17 = W*in
   wire signed [14:0] m229_17;
   assign m229_17 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_18 = W*in
   wire signed [14:0] m229_18;
   assign m229_18 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_19 = W*in
   wire signed [14:0] m229_19;
   assign m229_19 ={ {3{in229[14]}} , in229[14:3] };

   // m229_20 = W*in
   wire signed [14:0] m229_20;
   assign m229_20 ={ {4{neg229[14]}} , neg229[14:4] };

   // m229_21 = W*in
   wire signed [14:0] m229_21;
   assign m229_21 =15'b0;

   // m229_22 = W*in
   wire signed [14:0] m229_22;
   assign m229_22 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_23 = W*in
   wire signed [14:0] m229_23;
   assign m229_23 =15'b0;

   // m229_24 = W*in
   wire signed [14:0] m229_24;
   assign m229_24 ={ {3{in229[14]}} , in229[14:3] };

   // m229_25 = W*in
   wire signed [14:0] m229_25;
   assign m229_25 =15'b0;

   // m229_26 = W*in
   wire signed [14:0] m229_26;
   assign m229_26 ={ {4{in229[14]}} , in229[14:4] };

   // m229_27 = W*in
   wire signed [14:0] m229_27;
   assign m229_27 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_28 = W*in
   wire signed [14:0] m229_28;
   assign m229_28 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_29 = W*in
   wire signed [14:0] m229_29;
   assign m229_29 ={ {3{in229[14]}} , in229[14:3] };

   // m229_30 = W*in
   wire signed [14:0] m229_30;
   assign m229_30 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_31 = W*in
   wire signed [14:0] m229_31;
   assign m229_31 ={ {4{in229[14]}} , in229[14:4] };

   // m229_32 = W*in
   wire signed [14:0] m229_32;
   assign m229_32 =15'b0;

   // m229_33 = W*in
   wire signed [14:0] m229_33;
   assign m229_33 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_34 = W*in
   wire signed [14:0] m229_34;
   assign m229_34 ={ {3{in229[14]}} , in229[14:3] };

   // m229_35 = W*in
   wire signed [14:0] m229_35;
   assign m229_35 =15'b0;

   // m229_36 = W*in
   wire signed [14:0] m229_36;
   assign m229_36 =15'b0;

   // m229_37 = W*in
   wire signed [14:0] m229_37;
   assign m229_37 =15'b0;

   // m229_38 = W*in
   wire signed [14:0] m229_38;
   assign m229_38 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_39 = W*in
   wire signed [14:0] m229_39;
   assign m229_39 =15'b0;

   // m229_40 = W*in
   wire signed [14:0] m229_40;
   assign m229_40 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_41 = W*in
   wire signed [14:0] m229_41;
   assign m229_41 =15'b0;

   // m229_42 = W*in
   wire signed [14:0] m229_42;
   assign m229_42 =15'b0;

   // m229_43 = W*in
   wire signed [14:0] m229_43;
   assign m229_43 =15'b0;

   // m229_44 = W*in
   wire signed [14:0] m229_44;
   assign m229_44 =15'b0;

   // m229_45 = W*in
   wire signed [14:0] m229_45;
   assign m229_45 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_46 = W*in
   wire signed [14:0] m229_46;
   assign m229_46 =15'b0;

   // m229_47 = W*in
   wire signed [14:0] m229_47;
   assign m229_47 ={ {2{in229[14]}} , in229[14:2] };

   // m229_48 = W*in
   wire signed [14:0] m229_48;
   assign m229_48 =15'b0;

   // m229_49 = W*in
   wire signed [14:0] m229_49;
   assign m229_49 =15'b0;

   // m229_50 = W*in
   wire signed [14:0] m229_50;
   assign m229_50 =15'b0;

   // m229_51 = W*in
   wire signed [14:0] m229_51;
   assign m229_51 =15'b0;

   // m229_52 = W*in
   wire signed [14:0] m229_52;
   assign m229_52 ={ {3{in229[14]}} , in229[14:3] };

   // m229_53 = W*in
   wire signed [14:0] m229_53;
   assign m229_53 =15'b0;

   // m229_54 = W*in
   wire signed [14:0] m229_54;
   assign m229_54 =15'b0;

   // m229_55 = W*in
   wire signed [14:0] m229_55;
   assign m229_55 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_56 = W*in
   wire signed [14:0] m229_56;
   assign m229_56 =15'b0;

   // m229_57 = W*in
   wire signed [14:0] m229_57;
   assign m229_57 =15'b0;

   // m229_58 = W*in
   wire signed [14:0] m229_58;
   assign m229_58 =15'b0;

   // m229_59 = W*in
   wire signed [14:0] m229_59;
   assign m229_59 ={ {4{in229[14]}} , in229[14:4] };

   // m229_60 = W*in
   wire signed [14:0] m229_60;
   assign m229_60 =15'b0;

   // m229_61 = W*in
   wire signed [14:0] m229_61;
   assign m229_61 =15'b0;

   // m229_62 = W*in
   wire signed [14:0] m229_62;
   assign m229_62 =15'b0;

   // m229_63 = W*in
   wire signed [14:0] m229_63;
   assign m229_63 =15'b0;

   // m229_64 = W*in
   wire signed [14:0] m229_64;
   assign m229_64 =15'b0;

   // m229_65 = W*in
   wire signed [14:0] m229_65;
   assign m229_65 =15'b0;

   // m229_66 = W*in
   wire signed [14:0] m229_66;
   assign m229_66 =15'b0;

   // m229_67 = W*in
   wire signed [14:0] m229_67;
   assign m229_67 =15'b0;

   // m229_68 = W*in
   wire signed [14:0] m229_68;
   assign m229_68 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_69 = W*in
   wire signed [14:0] m229_69;
   assign m229_69 =15'b0;

   // m229_70 = W*in
   wire signed [14:0] m229_70;
   assign m229_70 =15'b0;

   // m229_71 = W*in
   wire signed [14:0] m229_71;
   assign m229_71 =15'b0;

   // m229_72 = W*in
   wire signed [14:0] m229_72;
   assign m229_72 =15'b0;

   // m229_73 = W*in
   wire signed [14:0] m229_73;
   assign m229_73 ={ {3{in229[14]}} , in229[14:3] };

   // m229_74 = W*in
   wire signed [14:0] m229_74;
   assign m229_74 =15'b0;

   // m229_75 = W*in
   wire signed [14:0] m229_75;
   assign m229_75 =15'b0;

   // m229_76 = W*in
   wire signed [14:0] m229_76;
   assign m229_76 =15'b0;

   // m229_77 = W*in
   wire signed [14:0] m229_77;
   assign m229_77 =15'b0;

   // m229_78 = W*in
   wire signed [14:0] m229_78;
   assign m229_78 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_79 = W*in
   wire signed [14:0] m229_79;
   assign m229_79 ={ {2{in229[14]}} , in229[14:2] };

   // m229_80 = W*in
   wire signed [14:0] m229_80;
   assign m229_80 =15'b0;

   // m229_81 = W*in
   wire signed [14:0] m229_81;
   assign m229_81 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_82 = W*in
   wire signed [14:0] m229_82;
   assign m229_82 =15'b0;

   // m229_83 = W*in
   wire signed [14:0] m229_83;
   assign m229_83 =15'b0;

   // m229_84 = W*in
   wire signed [14:0] m229_84;
   assign m229_84 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_85 = W*in
   wire signed [14:0] m229_85;
   assign m229_85 =15'b0;

   // m229_86 = W*in
   wire signed [14:0] m229_86;
   assign m229_86 =15'b0;

   // m229_87 = W*in
   wire signed [14:0] m229_87;
   assign m229_87 =15'b0;

   // m229_88 = W*in
   wire signed [14:0] m229_88;
   assign m229_88 ={ {3{in229[14]}} , in229[14:3] };

   // m229_89 = W*in
   wire signed [14:0] m229_89;
   assign m229_89 =15'b0;

   // m229_90 = W*in
   wire signed [14:0] m229_90;
   assign m229_90 =15'b0;

   // m229_91 = W*in
   wire signed [14:0] m229_91;
   assign m229_91 =15'b0;

   // m229_92 = W*in
   wire signed [14:0] m229_92;
   assign m229_92 =15'b0;

   // m229_93 = W*in
   wire signed [14:0] m229_93;
   assign m229_93 =15'b0;

   // m229_94 = W*in
   wire signed [14:0] m229_94;
   assign m229_94 =15'b0;

   // m229_95 = W*in
   wire signed [14:0] m229_95;
   assign m229_95 =15'b0;

   // m229_96 = W*in
   wire signed [14:0] m229_96;
   assign m229_96 ={ {3{in229[14]}} , in229[14:3] };

   // m229_97 = W*in
   wire signed [14:0] m229_97;
   assign m229_97 ={ {3{neg229[14]}} , neg229[14:3] };

   // m229_98 = W*in
   wire signed [14:0] m229_98;
   assign m229_98 =15'b0;

   // m229_99 = W*in
   wire signed [14:0] m229_99;
   assign m229_99 =15'b0;

   // m229_100 = W*in
   wire signed [14:0] m229_100;
   assign m229_100 =15'b0;

   // m230_1 = W*in
   wire signed [14:0] m230_1;
   assign m230_1 =15'b0;

   // m230_2 = W*in
   wire signed [14:0] m230_2;
   assign m230_2 =15'b0;

   // m230_3 = W*in
   wire signed [14:0] m230_3;
   assign m230_3 =15'b0;

   // m230_4 = W*in
   wire signed [14:0] m230_4;
   assign m230_4 =15'b0;

   // m230_5 = W*in
   wire signed [14:0] m230_5;
   assign m230_5 ={ {4{in230[14]}} , in230[14:4] };

   // m230_6 = W*in
   wire signed [14:0] m230_6;
   assign m230_6 =15'b0;

   // m230_7 = W*in
   wire signed [14:0] m230_7;
   assign m230_7 =15'b0;

   // m230_8 = W*in
   wire signed [14:0] m230_8;
   assign m230_8 =15'b0;

   // m230_9 = W*in
   wire signed [14:0] m230_9;
   assign m230_9 =15'b0;

   // m230_10 = W*in
   wire signed [14:0] m230_10;
   assign m230_10 =15'b0;

   // m230_11 = W*in
   wire signed [14:0] m230_11;
   assign m230_11 =15'b0;

   // m230_12 = W*in
   wire signed [14:0] m230_12;
   assign m230_12 =15'b0;

   // m230_13 = W*in
   wire signed [14:0] m230_13;
   assign m230_13 =15'b0;

   // m230_14 = W*in
   wire signed [14:0] m230_14;
   assign m230_14 =15'b0;

   // m230_15 = W*in
   wire signed [14:0] m230_15;
   assign m230_15 ={ {3{in230[14]}} , in230[14:3] };

   // m230_16 = W*in
   wire signed [14:0] m230_16;
   assign m230_16 =15'b0;

   // m230_17 = W*in
   wire signed [14:0] m230_17;
   assign m230_17 =15'b0;

   // m230_18 = W*in
   wire signed [14:0] m230_18;
   assign m230_18 =15'b0;

   // m230_19 = W*in
   wire signed [14:0] m230_19;
   assign m230_19 =15'b0;

   // m230_20 = W*in
   wire signed [14:0] m230_20;
   assign m230_20 =15'b0;

   // m230_21 = W*in
   wire signed [14:0] m230_21;
   assign m230_21 =15'b0;

   // m230_22 = W*in
   wire signed [14:0] m230_22;
   assign m230_22 =15'b0;

   // m230_23 = W*in
   wire signed [14:0] m230_23;
   assign m230_23 =15'b0;

   // m230_24 = W*in
   wire signed [14:0] m230_24;
   assign m230_24 =15'b0;

   // m230_25 = W*in
   wire signed [14:0] m230_25;
   assign m230_25 ={ {4{neg230[14]}} , neg230[14:4] };

   // m230_26 = W*in
   wire signed [14:0] m230_26;
   assign m230_26 ={ {4{neg230[14]}} , neg230[14:4] };

   // m230_27 = W*in
   wire signed [14:0] m230_27;
   assign m230_27 ={ {4{in230[14]}} , in230[14:4] };

   // m230_28 = W*in
   wire signed [14:0] m230_28;
   assign m230_28 ={ {4{in230[14]}} , in230[14:4] };

   // m230_29 = W*in
   wire signed [14:0] m230_29;
   assign m230_29 ={ {4{neg230[14]}} , neg230[14:4] };

   // m230_30 = W*in
   wire signed [14:0] m230_30;
   assign m230_30 =15'b0;

   // m230_31 = W*in
   wire signed [14:0] m230_31;
   assign m230_31 ={ {4{neg230[14]}} , neg230[14:4] };

   // m230_32 = W*in
   wire signed [14:0] m230_32;
   assign m230_32 =15'b0;

   // m230_33 = W*in
   wire signed [14:0] m230_33;
   assign m230_33 =15'b0;

   // m230_34 = W*in
   wire signed [14:0] m230_34;
   assign m230_34 ={ {3{neg230[14]}} , neg230[14:3] };

   // m230_35 = W*in
   wire signed [14:0] m230_35;
   assign m230_35 =15'b0;

   // m230_36 = W*in
   wire signed [14:0] m230_36;
   assign m230_36 =15'b0;

   // m230_37 = W*in
   wire signed [14:0] m230_37;
   assign m230_37 =15'b0;

   // m230_38 = W*in
   wire signed [14:0] m230_38;
   assign m230_38 =15'b0;

   // m230_39 = W*in
   wire signed [14:0] m230_39;
   assign m230_39 =15'b0;

   // m230_40 = W*in
   wire signed [14:0] m230_40;
   assign m230_40 ={ {4{in230[14]}} , in230[14:4] };

   // m230_41 = W*in
   wire signed [14:0] m230_41;
   assign m230_41 =15'b0;

   // m230_42 = W*in
   wire signed [14:0] m230_42;
   assign m230_42 =15'b0;

   // m230_43 = W*in
   wire signed [14:0] m230_43;
   assign m230_43 =15'b0;

   // m230_44 = W*in
   wire signed [14:0] m230_44;
   assign m230_44 =15'b0;

   // m230_45 = W*in
   wire signed [14:0] m230_45;
   assign m230_45 =15'b0;

   // m230_46 = W*in
   wire signed [14:0] m230_46;
   assign m230_46 =15'b0;

   // m230_47 = W*in
   wire signed [14:0] m230_47;
   assign m230_47 =15'b0;

   // m230_48 = W*in
   wire signed [14:0] m230_48;
   assign m230_48 =15'b0;

   // m230_49 = W*in
   wire signed [14:0] m230_49;
   assign m230_49 =15'b0;

   // m230_50 = W*in
   wire signed [14:0] m230_50;
   assign m230_50 =15'b0;

   // m230_51 = W*in
   wire signed [14:0] m230_51;
   assign m230_51 =15'b0;

   // m230_52 = W*in
   wire signed [14:0] m230_52;
   assign m230_52 =15'b0;

   // m230_53 = W*in
   wire signed [14:0] m230_53;
   assign m230_53 =15'b0;

   // m230_54 = W*in
   wire signed [14:0] m230_54;
   assign m230_54 =15'b0;

   // m230_55 = W*in
   wire signed [14:0] m230_55;
   assign m230_55 =15'b0;

   // m230_56 = W*in
   wire signed [14:0] m230_56;
   assign m230_56 =15'b0;

   // m230_57 = W*in
   wire signed [14:0] m230_57;
   assign m230_57 =15'b0;

   // m230_58 = W*in
   wire signed [14:0] m230_58;
   assign m230_58 =15'b0;

   // m230_59 = W*in
   wire signed [14:0] m230_59;
   assign m230_59 =15'b0;

   // m230_60 = W*in
   wire signed [14:0] m230_60;
   assign m230_60 ={ {3{neg230[14]}} , neg230[14:3] };

   // m230_61 = W*in
   wire signed [14:0] m230_61;
   assign m230_61 =15'b0;

   // m230_62 = W*in
   wire signed [14:0] m230_62;
   assign m230_62 =15'b0;

   // m230_63 = W*in
   wire signed [14:0] m230_63;
   assign m230_63 ={ {3{in230[14]}} , in230[14:3] };

   // m230_64 = W*in
   wire signed [14:0] m230_64;
   assign m230_64 =15'b0;

   // m230_65 = W*in
   wire signed [14:0] m230_65;
   assign m230_65 =15'b0;

   // m230_66 = W*in
   wire signed [14:0] m230_66;
   assign m230_66 =15'b0;

   // m230_67 = W*in
   wire signed [14:0] m230_67;
   assign m230_67 =15'b0;

   // m230_68 = W*in
   wire signed [14:0] m230_68;
   assign m230_68 =15'b0;

   // m230_69 = W*in
   wire signed [14:0] m230_69;
   assign m230_69 ={ {4{neg230[14]}} , neg230[14:4] };

   // m230_70 = W*in
   wire signed [14:0] m230_70;
   assign m230_70 ={ {4{in230[14]}} , in230[14:4] };

   // m230_71 = W*in
   wire signed [14:0] m230_71;
   assign m230_71 =15'b0;

   // m230_72 = W*in
   wire signed [14:0] m230_72;
   assign m230_72 =15'b0;

   // m230_73 = W*in
   wire signed [14:0] m230_73;
   assign m230_73 =15'b0;

   // m230_74 = W*in
   wire signed [14:0] m230_74;
   assign m230_74 =15'b0;

   // m230_75 = W*in
   wire signed [14:0] m230_75;
   assign m230_75 =15'b0;

   // m230_76 = W*in
   wire signed [14:0] m230_76;
   assign m230_76 =15'b0;

   // m230_77 = W*in
   wire signed [14:0] m230_77;
   assign m230_77 =15'b0;

   // m230_78 = W*in
   wire signed [14:0] m230_78;
   assign m230_78 =15'b0;

   // m230_79 = W*in
   wire signed [14:0] m230_79;
   assign m230_79 =15'b0;

   // m230_80 = W*in
   wire signed [14:0] m230_80;
   assign m230_80 =15'b0;

   // m230_81 = W*in
   wire signed [14:0] m230_81;
   assign m230_81 =15'b0;

   // m230_82 = W*in
   wire signed [14:0] m230_82;
   assign m230_82 =15'b0;

   // m230_83 = W*in
   wire signed [14:0] m230_83;
   assign m230_83 =15'b0;

   // m230_84 = W*in
   wire signed [14:0] m230_84;
   assign m230_84 =15'b0;

   // m230_85 = W*in
   wire signed [14:0] m230_85;
   assign m230_85 =15'b0;

   // m230_86 = W*in
   wire signed [14:0] m230_86;
   assign m230_86 =15'b0;

   // m230_87 = W*in
   wire signed [14:0] m230_87;
   assign m230_87 =15'b0;

   // m230_88 = W*in
   wire signed [14:0] m230_88;
   assign m230_88 =15'b0;

   // m230_89 = W*in
   wire signed [14:0] m230_89;
   assign m230_89 =15'b0;

   // m230_90 = W*in
   wire signed [14:0] m230_90;
   assign m230_90 =15'b0;

   // m230_91 = W*in
   wire signed [14:0] m230_91;
   assign m230_91 =15'b0;

   // m230_92 = W*in
   wire signed [14:0] m230_92;
   assign m230_92 =15'b0;

   // m230_93 = W*in
   wire signed [14:0] m230_93;
   assign m230_93 =15'b0;

   // m230_94 = W*in
   wire signed [14:0] m230_94;
   assign m230_94 =15'b0;

   // m230_95 = W*in
   wire signed [14:0] m230_95;
   assign m230_95 =15'b0;

   // m230_96 = W*in
   wire signed [14:0] m230_96;
   assign m230_96 =15'b0;

   // m230_97 = W*in
   wire signed [14:0] m230_97;
   assign m230_97 =15'b0;

   // m230_98 = W*in
   wire signed [14:0] m230_98;
   assign m230_98 =15'b0;

   // m230_99 = W*in
   wire signed [14:0] m230_99;
   assign m230_99 =15'b0;

   // m230_100 = W*in
   wire signed [14:0] m230_100;
   assign m230_100 =15'b0;

   // m231_1 = W*in
   wire signed [14:0] m231_1;
   assign m231_1 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_2 = W*in
   wire signed [14:0] m231_2;
   assign m231_2 =15'b0;

   // m231_3 = W*in
   wire signed [14:0] m231_3;
   assign m231_3 =15'b0;

   // m231_4 = W*in
   wire signed [14:0] m231_4;
   assign m231_4 =15'b0;

   // m231_5 = W*in
   wire signed [14:0] m231_5;
   assign m231_5 ={ {3{in231[14]}} , in231[14:3] };

   // m231_6 = W*in
   wire signed [14:0] m231_6;
   assign m231_6 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_7 = W*in
   wire signed [14:0] m231_7;
   assign m231_7 =15'b0;

   // m231_8 = W*in
   wire signed [14:0] m231_8;
   assign m231_8 =15'b0;

   // m231_9 = W*in
   wire signed [14:0] m231_9;
   assign m231_9 =15'b0;

   // m231_10 = W*in
   wire signed [14:0] m231_10;
   assign m231_10 ={ {3{in231[14]}} , in231[14:3] };

   // m231_11 = W*in
   wire signed [14:0] m231_11;
   assign m231_11 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_12 = W*in
   wire signed [14:0] m231_12;
   assign m231_12 =15'b0;

   // m231_13 = W*in
   wire signed [14:0] m231_13;
   assign m231_13 =15'b0;

   // m231_14 = W*in
   wire signed [14:0] m231_14;
   assign m231_14 ={ {3{in231[14]}} , in231[14:3] };

   // m231_15 = W*in
   wire signed [14:0] m231_15;
   assign m231_15 ={ {4{in231[14]}} , in231[14:4] };

   // m231_16 = W*in
   wire signed [14:0] m231_16;
   assign m231_16 ={ {4{in231[14]}} , in231[14:4] };

   // m231_17 = W*in
   wire signed [14:0] m231_17;
   assign m231_17 =15'b0;

   // m231_18 = W*in
   wire signed [14:0] m231_18;
   assign m231_18 =15'b0;

   // m231_19 = W*in
   wire signed [14:0] m231_19;
   assign m231_19 =15'b0;

   // m231_20 = W*in
   wire signed [14:0] m231_20;
   assign m231_20 ={ {4{neg231[14]}} , neg231[14:4] };

   // m231_21 = W*in
   wire signed [14:0] m231_21;
   assign m231_21 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_22 = W*in
   wire signed [14:0] m231_22;
   assign m231_22 =15'b0;

   // m231_23 = W*in
   wire signed [14:0] m231_23;
   assign m231_23 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_24 = W*in
   wire signed [14:0] m231_24;
   assign m231_24 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_25 = W*in
   wire signed [14:0] m231_25;
   assign m231_25 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_26 = W*in
   wire signed [14:0] m231_26;
   assign m231_26 =15'b0;

   // m231_27 = W*in
   wire signed [14:0] m231_27;
   assign m231_27 =15'b0;

   // m231_28 = W*in
   wire signed [14:0] m231_28;
   assign m231_28 =15'b0;

   // m231_29 = W*in
   wire signed [14:0] m231_29;
   assign m231_29 =15'b0;

   // m231_30 = W*in
   wire signed [14:0] m231_30;
   assign m231_30 =15'b0;

   // m231_31 = W*in
   wire signed [14:0] m231_31;
   assign m231_31 ={ {3{in231[14]}} , in231[14:3] };

   // m231_32 = W*in
   wire signed [14:0] m231_32;
   assign m231_32 =15'b0;

   // m231_33 = W*in
   wire signed [14:0] m231_33;
   assign m231_33 =15'b0;

   // m231_34 = W*in
   wire signed [14:0] m231_34;
   assign m231_34 =15'b0;

   // m231_35 = W*in
   wire signed [14:0] m231_35;
   assign m231_35 =15'b0;

   // m231_36 = W*in
   wire signed [14:0] m231_36;
   assign m231_36 =15'b0;

   // m231_37 = W*in
   wire signed [14:0] m231_37;
   assign m231_37 =15'b0;

   // m231_38 = W*in
   wire signed [14:0] m231_38;
   assign m231_38 =15'b0;

   // m231_39 = W*in
   wire signed [14:0] m231_39;
   assign m231_39 =15'b0;

   // m231_40 = W*in
   wire signed [14:0] m231_40;
   assign m231_40 ={ {4{in231[14]}} , in231[14:4] };

   // m231_41 = W*in
   wire signed [14:0] m231_41;
   assign m231_41 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_42 = W*in
   wire signed [14:0] m231_42;
   assign m231_42 =15'b0;

   // m231_43 = W*in
   wire signed [14:0] m231_43;
   assign m231_43 =15'b0;

   // m231_44 = W*in
   wire signed [14:0] m231_44;
   assign m231_44 =15'b0;

   // m231_45 = W*in
   wire signed [14:0] m231_45;
   assign m231_45 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_46 = W*in
   wire signed [14:0] m231_46;
   assign m231_46 ={ {3{in231[14]}} , in231[14:3] };

   // m231_47 = W*in
   wire signed [14:0] m231_47;
   assign m231_47 =15'b0;

   // m231_48 = W*in
   wire signed [14:0] m231_48;
   assign m231_48 ={ {3{in231[14]}} , in231[14:3] };

   // m231_49 = W*in
   wire signed [14:0] m231_49;
   assign m231_49 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_50 = W*in
   wire signed [14:0] m231_50;
   assign m231_50 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_51 = W*in
   wire signed [14:0] m231_51;
   assign m231_51 =15'b0;

   // m231_52 = W*in
   wire signed [14:0] m231_52;
   assign m231_52 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_53 = W*in
   wire signed [14:0] m231_53;
   assign m231_53 =15'b0;

   // m231_54 = W*in
   wire signed [14:0] m231_54;
   assign m231_54 =15'b0;

   // m231_55 = W*in
   wire signed [14:0] m231_55;
   assign m231_55 ={ {3{in231[14]}} , in231[14:3] };

   // m231_56 = W*in
   wire signed [14:0] m231_56;
   assign m231_56 =15'b0;

   // m231_57 = W*in
   wire signed [14:0] m231_57;
   assign m231_57 ={ {2{in231[14]}} , in231[14:2] };

   // m231_58 = W*in
   wire signed [14:0] m231_58;
   assign m231_58 =15'b0;

   // m231_59 = W*in
   wire signed [14:0] m231_59;
   assign m231_59 =15'b0;

   // m231_60 = W*in
   wire signed [14:0] m231_60;
   assign m231_60 =15'b0;

   // m231_61 = W*in
   wire signed [14:0] m231_61;
   assign m231_61 ={ {3{in231[14]}} , in231[14:3] };

   // m231_62 = W*in
   wire signed [14:0] m231_62;
   assign m231_62 =15'b0;

   // m231_63 = W*in
   wire signed [14:0] m231_63;
   assign m231_63 ={ {2{in231[14]}} , in231[14:2] };

   // m231_64 = W*in
   wire signed [14:0] m231_64;
   assign m231_64 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_65 = W*in
   wire signed [14:0] m231_65;
   assign m231_65 =15'b0;

   // m231_66 = W*in
   wire signed [14:0] m231_66;
   assign m231_66 =15'b0;

   // m231_67 = W*in
   wire signed [14:0] m231_67;
   assign m231_67 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_68 = W*in
   wire signed [14:0] m231_68;
   assign m231_68 ={ {4{in231[14]}} , in231[14:4] };

   // m231_69 = W*in
   wire signed [14:0] m231_69;
   assign m231_69 =15'b0;

   // m231_70 = W*in
   wire signed [14:0] m231_70;
   assign m231_70 =15'b0;

   // m231_71 = W*in
   wire signed [14:0] m231_71;
   assign m231_71 ={ {3{in231[14]}} , in231[14:3] };

   // m231_72 = W*in
   wire signed [14:0] m231_72;
   assign m231_72 =15'b0;

   // m231_73 = W*in
   wire signed [14:0] m231_73;
   assign m231_73 =15'b0;

   // m231_74 = W*in
   wire signed [14:0] m231_74;
   assign m231_74 =15'b0;

   // m231_75 = W*in
   wire signed [14:0] m231_75;
   assign m231_75 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_76 = W*in
   wire signed [14:0] m231_76;
   assign m231_76 =15'b0;

   // m231_77 = W*in
   wire signed [14:0] m231_77;
   assign m231_77 =15'b0;

   // m231_78 = W*in
   wire signed [14:0] m231_78;
   assign m231_78 =15'b0;

   // m231_79 = W*in
   wire signed [14:0] m231_79;
   assign m231_79 =15'b0;

   // m231_80 = W*in
   wire signed [14:0] m231_80;
   assign m231_80 =15'b0;

   // m231_81 = W*in
   wire signed [14:0] m231_81;
   assign m231_81 =15'b0;

   // m231_82 = W*in
   wire signed [14:0] m231_82;
   assign m231_82 ={ {3{in231[14]}} , in231[14:3] };

   // m231_83 = W*in
   wire signed [14:0] m231_83;
   assign m231_83 ={ {3{in231[14]}} , in231[14:3] };

   // m231_84 = W*in
   wire signed [14:0] m231_84;
   assign m231_84 =15'b0;

   // m231_85 = W*in
   wire signed [14:0] m231_85;
   assign m231_85 =15'b0;

   // m231_86 = W*in
   wire signed [14:0] m231_86;
   assign m231_86 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_87 = W*in
   wire signed [14:0] m231_87;
   assign m231_87 =15'b0;

   // m231_88 = W*in
   wire signed [14:0] m231_88;
   assign m231_88 =15'b0;

   // m231_89 = W*in
   wire signed [14:0] m231_89;
   assign m231_89 ={ {3{in231[14]}} , in231[14:3] };

   // m231_90 = W*in
   wire signed [14:0] m231_90;
   assign m231_90 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_91 = W*in
   wire signed [14:0] m231_91;
   assign m231_91 =15'b0;

   // m231_92 = W*in
   wire signed [14:0] m231_92;
   assign m231_92 =15'b0;

   // m231_93 = W*in
   wire signed [14:0] m231_93;
   assign m231_93 =15'b0;

   // m231_94 = W*in
   wire signed [14:0] m231_94;
   assign m231_94 =15'b0;

   // m231_95 = W*in
   wire signed [14:0] m231_95;
   assign m231_95 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_96 = W*in
   wire signed [14:0] m231_96;
   assign m231_96 ={ {3{neg231[14]}} , neg231[14:3] };

   // m231_97 = W*in
   wire signed [14:0] m231_97;
   assign m231_97 =15'b0;

   // m231_98 = W*in
   wire signed [14:0] m231_98;
   assign m231_98 =15'b0;

   // m231_99 = W*in
   wire signed [14:0] m231_99;
   assign m231_99 =15'b0;

   // m231_100 = W*in
   wire signed [14:0] m231_100;
   assign m231_100 ={ {3{in231[14]}} , in231[14:3] };

   // m232_1 = W*in
   wire signed [14:0] m232_1;
   assign m232_1 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_2 = W*in
   wire signed [14:0] m232_2;
   assign m232_2 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_3 = W*in
   wire signed [14:0] m232_3;
   assign m232_3 ={ {3{in232[14]}} , in232[14:3] };

   // m232_4 = W*in
   wire signed [14:0] m232_4;
   assign m232_4 =15'b0;

   // m232_5 = W*in
   wire signed [14:0] m232_5;
   assign m232_5 ={ {4{neg232[14]}} , neg232[14:4] };

   // m232_6 = W*in
   wire signed [14:0] m232_6;
   assign m232_6 =15'b0;

   // m232_7 = W*in
   wire signed [14:0] m232_7;
   assign m232_7 =15'b0;

   // m232_8 = W*in
   wire signed [14:0] m232_8;
   assign m232_8 ={ {3{in232[14]}} , in232[14:3] };

   // m232_9 = W*in
   wire signed [14:0] m232_9;
   assign m232_9 =15'b0;

   // m232_10 = W*in
   wire signed [14:0] m232_10;
   assign m232_10 ={ {3{in232[14]}} , in232[14:3] };

   // m232_11 = W*in
   wire signed [14:0] m232_11;
   assign m232_11 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_12 = W*in
   wire signed [14:0] m232_12;
   assign m232_12 =15'b0;

   // m232_13 = W*in
   wire signed [14:0] m232_13;
   assign m232_13 =15'b0;

   // m232_14 = W*in
   wire signed [14:0] m232_14;
   assign m232_14 =15'b0;

   // m232_15 = W*in
   wire signed [14:0] m232_15;
   assign m232_15 ={ {3{in232[14]}} , in232[14:3] };

   // m232_16 = W*in
   wire signed [14:0] m232_16;
   assign m232_16 =15'b0;

   // m232_17 = W*in
   wire signed [14:0] m232_17;
   assign m232_17 =15'b0;

   // m232_18 = W*in
   wire signed [14:0] m232_18;
   assign m232_18 =15'b0;

   // m232_19 = W*in
   wire signed [14:0] m232_19;
   assign m232_19 =15'b0;

   // m232_20 = W*in
   wire signed [14:0] m232_20;
   assign m232_20 =15'b0;

   // m232_21 = W*in
   wire signed [14:0] m232_21;
   assign m232_21 ={ {4{neg232[14]}} , neg232[14:4] };

   // m232_22 = W*in
   wire signed [14:0] m232_22;
   assign m232_22 =15'b0;

   // m232_23 = W*in
   wire signed [14:0] m232_23;
   assign m232_23 =15'b0;

   // m232_24 = W*in
   wire signed [14:0] m232_24;
   assign m232_24 =15'b0;

   // m232_25 = W*in
   wire signed [14:0] m232_25;
   assign m232_25 ={ {4{neg232[14]}} , neg232[14:4] };

   // m232_26 = W*in
   wire signed [14:0] m232_26;
   assign m232_26 =15'b0;

   // m232_27 = W*in
   wire signed [14:0] m232_27;
   assign m232_27 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_28 = W*in
   wire signed [14:0] m232_28;
   assign m232_28 =15'b0;

   // m232_29 = W*in
   wire signed [14:0] m232_29;
   assign m232_29 =15'b0;

   // m232_30 = W*in
   wire signed [14:0] m232_30;
   assign m232_30 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_31 = W*in
   wire signed [14:0] m232_31;
   assign m232_31 =15'b0;

   // m232_32 = W*in
   wire signed [14:0] m232_32;
   assign m232_32 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_33 = W*in
   wire signed [14:0] m232_33;
   assign m232_33 =15'b0;

   // m232_34 = W*in
   wire signed [14:0] m232_34;
   assign m232_34 =15'b0;

   // m232_35 = W*in
   wire signed [14:0] m232_35;
   assign m232_35 =15'b0;

   // m232_36 = W*in
   wire signed [14:0] m232_36;
   assign m232_36 =15'b0;

   // m232_37 = W*in
   wire signed [14:0] m232_37;
   assign m232_37 =15'b0;

   // m232_38 = W*in
   wire signed [14:0] m232_38;
   assign m232_38 =15'b0;

   // m232_39 = W*in
   wire signed [14:0] m232_39;
   assign m232_39 =15'b0;

   // m232_40 = W*in
   wire signed [14:0] m232_40;
   assign m232_40 =15'b0;

   // m232_41 = W*in
   wire signed [14:0] m232_41;
   assign m232_41 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_42 = W*in
   wire signed [14:0] m232_42;
   assign m232_42 =15'b0;

   // m232_43 = W*in
   wire signed [14:0] m232_43;
   assign m232_43 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_44 = W*in
   wire signed [14:0] m232_44;
   assign m232_44 =15'b0;

   // m232_45 = W*in
   wire signed [14:0] m232_45;
   assign m232_45 =15'b0;

   // m232_46 = W*in
   wire signed [14:0] m232_46;
   assign m232_46 =15'b0;

   // m232_47 = W*in
   wire signed [14:0] m232_47;
   assign m232_47 =15'b0;

   // m232_48 = W*in
   wire signed [14:0] m232_48;
   assign m232_48 ={ {3{in232[14]}} , in232[14:3] };

   // m232_49 = W*in
   wire signed [14:0] m232_49;
   assign m232_49 ={ {3{in232[14]}} , in232[14:3] };

   // m232_50 = W*in
   wire signed [14:0] m232_50;
   assign m232_50 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_51 = W*in
   wire signed [14:0] m232_51;
   assign m232_51 =15'b0;

   // m232_52 = W*in
   wire signed [14:0] m232_52;
   assign m232_52 =15'b0;

   // m232_53 = W*in
   wire signed [14:0] m232_53;
   assign m232_53 ={ {3{in232[14]}} , in232[14:3] };

   // m232_54 = W*in
   wire signed [14:0] m232_54;
   assign m232_54 =15'b0;

   // m232_55 = W*in
   wire signed [14:0] m232_55;
   assign m232_55 =15'b0;

   // m232_56 = W*in
   wire signed [14:0] m232_56;
   assign m232_56 =15'b0;

   // m232_57 = W*in
   wire signed [14:0] m232_57;
   assign m232_57 =15'b0;

   // m232_58 = W*in
   wire signed [14:0] m232_58;
   assign m232_58 ={ {3{in232[14]}} , in232[14:3] };

   // m232_59 = W*in
   wire signed [14:0] m232_59;
   assign m232_59 =15'b0;

   // m232_60 = W*in
   wire signed [14:0] m232_60;
   assign m232_60 =15'b0;

   // m232_61 = W*in
   wire signed [14:0] m232_61;
   assign m232_61 ={ {3{in232[14]}} , in232[14:3] };

   // m232_62 = W*in
   wire signed [14:0] m232_62;
   assign m232_62 =15'b0;

   // m232_63 = W*in
   wire signed [14:0] m232_63;
   assign m232_63 ={ {2{in232[14]}} , in232[14:2] };

   // m232_64 = W*in
   wire signed [14:0] m232_64;
   assign m232_64 =15'b0;

   // m232_65 = W*in
   wire signed [14:0] m232_65;
   assign m232_65 =15'b0;

   // m232_66 = W*in
   wire signed [14:0] m232_66;
   assign m232_66 =15'b0;

   // m232_67 = W*in
   wire signed [14:0] m232_67;
   assign m232_67 =15'b0;

   // m232_68 = W*in
   wire signed [14:0] m232_68;
   assign m232_68 =15'b0;

   // m232_69 = W*in
   wire signed [14:0] m232_69;
   assign m232_69 =15'b0;

   // m232_70 = W*in
   wire signed [14:0] m232_70;
   assign m232_70 =15'b0;

   // m232_71 = W*in
   wire signed [14:0] m232_71;
   assign m232_71 ={ {3{in232[14]}} , in232[14:3] };

   // m232_72 = W*in
   wire signed [14:0] m232_72;
   assign m232_72 =15'b0;

   // m232_73 = W*in
   wire signed [14:0] m232_73;
   assign m232_73 =15'b0;

   // m232_74 = W*in
   wire signed [14:0] m232_74;
   assign m232_74 =15'b0;

   // m232_75 = W*in
   wire signed [14:0] m232_75;
   assign m232_75 =15'b0;

   // m232_76 = W*in
   wire signed [14:0] m232_76;
   assign m232_76 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_77 = W*in
   wire signed [14:0] m232_77;
   assign m232_77 =15'b0;

   // m232_78 = W*in
   wire signed [14:0] m232_78;
   assign m232_78 =15'b0;

   // m232_79 = W*in
   wire signed [14:0] m232_79;
   assign m232_79 =15'b0;

   // m232_80 = W*in
   wire signed [14:0] m232_80;
   assign m232_80 =15'b0;

   // m232_81 = W*in
   wire signed [14:0] m232_81;
   assign m232_81 =15'b0;

   // m232_82 = W*in
   wire signed [14:0] m232_82;
   assign m232_82 =15'b0;

   // m232_83 = W*in
   wire signed [14:0] m232_83;
   assign m232_83 =15'b0;

   // m232_84 = W*in
   wire signed [14:0] m232_84;
   assign m232_84 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_85 = W*in
   wire signed [14:0] m232_85;
   assign m232_85 =15'b0;

   // m232_86 = W*in
   wire signed [14:0] m232_86;
   assign m232_86 =15'b0;

   // m232_87 = W*in
   wire signed [14:0] m232_87;
   assign m232_87 =15'b0;

   // m232_88 = W*in
   wire signed [14:0] m232_88;
   assign m232_88 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_89 = W*in
   wire signed [14:0] m232_89;
   assign m232_89 =15'b0;

   // m232_90 = W*in
   wire signed [14:0] m232_90;
   assign m232_90 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_91 = W*in
   wire signed [14:0] m232_91;
   assign m232_91 ={ {3{in232[14]}} , in232[14:3] };

   // m232_92 = W*in
   wire signed [14:0] m232_92;
   assign m232_92 =15'b0;

   // m232_93 = W*in
   wire signed [14:0] m232_93;
   assign m232_93 =15'b0;

   // m232_94 = W*in
   wire signed [14:0] m232_94;
   assign m232_94 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_95 = W*in
   wire signed [14:0] m232_95;
   assign m232_95 ={ {3{neg232[14]}} , neg232[14:3] };

   // m232_96 = W*in
   wire signed [14:0] m232_96;
   assign m232_96 =15'b0;

   // m232_97 = W*in
   wire signed [14:0] m232_97;
   assign m232_97 =15'b0;

   // m232_98 = W*in
   wire signed [14:0] m232_98;
   assign m232_98 =15'b0;

   // m232_99 = W*in
   wire signed [14:0] m232_99;
   assign m232_99 =15'b0;

   // m232_100 = W*in
   wire signed [14:0] m232_100;
   assign m232_100 =15'b0;

   // m233_1 = W*in
   wire signed [14:0] m233_1;
   assign m233_1 =15'b0;

   // m233_2 = W*in
   wire signed [14:0] m233_2;
   assign m233_2 =15'b0;

   // m233_3 = W*in
   wire signed [14:0] m233_3;
   assign m233_3 =15'b0;

   // m233_4 = W*in
   wire signed [14:0] m233_4;
   assign m233_4 ={ {2{neg233[14]}} , neg233[14:2] };

   // m233_5 = W*in
   wire signed [14:0] m233_5;
   assign m233_5 =15'b0;

   // m233_6 = W*in
   wire signed [14:0] m233_6;
   assign m233_6 =15'b0;

   // m233_7 = W*in
   wire signed [14:0] m233_7;
   assign m233_7 =15'b0;

   // m233_8 = W*in
   wire signed [14:0] m233_8;
   assign m233_8 =15'b0;

   // m233_9 = W*in
   wire signed [14:0] m233_9;
   assign m233_9 ={ {3{in233[14]}} , in233[14:3] };

   // m233_10 = W*in
   wire signed [14:0] m233_10;
   assign m233_10 =15'b0;

   // m233_11 = W*in
   wire signed [14:0] m233_11;
   assign m233_11 =15'b0;

   // m233_12 = W*in
   wire signed [14:0] m233_12;
   assign m233_12 =15'b0;

   // m233_13 = W*in
   wire signed [14:0] m233_13;
   assign m233_13 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_14 = W*in
   wire signed [14:0] m233_14;
   assign m233_14 =15'b0;

   // m233_15 = W*in
   wire signed [14:0] m233_15;
   assign m233_15 =15'b0;

   // m233_16 = W*in
   wire signed [14:0] m233_16;
   assign m233_16 =15'b0;

   // m233_17 = W*in
   wire signed [14:0] m233_17;
   assign m233_17 =15'b0;

   // m233_18 = W*in
   wire signed [14:0] m233_18;
   assign m233_18 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_19 = W*in
   wire signed [14:0] m233_19;
   assign m233_19 =15'b0;

   // m233_20 = W*in
   wire signed [14:0] m233_20;
   assign m233_20 =15'b0;

   // m233_21 = W*in
   wire signed [14:0] m233_21;
   assign m233_21 ={ {4{neg233[14]}} , neg233[14:4] };

   // m233_22 = W*in
   wire signed [14:0] m233_22;
   assign m233_22 =15'b0;

   // m233_23 = W*in
   wire signed [14:0] m233_23;
   assign m233_23 =15'b0;

   // m233_24 = W*in
   wire signed [14:0] m233_24;
   assign m233_24 =15'b0;

   // m233_25 = W*in
   wire signed [14:0] m233_25;
   assign m233_25 =15'b0;

   // m233_26 = W*in
   wire signed [14:0] m233_26;
   assign m233_26 ={ {3{in233[14]}} , in233[14:3] };

   // m233_27 = W*in
   wire signed [14:0] m233_27;
   assign m233_27 =15'b0;

   // m233_28 = W*in
   wire signed [14:0] m233_28;
   assign m233_28 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_29 = W*in
   wire signed [14:0] m233_29;
   assign m233_29 =15'b0;

   // m233_30 = W*in
   wire signed [14:0] m233_30;
   assign m233_30 =15'b0;

   // m233_31 = W*in
   wire signed [14:0] m233_31;
   assign m233_31 ={ {3{in233[14]}} , in233[14:3] };

   // m233_32 = W*in
   wire signed [14:0] m233_32;
   assign m233_32 =15'b0;

   // m233_33 = W*in
   wire signed [14:0] m233_33;
   assign m233_33 =15'b0;

   // m233_34 = W*in
   wire signed [14:0] m233_34;
   assign m233_34 =15'b0;

   // m233_35 = W*in
   wire signed [14:0] m233_35;
   assign m233_35 ={ {3{in233[14]}} , in233[14:3] };

   // m233_36 = W*in
   wire signed [14:0] m233_36;
   assign m233_36 =15'b0;

   // m233_37 = W*in
   wire signed [14:0] m233_37;
   assign m233_37 =15'b0;

   // m233_38 = W*in
   wire signed [14:0] m233_38;
   assign m233_38 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_39 = W*in
   wire signed [14:0] m233_39;
   assign m233_39 =15'b0;

   // m233_40 = W*in
   wire signed [14:0] m233_40;
   assign m233_40 ={ {3{in233[14]}} , in233[14:3] };

   // m233_41 = W*in
   wire signed [14:0] m233_41;
   assign m233_41 =15'b0;

   // m233_42 = W*in
   wire signed [14:0] m233_42;
   assign m233_42 ={ {3{in233[14]}} , in233[14:3] };

   // m233_43 = W*in
   wire signed [14:0] m233_43;
   assign m233_43 =15'b0;

   // m233_44 = W*in
   wire signed [14:0] m233_44;
   assign m233_44 =15'b0;

   // m233_45 = W*in
   wire signed [14:0] m233_45;
   assign m233_45 =15'b0;

   // m233_46 = W*in
   wire signed [14:0] m233_46;
   assign m233_46 =15'b0;

   // m233_47 = W*in
   wire signed [14:0] m233_47;
   assign m233_47 ={ {3{in233[14]}} , in233[14:3] };

   // m233_48 = W*in
   wire signed [14:0] m233_48;
   assign m233_48 ={ {3{in233[14]}} , in233[14:3] };

   // m233_49 = W*in
   wire signed [14:0] m233_49;
   assign m233_49 =15'b0;

   // m233_50 = W*in
   wire signed [14:0] m233_50;
   assign m233_50 =15'b0;

   // m233_51 = W*in
   wire signed [14:0] m233_51;
   assign m233_51 ={ {3{in233[14]}} , in233[14:3] };

   // m233_52 = W*in
   wire signed [14:0] m233_52;
   assign m233_52 =15'b0;

   // m233_53 = W*in
   wire signed [14:0] m233_53;
   assign m233_53 =15'b0;

   // m233_54 = W*in
   wire signed [14:0] m233_54;
   assign m233_54 =15'b0;

   // m233_55 = W*in
   wire signed [14:0] m233_55;
   assign m233_55 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_56 = W*in
   wire signed [14:0] m233_56;
   assign m233_56 =15'b0;

   // m233_57 = W*in
   wire signed [14:0] m233_57;
   assign m233_57 ={ {3{in233[14]}} , in233[14:3] };

   // m233_58 = W*in
   wire signed [14:0] m233_58;
   assign m233_58 =15'b0;

   // m233_59 = W*in
   wire signed [14:0] m233_59;
   assign m233_59 =15'b0;

   // m233_60 = W*in
   wire signed [14:0] m233_60;
   assign m233_60 =15'b0;

   // m233_61 = W*in
   wire signed [14:0] m233_61;
   assign m233_61 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_62 = W*in
   wire signed [14:0] m233_62;
   assign m233_62 =15'b0;

   // m233_63 = W*in
   wire signed [14:0] m233_63;
   assign m233_63 =15'b0;

   // m233_64 = W*in
   wire signed [14:0] m233_64;
   assign m233_64 =15'b0;

   // m233_65 = W*in
   wire signed [14:0] m233_65;
   assign m233_65 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_66 = W*in
   wire signed [14:0] m233_66;
   assign m233_66 ={ {3{in233[14]}} , in233[14:3] };

   // m233_67 = W*in
   wire signed [14:0] m233_67;
   assign m233_67 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_68 = W*in
   wire signed [14:0] m233_68;
   assign m233_68 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_69 = W*in
   wire signed [14:0] m233_69;
   assign m233_69 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_70 = W*in
   wire signed [14:0] m233_70;
   assign m233_70 ={ {3{in233[14]}} , in233[14:3] };

   // m233_71 = W*in
   wire signed [14:0] m233_71;
   assign m233_71 =15'b0;

   // m233_72 = W*in
   wire signed [14:0] m233_72;
   assign m233_72 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_73 = W*in
   wire signed [14:0] m233_73;
   assign m233_73 =15'b0;

   // m233_74 = W*in
   wire signed [14:0] m233_74;
   assign m233_74 ={ {4{in233[14]}} , in233[14:4] };

   // m233_75 = W*in
   wire signed [14:0] m233_75;
   assign m233_75 =15'b0;

   // m233_76 = W*in
   wire signed [14:0] m233_76;
   assign m233_76 =15'b0;

   // m233_77 = W*in
   wire signed [14:0] m233_77;
   assign m233_77 =15'b0;

   // m233_78 = W*in
   wire signed [14:0] m233_78;
   assign m233_78 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_79 = W*in
   wire signed [14:0] m233_79;
   assign m233_79 ={ {3{in233[14]}} , in233[14:3] };

   // m233_80 = W*in
   wire signed [14:0] m233_80;
   assign m233_80 =15'b0;

   // m233_81 = W*in
   wire signed [14:0] m233_81;
   assign m233_81 =15'b0;

   // m233_82 = W*in
   wire signed [14:0] m233_82;
   assign m233_82 =15'b0;

   // m233_83 = W*in
   wire signed [14:0] m233_83;
   assign m233_83 =15'b0;

   // m233_84 = W*in
   wire signed [14:0] m233_84;
   assign m233_84 =15'b0;

   // m233_85 = W*in
   wire signed [14:0] m233_85;
   assign m233_85 =15'b0;

   // m233_86 = W*in
   wire signed [14:0] m233_86;
   assign m233_86 =15'b0;

   // m233_87 = W*in
   wire signed [14:0] m233_87;
   assign m233_87 =15'b0;

   // m233_88 = W*in
   wire signed [14:0] m233_88;
   assign m233_88 =15'b0;

   // m233_89 = W*in
   wire signed [14:0] m233_89;
   assign m233_89 =15'b0;

   // m233_90 = W*in
   wire signed [14:0] m233_90;
   assign m233_90 =15'b0;

   // m233_91 = W*in
   wire signed [14:0] m233_91;
   assign m233_91 ={ {3{in233[14]}} , in233[14:3] };

   // m233_92 = W*in
   wire signed [14:0] m233_92;
   assign m233_92 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_93 = W*in
   wire signed [14:0] m233_93;
   assign m233_93 =15'b0;

   // m233_94 = W*in
   wire signed [14:0] m233_94;
   assign m233_94 ={ {4{in233[14]}} , in233[14:4] };

   // m233_95 = W*in
   wire signed [14:0] m233_95;
   assign m233_95 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_96 = W*in
   wire signed [14:0] m233_96;
   assign m233_96 =15'b0;

   // m233_97 = W*in
   wire signed [14:0] m233_97;
   assign m233_97 ={ {3{neg233[14]}} , neg233[14:3] };

   // m233_98 = W*in
   wire signed [14:0] m233_98;
   assign m233_98 =15'b0;

   // m233_99 = W*in
   wire signed [14:0] m233_99;
   assign m233_99 ={ {4{neg233[14]}} , neg233[14:4] };

   // m233_100 = W*in
   wire signed [14:0] m233_100;
   assign m233_100 ={ {3{in233[14]}} , in233[14:3] };

   // m234_1 = W*in
   wire signed [14:0] m234_1;
   assign m234_1 =15'b0;

   // m234_2 = W*in
   wire signed [14:0] m234_2;
   assign m234_2 =15'b0;

   // m234_3 = W*in
   wire signed [14:0] m234_3;
   assign m234_3 =15'b0;

   // m234_4 = W*in
   wire signed [14:0] m234_4;
   assign m234_4 =15'b0;

   // m234_5 = W*in
   wire signed [14:0] m234_5;
   assign m234_5 ={ {4{neg234[14]}} , neg234[14:4] };

   // m234_6 = W*in
   wire signed [14:0] m234_6;
   assign m234_6 =15'b0;

   // m234_7 = W*in
   wire signed [14:0] m234_7;
   assign m234_7 =15'b0;

   // m234_8 = W*in
   wire signed [14:0] m234_8;
   assign m234_8 =15'b0;

   // m234_9 = W*in
   wire signed [14:0] m234_9;
   assign m234_9 ={ {3{in234[14]}} , in234[14:3] };

   // m234_10 = W*in
   wire signed [14:0] m234_10;
   assign m234_10 =15'b0;

   // m234_11 = W*in
   wire signed [14:0] m234_11;
   assign m234_11 =15'b0;

   // m234_12 = W*in
   wire signed [14:0] m234_12;
   assign m234_12 =15'b0;

   // m234_13 = W*in
   wire signed [14:0] m234_13;
   assign m234_13 =15'b0;

   // m234_14 = W*in
   wire signed [14:0] m234_14;
   assign m234_14 =15'b0;

   // m234_15 = W*in
   wire signed [14:0] m234_15;
   assign m234_15 =15'b0;

   // m234_16 = W*in
   wire signed [14:0] m234_16;
   assign m234_16 ={ {4{in234[14]}} , in234[14:4] };

   // m234_17 = W*in
   wire signed [14:0] m234_17;
   assign m234_17 =15'b0;

   // m234_18 = W*in
   wire signed [14:0] m234_18;
   assign m234_18 =15'b0;

   // m234_19 = W*in
   wire signed [14:0] m234_19;
   assign m234_19 =15'b0;

   // m234_20 = W*in
   wire signed [14:0] m234_20;
   assign m234_20 =15'b0;

   // m234_21 = W*in
   wire signed [14:0] m234_21;
   assign m234_21 ={ {4{neg234[14]}} , neg234[14:4] };

   // m234_22 = W*in
   wire signed [14:0] m234_22;
   assign m234_22 =15'b0;

   // m234_23 = W*in
   wire signed [14:0] m234_23;
   assign m234_23 =15'b0;

   // m234_24 = W*in
   wire signed [14:0] m234_24;
   assign m234_24 ={ {3{in234[14]}} , in234[14:3] };

   // m234_25 = W*in
   wire signed [14:0] m234_25;
   assign m234_25 ={ {4{neg234[14]}} , neg234[14:4] };

   // m234_26 = W*in
   wire signed [14:0] m234_26;
   assign m234_26 =15'b0;

   // m234_27 = W*in
   wire signed [14:0] m234_27;
   assign m234_27 =15'b0;

   // m234_28 = W*in
   wire signed [14:0] m234_28;
   assign m234_28 =15'b0;

   // m234_29 = W*in
   wire signed [14:0] m234_29;
   assign m234_29 =15'b0;

   // m234_30 = W*in
   wire signed [14:0] m234_30;
   assign m234_30 =15'b0;

   // m234_31 = W*in
   wire signed [14:0] m234_31;
   assign m234_31 ={ {3{in234[14]}} , in234[14:3] };

   // m234_32 = W*in
   wire signed [14:0] m234_32;
   assign m234_32 ={ {3{in234[14]}} , in234[14:3] };

   // m234_33 = W*in
   wire signed [14:0] m234_33;
   assign m234_33 =15'b0;

   // m234_34 = W*in
   wire signed [14:0] m234_34;
   assign m234_34 =15'b0;

   // m234_35 = W*in
   wire signed [14:0] m234_35;
   assign m234_35 ={ {3{in234[14]}} , in234[14:3] };

   // m234_36 = W*in
   wire signed [14:0] m234_36;
   assign m234_36 =15'b0;

   // m234_37 = W*in
   wire signed [14:0] m234_37;
   assign m234_37 =15'b0;

   // m234_38 = W*in
   wire signed [14:0] m234_38;
   assign m234_38 =15'b0;

   // m234_39 = W*in
   wire signed [14:0] m234_39;
   assign m234_39 =15'b0;

   // m234_40 = W*in
   wire signed [14:0] m234_40;
   assign m234_40 ={ {3{in234[14]}} , in234[14:3] };

   // m234_41 = W*in
   wire signed [14:0] m234_41;
   assign m234_41 =15'b0;

   // m234_42 = W*in
   wire signed [14:0] m234_42;
   assign m234_42 =15'b0;

   // m234_43 = W*in
   wire signed [14:0] m234_43;
   assign m234_43 =15'b0;

   // m234_44 = W*in
   wire signed [14:0] m234_44;
   assign m234_44 =15'b0;

   // m234_45 = W*in
   wire signed [14:0] m234_45;
   assign m234_45 =15'b0;

   // m234_46 = W*in
   wire signed [14:0] m234_46;
   assign m234_46 =15'b0;

   // m234_47 = W*in
   wire signed [14:0] m234_47;
   assign m234_47 ={ {3{in234[14]}} , in234[14:3] };

   // m234_48 = W*in
   wire signed [14:0] m234_48;
   assign m234_48 =15'b0;

   // m234_49 = W*in
   wire signed [14:0] m234_49;
   assign m234_49 =15'b0;

   // m234_50 = W*in
   wire signed [14:0] m234_50;
   assign m234_50 =15'b0;

   // m234_51 = W*in
   wire signed [14:0] m234_51;
   assign m234_51 =15'b0;

   // m234_52 = W*in
   wire signed [14:0] m234_52;
   assign m234_52 ={ {3{neg234[14]}} , neg234[14:3] };

   // m234_53 = W*in
   wire signed [14:0] m234_53;
   assign m234_53 ={ {3{neg234[14]}} , neg234[14:3] };

   // m234_54 = W*in
   wire signed [14:0] m234_54;
   assign m234_54 =15'b0;

   // m234_55 = W*in
   wire signed [14:0] m234_55;
   assign m234_55 =15'b0;

   // m234_56 = W*in
   wire signed [14:0] m234_56;
   assign m234_56 =15'b0;

   // m234_57 = W*in
   wire signed [14:0] m234_57;
   assign m234_57 =15'b0;

   // m234_58 = W*in
   wire signed [14:0] m234_58;
   assign m234_58 =15'b0;

   // m234_59 = W*in
   wire signed [14:0] m234_59;
   assign m234_59 =15'b0;

   // m234_60 = W*in
   wire signed [14:0] m234_60;
   assign m234_60 =15'b0;

   // m234_61 = W*in
   wire signed [14:0] m234_61;
   assign m234_61 =15'b0;

   // m234_62 = W*in
   wire signed [14:0] m234_62;
   assign m234_62 =15'b0;

   // m234_63 = W*in
   wire signed [14:0] m234_63;
   assign m234_63 =15'b0;

   // m234_64 = W*in
   wire signed [14:0] m234_64;
   assign m234_64 ={ {3{neg234[14]}} , neg234[14:3] };

   // m234_65 = W*in
   wire signed [14:0] m234_65;
   assign m234_65 =15'b0;

   // m234_66 = W*in
   wire signed [14:0] m234_66;
   assign m234_66 =15'b0;

   // m234_67 = W*in
   wire signed [14:0] m234_67;
   assign m234_67 =15'b0;

   // m234_68 = W*in
   wire signed [14:0] m234_68;
   assign m234_68 =15'b0;

   // m234_69 = W*in
   wire signed [14:0] m234_69;
   assign m234_69 =15'b0;

   // m234_70 = W*in
   wire signed [14:0] m234_70;
   assign m234_70 ={ {3{in234[14]}} , in234[14:3] };

   // m234_71 = W*in
   wire signed [14:0] m234_71;
   assign m234_71 =15'b0;

   // m234_72 = W*in
   wire signed [14:0] m234_72;
   assign m234_72 =15'b0;

   // m234_73 = W*in
   wire signed [14:0] m234_73;
   assign m234_73 =15'b0;

   // m234_74 = W*in
   wire signed [14:0] m234_74;
   assign m234_74 ={ {3{in234[14]}} , in234[14:3] };

   // m234_75 = W*in
   wire signed [14:0] m234_75;
   assign m234_75 =15'b0;

   // m234_76 = W*in
   wire signed [14:0] m234_76;
   assign m234_76 =15'b0;

   // m234_77 = W*in
   wire signed [14:0] m234_77;
   assign m234_77 =15'b0;

   // m234_78 = W*in
   wire signed [14:0] m234_78;
   assign m234_78 ={ {3{neg234[14]}} , neg234[14:3] };

   // m234_79 = W*in
   wire signed [14:0] m234_79;
   assign m234_79 =15'b0;

   // m234_80 = W*in
   wire signed [14:0] m234_80;
   assign m234_80 =15'b0;

   // m234_81 = W*in
   wire signed [14:0] m234_81;
   assign m234_81 =15'b0;

   // m234_82 = W*in
   wire signed [14:0] m234_82;
   assign m234_82 =15'b0;

   // m234_83 = W*in
   wire signed [14:0] m234_83;
   assign m234_83 =15'b0;

   // m234_84 = W*in
   wire signed [14:0] m234_84;
   assign m234_84 =15'b0;

   // m234_85 = W*in
   wire signed [14:0] m234_85;
   assign m234_85 =15'b0;

   // m234_86 = W*in
   wire signed [14:0] m234_86;
   assign m234_86 =15'b0;

   // m234_87 = W*in
   wire signed [14:0] m234_87;
   assign m234_87 =15'b0;

   // m234_88 = W*in
   wire signed [14:0] m234_88;
   assign m234_88 =15'b0;

   // m234_89 = W*in
   wire signed [14:0] m234_89;
   assign m234_89 =15'b0;

   // m234_90 = W*in
   wire signed [14:0] m234_90;
   assign m234_90 ={ {3{neg234[14]}} , neg234[14:3] };

   // m234_91 = W*in
   wire signed [14:0] m234_91;
   assign m234_91 =15'b0;

   // m234_92 = W*in
   wire signed [14:0] m234_92;
   assign m234_92 =15'b0;

   // m234_93 = W*in
   wire signed [14:0] m234_93;
   assign m234_93 =15'b0;

   // m234_94 = W*in
   wire signed [14:0] m234_94;
   assign m234_94 =15'b0;

   // m234_95 = W*in
   wire signed [14:0] m234_95;
   assign m234_95 =15'b0;

   // m234_96 = W*in
   wire signed [14:0] m234_96;
   assign m234_96 =15'b0;

   // m234_97 = W*in
   wire signed [14:0] m234_97;
   assign m234_97 =15'b0;

   // m234_98 = W*in
   wire signed [14:0] m234_98;
   assign m234_98 =15'b0;

   // m234_99 = W*in
   wire signed [14:0] m234_99;
   assign m234_99 =15'b0;

   // m234_100 = W*in
   wire signed [14:0] m234_100;
   assign m234_100 =15'b0;

   // m235_1 = W*in
   wire signed [14:0] m235_1;
   assign m235_1 =15'b0;

   // m235_2 = W*in
   wire signed [14:0] m235_2;
   assign m235_2 =15'b0;

   // m235_3 = W*in
   wire signed [14:0] m235_3;
   assign m235_3 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_4 = W*in
   wire signed [14:0] m235_4;
   assign m235_4 ={ {3{in235[14]}} , in235[14:3] };

   // m235_5 = W*in
   wire signed [14:0] m235_5;
   assign m235_5 =15'b0;

   // m235_6 = W*in
   wire signed [14:0] m235_6;
   assign m235_6 =15'b0;

   // m235_7 = W*in
   wire signed [14:0] m235_7;
   assign m235_7 =15'b0;

   // m235_8 = W*in
   wire signed [14:0] m235_8;
   assign m235_8 =15'b0;

   // m235_9 = W*in
   wire signed [14:0] m235_9;
   assign m235_9 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_10 = W*in
   wire signed [14:0] m235_10;
   assign m235_10 =15'b0;

   // m235_11 = W*in
   wire signed [14:0] m235_11;
   assign m235_11 =15'b0;

   // m235_12 = W*in
   wire signed [14:0] m235_12;
   assign m235_12 =15'b0;

   // m235_13 = W*in
   wire signed [14:0] m235_13;
   assign m235_13 =15'b0;

   // m235_14 = W*in
   wire signed [14:0] m235_14;
   assign m235_14 =15'b0;

   // m235_15 = W*in
   wire signed [14:0] m235_15;
   assign m235_15 ={ {2{in235[14]}} , in235[14:2] };

   // m235_16 = W*in
   wire signed [14:0] m235_16;
   assign m235_16 =15'b0;

   // m235_17 = W*in
   wire signed [14:0] m235_17;
   assign m235_17 =15'b0;

   // m235_18 = W*in
   wire signed [14:0] m235_18;
   assign m235_18 ={ {4{in235[14]}} , in235[14:4] };

   // m235_19 = W*in
   wire signed [14:0] m235_19;
   assign m235_19 =15'b0;

   // m235_20 = W*in
   wire signed [14:0] m235_20;
   assign m235_20 ={ {4{neg235[14]}} , neg235[14:4] };

   // m235_21 = W*in
   wire signed [14:0] m235_21;
   assign m235_21 ={ {4{in235[14]}} , in235[14:4] };

   // m235_22 = W*in
   wire signed [14:0] m235_22;
   assign m235_22 ={ {2{neg235[14]}} , neg235[14:2] };

   // m235_23 = W*in
   wire signed [14:0] m235_23;
   assign m235_23 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_24 = W*in
   wire signed [14:0] m235_24;
   assign m235_24 =15'b0;

   // m235_25 = W*in
   wire signed [14:0] m235_25;
   assign m235_25 ={ {4{neg235[14]}} , neg235[14:4] };

   // m235_26 = W*in
   wire signed [14:0] m235_26;
   assign m235_26 =15'b0;

   // m235_27 = W*in
   wire signed [14:0] m235_27;
   assign m235_27 =15'b0;

   // m235_28 = W*in
   wire signed [14:0] m235_28;
   assign m235_28 ={ {3{in235[14]}} , in235[14:3] };

   // m235_29 = W*in
   wire signed [14:0] m235_29;
   assign m235_29 =15'b0;

   // m235_30 = W*in
   wire signed [14:0] m235_30;
   assign m235_30 ={ {3{in235[14]}} , in235[14:3] };

   // m235_31 = W*in
   wire signed [14:0] m235_31;
   assign m235_31 =15'b0;

   // m235_32 = W*in
   wire signed [14:0] m235_32;
   assign m235_32 =15'b0;

   // m235_33 = W*in
   wire signed [14:0] m235_33;
   assign m235_33 =15'b0;

   // m235_34 = W*in
   wire signed [14:0] m235_34;
   assign m235_34 =15'b0;

   // m235_35 = W*in
   wire signed [14:0] m235_35;
   assign m235_35 =15'b0;

   // m235_36 = W*in
   wire signed [14:0] m235_36;
   assign m235_36 =15'b0;

   // m235_37 = W*in
   wire signed [14:0] m235_37;
   assign m235_37 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_38 = W*in
   wire signed [14:0] m235_38;
   assign m235_38 =15'b0;

   // m235_39 = W*in
   wire signed [14:0] m235_39;
   assign m235_39 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_40 = W*in
   wire signed [14:0] m235_40;
   assign m235_40 =15'b0;

   // m235_41 = W*in
   wire signed [14:0] m235_41;
   assign m235_41 =15'b0;

   // m235_42 = W*in
   wire signed [14:0] m235_42;
   assign m235_42 =15'b0;

   // m235_43 = W*in
   wire signed [14:0] m235_43;
   assign m235_43 =15'b0;

   // m235_44 = W*in
   wire signed [14:0] m235_44;
   assign m235_44 =15'b0;

   // m235_45 = W*in
   wire signed [14:0] m235_45;
   assign m235_45 =15'b0;

   // m235_46 = W*in
   wire signed [14:0] m235_46;
   assign m235_46 =15'b0;

   // m235_47 = W*in
   wire signed [14:0] m235_47;
   assign m235_47 =15'b0;

   // m235_48 = W*in
   wire signed [14:0] m235_48;
   assign m235_48 ={ {2{in235[14]}} , in235[14:2] };

   // m235_49 = W*in
   wire signed [14:0] m235_49;
   assign m235_49 ={ {3{in235[14]}} , in235[14:3] };

   // m235_50 = W*in
   wire signed [14:0] m235_50;
   assign m235_50 =15'b0;

   // m235_51 = W*in
   wire signed [14:0] m235_51;
   assign m235_51 =15'b0;

   // m235_52 = W*in
   wire signed [14:0] m235_52;
   assign m235_52 =15'b0;

   // m235_53 = W*in
   wire signed [14:0] m235_53;
   assign m235_53 =15'b0;

   // m235_54 = W*in
   wire signed [14:0] m235_54;
   assign m235_54 =15'b0;

   // m235_55 = W*in
   wire signed [14:0] m235_55;
   assign m235_55 =15'b0;

   // m235_56 = W*in
   wire signed [14:0] m235_56;
   assign m235_56 =15'b0;

   // m235_57 = W*in
   wire signed [14:0] m235_57;
   assign m235_57 =15'b0;

   // m235_58 = W*in
   wire signed [14:0] m235_58;
   assign m235_58 =15'b0;

   // m235_59 = W*in
   wire signed [14:0] m235_59;
   assign m235_59 =15'b0;

   // m235_60 = W*in
   wire signed [14:0] m235_60;
   assign m235_60 =15'b0;

   // m235_61 = W*in
   wire signed [14:0] m235_61;
   assign m235_61 ={ {3{in235[14]}} , in235[14:3] };

   // m235_62 = W*in
   wire signed [14:0] m235_62;
   assign m235_62 =15'b0;

   // m235_63 = W*in
   wire signed [14:0] m235_63;
   assign m235_63 =15'b0;

   // m235_64 = W*in
   wire signed [14:0] m235_64;
   assign m235_64 =15'b0;

   // m235_65 = W*in
   wire signed [14:0] m235_65;
   assign m235_65 ={ {3{in235[14]}} , in235[14:3] };

   // m235_66 = W*in
   wire signed [14:0] m235_66;
   assign m235_66 =15'b0;

   // m235_67 = W*in
   wire signed [14:0] m235_67;
   assign m235_67 ={ {2{in235[14]}} , in235[14:2] };

   // m235_68 = W*in
   wire signed [14:0] m235_68;
   assign m235_68 =15'b0;

   // m235_69 = W*in
   wire signed [14:0] m235_69;
   assign m235_69 ={ {4{in235[14]}} , in235[14:4] };

   // m235_70 = W*in
   wire signed [14:0] m235_70;
   assign m235_70 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_71 = W*in
   wire signed [14:0] m235_71;
   assign m235_71 =15'b0;

   // m235_72 = W*in
   wire signed [14:0] m235_72;
   assign m235_72 =15'b0;

   // m235_73 = W*in
   wire signed [14:0] m235_73;
   assign m235_73 =15'b0;

   // m235_74 = W*in
   wire signed [14:0] m235_74;
   assign m235_74 ={ {4{neg235[14]}} , neg235[14:4] };

   // m235_75 = W*in
   wire signed [14:0] m235_75;
   assign m235_75 =15'b0;

   // m235_76 = W*in
   wire signed [14:0] m235_76;
   assign m235_76 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_77 = W*in
   wire signed [14:0] m235_77;
   assign m235_77 =15'b0;

   // m235_78 = W*in
   wire signed [14:0] m235_78;
   assign m235_78 ={ {3{in235[14]}} , in235[14:3] };

   // m235_79 = W*in
   wire signed [14:0] m235_79;
   assign m235_79 =15'b0;

   // m235_80 = W*in
   wire signed [14:0] m235_80;
   assign m235_80 =15'b0;

   // m235_81 = W*in
   wire signed [14:0] m235_81;
   assign m235_81 ={ {3{in235[14]}} , in235[14:3] };

   // m235_82 = W*in
   wire signed [14:0] m235_82;
   assign m235_82 =15'b0;

   // m235_83 = W*in
   wire signed [14:0] m235_83;
   assign m235_83 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_84 = W*in
   wire signed [14:0] m235_84;
   assign m235_84 ={ {3{in235[14]}} , in235[14:3] };

   // m235_85 = W*in
   wire signed [14:0] m235_85;
   assign m235_85 =15'b0;

   // m235_86 = W*in
   wire signed [14:0] m235_86;
   assign m235_86 =15'b0;

   // m235_87 = W*in
   wire signed [14:0] m235_87;
   assign m235_87 =15'b0;

   // m235_88 = W*in
   wire signed [14:0] m235_88;
   assign m235_88 =15'b0;

   // m235_89 = W*in
   wire signed [14:0] m235_89;
   assign m235_89 =15'b0;

   // m235_90 = W*in
   wire signed [14:0] m235_90;
   assign m235_90 =15'b0;

   // m235_91 = W*in
   wire signed [14:0] m235_91;
   assign m235_91 =15'b0;

   // m235_92 = W*in
   wire signed [14:0] m235_92;
   assign m235_92 ={ {4{in235[14]}} , in235[14:4] };

   // m235_93 = W*in
   wire signed [14:0] m235_93;
   assign m235_93 =15'b0;

   // m235_94 = W*in
   wire signed [14:0] m235_94;
   assign m235_94 ={ {3{neg235[14]}} , neg235[14:3] };

   // m235_95 = W*in
   wire signed [14:0] m235_95;
   assign m235_95 =15'b0;

   // m235_96 = W*in
   wire signed [14:0] m235_96;
   assign m235_96 =15'b0;

   // m235_97 = W*in
   wire signed [14:0] m235_97;
   assign m235_97 =15'b0;

   // m235_98 = W*in
   wire signed [14:0] m235_98;
   assign m235_98 ={ {3{in235[14]}} , in235[14:3] };

   // m235_99 = W*in
   wire signed [14:0] m235_99;
   assign m235_99 =15'b0;

   // m235_100 = W*in
   wire signed [14:0] m235_100;
   assign m235_100 ={ {3{neg235[14]}} , neg235[14:3] };

   // m236_1 = W*in
   wire signed [14:0] m236_1;
   assign m236_1 =15'b0;

   // m236_2 = W*in
   wire signed [14:0] m236_2;
   assign m236_2 =15'b0;

   // m236_3 = W*in
   wire signed [14:0] m236_3;
   assign m236_3 =15'b0;

   // m236_4 = W*in
   wire signed [14:0] m236_4;
   assign m236_4 =15'b0;

   // m236_5 = W*in
   wire signed [14:0] m236_5;
   assign m236_5 =15'b0;

   // m236_6 = W*in
   wire signed [14:0] m236_6;
   assign m236_6 =15'b0;

   // m236_7 = W*in
   wire signed [14:0] m236_7;
   assign m236_7 =15'b0;

   // m236_8 = W*in
   wire signed [14:0] m236_8;
   assign m236_8 =15'b0;

   // m236_9 = W*in
   wire signed [14:0] m236_9;
   assign m236_9 =15'b0;

   // m236_10 = W*in
   wire signed [14:0] m236_10;
   assign m236_10 ={ {4{neg236[14]}} , neg236[14:4] };

   // m236_11 = W*in
   wire signed [14:0] m236_11;
   assign m236_11 =15'b0;

   // m236_12 = W*in
   wire signed [14:0] m236_12;
   assign m236_12 =15'b0;

   // m236_13 = W*in
   wire signed [14:0] m236_13;
   assign m236_13 =15'b0;

   // m236_14 = W*in
   wire signed [14:0] m236_14;
   assign m236_14 =15'b0;

   // m236_15 = W*in
   wire signed [14:0] m236_15;
   assign m236_15 =15'b0;

   // m236_16 = W*in
   wire signed [14:0] m236_16;
   assign m236_16 =15'b0;

   // m236_17 = W*in
   wire signed [14:0] m236_17;
   assign m236_17 =15'b0;

   // m236_18 = W*in
   wire signed [14:0] m236_18;
   assign m236_18 =15'b0;

   // m236_19 = W*in
   wire signed [14:0] m236_19;
   assign m236_19 =15'b0;

   // m236_20 = W*in
   wire signed [14:0] m236_20;
   assign m236_20 ={ {3{in236[14]}} , in236[14:3] };

   // m236_21 = W*in
   wire signed [14:0] m236_21;
   assign m236_21 ={ {3{in236[14]}} , in236[14:3] };

   // m236_22 = W*in
   wire signed [14:0] m236_22;
   assign m236_22 =15'b0;

   // m236_23 = W*in
   wire signed [14:0] m236_23;
   assign m236_23 =15'b0;

   // m236_24 = W*in
   wire signed [14:0] m236_24;
   assign m236_24 =15'b0;

   // m236_25 = W*in
   wire signed [14:0] m236_25;
   assign m236_25 =15'b0;

   // m236_26 = W*in
   wire signed [14:0] m236_26;
   assign m236_26 =15'b0;

   // m236_27 = W*in
   wire signed [14:0] m236_27;
   assign m236_27 =15'b0;

   // m236_28 = W*in
   wire signed [14:0] m236_28;
   assign m236_28 =15'b0;

   // m236_29 = W*in
   wire signed [14:0] m236_29;
   assign m236_29 =15'b0;

   // m236_30 = W*in
   wire signed [14:0] m236_30;
   assign m236_30 =15'b0;

   // m236_31 = W*in
   wire signed [14:0] m236_31;
   assign m236_31 =15'b0;

   // m236_32 = W*in
   wire signed [14:0] m236_32;
   assign m236_32 =15'b0;

   // m236_33 = W*in
   wire signed [14:0] m236_33;
   assign m236_33 =15'b0;

   // m236_34 = W*in
   wire signed [14:0] m236_34;
   assign m236_34 =15'b0;

   // m236_35 = W*in
   wire signed [14:0] m236_35;
   assign m236_35 =15'b0;

   // m236_36 = W*in
   wire signed [14:0] m236_36;
   assign m236_36 =15'b0;

   // m236_37 = W*in
   wire signed [14:0] m236_37;
   assign m236_37 =15'b0;

   // m236_38 = W*in
   wire signed [14:0] m236_38;
   assign m236_38 =15'b0;

   // m236_39 = W*in
   wire signed [14:0] m236_39;
   assign m236_39 =15'b0;

   // m236_40 = W*in
   wire signed [14:0] m236_40;
   assign m236_40 =15'b0;

   // m236_41 = W*in
   wire signed [14:0] m236_41;
   assign m236_41 =15'b0;

   // m236_42 = W*in
   wire signed [14:0] m236_42;
   assign m236_42 =15'b0;

   // m236_43 = W*in
   wire signed [14:0] m236_43;
   assign m236_43 ={ {3{in236[14]}} , in236[14:3] };

   // m236_44 = W*in
   wire signed [14:0] m236_44;
   assign m236_44 =15'b0;

   // m236_45 = W*in
   wire signed [14:0] m236_45;
   assign m236_45 =15'b0;

   // m236_46 = W*in
   wire signed [14:0] m236_46;
   assign m236_46 =15'b0;

   // m236_47 = W*in
   wire signed [14:0] m236_47;
   assign m236_47 =15'b0;

   // m236_48 = W*in
   wire signed [14:0] m236_48;
   assign m236_48 =15'b0;

   // m236_49 = W*in
   wire signed [14:0] m236_49;
   assign m236_49 =15'b0;

   // m236_50 = W*in
   wire signed [14:0] m236_50;
   assign m236_50 ={ {3{neg236[14]}} , neg236[14:3] };

   // m236_51 = W*in
   wire signed [14:0] m236_51;
   assign m236_51 =15'b0;

   // m236_52 = W*in
   wire signed [14:0] m236_52;
   assign m236_52 =15'b0;

   // m236_53 = W*in
   wire signed [14:0] m236_53;
   assign m236_53 =15'b0;

   // m236_54 = W*in
   wire signed [14:0] m236_54;
   assign m236_54 =15'b0;

   // m236_55 = W*in
   wire signed [14:0] m236_55;
   assign m236_55 =15'b0;

   // m236_56 = W*in
   wire signed [14:0] m236_56;
   assign m236_56 =15'b0;

   // m236_57 = W*in
   wire signed [14:0] m236_57;
   assign m236_57 =15'b0;

   // m236_58 = W*in
   wire signed [14:0] m236_58;
   assign m236_58 =15'b0;

   // m236_59 = W*in
   wire signed [14:0] m236_59;
   assign m236_59 ={ {3{in236[14]}} , in236[14:3] };

   // m236_60 = W*in
   wire signed [14:0] m236_60;
   assign m236_60 =15'b0;

   // m236_61 = W*in
   wire signed [14:0] m236_61;
   assign m236_61 =15'b0;

   // m236_62 = W*in
   wire signed [14:0] m236_62;
   assign m236_62 ={ {3{in236[14]}} , in236[14:3] };

   // m236_63 = W*in
   wire signed [14:0] m236_63;
   assign m236_63 =15'b0;

   // m236_64 = W*in
   wire signed [14:0] m236_64;
   assign m236_64 =15'b0;

   // m236_65 = W*in
   wire signed [14:0] m236_65;
   assign m236_65 =15'b0;

   // m236_66 = W*in
   wire signed [14:0] m236_66;
   assign m236_66 =15'b0;

   // m236_67 = W*in
   wire signed [14:0] m236_67;
   assign m236_67 =15'b0;

   // m236_68 = W*in
   wire signed [14:0] m236_68;
   assign m236_68 =15'b0;

   // m236_69 = W*in
   wire signed [14:0] m236_69;
   assign m236_69 =15'b0;

   // m236_70 = W*in
   wire signed [14:0] m236_70;
   assign m236_70 =15'b0;

   // m236_71 = W*in
   wire signed [14:0] m236_71;
   assign m236_71 =15'b0;

   // m236_72 = W*in
   wire signed [14:0] m236_72;
   assign m236_72 =15'b0;

   // m236_73 = W*in
   wire signed [14:0] m236_73;
   assign m236_73 =15'b0;

   // m236_74 = W*in
   wire signed [14:0] m236_74;
   assign m236_74 =15'b0;

   // m236_75 = W*in
   wire signed [14:0] m236_75;
   assign m236_75 ={ {4{in236[14]}} , in236[14:4] };

   // m236_76 = W*in
   wire signed [14:0] m236_76;
   assign m236_76 ={ {4{neg236[14]}} , neg236[14:4] };

   // m236_77 = W*in
   wire signed [14:0] m236_77;
   assign m236_77 =15'b0;

   // m236_78 = W*in
   wire signed [14:0] m236_78;
   assign m236_78 =15'b0;

   // m236_79 = W*in
   wire signed [14:0] m236_79;
   assign m236_79 =15'b0;

   // m236_80 = W*in
   wire signed [14:0] m236_80;
   assign m236_80 =15'b0;

   // m236_81 = W*in
   wire signed [14:0] m236_81;
   assign m236_81 ={ {3{neg236[14]}} , neg236[14:3] };

   // m236_82 = W*in
   wire signed [14:0] m236_82;
   assign m236_82 =15'b0;

   // m236_83 = W*in
   wire signed [14:0] m236_83;
   assign m236_83 =15'b0;

   // m236_84 = W*in
   wire signed [14:0] m236_84;
   assign m236_84 =15'b0;

   // m236_85 = W*in
   wire signed [14:0] m236_85;
   assign m236_85 ={ {3{neg236[14]}} , neg236[14:3] };

   // m236_86 = W*in
   wire signed [14:0] m236_86;
   assign m236_86 =15'b0;

   // m236_87 = W*in
   wire signed [14:0] m236_87;
   assign m236_87 =15'b0;

   // m236_88 = W*in
   wire signed [14:0] m236_88;
   assign m236_88 =15'b0;

   // m236_89 = W*in
   wire signed [14:0] m236_89;
   assign m236_89 =15'b0;

   // m236_90 = W*in
   wire signed [14:0] m236_90;
   assign m236_90 =15'b0;

   // m236_91 = W*in
   wire signed [14:0] m236_91;
   assign m236_91 =15'b0;

   // m236_92 = W*in
   wire signed [14:0] m236_92;
   assign m236_92 =15'b0;

   // m236_93 = W*in
   wire signed [14:0] m236_93;
   assign m236_93 =15'b0;

   // m236_94 = W*in
   wire signed [14:0] m236_94;
   assign m236_94 =15'b0;

   // m236_95 = W*in
   wire signed [14:0] m236_95;
   assign m236_95 ={ {4{in236[14]}} , in236[14:4] };

   // m236_96 = W*in
   wire signed [14:0] m236_96;
   assign m236_96 =15'b0;

   // m236_97 = W*in
   wire signed [14:0] m236_97;
   assign m236_97 =15'b0;

   // m236_98 = W*in
   wire signed [14:0] m236_98;
   assign m236_98 =15'b0;

   // m236_99 = W*in
   wire signed [14:0] m236_99;
   assign m236_99 =15'b0;

   // m236_100 = W*in
   wire signed [14:0] m236_100;
   assign m236_100 =15'b0;

   // m237_1 = W*in
   wire signed [14:0] m237_1;
   assign m237_1 =15'b0;

   // m237_2 = W*in
   wire signed [14:0] m237_2;
   assign m237_2 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_3 = W*in
   wire signed [14:0] m237_3;
   assign m237_3 =15'b0;

   // m237_4 = W*in
   wire signed [14:0] m237_4;
   assign m237_4 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_5 = W*in
   wire signed [14:0] m237_5;
   assign m237_5 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_6 = W*in
   wire signed [14:0] m237_6;
   assign m237_6 =15'b0;

   // m237_7 = W*in
   wire signed [14:0] m237_7;
   assign m237_7 =15'b0;

   // m237_8 = W*in
   wire signed [14:0] m237_8;
   assign m237_8 =15'b0;

   // m237_9 = W*in
   wire signed [14:0] m237_9;
   assign m237_9 =15'b0;

   // m237_10 = W*in
   wire signed [14:0] m237_10;
   assign m237_10 =15'b0;

   // m237_11 = W*in
   wire signed [14:0] m237_11;
   assign m237_11 ={ {3{in237[14]}} , in237[14:3] };

   // m237_12 = W*in
   wire signed [14:0] m237_12;
   assign m237_12 =15'b0;

   // m237_13 = W*in
   wire signed [14:0] m237_13;
   assign m237_13 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_14 = W*in
   wire signed [14:0] m237_14;
   assign m237_14 =15'b0;

   // m237_15 = W*in
   wire signed [14:0] m237_15;
   assign m237_15 =15'b0;

   // m237_16 = W*in
   wire signed [14:0] m237_16;
   assign m237_16 =15'b0;

   // m237_17 = W*in
   wire signed [14:0] m237_17;
   assign m237_17 =15'b0;

   // m237_18 = W*in
   wire signed [14:0] m237_18;
   assign m237_18 =15'b0;

   // m237_19 = W*in
   wire signed [14:0] m237_19;
   assign m237_19 =15'b0;

   // m237_20 = W*in
   wire signed [14:0] m237_20;
   assign m237_20 =15'b0;

   // m237_21 = W*in
   wire signed [14:0] m237_21;
   assign m237_21 =15'b0;

   // m237_22 = W*in
   wire signed [14:0] m237_22;
   assign m237_22 =15'b0;

   // m237_23 = W*in
   wire signed [14:0] m237_23;
   assign m237_23 =15'b0;

   // m237_24 = W*in
   wire signed [14:0] m237_24;
   assign m237_24 =15'b0;

   // m237_25 = W*in
   wire signed [14:0] m237_25;
   assign m237_25 =15'b0;

   // m237_26 = W*in
   wire signed [14:0] m237_26;
   assign m237_26 =15'b0;

   // m237_27 = W*in
   wire signed [14:0] m237_27;
   assign m237_27 =15'b0;

   // m237_28 = W*in
   wire signed [14:0] m237_28;
   assign m237_28 =15'b0;

   // m237_29 = W*in
   wire signed [14:0] m237_29;
   assign m237_29 =15'b0;

   // m237_30 = W*in
   wire signed [14:0] m237_30;
   assign m237_30 =15'b0;

   // m237_31 = W*in
   wire signed [14:0] m237_31;
   assign m237_31 ={ {3{in237[14]}} , in237[14:3] };

   // m237_32 = W*in
   wire signed [14:0] m237_32;
   assign m237_32 =15'b0;

   // m237_33 = W*in
   wire signed [14:0] m237_33;
   assign m237_33 =15'b0;

   // m237_34 = W*in
   wire signed [14:0] m237_34;
   assign m237_34 =15'b0;

   // m237_35 = W*in
   wire signed [14:0] m237_35;
   assign m237_35 =15'b0;

   // m237_36 = W*in
   wire signed [14:0] m237_36;
   assign m237_36 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_37 = W*in
   wire signed [14:0] m237_37;
   assign m237_37 =15'b0;

   // m237_38 = W*in
   wire signed [14:0] m237_38;
   assign m237_38 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_39 = W*in
   wire signed [14:0] m237_39;
   assign m237_39 ={ {3{in237[14]}} , in237[14:3] };

   // m237_40 = W*in
   wire signed [14:0] m237_40;
   assign m237_40 =15'b0;

   // m237_41 = W*in
   wire signed [14:0] m237_41;
   assign m237_41 ={ {3{in237[14]}} , in237[14:3] };

   // m237_42 = W*in
   wire signed [14:0] m237_42;
   assign m237_42 =15'b0;

   // m237_43 = W*in
   wire signed [14:0] m237_43;
   assign m237_43 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_44 = W*in
   wire signed [14:0] m237_44;
   assign m237_44 =15'b0;

   // m237_45 = W*in
   wire signed [14:0] m237_45;
   assign m237_45 =15'b0;

   // m237_46 = W*in
   wire signed [14:0] m237_46;
   assign m237_46 =15'b0;

   // m237_47 = W*in
   wire signed [14:0] m237_47;
   assign m237_47 =15'b0;

   // m237_48 = W*in
   wire signed [14:0] m237_48;
   assign m237_48 =15'b0;

   // m237_49 = W*in
   wire signed [14:0] m237_49;
   assign m237_49 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_50 = W*in
   wire signed [14:0] m237_50;
   assign m237_50 =15'b0;

   // m237_51 = W*in
   wire signed [14:0] m237_51;
   assign m237_51 =15'b0;

   // m237_52 = W*in
   wire signed [14:0] m237_52;
   assign m237_52 ={ {3{in237[14]}} , in237[14:3] };

   // m237_53 = W*in
   wire signed [14:0] m237_53;
   assign m237_53 ={ {3{in237[14]}} , in237[14:3] };

   // m237_54 = W*in
   wire signed [14:0] m237_54;
   assign m237_54 =15'b0;

   // m237_55 = W*in
   wire signed [14:0] m237_55;
   assign m237_55 =15'b0;

   // m237_56 = W*in
   wire signed [14:0] m237_56;
   assign m237_56 ={ {3{in237[14]}} , in237[14:3] };

   // m237_57 = W*in
   wire signed [14:0] m237_57;
   assign m237_57 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_58 = W*in
   wire signed [14:0] m237_58;
   assign m237_58 =15'b0;

   // m237_59 = W*in
   wire signed [14:0] m237_59;
   assign m237_59 =15'b0;

   // m237_60 = W*in
   wire signed [14:0] m237_60;
   assign m237_60 =15'b0;

   // m237_61 = W*in
   wire signed [14:0] m237_61;
   assign m237_61 =15'b0;

   // m237_62 = W*in
   wire signed [14:0] m237_62;
   assign m237_62 =15'b0;

   // m237_63 = W*in
   wire signed [14:0] m237_63;
   assign m237_63 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_64 = W*in
   wire signed [14:0] m237_64;
   assign m237_64 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_65 = W*in
   wire signed [14:0] m237_65;
   assign m237_65 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_66 = W*in
   wire signed [14:0] m237_66;
   assign m237_66 =15'b0;

   // m237_67 = W*in
   wire signed [14:0] m237_67;
   assign m237_67 =15'b0;

   // m237_68 = W*in
   wire signed [14:0] m237_68;
   assign m237_68 =15'b0;

   // m237_69 = W*in
   wire signed [14:0] m237_69;
   assign m237_69 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_70 = W*in
   wire signed [14:0] m237_70;
   assign m237_70 ={ {3{in237[14]}} , in237[14:3] };

   // m237_71 = W*in
   wire signed [14:0] m237_71;
   assign m237_71 ={ {3{in237[14]}} , in237[14:3] };

   // m237_72 = W*in
   wire signed [14:0] m237_72;
   assign m237_72 =15'b0;

   // m237_73 = W*in
   wire signed [14:0] m237_73;
   assign m237_73 =15'b0;

   // m237_74 = W*in
   wire signed [14:0] m237_74;
   assign m237_74 ={ {4{in237[14]}} , in237[14:4] };

   // m237_75 = W*in
   wire signed [14:0] m237_75;
   assign m237_75 =15'b0;

   // m237_76 = W*in
   wire signed [14:0] m237_76;
   assign m237_76 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_77 = W*in
   wire signed [14:0] m237_77;
   assign m237_77 =15'b0;

   // m237_78 = W*in
   wire signed [14:0] m237_78;
   assign m237_78 =15'b0;

   // m237_79 = W*in
   wire signed [14:0] m237_79;
   assign m237_79 =15'b0;

   // m237_80 = W*in
   wire signed [14:0] m237_80;
   assign m237_80 =15'b0;

   // m237_81 = W*in
   wire signed [14:0] m237_81;
   assign m237_81 =15'b0;

   // m237_82 = W*in
   wire signed [14:0] m237_82;
   assign m237_82 ={ {4{neg237[14]}} , neg237[14:4] };

   // m237_83 = W*in
   wire signed [14:0] m237_83;
   assign m237_83 =15'b0;

   // m237_84 = W*in
   wire signed [14:0] m237_84;
   assign m237_84 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_85 = W*in
   wire signed [14:0] m237_85;
   assign m237_85 ={ {3{in237[14]}} , in237[14:3] };

   // m237_86 = W*in
   wire signed [14:0] m237_86;
   assign m237_86 ={ {3{neg237[14]}} , neg237[14:3] };

   // m237_87 = W*in
   wire signed [14:0] m237_87;
   assign m237_87 =15'b0;

   // m237_88 = W*in
   wire signed [14:0] m237_88;
   assign m237_88 =15'b0;

   // m237_89 = W*in
   wire signed [14:0] m237_89;
   assign m237_89 =15'b0;

   // m237_90 = W*in
   wire signed [14:0] m237_90;
   assign m237_90 =15'b0;

   // m237_91 = W*in
   wire signed [14:0] m237_91;
   assign m237_91 ={ {3{in237[14]}} , in237[14:3] };

   // m237_92 = W*in
   wire signed [14:0] m237_92;
   assign m237_92 =15'b0;

   // m237_93 = W*in
   wire signed [14:0] m237_93;
   assign m237_93 =15'b0;

   // m237_94 = W*in
   wire signed [14:0] m237_94;
   assign m237_94 =15'b0;

   // m237_95 = W*in
   wire signed [14:0] m237_95;
   assign m237_95 =15'b0;

   // m237_96 = W*in
   wire signed [14:0] m237_96;
   assign m237_96 =15'b0;

   // m237_97 = W*in
   wire signed [14:0] m237_97;
   assign m237_97 =15'b0;

   // m237_98 = W*in
   wire signed [14:0] m237_98;
   assign m237_98 =15'b0;

   // m237_99 = W*in
   wire signed [14:0] m237_99;
   assign m237_99 ={ {3{in237[14]}} , in237[14:3] };

   // m237_100 = W*in
   wire signed [14:0] m237_100;
   assign m237_100 =15'b0;

   // m238_1 = W*in
   wire signed [14:0] m238_1;
   assign m238_1 =15'b0;

   // m238_2 = W*in
   wire signed [14:0] m238_2;
   assign m238_2 =15'b0;

   // m238_3 = W*in
   wire signed [14:0] m238_3;
   assign m238_3 =15'b0;

   // m238_4 = W*in
   wire signed [14:0] m238_4;
   assign m238_4 =15'b0;

   // m238_5 = W*in
   wire signed [14:0] m238_5;
   assign m238_5 =15'b0;

   // m238_6 = W*in
   wire signed [14:0] m238_6;
   assign m238_6 =15'b0;

   // m238_7 = W*in
   wire signed [14:0] m238_7;
   assign m238_7 =15'b0;

   // m238_8 = W*in
   wire signed [14:0] m238_8;
   assign m238_8 =15'b0;

   // m238_9 = W*in
   wire signed [14:0] m238_9;
   assign m238_9 ={ {3{neg238[14]}} , neg238[14:3] };

   // m238_10 = W*in
   wire signed [14:0] m238_10;
   assign m238_10 =15'b0;

   // m238_11 = W*in
   wire signed [14:0] m238_11;
   assign m238_11 =15'b0;

   // m238_12 = W*in
   wire signed [14:0] m238_12;
   assign m238_12 =15'b0;

   // m238_13 = W*in
   wire signed [14:0] m238_13;
   assign m238_13 =15'b0;

   // m238_14 = W*in
   wire signed [14:0] m238_14;
   assign m238_14 ={ {4{neg238[14]}} , neg238[14:4] };

   // m238_15 = W*in
   wire signed [14:0] m238_15;
   assign m238_15 =15'b0;

   // m238_16 = W*in
   wire signed [14:0] m238_16;
   assign m238_16 =15'b0;

   // m238_17 = W*in
   wire signed [14:0] m238_17;
   assign m238_17 =15'b0;

   // m238_18 = W*in
   wire signed [14:0] m238_18;
   assign m238_18 =15'b0;

   // m238_19 = W*in
   wire signed [14:0] m238_19;
   assign m238_19 =15'b0;

   // m238_20 = W*in
   wire signed [14:0] m238_20;
   assign m238_20 =15'b0;

   // m238_21 = W*in
   wire signed [14:0] m238_21;
   assign m238_21 =15'b0;

   // m238_22 = W*in
   wire signed [14:0] m238_22;
   assign m238_22 =15'b0;

   // m238_23 = W*in
   wire signed [14:0] m238_23;
   assign m238_23 =15'b0;

   // m238_24 = W*in
   wire signed [14:0] m238_24;
   assign m238_24 ={ {3{in238[14]}} , in238[14:3] };

   // m238_25 = W*in
   wire signed [14:0] m238_25;
   assign m238_25 =15'b0;

   // m238_26 = W*in
   wire signed [14:0] m238_26;
   assign m238_26 ={ {3{neg238[14]}} , neg238[14:3] };

   // m238_27 = W*in
   wire signed [14:0] m238_27;
   assign m238_27 =15'b0;

   // m238_28 = W*in
   wire signed [14:0] m238_28;
   assign m238_28 =15'b0;

   // m238_29 = W*in
   wire signed [14:0] m238_29;
   assign m238_29 =15'b0;

   // m238_30 = W*in
   wire signed [14:0] m238_30;
   assign m238_30 ={ {3{neg238[14]}} , neg238[14:3] };

   // m238_31 = W*in
   wire signed [14:0] m238_31;
   assign m238_31 =15'b0;

   // m238_32 = W*in
   wire signed [14:0] m238_32;
   assign m238_32 =15'b0;

   // m238_33 = W*in
   wire signed [14:0] m238_33;
   assign m238_33 ={ {3{neg238[14]}} , neg238[14:3] };

   // m238_34 = W*in
   wire signed [14:0] m238_34;
   assign m238_34 =15'b0;

   // m238_35 = W*in
   wire signed [14:0] m238_35;
   assign m238_35 =15'b0;

   // m238_36 = W*in
   wire signed [14:0] m238_36;
   assign m238_36 ={ {3{neg238[14]}} , neg238[14:3] };

   // m238_37 = W*in
   wire signed [14:0] m238_37;
   assign m238_37 ={ {3{in238[14]}} , in238[14:3] };

   // m238_38 = W*in
   wire signed [14:0] m238_38;
   assign m238_38 =15'b0;

   // m238_39 = W*in
   wire signed [14:0] m238_39;
   assign m238_39 =15'b0;

   // m238_40 = W*in
   wire signed [14:0] m238_40;
   assign m238_40 =15'b0;

   // m238_41 = W*in
   wire signed [14:0] m238_41;
   assign m238_41 =15'b0;

   // m238_42 = W*in
   wire signed [14:0] m238_42;
   assign m238_42 =15'b0;

   // m238_43 = W*in
   wire signed [14:0] m238_43;
   assign m238_43 =15'b0;

   // m238_44 = W*in
   wire signed [14:0] m238_44;
   assign m238_44 =15'b0;

   // m238_45 = W*in
   wire signed [14:0] m238_45;
   assign m238_45 =15'b0;

   // m238_46 = W*in
   wire signed [14:0] m238_46;
   assign m238_46 =15'b0;

   // m238_47 = W*in
   wire signed [14:0] m238_47;
   assign m238_47 =15'b0;

   // m238_48 = W*in
   wire signed [14:0] m238_48;
   assign m238_48 =15'b0;

   // m238_49 = W*in
   wire signed [14:0] m238_49;
   assign m238_49 =15'b0;

   // m238_50 = W*in
   wire signed [14:0] m238_50;
   assign m238_50 =15'b0;

   // m238_51 = W*in
   wire signed [14:0] m238_51;
   assign m238_51 =15'b0;

   // m238_52 = W*in
   wire signed [14:0] m238_52;
   assign m238_52 =15'b0;

   // m238_53 = W*in
   wire signed [14:0] m238_53;
   assign m238_53 =15'b0;

   // m238_54 = W*in
   wire signed [14:0] m238_54;
   assign m238_54 =15'b0;

   // m238_55 = W*in
   wire signed [14:0] m238_55;
   assign m238_55 =15'b0;

   // m238_56 = W*in
   wire signed [14:0] m238_56;
   assign m238_56 =15'b0;

   // m238_57 = W*in
   wire signed [14:0] m238_57;
   assign m238_57 =15'b0;

   // m238_58 = W*in
   wire signed [14:0] m238_58;
   assign m238_58 =15'b0;

   // m238_59 = W*in
   wire signed [14:0] m238_59;
   assign m238_59 =15'b0;

   // m238_60 = W*in
   wire signed [14:0] m238_60;
   assign m238_60 =15'b0;

   // m238_61 = W*in
   wire signed [14:0] m238_61;
   assign m238_61 =15'b0;

   // m238_62 = W*in
   wire signed [14:0] m238_62;
   assign m238_62 =15'b0;

   // m238_63 = W*in
   wire signed [14:0] m238_63;
   assign m238_63 ={ {3{in238[14]}} , in238[14:3] };

   // m238_64 = W*in
   wire signed [14:0] m238_64;
   assign m238_64 =15'b0;

   // m238_65 = W*in
   wire signed [14:0] m238_65;
   assign m238_65 =15'b0;

   // m238_66 = W*in
   wire signed [14:0] m238_66;
   assign m238_66 =15'b0;

   // m238_67 = W*in
   wire signed [14:0] m238_67;
   assign m238_67 =15'b0;

   // m238_68 = W*in
   wire signed [14:0] m238_68;
   assign m238_68 =15'b0;

   // m238_69 = W*in
   wire signed [14:0] m238_69;
   assign m238_69 =15'b0;

   // m238_70 = W*in
   wire signed [14:0] m238_70;
   assign m238_70 =15'b0;

   // m238_71 = W*in
   wire signed [14:0] m238_71;
   assign m238_71 =15'b0;

   // m238_72 = W*in
   wire signed [14:0] m238_72;
   assign m238_72 =15'b0;

   // m238_73 = W*in
   wire signed [14:0] m238_73;
   assign m238_73 =15'b0;

   // m238_74 = W*in
   wire signed [14:0] m238_74;
   assign m238_74 =15'b0;

   // m238_75 = W*in
   wire signed [14:0] m238_75;
   assign m238_75 =15'b0;

   // m238_76 = W*in
   wire signed [14:0] m238_76;
   assign m238_76 ={ {4{neg238[14]}} , neg238[14:4] };

   // m238_77 = W*in
   wire signed [14:0] m238_77;
   assign m238_77 =15'b0;

   // m238_78 = W*in
   wire signed [14:0] m238_78;
   assign m238_78 =15'b0;

   // m238_79 = W*in
   wire signed [14:0] m238_79;
   assign m238_79 =15'b0;

   // m238_80 = W*in
   wire signed [14:0] m238_80;
   assign m238_80 =15'b0;

   // m238_81 = W*in
   wire signed [14:0] m238_81;
   assign m238_81 =15'b0;

   // m238_82 = W*in
   wire signed [14:0] m238_82;
   assign m238_82 =15'b0;

   // m238_83 = W*in
   wire signed [14:0] m238_83;
   assign m238_83 ={ {2{in238[14]}} , in238[14:2] };

   // m238_84 = W*in
   wire signed [14:0] m238_84;
   assign m238_84 =15'b0;

   // m238_85 = W*in
   wire signed [14:0] m238_85;
   assign m238_85 =15'b0;

   // m238_86 = W*in
   wire signed [14:0] m238_86;
   assign m238_86 ={ {3{neg238[14]}} , neg238[14:3] };

   // m238_87 = W*in
   wire signed [14:0] m238_87;
   assign m238_87 =15'b0;

   // m238_88 = W*in
   wire signed [14:0] m238_88;
   assign m238_88 =15'b0;

   // m238_89 = W*in
   wire signed [14:0] m238_89;
   assign m238_89 =15'b0;

   // m238_90 = W*in
   wire signed [14:0] m238_90;
   assign m238_90 =15'b0;

   // m238_91 = W*in
   wire signed [14:0] m238_91;
   assign m238_91 ={ {3{in238[14]}} , in238[14:3] };

   // m238_92 = W*in
   wire signed [14:0] m238_92;
   assign m238_92 =15'b0;

   // m238_93 = W*in
   wire signed [14:0] m238_93;
   assign m238_93 =15'b0;

   // m238_94 = W*in
   wire signed [14:0] m238_94;
   assign m238_94 =15'b0;

   // m238_95 = W*in
   wire signed [14:0] m238_95;
   assign m238_95 =15'b0;

   // m238_96 = W*in
   wire signed [14:0] m238_96;
   assign m238_96 =15'b0;

   // m238_97 = W*in
   wire signed [14:0] m238_97;
   assign m238_97 =15'b0;

   // m238_98 = W*in
   wire signed [14:0] m238_98;
   assign m238_98 =15'b0;

   // m238_99 = W*in
   wire signed [14:0] m238_99;
   assign m238_99 =15'b0;

   // m238_100 = W*in
   wire signed [14:0] m238_100;
   assign m238_100 =15'b0;

   // m239_1 = W*in
   wire signed [14:0] m239_1;
   assign m239_1 =15'b0;

   // m239_2 = W*in
   wire signed [14:0] m239_2;
   assign m239_2 =15'b0;

   // m239_3 = W*in
   wire signed [14:0] m239_3;
   assign m239_3 =15'b0;

   // m239_4 = W*in
   wire signed [14:0] m239_4;
   assign m239_4 =15'b0;

   // m239_5 = W*in
   wire signed [14:0] m239_5;
   assign m239_5 =15'b0;

   // m239_6 = W*in
   wire signed [14:0] m239_6;
   assign m239_6 =15'b0;

   // m239_7 = W*in
   wire signed [14:0] m239_7;
   assign m239_7 =15'b0;

   // m239_8 = W*in
   wire signed [14:0] m239_8;
   assign m239_8 =15'b0;

   // m239_9 = W*in
   wire signed [14:0] m239_9;
   assign m239_9 =15'b0;

   // m239_10 = W*in
   wire signed [14:0] m239_10;
   assign m239_10 ={ {3{in239[14]}} , in239[14:3] };

   // m239_11 = W*in
   wire signed [14:0] m239_11;
   assign m239_11 =15'b0;

   // m239_12 = W*in
   wire signed [14:0] m239_12;
   assign m239_12 =15'b0;

   // m239_13 = W*in
   wire signed [14:0] m239_13;
   assign m239_13 =15'b0;

   // m239_14 = W*in
   wire signed [14:0] m239_14;
   assign m239_14 =15'b0;

   // m239_15 = W*in
   wire signed [14:0] m239_15;
   assign m239_15 =15'b0;

   // m239_16 = W*in
   wire signed [14:0] m239_16;
   assign m239_16 =15'b0;

   // m239_17 = W*in
   wire signed [14:0] m239_17;
   assign m239_17 =15'b0;

   // m239_18 = W*in
   wire signed [14:0] m239_18;
   assign m239_18 =15'b0;

   // m239_19 = W*in
   wire signed [14:0] m239_19;
   assign m239_19 =15'b0;

   // m239_20 = W*in
   wire signed [14:0] m239_20;
   assign m239_20 =15'b0;

   // m239_21 = W*in
   wire signed [14:0] m239_21;
   assign m239_21 =15'b0;

   // m239_22 = W*in
   wire signed [14:0] m239_22;
   assign m239_22 =15'b0;

   // m239_23 = W*in
   wire signed [14:0] m239_23;
   assign m239_23 =15'b0;

   // m239_24 = W*in
   wire signed [14:0] m239_24;
   assign m239_24 =15'b0;

   // m239_25 = W*in
   wire signed [14:0] m239_25;
   assign m239_25 ={ {3{in239[14]}} , in239[14:3] };

   // m239_26 = W*in
   wire signed [14:0] m239_26;
   assign m239_26 ={ {3{neg239[14]}} , neg239[14:3] };

   // m239_27 = W*in
   wire signed [14:0] m239_27;
   assign m239_27 =15'b0;

   // m239_28 = W*in
   wire signed [14:0] m239_28;
   assign m239_28 =15'b0;

   // m239_29 = W*in
   wire signed [14:0] m239_29;
   assign m239_29 =15'b0;

   // m239_30 = W*in
   wire signed [14:0] m239_30;
   assign m239_30 =15'b0;

   // m239_31 = W*in
   wire signed [14:0] m239_31;
   assign m239_31 ={ {3{neg239[14]}} , neg239[14:3] };

   // m239_32 = W*in
   wire signed [14:0] m239_32;
   assign m239_32 =15'b0;

   // m239_33 = W*in
   wire signed [14:0] m239_33;
   assign m239_33 =15'b0;

   // m239_34 = W*in
   wire signed [14:0] m239_34;
   assign m239_34 =15'b0;

   // m239_35 = W*in
   wire signed [14:0] m239_35;
   assign m239_35 =15'b0;

   // m239_36 = W*in
   wire signed [14:0] m239_36;
   assign m239_36 =15'b0;

   // m239_37 = W*in
   wire signed [14:0] m239_37;
   assign m239_37 =15'b0;

   // m239_38 = W*in
   wire signed [14:0] m239_38;
   assign m239_38 =15'b0;

   // m239_39 = W*in
   wire signed [14:0] m239_39;
   assign m239_39 =15'b0;

   // m239_40 = W*in
   wire signed [14:0] m239_40;
   assign m239_40 =15'b0;

   // m239_41 = W*in
   wire signed [14:0] m239_41;
   assign m239_41 =15'b0;

   // m239_42 = W*in
   wire signed [14:0] m239_42;
   assign m239_42 =15'b0;

   // m239_43 = W*in
   wire signed [14:0] m239_43;
   assign m239_43 =15'b0;

   // m239_44 = W*in
   wire signed [14:0] m239_44;
   assign m239_44 =15'b0;

   // m239_45 = W*in
   wire signed [14:0] m239_45;
   assign m239_45 =15'b0;

   // m239_46 = W*in
   wire signed [14:0] m239_46;
   assign m239_46 ={ {3{in239[14]}} , in239[14:3] };

   // m239_47 = W*in
   wire signed [14:0] m239_47;
   assign m239_47 =15'b0;

   // m239_48 = W*in
   wire signed [14:0] m239_48;
   assign m239_48 =15'b0;

   // m239_49 = W*in
   wire signed [14:0] m239_49;
   assign m239_49 =15'b0;

   // m239_50 = W*in
   wire signed [14:0] m239_50;
   assign m239_50 =15'b0;

   // m239_51 = W*in
   wire signed [14:0] m239_51;
   assign m239_51 =15'b0;

   // m239_52 = W*in
   wire signed [14:0] m239_52;
   assign m239_52 =15'b0;

   // m239_53 = W*in
   wire signed [14:0] m239_53;
   assign m239_53 =15'b0;

   // m239_54 = W*in
   wire signed [14:0] m239_54;
   assign m239_54 =15'b0;

   // m239_55 = W*in
   wire signed [14:0] m239_55;
   assign m239_55 =15'b0;

   // m239_56 = W*in
   wire signed [14:0] m239_56;
   assign m239_56 =15'b0;

   // m239_57 = W*in
   wire signed [14:0] m239_57;
   assign m239_57 =15'b0;

   // m239_58 = W*in
   wire signed [14:0] m239_58;
   assign m239_58 ={ {3{neg239[14]}} , neg239[14:3] };

   // m239_59 = W*in
   wire signed [14:0] m239_59;
   assign m239_59 =15'b0;

   // m239_60 = W*in
   wire signed [14:0] m239_60;
   assign m239_60 =15'b0;

   // m239_61 = W*in
   wire signed [14:0] m239_61;
   assign m239_61 =15'b0;

   // m239_62 = W*in
   wire signed [14:0] m239_62;
   assign m239_62 =15'b0;

   // m239_63 = W*in
   wire signed [14:0] m239_63;
   assign m239_63 =15'b0;

   // m239_64 = W*in
   wire signed [14:0] m239_64;
   assign m239_64 =15'b0;

   // m239_65 = W*in
   wire signed [14:0] m239_65;
   assign m239_65 =15'b0;

   // m239_66 = W*in
   wire signed [14:0] m239_66;
   assign m239_66 =15'b0;

   // m239_67 = W*in
   wire signed [14:0] m239_67;
   assign m239_67 =15'b0;

   // m239_68 = W*in
   wire signed [14:0] m239_68;
   assign m239_68 ={ {4{neg239[14]}} , neg239[14:4] };

   // m239_69 = W*in
   wire signed [14:0] m239_69;
   assign m239_69 =15'b0;

   // m239_70 = W*in
   wire signed [14:0] m239_70;
   assign m239_70 =15'b0;

   // m239_71 = W*in
   wire signed [14:0] m239_71;
   assign m239_71 =15'b0;

   // m239_72 = W*in
   wire signed [14:0] m239_72;
   assign m239_72 ={ {3{in239[14]}} , in239[14:3] };

   // m239_73 = W*in
   wire signed [14:0] m239_73;
   assign m239_73 =15'b0;

   // m239_74 = W*in
   wire signed [14:0] m239_74;
   assign m239_74 =15'b0;

   // m239_75 = W*in
   wire signed [14:0] m239_75;
   assign m239_75 =15'b0;

   // m239_76 = W*in
   wire signed [14:0] m239_76;
   assign m239_76 =15'b0;

   // m239_77 = W*in
   wire signed [14:0] m239_77;
   assign m239_77 =15'b0;

   // m239_78 = W*in
   wire signed [14:0] m239_78;
   assign m239_78 =15'b0;

   // m239_79 = W*in
   wire signed [14:0] m239_79;
   assign m239_79 =15'b0;

   // m239_80 = W*in
   wire signed [14:0] m239_80;
   assign m239_80 ={ {3{in239[14]}} , in239[14:3] };

   // m239_81 = W*in
   wire signed [14:0] m239_81;
   assign m239_81 =15'b0;

   // m239_82 = W*in
   wire signed [14:0] m239_82;
   assign m239_82 =15'b0;

   // m239_83 = W*in
   wire signed [14:0] m239_83;
   assign m239_83 =15'b0;

   // m239_84 = W*in
   wire signed [14:0] m239_84;
   assign m239_84 =15'b0;

   // m239_85 = W*in
   wire signed [14:0] m239_85;
   assign m239_85 =15'b0;

   // m239_86 = W*in
   wire signed [14:0] m239_86;
   assign m239_86 =15'b0;

   // m239_87 = W*in
   wire signed [14:0] m239_87;
   assign m239_87 =15'b0;

   // m239_88 = W*in
   wire signed [14:0] m239_88;
   assign m239_88 =15'b0;

   // m239_89 = W*in
   wire signed [14:0] m239_89;
   assign m239_89 =15'b0;

   // m239_90 = W*in
   wire signed [14:0] m239_90;
   assign m239_90 =15'b0;

   // m239_91 = W*in
   wire signed [14:0] m239_91;
   assign m239_91 =15'b0;

   // m239_92 = W*in
   wire signed [14:0] m239_92;
   assign m239_92 ={ {3{neg239[14]}} , neg239[14:3] };

   // m239_93 = W*in
   wire signed [14:0] m239_93;
   assign m239_93 ={ {3{in239[14]}} , in239[14:3] };

   // m239_94 = W*in
   wire signed [14:0] m239_94;
   assign m239_94 =15'b0;

   // m239_95 = W*in
   wire signed [14:0] m239_95;
   assign m239_95 ={ {3{in239[14]}} , in239[14:3] };

   // m239_96 = W*in
   wire signed [14:0] m239_96;
   assign m239_96 ={ {3{in239[14]}} , in239[14:3] };

   // m239_97 = W*in
   wire signed [14:0] m239_97;
   assign m239_97 =15'b0;

   // m239_98 = W*in
   wire signed [14:0] m239_98;
   assign m239_98 =15'b0;

   // m239_99 = W*in
   wire signed [14:0] m239_99;
   assign m239_99 =15'b0;

   // m239_100 = W*in
   wire signed [14:0] m239_100;
   assign m239_100 =15'b0;

   // m240_1 = W*in
   wire signed [14:0] m240_1;
   assign m240_1 =15'b0;

   // m240_2 = W*in
   wire signed [14:0] m240_2;
   assign m240_2 =15'b0;

   // m240_3 = W*in
   wire signed [14:0] m240_3;
   assign m240_3 =15'b0;

   // m240_4 = W*in
   wire signed [14:0] m240_4;
   assign m240_4 =15'b0;

   // m240_5 = W*in
   wire signed [14:0] m240_5;
   assign m240_5 ={ {3{neg240[14]}} , neg240[14:3] };

   // m240_6 = W*in
   wire signed [14:0] m240_6;
   assign m240_6 =15'b0;

   // m240_7 = W*in
   wire signed [14:0] m240_7;
   assign m240_7 =15'b0;

   // m240_8 = W*in
   wire signed [14:0] m240_8;
   assign m240_8 ={ {4{neg240[14]}} , neg240[14:4] };

   // m240_9 = W*in
   wire signed [14:0] m240_9;
   assign m240_9 =15'b0;

   // m240_10 = W*in
   wire signed [14:0] m240_10;
   assign m240_10 =15'b0;

   // m240_11 = W*in
   wire signed [14:0] m240_11;
   assign m240_11 =15'b0;

   // m240_12 = W*in
   wire signed [14:0] m240_12;
   assign m240_12 =15'b0;

   // m240_13 = W*in
   wire signed [14:0] m240_13;
   assign m240_13 =15'b0;

   // m240_14 = W*in
   wire signed [14:0] m240_14;
   assign m240_14 ={ {3{neg240[14]}} , neg240[14:3] };

   // m240_15 = W*in
   wire signed [14:0] m240_15;
   assign m240_15 =15'b0;

   // m240_16 = W*in
   wire signed [14:0] m240_16;
   assign m240_16 ={ {3{neg240[14]}} , neg240[14:3] };

   // m240_17 = W*in
   wire signed [14:0] m240_17;
   assign m240_17 =15'b0;

   // m240_18 = W*in
   wire signed [14:0] m240_18;
   assign m240_18 =15'b0;

   // m240_19 = W*in
   wire signed [14:0] m240_19;
   assign m240_19 =15'b0;

   // m240_20 = W*in
   wire signed [14:0] m240_20;
   assign m240_20 ={ {3{neg240[14]}} , neg240[14:3] };

   // m240_21 = W*in
   wire signed [14:0] m240_21;
   assign m240_21 =15'b0;

   // m240_22 = W*in
   wire signed [14:0] m240_22;
   assign m240_22 =15'b0;

   // m240_23 = W*in
   wire signed [14:0] m240_23;
   assign m240_23 =15'b0;

   // m240_24 = W*in
   wire signed [14:0] m240_24;
   assign m240_24 =15'b0;

   // m240_25 = W*in
   wire signed [14:0] m240_25;
   assign m240_25 =15'b0;

   // m240_26 = W*in
   wire signed [14:0] m240_26;
   assign m240_26 =15'b0;

   // m240_27 = W*in
   wire signed [14:0] m240_27;
   assign m240_27 ={ {3{in240[14]}} , in240[14:3] };

   // m240_28 = W*in
   wire signed [14:0] m240_28;
   assign m240_28 =15'b0;

   // m240_29 = W*in
   wire signed [14:0] m240_29;
   assign m240_29 =15'b0;

   // m240_30 = W*in
   wire signed [14:0] m240_30;
   assign m240_30 =15'b0;

   // m240_31 = W*in
   wire signed [14:0] m240_31;
   assign m240_31 =15'b0;

   // m240_32 = W*in
   wire signed [14:0] m240_32;
   assign m240_32 =15'b0;

   // m240_33 = W*in
   wire signed [14:0] m240_33;
   assign m240_33 =15'b0;

   // m240_34 = W*in
   wire signed [14:0] m240_34;
   assign m240_34 =15'b0;

   // m240_35 = W*in
   wire signed [14:0] m240_35;
   assign m240_35 =15'b0;

   // m240_36 = W*in
   wire signed [14:0] m240_36;
   assign m240_36 =15'b0;

   // m240_37 = W*in
   wire signed [14:0] m240_37;
   assign m240_37 =15'b0;

   // m240_38 = W*in
   wire signed [14:0] m240_38;
   assign m240_38 =15'b0;

   // m240_39 = W*in
   wire signed [14:0] m240_39;
   assign m240_39 =15'b0;

   // m240_40 = W*in
   wire signed [14:0] m240_40;
   assign m240_40 ={ {4{neg240[14]}} , neg240[14:4] };

   // m240_41 = W*in
   wire signed [14:0] m240_41;
   assign m240_41 =15'b0;

   // m240_42 = W*in
   wire signed [14:0] m240_42;
   assign m240_42 =15'b0;

   // m240_43 = W*in
   wire signed [14:0] m240_43;
   assign m240_43 =15'b0;

   // m240_44 = W*in
   wire signed [14:0] m240_44;
   assign m240_44 =15'b0;

   // m240_45 = W*in
   wire signed [14:0] m240_45;
   assign m240_45 =15'b0;

   // m240_46 = W*in
   wire signed [14:0] m240_46;
   assign m240_46 =15'b0;

   // m240_47 = W*in
   wire signed [14:0] m240_47;
   assign m240_47 =15'b0;

   // m240_48 = W*in
   wire signed [14:0] m240_48;
   assign m240_48 =15'b0;

   // m240_49 = W*in
   wire signed [14:0] m240_49;
   assign m240_49 =15'b0;

   // m240_50 = W*in
   wire signed [14:0] m240_50;
   assign m240_50 =15'b0;

   // m240_51 = W*in
   wire signed [14:0] m240_51;
   assign m240_51 =15'b0;

   // m240_52 = W*in
   wire signed [14:0] m240_52;
   assign m240_52 =15'b0;

   // m240_53 = W*in
   wire signed [14:0] m240_53;
   assign m240_53 =15'b0;

   // m240_54 = W*in
   wire signed [14:0] m240_54;
   assign m240_54 =15'b0;

   // m240_55 = W*in
   wire signed [14:0] m240_55;
   assign m240_55 =15'b0;

   // m240_56 = W*in
   wire signed [14:0] m240_56;
   assign m240_56 =15'b0;

   // m240_57 = W*in
   wire signed [14:0] m240_57;
   assign m240_57 =15'b0;

   // m240_58 = W*in
   wire signed [14:0] m240_58;
   assign m240_58 =15'b0;

   // m240_59 = W*in
   wire signed [14:0] m240_59;
   assign m240_59 =15'b0;

   // m240_60 = W*in
   wire signed [14:0] m240_60;
   assign m240_60 =15'b0;

   // m240_61 = W*in
   wire signed [14:0] m240_61;
   assign m240_61 ={ {4{neg240[14]}} , neg240[14:4] };

   // m240_62 = W*in
   wire signed [14:0] m240_62;
   assign m240_62 =15'b0;

   // m240_63 = W*in
   wire signed [14:0] m240_63;
   assign m240_63 =15'b0;

   // m240_64 = W*in
   wire signed [14:0] m240_64;
   assign m240_64 =15'b0;

   // m240_65 = W*in
   wire signed [14:0] m240_65;
   assign m240_65 =15'b0;

   // m240_66 = W*in
   wire signed [14:0] m240_66;
   assign m240_66 =15'b0;

   // m240_67 = W*in
   wire signed [14:0] m240_67;
   assign m240_67 =15'b0;

   // m240_68 = W*in
   wire signed [14:0] m240_68;
   assign m240_68 =15'b0;

   // m240_69 = W*in
   wire signed [14:0] m240_69;
   assign m240_69 ={ {4{in240[14]}} , in240[14:4] };

   // m240_70 = W*in
   wire signed [14:0] m240_70;
   assign m240_70 =15'b0;

   // m240_71 = W*in
   wire signed [14:0] m240_71;
   assign m240_71 =15'b0;

   // m240_72 = W*in
   wire signed [14:0] m240_72;
   assign m240_72 ={ {2{in240[14]}} , in240[14:2] };

   // m240_73 = W*in
   wire signed [14:0] m240_73;
   assign m240_73 =15'b0;

   // m240_74 = W*in
   wire signed [14:0] m240_74;
   assign m240_74 =15'b0;

   // m240_75 = W*in
   wire signed [14:0] m240_75;
   assign m240_75 =15'b0;

   // m240_76 = W*in
   wire signed [14:0] m240_76;
   assign m240_76 ={ {4{neg240[14]}} , neg240[14:4] };

   // m240_77 = W*in
   wire signed [14:0] m240_77;
   assign m240_77 ={ {3{neg240[14]}} , neg240[14:3] };

   // m240_78 = W*in
   wire signed [14:0] m240_78;
   assign m240_78 =15'b0;

   // m240_79 = W*in
   wire signed [14:0] m240_79;
   assign m240_79 =15'b0;

   // m240_80 = W*in
   wire signed [14:0] m240_80;
   assign m240_80 =15'b0;

   // m240_81 = W*in
   wire signed [14:0] m240_81;
   assign m240_81 =15'b0;

   // m240_82 = W*in
   wire signed [14:0] m240_82;
   assign m240_82 ={ {4{neg240[14]}} , neg240[14:4] };

   // m240_83 = W*in
   wire signed [14:0] m240_83;
   assign m240_83 =15'b0;

   // m240_84 = W*in
   wire signed [14:0] m240_84;
   assign m240_84 =15'b0;

   // m240_85 = W*in
   wire signed [14:0] m240_85;
   assign m240_85 =15'b0;

   // m240_86 = W*in
   wire signed [14:0] m240_86;
   assign m240_86 =15'b0;

   // m240_87 = W*in
   wire signed [14:0] m240_87;
   assign m240_87 =15'b0;

   // m240_88 = W*in
   wire signed [14:0] m240_88;
   assign m240_88 =15'b0;

   // m240_89 = W*in
   wire signed [14:0] m240_89;
   assign m240_89 =15'b0;

   // m240_90 = W*in
   wire signed [14:0] m240_90;
   assign m240_90 =15'b0;

   // m240_91 = W*in
   wire signed [14:0] m240_91;
   assign m240_91 =15'b0;

   // m240_92 = W*in
   wire signed [14:0] m240_92;
   assign m240_92 =15'b0;

   // m240_93 = W*in
   wire signed [14:0] m240_93;
   assign m240_93 =15'b0;

   // m240_94 = W*in
   wire signed [14:0] m240_94;
   assign m240_94 =15'b0;

   // m240_95 = W*in
   wire signed [14:0] m240_95;
   assign m240_95 =15'b0;

   // m240_96 = W*in
   wire signed [14:0] m240_96;
   assign m240_96 =15'b0;

   // m240_97 = W*in
   wire signed [14:0] m240_97;
   assign m240_97 =15'b0;

   // m240_98 = W*in
   wire signed [14:0] m240_98;
   assign m240_98 =15'b0;

   // m240_99 = W*in
   wire signed [14:0] m240_99;
   assign m240_99 =15'b0;

   // m240_100 = W*in
   wire signed [14:0] m240_100;
   assign m240_100 =15'b0;

   // m241_1 = W*in
   wire signed [14:0] m241_1;
   assign m241_1 =15'b0;

   // m241_2 = W*in
   wire signed [14:0] m241_2;
   assign m241_2 ={ {4{in241[14]}} , in241[14:4] };

   // m241_3 = W*in
   wire signed [14:0] m241_3;
   assign m241_3 =15'b0;

   // m241_4 = W*in
   wire signed [14:0] m241_4;
   assign m241_4 ={ {4{neg241[14]}} , neg241[14:4] };

   // m241_5 = W*in
   wire signed [14:0] m241_5;
   assign m241_5 =15'b0;

   // m241_6 = W*in
   wire signed [14:0] m241_6;
   assign m241_6 =15'b0;

   // m241_7 = W*in
   wire signed [14:0] m241_7;
   assign m241_7 =15'b0;

   // m241_8 = W*in
   wire signed [14:0] m241_8;
   assign m241_8 =15'b0;

   // m241_9 = W*in
   wire signed [14:0] m241_9;
   assign m241_9 ={ {4{in241[14]}} , in241[14:4] };

   // m241_10 = W*in
   wire signed [14:0] m241_10;
   assign m241_10 =15'b0;

   // m241_11 = W*in
   wire signed [14:0] m241_11;
   assign m241_11 =15'b0;

   // m241_12 = W*in
   wire signed [14:0] m241_12;
   assign m241_12 =15'b0;

   // m241_13 = W*in
   wire signed [14:0] m241_13;
   assign m241_13 =15'b0;

   // m241_14 = W*in
   wire signed [14:0] m241_14;
   assign m241_14 =15'b0;

   // m241_15 = W*in
   wire signed [14:0] m241_15;
   assign m241_15 =15'b0;

   // m241_16 = W*in
   wire signed [14:0] m241_16;
   assign m241_16 =15'b0;

   // m241_17 = W*in
   wire signed [14:0] m241_17;
   assign m241_17 =15'b0;

   // m241_18 = W*in
   wire signed [14:0] m241_18;
   assign m241_18 =15'b0;

   // m241_19 = W*in
   wire signed [14:0] m241_19;
   assign m241_19 =15'b0;

   // m241_20 = W*in
   wire signed [14:0] m241_20;
   assign m241_20 =15'b0;

   // m241_21 = W*in
   wire signed [14:0] m241_21;
   assign m241_21 =15'b0;

   // m241_22 = W*in
   wire signed [14:0] m241_22;
   assign m241_22 =15'b0;

   // m241_23 = W*in
   wire signed [14:0] m241_23;
   assign m241_23 =15'b0;

   // m241_24 = W*in
   wire signed [14:0] m241_24;
   assign m241_24 =15'b0;

   // m241_25 = W*in
   wire signed [14:0] m241_25;
   assign m241_25 =15'b0;

   // m241_26 = W*in
   wire signed [14:0] m241_26;
   assign m241_26 =15'b0;

   // m241_27 = W*in
   wire signed [14:0] m241_27;
   assign m241_27 =15'b0;

   // m241_28 = W*in
   wire signed [14:0] m241_28;
   assign m241_28 =15'b0;

   // m241_29 = W*in
   wire signed [14:0] m241_29;
   assign m241_29 =15'b0;

   // m241_30 = W*in
   wire signed [14:0] m241_30;
   assign m241_30 =15'b0;

   // m241_31 = W*in
   wire signed [14:0] m241_31;
   assign m241_31 =15'b0;

   // m241_32 = W*in
   wire signed [14:0] m241_32;
   assign m241_32 =15'b0;

   // m241_33 = W*in
   wire signed [14:0] m241_33;
   assign m241_33 =15'b0;

   // m241_34 = W*in
   wire signed [14:0] m241_34;
   assign m241_34 =15'b0;

   // m241_35 = W*in
   wire signed [14:0] m241_35;
   assign m241_35 =15'b0;

   // m241_36 = W*in
   wire signed [14:0] m241_36;
   assign m241_36 =15'b0;

   // m241_37 = W*in
   wire signed [14:0] m241_37;
   assign m241_37 =15'b0;

   // m241_38 = W*in
   wire signed [14:0] m241_38;
   assign m241_38 =15'b0;

   // m241_39 = W*in
   wire signed [14:0] m241_39;
   assign m241_39 =15'b0;

   // m241_40 = W*in
   wire signed [14:0] m241_40;
   assign m241_40 =15'b0;

   // m241_41 = W*in
   wire signed [14:0] m241_41;
   assign m241_41 =15'b0;

   // m241_42 = W*in
   wire signed [14:0] m241_42;
   assign m241_42 =15'b0;

   // m241_43 = W*in
   wire signed [14:0] m241_43;
   assign m241_43 =15'b0;

   // m241_44 = W*in
   wire signed [14:0] m241_44;
   assign m241_44 ={ {4{neg241[14]}} , neg241[14:4] };

   // m241_45 = W*in
   wire signed [14:0] m241_45;
   assign m241_45 =15'b0;

   // m241_46 = W*in
   wire signed [14:0] m241_46;
   assign m241_46 ={ {4{neg241[14]}} , neg241[14:4] };

   // m241_47 = W*in
   wire signed [14:0] m241_47;
   assign m241_47 =15'b0;

   // m241_48 = W*in
   wire signed [14:0] m241_48;
   assign m241_48 ={ {4{neg241[14]}} , neg241[14:4] };

   // m241_49 = W*in
   wire signed [14:0] m241_49;
   assign m241_49 =15'b0;

   // m241_50 = W*in
   wire signed [14:0] m241_50;
   assign m241_50 =15'b0;

   // m241_51 = W*in
   wire signed [14:0] m241_51;
   assign m241_51 =15'b0;

   // m241_52 = W*in
   wire signed [14:0] m241_52;
   assign m241_52 ={ {3{in241[14]}} , in241[14:3] };

   // m241_53 = W*in
   wire signed [14:0] m241_53;
   assign m241_53 =15'b0;

   // m241_54 = W*in
   wire signed [14:0] m241_54;
   assign m241_54 =15'b0;

   // m241_55 = W*in
   wire signed [14:0] m241_55;
   assign m241_55 =15'b0;

   // m241_56 = W*in
   wire signed [14:0] m241_56;
   assign m241_56 =15'b0;

   // m241_57 = W*in
   wire signed [14:0] m241_57;
   assign m241_57 =15'b0;

   // m241_58 = W*in
   wire signed [14:0] m241_58;
   assign m241_58 ={ {4{in241[14]}} , in241[14:4] };

   // m241_59 = W*in
   wire signed [14:0] m241_59;
   assign m241_59 =15'b0;

   // m241_60 = W*in
   wire signed [14:0] m241_60;
   assign m241_60 ={ {3{neg241[14]}} , neg241[14:3] };

   // m241_61 = W*in
   wire signed [14:0] m241_61;
   assign m241_61 =15'b0;

   // m241_62 = W*in
   wire signed [14:0] m241_62;
   assign m241_62 =15'b0;

   // m241_63 = W*in
   wire signed [14:0] m241_63;
   assign m241_63 =15'b0;

   // m241_64 = W*in
   wire signed [14:0] m241_64;
   assign m241_64 =15'b0;

   // m241_65 = W*in
   wire signed [14:0] m241_65;
   assign m241_65 =15'b0;

   // m241_66 = W*in
   wire signed [14:0] m241_66;
   assign m241_66 =15'b0;

   // m241_67 = W*in
   wire signed [14:0] m241_67;
   assign m241_67 ={ {4{in241[14]}} , in241[14:4] };

   // m241_68 = W*in
   wire signed [14:0] m241_68;
   assign m241_68 =15'b0;

   // m241_69 = W*in
   wire signed [14:0] m241_69;
   assign m241_69 =15'b0;

   // m241_70 = W*in
   wire signed [14:0] m241_70;
   assign m241_70 =15'b0;

   // m241_71 = W*in
   wire signed [14:0] m241_71;
   assign m241_71 =15'b0;

   // m241_72 = W*in
   wire signed [14:0] m241_72;
   assign m241_72 =15'b0;

   // m241_73 = W*in
   wire signed [14:0] m241_73;
   assign m241_73 =15'b0;

   // m241_74 = W*in
   wire signed [14:0] m241_74;
   assign m241_74 ={ {3{neg241[14]}} , neg241[14:3] };

   // m241_75 = W*in
   wire signed [14:0] m241_75;
   assign m241_75 =15'b0;

   // m241_76 = W*in
   wire signed [14:0] m241_76;
   assign m241_76 ={ {3{neg241[14]}} , neg241[14:3] };

   // m241_77 = W*in
   wire signed [14:0] m241_77;
   assign m241_77 ={ {3{neg241[14]}} , neg241[14:3] };

   // m241_78 = W*in
   wire signed [14:0] m241_78;
   assign m241_78 =15'b0;

   // m241_79 = W*in
   wire signed [14:0] m241_79;
   assign m241_79 =15'b0;

   // m241_80 = W*in
   wire signed [14:0] m241_80;
   assign m241_80 =15'b0;

   // m241_81 = W*in
   wire signed [14:0] m241_81;
   assign m241_81 =15'b0;

   // m241_82 = W*in
   wire signed [14:0] m241_82;
   assign m241_82 =15'b0;

   // m241_83 = W*in
   wire signed [14:0] m241_83;
   assign m241_83 =15'b0;

   // m241_84 = W*in
   wire signed [14:0] m241_84;
   assign m241_84 =15'b0;

   // m241_85 = W*in
   wire signed [14:0] m241_85;
   assign m241_85 ={ {4{in241[14]}} , in241[14:4] };

   // m241_86 = W*in
   wire signed [14:0] m241_86;
   assign m241_86 =15'b0;

   // m241_87 = W*in
   wire signed [14:0] m241_87;
   assign m241_87 =15'b0;

   // m241_88 = W*in
   wire signed [14:0] m241_88;
   assign m241_88 =15'b0;

   // m241_89 = W*in
   wire signed [14:0] m241_89;
   assign m241_89 =15'b0;

   // m241_90 = W*in
   wire signed [14:0] m241_90;
   assign m241_90 =15'b0;

   // m241_91 = W*in
   wire signed [14:0] m241_91;
   assign m241_91 =15'b0;

   // m241_92 = W*in
   wire signed [14:0] m241_92;
   assign m241_92 =15'b0;

   // m241_93 = W*in
   wire signed [14:0] m241_93;
   assign m241_93 =15'b0;

   // m241_94 = W*in
   wire signed [14:0] m241_94;
   assign m241_94 =15'b0;

   // m241_95 = W*in
   wire signed [14:0] m241_95;
   assign m241_95 =15'b0;

   // m241_96 = W*in
   wire signed [14:0] m241_96;
   assign m241_96 =15'b0;

   // m241_97 = W*in
   wire signed [14:0] m241_97;
   assign m241_97 =15'b0;

   // m241_98 = W*in
   wire signed [14:0] m241_98;
   assign m241_98 =15'b0;

   // m241_99 = W*in
   wire signed [14:0] m241_99;
   assign m241_99 =15'b0;

   // m241_100 = W*in
   wire signed [14:0] m241_100;
   assign m241_100 =15'b0;

   // m242_1 = W*in
   wire signed [14:0] m242_1;
   assign m242_1 =15'b0;

   // m242_2 = W*in
   wire signed [14:0] m242_2;
   assign m242_2 =15'b0;

   // m242_3 = W*in
   wire signed [14:0] m242_3;
   assign m242_3 =15'b0;

   // m242_4 = W*in
   wire signed [14:0] m242_4;
   assign m242_4 =15'b0;

   // m242_5 = W*in
   wire signed [14:0] m242_5;
   assign m242_5 =15'b0;

   // m242_6 = W*in
   wire signed [14:0] m242_6;
   assign m242_6 =15'b0;

   // m242_7 = W*in
   wire signed [14:0] m242_7;
   assign m242_7 =15'b0;

   // m242_8 = W*in
   wire signed [14:0] m242_8;
   assign m242_8 =15'b0;

   // m242_9 = W*in
   wire signed [14:0] m242_9;
   assign m242_9 =15'b0;

   // m242_10 = W*in
   wire signed [14:0] m242_10;
   assign m242_10 =15'b0;

   // m242_11 = W*in
   wire signed [14:0] m242_11;
   assign m242_11 =15'b0;

   // m242_12 = W*in
   wire signed [14:0] m242_12;
   assign m242_12 =15'b0;

   // m242_13 = W*in
   wire signed [14:0] m242_13;
   assign m242_13 ={ {3{neg242[14]}} , neg242[14:3] };

   // m242_14 = W*in
   wire signed [14:0] m242_14;
   assign m242_14 =15'b0;

   // m242_15 = W*in
   wire signed [14:0] m242_15;
   assign m242_15 ={ {3{in242[14]}} , in242[14:3] };

   // m242_16 = W*in
   wire signed [14:0] m242_16;
   assign m242_16 =15'b0;

   // m242_17 = W*in
   wire signed [14:0] m242_17;
   assign m242_17 =15'b0;

   // m242_18 = W*in
   wire signed [14:0] m242_18;
   assign m242_18 =15'b0;

   // m242_19 = W*in
   wire signed [14:0] m242_19;
   assign m242_19 =15'b0;

   // m242_20 = W*in
   wire signed [14:0] m242_20;
   assign m242_20 ={ {3{neg242[14]}} , neg242[14:3] };

   // m242_21 = W*in
   wire signed [14:0] m242_21;
   assign m242_21 ={ {4{neg242[14]}} , neg242[14:4] };

   // m242_22 = W*in
   wire signed [14:0] m242_22;
   assign m242_22 =15'b0;

   // m242_23 = W*in
   wire signed [14:0] m242_23;
   assign m242_23 =15'b0;

   // m242_24 = W*in
   wire signed [14:0] m242_24;
   assign m242_24 =15'b0;

   // m242_25 = W*in
   wire signed [14:0] m242_25;
   assign m242_25 =15'b0;

   // m242_26 = W*in
   wire signed [14:0] m242_26;
   assign m242_26 =15'b0;

   // m242_27 = W*in
   wire signed [14:0] m242_27;
   assign m242_27 =15'b0;

   // m242_28 = W*in
   wire signed [14:0] m242_28;
   assign m242_28 =15'b0;

   // m242_29 = W*in
   wire signed [14:0] m242_29;
   assign m242_29 =15'b0;

   // m242_30 = W*in
   wire signed [14:0] m242_30;
   assign m242_30 ={ {3{in242[14]}} , in242[14:3] };

   // m242_31 = W*in
   wire signed [14:0] m242_31;
   assign m242_31 =15'b0;

   // m242_32 = W*in
   wire signed [14:0] m242_32;
   assign m242_32 ={ {4{neg242[14]}} , neg242[14:4] };

   // m242_33 = W*in
   wire signed [14:0] m242_33;
   assign m242_33 =15'b0;

   // m242_34 = W*in
   wire signed [14:0] m242_34;
   assign m242_34 =15'b0;

   // m242_35 = W*in
   wire signed [14:0] m242_35;
   assign m242_35 =15'b0;

   // m242_36 = W*in
   wire signed [14:0] m242_36;
   assign m242_36 =15'b0;

   // m242_37 = W*in
   wire signed [14:0] m242_37;
   assign m242_37 =15'b0;

   // m242_38 = W*in
   wire signed [14:0] m242_38;
   assign m242_38 =15'b0;

   // m242_39 = W*in
   wire signed [14:0] m242_39;
   assign m242_39 =15'b0;

   // m242_40 = W*in
   wire signed [14:0] m242_40;
   assign m242_40 =15'b0;

   // m242_41 = W*in
   wire signed [14:0] m242_41;
   assign m242_41 ={ {3{in242[14]}} , in242[14:3] };

   // m242_42 = W*in
   wire signed [14:0] m242_42;
   assign m242_42 =15'b0;

   // m242_43 = W*in
   wire signed [14:0] m242_43;
   assign m242_43 =15'b0;

   // m242_44 = W*in
   wire signed [14:0] m242_44;
   assign m242_44 =15'b0;

   // m242_45 = W*in
   wire signed [14:0] m242_45;
   assign m242_45 =15'b0;

   // m242_46 = W*in
   wire signed [14:0] m242_46;
   assign m242_46 =15'b0;

   // m242_47 = W*in
   wire signed [14:0] m242_47;
   assign m242_47 =15'b0;

   // m242_48 = W*in
   wire signed [14:0] m242_48;
   assign m242_48 =15'b0;

   // m242_49 = W*in
   wire signed [14:0] m242_49;
   assign m242_49 =15'b0;

   // m242_50 = W*in
   wire signed [14:0] m242_50;
   assign m242_50 ={ {3{in242[14]}} , in242[14:3] };

   // m242_51 = W*in
   wire signed [14:0] m242_51;
   assign m242_51 =15'b0;

   // m242_52 = W*in
   wire signed [14:0] m242_52;
   assign m242_52 =15'b0;

   // m242_53 = W*in
   wire signed [14:0] m242_53;
   assign m242_53 =15'b0;

   // m242_54 = W*in
   wire signed [14:0] m242_54;
   assign m242_54 =15'b0;

   // m242_55 = W*in
   wire signed [14:0] m242_55;
   assign m242_55 =15'b0;

   // m242_56 = W*in
   wire signed [14:0] m242_56;
   assign m242_56 =15'b0;

   // m242_57 = W*in
   wire signed [14:0] m242_57;
   assign m242_57 ={ {3{neg242[14]}} , neg242[14:3] };

   // m242_58 = W*in
   wire signed [14:0] m242_58;
   assign m242_58 =15'b0;

   // m242_59 = W*in
   wire signed [14:0] m242_59;
   assign m242_59 =15'b0;

   // m242_60 = W*in
   wire signed [14:0] m242_60;
   assign m242_60 =15'b0;

   // m242_61 = W*in
   wire signed [14:0] m242_61;
   assign m242_61 =15'b0;

   // m242_62 = W*in
   wire signed [14:0] m242_62;
   assign m242_62 ={ {3{neg242[14]}} , neg242[14:3] };

   // m242_63 = W*in
   wire signed [14:0] m242_63;
   assign m242_63 =15'b0;

   // m242_64 = W*in
   wire signed [14:0] m242_64;
   assign m242_64 ={ {4{neg242[14]}} , neg242[14:4] };

   // m242_65 = W*in
   wire signed [14:0] m242_65;
   assign m242_65 =15'b0;

   // m242_66 = W*in
   wire signed [14:0] m242_66;
   assign m242_66 =15'b0;

   // m242_67 = W*in
   wire signed [14:0] m242_67;
   assign m242_67 ={ {3{in242[14]}} , in242[14:3] };

   // m242_68 = W*in
   wire signed [14:0] m242_68;
   assign m242_68 =15'b0;

   // m242_69 = W*in
   wire signed [14:0] m242_69;
   assign m242_69 =15'b0;

   // m242_70 = W*in
   wire signed [14:0] m242_70;
   assign m242_70 =15'b0;

   // m242_71 = W*in
   wire signed [14:0] m242_71;
   assign m242_71 =15'b0;

   // m242_72 = W*in
   wire signed [14:0] m242_72;
   assign m242_72 =15'b0;

   // m242_73 = W*in
   wire signed [14:0] m242_73;
   assign m242_73 =15'b0;

   // m242_74 = W*in
   wire signed [14:0] m242_74;
   assign m242_74 ={ {3{neg242[14]}} , neg242[14:3] };

   // m242_75 = W*in
   wire signed [14:0] m242_75;
   assign m242_75 =15'b0;

   // m242_76 = W*in
   wire signed [14:0] m242_76;
   assign m242_76 =15'b0;

   // m242_77 = W*in
   wire signed [14:0] m242_77;
   assign m242_77 ={ {3{in242[14]}} , in242[14:3] };

   // m242_78 = W*in
   wire signed [14:0] m242_78;
   assign m242_78 ={ {3{in242[14]}} , in242[14:3] };

   // m242_79 = W*in
   wire signed [14:0] m242_79;
   assign m242_79 =15'b0;

   // m242_80 = W*in
   wire signed [14:0] m242_80;
   assign m242_80 ={ {3{in242[14]}} , in242[14:3] };

   // m242_81 = W*in
   wire signed [14:0] m242_81;
   assign m242_81 =15'b0;

   // m242_82 = W*in
   wire signed [14:0] m242_82;
   assign m242_82 =15'b0;

   // m242_83 = W*in
   wire signed [14:0] m242_83;
   assign m242_83 =15'b0;

   // m242_84 = W*in
   wire signed [14:0] m242_84;
   assign m242_84 =15'b0;

   // m242_85 = W*in
   wire signed [14:0] m242_85;
   assign m242_85 =15'b0;

   // m242_86 = W*in
   wire signed [14:0] m242_86;
   assign m242_86 =15'b0;

   // m242_87 = W*in
   wire signed [14:0] m242_87;
   assign m242_87 ={ {3{neg242[14]}} , neg242[14:3] };

   // m242_88 = W*in
   wire signed [14:0] m242_88;
   assign m242_88 =15'b0;

   // m242_89 = W*in
   wire signed [14:0] m242_89;
   assign m242_89 =15'b0;

   // m242_90 = W*in
   wire signed [14:0] m242_90;
   assign m242_90 =15'b0;

   // m242_91 = W*in
   wire signed [14:0] m242_91;
   assign m242_91 =15'b0;

   // m242_92 = W*in
   wire signed [14:0] m242_92;
   assign m242_92 =15'b0;

   // m242_93 = W*in
   wire signed [14:0] m242_93;
   assign m242_93 =15'b0;

   // m242_94 = W*in
   wire signed [14:0] m242_94;
   assign m242_94 =15'b0;

   // m242_95 = W*in
   wire signed [14:0] m242_95;
   assign m242_95 =15'b0;

   // m242_96 = W*in
   wire signed [14:0] m242_96;
   assign m242_96 =15'b0;

   // m242_97 = W*in
   wire signed [14:0] m242_97;
   assign m242_97 =15'b0;

   // m242_98 = W*in
   wire signed [14:0] m242_98;
   assign m242_98 =15'b0;

   // m242_99 = W*in
   wire signed [14:0] m242_99;
   assign m242_99 =15'b0;

   // m242_100 = W*in
   wire signed [14:0] m242_100;
   assign m242_100 =15'b0;

   // m243_1 = W*in
   wire signed [14:0] m243_1;
   assign m243_1 =15'b0;

   // m243_2 = W*in
   wire signed [14:0] m243_2;
   assign m243_2 ={ {3{in243[14]}} , in243[14:3] };

   // m243_3 = W*in
   wire signed [14:0] m243_3;
   assign m243_3 =15'b0;

   // m243_4 = W*in
   wire signed [14:0] m243_4;
   assign m243_4 =15'b0;

   // m243_5 = W*in
   wire signed [14:0] m243_5;
   assign m243_5 =15'b0;

   // m243_6 = W*in
   wire signed [14:0] m243_6;
   assign m243_6 =15'b0;

   // m243_7 = W*in
   wire signed [14:0] m243_7;
   assign m243_7 =15'b0;

   // m243_8 = W*in
   wire signed [14:0] m243_8;
   assign m243_8 =15'b0;

   // m243_9 = W*in
   wire signed [14:0] m243_9;
   assign m243_9 =15'b0;

   // m243_10 = W*in
   wire signed [14:0] m243_10;
   assign m243_10 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_11 = W*in
   wire signed [14:0] m243_11;
   assign m243_11 =15'b0;

   // m243_12 = W*in
   wire signed [14:0] m243_12;
   assign m243_12 =15'b0;

   // m243_13 = W*in
   wire signed [14:0] m243_13;
   assign m243_13 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_14 = W*in
   wire signed [14:0] m243_14;
   assign m243_14 =15'b0;

   // m243_15 = W*in
   wire signed [14:0] m243_15;
   assign m243_15 =15'b0;

   // m243_16 = W*in
   wire signed [14:0] m243_16;
   assign m243_16 =15'b0;

   // m243_17 = W*in
   wire signed [14:0] m243_17;
   assign m243_17 =15'b0;

   // m243_18 = W*in
   wire signed [14:0] m243_18;
   assign m243_18 =15'b0;

   // m243_19 = W*in
   wire signed [14:0] m243_19;
   assign m243_19 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_20 = W*in
   wire signed [14:0] m243_20;
   assign m243_20 =15'b0;

   // m243_21 = W*in
   wire signed [14:0] m243_21;
   assign m243_21 ={ {3{in243[14]}} , in243[14:3] };

   // m243_22 = W*in
   wire signed [14:0] m243_22;
   assign m243_22 =15'b0;

   // m243_23 = W*in
   wire signed [14:0] m243_23;
   assign m243_23 =15'b0;

   // m243_24 = W*in
   wire signed [14:0] m243_24;
   assign m243_24 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_25 = W*in
   wire signed [14:0] m243_25;
   assign m243_25 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_26 = W*in
   wire signed [14:0] m243_26;
   assign m243_26 =15'b0;

   // m243_27 = W*in
   wire signed [14:0] m243_27;
   assign m243_27 =15'b0;

   // m243_28 = W*in
   wire signed [14:0] m243_28;
   assign m243_28 =15'b0;

   // m243_29 = W*in
   wire signed [14:0] m243_29;
   assign m243_29 =15'b0;

   // m243_30 = W*in
   wire signed [14:0] m243_30;
   assign m243_30 =15'b0;

   // m243_31 = W*in
   wire signed [14:0] m243_31;
   assign m243_31 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_32 = W*in
   wire signed [14:0] m243_32;
   assign m243_32 =15'b0;

   // m243_33 = W*in
   wire signed [14:0] m243_33;
   assign m243_33 =15'b0;

   // m243_34 = W*in
   wire signed [14:0] m243_34;
   assign m243_34 =15'b0;

   // m243_35 = W*in
   wire signed [14:0] m243_35;
   assign m243_35 ={ {3{in243[14]}} , in243[14:3] };

   // m243_36 = W*in
   wire signed [14:0] m243_36;
   assign m243_36 =15'b0;

   // m243_37 = W*in
   wire signed [14:0] m243_37;
   assign m243_37 =15'b0;

   // m243_38 = W*in
   wire signed [14:0] m243_38;
   assign m243_38 =15'b0;

   // m243_39 = W*in
   wire signed [14:0] m243_39;
   assign m243_39 =15'b0;

   // m243_40 = W*in
   wire signed [14:0] m243_40;
   assign m243_40 ={ {2{in243[14]}} , in243[14:2] };

   // m243_41 = W*in
   wire signed [14:0] m243_41;
   assign m243_41 =15'b0;

   // m243_42 = W*in
   wire signed [14:0] m243_42;
   assign m243_42 =15'b0;

   // m243_43 = W*in
   wire signed [14:0] m243_43;
   assign m243_43 =15'b0;

   // m243_44 = W*in
   wire signed [14:0] m243_44;
   assign m243_44 =15'b0;

   // m243_45 = W*in
   wire signed [14:0] m243_45;
   assign m243_45 ={ {3{in243[14]}} , in243[14:3] };

   // m243_46 = W*in
   wire signed [14:0] m243_46;
   assign m243_46 ={ {4{neg243[14]}} , neg243[14:4] };

   // m243_47 = W*in
   wire signed [14:0] m243_47;
   assign m243_47 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_48 = W*in
   wire signed [14:0] m243_48;
   assign m243_48 =15'b0;

   // m243_49 = W*in
   wire signed [14:0] m243_49;
   assign m243_49 =15'b0;

   // m243_50 = W*in
   wire signed [14:0] m243_50;
   assign m243_50 =15'b0;

   // m243_51 = W*in
   wire signed [14:0] m243_51;
   assign m243_51 =15'b0;

   // m243_52 = W*in
   wire signed [14:0] m243_52;
   assign m243_52 =15'b0;

   // m243_53 = W*in
   wire signed [14:0] m243_53;
   assign m243_53 =15'b0;

   // m243_54 = W*in
   wire signed [14:0] m243_54;
   assign m243_54 =15'b0;

   // m243_55 = W*in
   wire signed [14:0] m243_55;
   assign m243_55 =15'b0;

   // m243_56 = W*in
   wire signed [14:0] m243_56;
   assign m243_56 =15'b0;

   // m243_57 = W*in
   wire signed [14:0] m243_57;
   assign m243_57 =15'b0;

   // m243_58 = W*in
   wire signed [14:0] m243_58;
   assign m243_58 =15'b0;

   // m243_59 = W*in
   wire signed [14:0] m243_59;
   assign m243_59 ={ {4{neg243[14]}} , neg243[14:4] };

   // m243_60 = W*in
   wire signed [14:0] m243_60;
   assign m243_60 =15'b0;

   // m243_61 = W*in
   wire signed [14:0] m243_61;
   assign m243_61 =15'b0;

   // m243_62 = W*in
   wire signed [14:0] m243_62;
   assign m243_62 =15'b0;

   // m243_63 = W*in
   wire signed [14:0] m243_63;
   assign m243_63 =15'b0;

   // m243_64 = W*in
   wire signed [14:0] m243_64;
   assign m243_64 =15'b0;

   // m243_65 = W*in
   wire signed [14:0] m243_65;
   assign m243_65 =15'b0;

   // m243_66 = W*in
   wire signed [14:0] m243_66;
   assign m243_66 =15'b0;

   // m243_67 = W*in
   wire signed [14:0] m243_67;
   assign m243_67 =15'b0;

   // m243_68 = W*in
   wire signed [14:0] m243_68;
   assign m243_68 =15'b0;

   // m243_69 = W*in
   wire signed [14:0] m243_69;
   assign m243_69 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_70 = W*in
   wire signed [14:0] m243_70;
   assign m243_70 =15'b0;

   // m243_71 = W*in
   wire signed [14:0] m243_71;
   assign m243_71 =15'b0;

   // m243_72 = W*in
   wire signed [14:0] m243_72;
   assign m243_72 =15'b0;

   // m243_73 = W*in
   wire signed [14:0] m243_73;
   assign m243_73 =15'b0;

   // m243_74 = W*in
   wire signed [14:0] m243_74;
   assign m243_74 ={ {3{in243[14]}} , in243[14:3] };

   // m243_75 = W*in
   wire signed [14:0] m243_75;
   assign m243_75 =15'b0;

   // m243_76 = W*in
   wire signed [14:0] m243_76;
   assign m243_76 =15'b0;

   // m243_77 = W*in
   wire signed [14:0] m243_77;
   assign m243_77 =15'b0;

   // m243_78 = W*in
   wire signed [14:0] m243_78;
   assign m243_78 ={ {3{in243[14]}} , in243[14:3] };

   // m243_79 = W*in
   wire signed [14:0] m243_79;
   assign m243_79 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_80 = W*in
   wire signed [14:0] m243_80;
   assign m243_80 =15'b0;

   // m243_81 = W*in
   wire signed [14:0] m243_81;
   assign m243_81 =15'b0;

   // m243_82 = W*in
   wire signed [14:0] m243_82;
   assign m243_82 =15'b0;

   // m243_83 = W*in
   wire signed [14:0] m243_83;
   assign m243_83 =15'b0;

   // m243_84 = W*in
   wire signed [14:0] m243_84;
   assign m243_84 =15'b0;

   // m243_85 = W*in
   wire signed [14:0] m243_85;
   assign m243_85 =15'b0;

   // m243_86 = W*in
   wire signed [14:0] m243_86;
   assign m243_86 =15'b0;

   // m243_87 = W*in
   wire signed [14:0] m243_87;
   assign m243_87 =15'b0;

   // m243_88 = W*in
   wire signed [14:0] m243_88;
   assign m243_88 =15'b0;

   // m243_89 = W*in
   wire signed [14:0] m243_89;
   assign m243_89 =15'b0;

   // m243_90 = W*in
   wire signed [14:0] m243_90;
   assign m243_90 ={ {3{in243[14]}} , in243[14:3] };

   // m243_91 = W*in
   wire signed [14:0] m243_91;
   assign m243_91 =15'b0;

   // m243_92 = W*in
   wire signed [14:0] m243_92;
   assign m243_92 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_93 = W*in
   wire signed [14:0] m243_93;
   assign m243_93 =15'b0;

   // m243_94 = W*in
   wire signed [14:0] m243_94;
   assign m243_94 ={ {3{neg243[14]}} , neg243[14:3] };

   // m243_95 = W*in
   wire signed [14:0] m243_95;
   assign m243_95 =15'b0;

   // m243_96 = W*in
   wire signed [14:0] m243_96;
   assign m243_96 =15'b0;

   // m243_97 = W*in
   wire signed [14:0] m243_97;
   assign m243_97 =15'b0;

   // m243_98 = W*in
   wire signed [14:0] m243_98;
   assign m243_98 =15'b0;

   // m243_99 = W*in
   wire signed [14:0] m243_99;
   assign m243_99 =15'b0;

   // m243_100 = W*in
   wire signed [14:0] m243_100;
   assign m243_100 =15'b0;

   // m244_1 = W*in
   wire signed [14:0] m244_1;
   assign m244_1 =15'b0;

   // m244_2 = W*in
   wire signed [14:0] m244_2;
   assign m244_2 =15'b0;

   // m244_3 = W*in
   wire signed [14:0] m244_3;
   assign m244_3 =15'b0;

   // m244_4 = W*in
   wire signed [14:0] m244_4;
   assign m244_4 =15'b0;

   // m244_5 = W*in
   wire signed [14:0] m244_5;
   assign m244_5 =15'b0;

   // m244_6 = W*in
   wire signed [14:0] m244_6;
   assign m244_6 =15'b0;

   // m244_7 = W*in
   wire signed [14:0] m244_7;
   assign m244_7 =15'b0;

   // m244_8 = W*in
   wire signed [14:0] m244_8;
   assign m244_8 =15'b0;

   // m244_9 = W*in
   wire signed [14:0] m244_9;
   assign m244_9 =15'b0;

   // m244_10 = W*in
   wire signed [14:0] m244_10;
   assign m244_10 =15'b0;

   // m244_11 = W*in
   wire signed [14:0] m244_11;
   assign m244_11 =15'b0;

   // m244_12 = W*in
   wire signed [14:0] m244_12;
   assign m244_12 =15'b0;

   // m244_13 = W*in
   wire signed [14:0] m244_13;
   assign m244_13 =15'b0;

   // m244_14 = W*in
   wire signed [14:0] m244_14;
   assign m244_14 =15'b0;

   // m244_15 = W*in
   wire signed [14:0] m244_15;
   assign m244_15 =15'b0;

   // m244_16 = W*in
   wire signed [14:0] m244_16;
   assign m244_16 =15'b0;

   // m244_17 = W*in
   wire signed [14:0] m244_17;
   assign m244_17 =15'b0;

   // m244_18 = W*in
   wire signed [14:0] m244_18;
   assign m244_18 =15'b0;

   // m244_19 = W*in
   wire signed [14:0] m244_19;
   assign m244_19 =15'b0;

   // m244_20 = W*in
   wire signed [14:0] m244_20;
   assign m244_20 ={ {4{in244[14]}} , in244[14:4] };

   // m244_21 = W*in
   wire signed [14:0] m244_21;
   assign m244_21 =15'b0;

   // m244_22 = W*in
   wire signed [14:0] m244_22;
   assign m244_22 =15'b0;

   // m244_23 = W*in
   wire signed [14:0] m244_23;
   assign m244_23 =15'b0;

   // m244_24 = W*in
   wire signed [14:0] m244_24;
   assign m244_24 =15'b0;

   // m244_25 = W*in
   wire signed [14:0] m244_25;
   assign m244_25 =15'b0;

   // m244_26 = W*in
   wire signed [14:0] m244_26;
   assign m244_26 =15'b0;

   // m244_27 = W*in
   wire signed [14:0] m244_27;
   assign m244_27 =15'b0;

   // m244_28 = W*in
   wire signed [14:0] m244_28;
   assign m244_28 =15'b0;

   // m244_29 = W*in
   wire signed [14:0] m244_29;
   assign m244_29 =15'b0;

   // m244_30 = W*in
   wire signed [14:0] m244_30;
   assign m244_30 =15'b0;

   // m244_31 = W*in
   wire signed [14:0] m244_31;
   assign m244_31 =15'b0;

   // m244_32 = W*in
   wire signed [14:0] m244_32;
   assign m244_32 =15'b0;

   // m244_33 = W*in
   wire signed [14:0] m244_33;
   assign m244_33 =15'b0;

   // m244_34 = W*in
   wire signed [14:0] m244_34;
   assign m244_34 =15'b0;

   // m244_35 = W*in
   wire signed [14:0] m244_35;
   assign m244_35 =15'b0;

   // m244_36 = W*in
   wire signed [14:0] m244_36;
   assign m244_36 =15'b0;

   // m244_37 = W*in
   wire signed [14:0] m244_37;
   assign m244_37 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_38 = W*in
   wire signed [14:0] m244_38;
   assign m244_38 =15'b0;

   // m244_39 = W*in
   wire signed [14:0] m244_39;
   assign m244_39 =15'b0;

   // m244_40 = W*in
   wire signed [14:0] m244_40;
   assign m244_40 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_41 = W*in
   wire signed [14:0] m244_41;
   assign m244_41 =15'b0;

   // m244_42 = W*in
   wire signed [14:0] m244_42;
   assign m244_42 =15'b0;

   // m244_43 = W*in
   wire signed [14:0] m244_43;
   assign m244_43 =15'b0;

   // m244_44 = W*in
   wire signed [14:0] m244_44;
   assign m244_44 =15'b0;

   // m244_45 = W*in
   wire signed [14:0] m244_45;
   assign m244_45 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_46 = W*in
   wire signed [14:0] m244_46;
   assign m244_46 =15'b0;

   // m244_47 = W*in
   wire signed [14:0] m244_47;
   assign m244_47 =15'b0;

   // m244_48 = W*in
   wire signed [14:0] m244_48;
   assign m244_48 =15'b0;

   // m244_49 = W*in
   wire signed [14:0] m244_49;
   assign m244_49 =15'b0;

   // m244_50 = W*in
   wire signed [14:0] m244_50;
   assign m244_50 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_51 = W*in
   wire signed [14:0] m244_51;
   assign m244_51 ={ {4{neg244[14]}} , neg244[14:4] };

   // m244_52 = W*in
   wire signed [14:0] m244_52;
   assign m244_52 =15'b0;

   // m244_53 = W*in
   wire signed [14:0] m244_53;
   assign m244_53 =15'b0;

   // m244_54 = W*in
   wire signed [14:0] m244_54;
   assign m244_54 =15'b0;

   // m244_55 = W*in
   wire signed [14:0] m244_55;
   assign m244_55 =15'b0;

   // m244_56 = W*in
   wire signed [14:0] m244_56;
   assign m244_56 =15'b0;

   // m244_57 = W*in
   wire signed [14:0] m244_57;
   assign m244_57 =15'b0;

   // m244_58 = W*in
   wire signed [14:0] m244_58;
   assign m244_58 ={ {3{in244[14]}} , in244[14:3] };

   // m244_59 = W*in
   wire signed [14:0] m244_59;
   assign m244_59 =15'b0;

   // m244_60 = W*in
   wire signed [14:0] m244_60;
   assign m244_60 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_61 = W*in
   wire signed [14:0] m244_61;
   assign m244_61 =15'b0;

   // m244_62 = W*in
   wire signed [14:0] m244_62;
   assign m244_62 =15'b0;

   // m244_63 = W*in
   wire signed [14:0] m244_63;
   assign m244_63 =15'b0;

   // m244_64 = W*in
   wire signed [14:0] m244_64;
   assign m244_64 =15'b0;

   // m244_65 = W*in
   wire signed [14:0] m244_65;
   assign m244_65 =15'b0;

   // m244_66 = W*in
   wire signed [14:0] m244_66;
   assign m244_66 =15'b0;

   // m244_67 = W*in
   wire signed [14:0] m244_67;
   assign m244_67 =15'b0;

   // m244_68 = W*in
   wire signed [14:0] m244_68;
   assign m244_68 =15'b0;

   // m244_69 = W*in
   wire signed [14:0] m244_69;
   assign m244_69 =15'b0;

   // m244_70 = W*in
   wire signed [14:0] m244_70;
   assign m244_70 =15'b0;

   // m244_71 = W*in
   wire signed [14:0] m244_71;
   assign m244_71 =15'b0;

   // m244_72 = W*in
   wire signed [14:0] m244_72;
   assign m244_72 =15'b0;

   // m244_73 = W*in
   wire signed [14:0] m244_73;
   assign m244_73 =15'b0;

   // m244_74 = W*in
   wire signed [14:0] m244_74;
   assign m244_74 ={ {4{in244[14]}} , in244[14:4] };

   // m244_75 = W*in
   wire signed [14:0] m244_75;
   assign m244_75 ={ {3{in244[14]}} , in244[14:3] };

   // m244_76 = W*in
   wire signed [14:0] m244_76;
   assign m244_76 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_77 = W*in
   wire signed [14:0] m244_77;
   assign m244_77 =15'b0;

   // m244_78 = W*in
   wire signed [14:0] m244_78;
   assign m244_78 =15'b0;

   // m244_79 = W*in
   wire signed [14:0] m244_79;
   assign m244_79 =15'b0;

   // m244_80 = W*in
   wire signed [14:0] m244_80;
   assign m244_80 =15'b0;

   // m244_81 = W*in
   wire signed [14:0] m244_81;
   assign m244_81 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_82 = W*in
   wire signed [14:0] m244_82;
   assign m244_82 =15'b0;

   // m244_83 = W*in
   wire signed [14:0] m244_83;
   assign m244_83 =15'b0;

   // m244_84 = W*in
   wire signed [14:0] m244_84;
   assign m244_84 =15'b0;

   // m244_85 = W*in
   wire signed [14:0] m244_85;
   assign m244_85 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_86 = W*in
   wire signed [14:0] m244_86;
   assign m244_86 =15'b0;

   // m244_87 = W*in
   wire signed [14:0] m244_87;
   assign m244_87 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_88 = W*in
   wire signed [14:0] m244_88;
   assign m244_88 ={ {3{in244[14]}} , in244[14:3] };

   // m244_89 = W*in
   wire signed [14:0] m244_89;
   assign m244_89 ={ {3{neg244[14]}} , neg244[14:3] };

   // m244_90 = W*in
   wire signed [14:0] m244_90;
   assign m244_90 =15'b0;

   // m244_91 = W*in
   wire signed [14:0] m244_91;
   assign m244_91 ={ {4{neg244[14]}} , neg244[14:4] };

   // m244_92 = W*in
   wire signed [14:0] m244_92;
   assign m244_92 =15'b0;

   // m244_93 = W*in
   wire signed [14:0] m244_93;
   assign m244_93 =15'b0;

   // m244_94 = W*in
   wire signed [14:0] m244_94;
   assign m244_94 =15'b0;

   // m244_95 = W*in
   wire signed [14:0] m244_95;
   assign m244_95 =15'b0;

   // m244_96 = W*in
   wire signed [14:0] m244_96;
   assign m244_96 =15'b0;

   // m244_97 = W*in
   wire signed [14:0] m244_97;
   assign m244_97 =15'b0;

   // m244_98 = W*in
   wire signed [14:0] m244_98;
   assign m244_98 =15'b0;

   // m244_99 = W*in
   wire signed [14:0] m244_99;
   assign m244_99 =15'b0;

   // m244_100 = W*in
   wire signed [14:0] m244_100;
   assign m244_100 =15'b0;

   // m245_1 = W*in
   wire signed [14:0] m245_1;
   assign m245_1 =15'b0;

   // m245_2 = W*in
   wire signed [14:0] m245_2;
   assign m245_2 =15'b0;

   // m245_3 = W*in
   wire signed [14:0] m245_3;
   assign m245_3 ={ {3{neg245[14]}} , neg245[14:3] };

   // m245_4 = W*in
   wire signed [14:0] m245_4;
   assign m245_4 =15'b0;

   // m245_5 = W*in
   wire signed [14:0] m245_5;
   assign m245_5 =15'b0;

   // m245_6 = W*in
   wire signed [14:0] m245_6;
   assign m245_6 ={ {4{neg245[14]}} , neg245[14:4] };

   // m245_7 = W*in
   wire signed [14:0] m245_7;
   assign m245_7 =15'b0;

   // m245_8 = W*in
   wire signed [14:0] m245_8;
   assign m245_8 =15'b0;

   // m245_9 = W*in
   wire signed [14:0] m245_9;
   assign m245_9 =15'b0;

   // m245_10 = W*in
   wire signed [14:0] m245_10;
   assign m245_10 =15'b0;

   // m245_11 = W*in
   wire signed [14:0] m245_11;
   assign m245_11 =15'b0;

   // m245_12 = W*in
   wire signed [14:0] m245_12;
   assign m245_12 =15'b0;

   // m245_13 = W*in
   wire signed [14:0] m245_13;
   assign m245_13 =15'b0;

   // m245_14 = W*in
   wire signed [14:0] m245_14;
   assign m245_14 =15'b0;

   // m245_15 = W*in
   wire signed [14:0] m245_15;
   assign m245_15 =15'b0;

   // m245_16 = W*in
   wire signed [14:0] m245_16;
   assign m245_16 =15'b0;

   // m245_17 = W*in
   wire signed [14:0] m245_17;
   assign m245_17 =15'b0;

   // m245_18 = W*in
   wire signed [14:0] m245_18;
   assign m245_18 =15'b0;

   // m245_19 = W*in
   wire signed [14:0] m245_19;
   assign m245_19 =15'b0;

   // m245_20 = W*in
   wire signed [14:0] m245_20;
   assign m245_20 ={ {4{neg245[14]}} , neg245[14:4] };

   // m245_21 = W*in
   wire signed [14:0] m245_21;
   assign m245_21 =15'b0;

   // m245_22 = W*in
   wire signed [14:0] m245_22;
   assign m245_22 =15'b0;

   // m245_23 = W*in
   wire signed [14:0] m245_23;
   assign m245_23 =15'b0;

   // m245_24 = W*in
   wire signed [14:0] m245_24;
   assign m245_24 =15'b0;

   // m245_25 = W*in
   wire signed [14:0] m245_25;
   assign m245_25 =15'b0;

   // m245_26 = W*in
   wire signed [14:0] m245_26;
   assign m245_26 ={ {4{neg245[14]}} , neg245[14:4] };

   // m245_27 = W*in
   wire signed [14:0] m245_27;
   assign m245_27 =15'b0;

   // m245_28 = W*in
   wire signed [14:0] m245_28;
   assign m245_28 =15'b0;

   // m245_29 = W*in
   wire signed [14:0] m245_29;
   assign m245_29 =15'b0;

   // m245_30 = W*in
   wire signed [14:0] m245_30;
   assign m245_30 =15'b0;

   // m245_31 = W*in
   wire signed [14:0] m245_31;
   assign m245_31 =15'b0;

   // m245_32 = W*in
   wire signed [14:0] m245_32;
   assign m245_32 =15'b0;

   // m245_33 = W*in
   wire signed [14:0] m245_33;
   assign m245_33 =15'b0;

   // m245_34 = W*in
   wire signed [14:0] m245_34;
   assign m245_34 =15'b0;

   // m245_35 = W*in
   wire signed [14:0] m245_35;
   assign m245_35 =15'b0;

   // m245_36 = W*in
   wire signed [14:0] m245_36;
   assign m245_36 =15'b0;

   // m245_37 = W*in
   wire signed [14:0] m245_37;
   assign m245_37 ={ {4{in245[14]}} , in245[14:4] };

   // m245_38 = W*in
   wire signed [14:0] m245_38;
   assign m245_38 ={ {4{neg245[14]}} , neg245[14:4] };

   // m245_39 = W*in
   wire signed [14:0] m245_39;
   assign m245_39 ={ {3{in245[14]}} , in245[14:3] };

   // m245_40 = W*in
   wire signed [14:0] m245_40;
   assign m245_40 =15'b0;

   // m245_41 = W*in
   wire signed [14:0] m245_41;
   assign m245_41 =15'b0;

   // m245_42 = W*in
   wire signed [14:0] m245_42;
   assign m245_42 =15'b0;

   // m245_43 = W*in
   wire signed [14:0] m245_43;
   assign m245_43 =15'b0;

   // m245_44 = W*in
   wire signed [14:0] m245_44;
   assign m245_44 =15'b0;

   // m245_45 = W*in
   wire signed [14:0] m245_45;
   assign m245_45 =15'b0;

   // m245_46 = W*in
   wire signed [14:0] m245_46;
   assign m245_46 =15'b0;

   // m245_47 = W*in
   wire signed [14:0] m245_47;
   assign m245_47 =15'b0;

   // m245_48 = W*in
   wire signed [14:0] m245_48;
   assign m245_48 =15'b0;

   // m245_49 = W*in
   wire signed [14:0] m245_49;
   assign m245_49 =15'b0;

   // m245_50 = W*in
   wire signed [14:0] m245_50;
   assign m245_50 =15'b0;

   // m245_51 = W*in
   wire signed [14:0] m245_51;
   assign m245_51 =15'b0;

   // m245_52 = W*in
   wire signed [14:0] m245_52;
   assign m245_52 =15'b0;

   // m245_53 = W*in
   wire signed [14:0] m245_53;
   assign m245_53 =15'b0;

   // m245_54 = W*in
   wire signed [14:0] m245_54;
   assign m245_54 =15'b0;

   // m245_55 = W*in
   wire signed [14:0] m245_55;
   assign m245_55 ={ {3{neg245[14]}} , neg245[14:3] };

   // m245_56 = W*in
   wire signed [14:0] m245_56;
   assign m245_56 =15'b0;

   // m245_57 = W*in
   wire signed [14:0] m245_57;
   assign m245_57 =15'b0;

   // m245_58 = W*in
   wire signed [14:0] m245_58;
   assign m245_58 =15'b0;

   // m245_59 = W*in
   wire signed [14:0] m245_59;
   assign m245_59 ={ {3{neg245[14]}} , neg245[14:3] };

   // m245_60 = W*in
   wire signed [14:0] m245_60;
   assign m245_60 =15'b0;

   // m245_61 = W*in
   wire signed [14:0] m245_61;
   assign m245_61 =15'b0;

   // m245_62 = W*in
   wire signed [14:0] m245_62;
   assign m245_62 =15'b0;

   // m245_63 = W*in
   wire signed [14:0] m245_63;
   assign m245_63 =15'b0;

   // m245_64 = W*in
   wire signed [14:0] m245_64;
   assign m245_64 =15'b0;

   // m245_65 = W*in
   wire signed [14:0] m245_65;
   assign m245_65 =15'b0;

   // m245_66 = W*in
   wire signed [14:0] m245_66;
   assign m245_66 =15'b0;

   // m245_67 = W*in
   wire signed [14:0] m245_67;
   assign m245_67 =15'b0;

   // m245_68 = W*in
   wire signed [14:0] m245_68;
   assign m245_68 =15'b0;

   // m245_69 = W*in
   wire signed [14:0] m245_69;
   assign m245_69 =15'b0;

   // m245_70 = W*in
   wire signed [14:0] m245_70;
   assign m245_70 =15'b0;

   // m245_71 = W*in
   wire signed [14:0] m245_71;
   assign m245_71 =15'b0;

   // m245_72 = W*in
   wire signed [14:0] m245_72;
   assign m245_72 =15'b0;

   // m245_73 = W*in
   wire signed [14:0] m245_73;
   assign m245_73 =15'b0;

   // m245_74 = W*in
   wire signed [14:0] m245_74;
   assign m245_74 =15'b0;

   // m245_75 = W*in
   wire signed [14:0] m245_75;
   assign m245_75 =15'b0;

   // m245_76 = W*in
   wire signed [14:0] m245_76;
   assign m245_76 ={ {4{neg245[14]}} , neg245[14:4] };

   // m245_77 = W*in
   wire signed [14:0] m245_77;
   assign m245_77 =15'b0;

   // m245_78 = W*in
   wire signed [14:0] m245_78;
   assign m245_78 =15'b0;

   // m245_79 = W*in
   wire signed [14:0] m245_79;
   assign m245_79 =15'b0;

   // m245_80 = W*in
   wire signed [14:0] m245_80;
   assign m245_80 =15'b0;

   // m245_81 = W*in
   wire signed [14:0] m245_81;
   assign m245_81 =15'b0;

   // m245_82 = W*in
   wire signed [14:0] m245_82;
   assign m245_82 =15'b0;

   // m245_83 = W*in
   wire signed [14:0] m245_83;
   assign m245_83 =15'b0;

   // m245_84 = W*in
   wire signed [14:0] m245_84;
   assign m245_84 =15'b0;

   // m245_85 = W*in
   wire signed [14:0] m245_85;
   assign m245_85 =15'b0;

   // m245_86 = W*in
   wire signed [14:0] m245_86;
   assign m245_86 =15'b0;

   // m245_87 = W*in
   wire signed [14:0] m245_87;
   assign m245_87 =15'b0;

   // m245_88 = W*in
   wire signed [14:0] m245_88;
   assign m245_88 =15'b0;

   // m245_89 = W*in
   wire signed [14:0] m245_89;
   assign m245_89 =15'b0;

   // m245_90 = W*in
   wire signed [14:0] m245_90;
   assign m245_90 =15'b0;

   // m245_91 = W*in
   wire signed [14:0] m245_91;
   assign m245_91 =15'b0;

   // m245_92 = W*in
   wire signed [14:0] m245_92;
   assign m245_92 =15'b0;

   // m245_93 = W*in
   wire signed [14:0] m245_93;
   assign m245_93 =15'b0;

   // m245_94 = W*in
   wire signed [14:0] m245_94;
   assign m245_94 =15'b0;

   // m245_95 = W*in
   wire signed [14:0] m245_95;
   assign m245_95 =15'b0;

   // m245_96 = W*in
   wire signed [14:0] m245_96;
   assign m245_96 =15'b0;

   // m245_97 = W*in
   wire signed [14:0] m245_97;
   assign m245_97 =15'b0;

   // m245_98 = W*in
   wire signed [14:0] m245_98;
   assign m245_98 ={ {3{in245[14]}} , in245[14:3] };

   // m245_99 = W*in
   wire signed [14:0] m245_99;
   assign m245_99 ={ {3{neg245[14]}} , neg245[14:3] };

   // m245_100 = W*in
   wire signed [14:0] m245_100;
   assign m245_100 =15'b0;

   // m246_1 = W*in
   wire signed [14:0] m246_1;
   assign m246_1 ={ {3{in246[14]}} , in246[14:3] };

   // m246_2 = W*in
   wire signed [14:0] m246_2;
   assign m246_2 =15'b0;

   // m246_3 = W*in
   wire signed [14:0] m246_3;
   assign m246_3 =15'b0;

   // m246_4 = W*in
   wire signed [14:0] m246_4;
   assign m246_4 ={ {4{neg246[14]}} , neg246[14:4] };

   // m246_5 = W*in
   wire signed [14:0] m246_5;
   assign m246_5 =15'b0;

   // m246_6 = W*in
   wire signed [14:0] m246_6;
   assign m246_6 ={ {3{in246[14]}} , in246[14:3] };

   // m246_7 = W*in
   wire signed [14:0] m246_7;
   assign m246_7 =15'b0;

   // m246_8 = W*in
   wire signed [14:0] m246_8;
   assign m246_8 ={ {3{in246[14]}} , in246[14:3] };

   // m246_9 = W*in
   wire signed [14:0] m246_9;
   assign m246_9 ={ {3{in246[14]}} , in246[14:3] };

   // m246_10 = W*in
   wire signed [14:0] m246_10;
   assign m246_10 =15'b0;

   // m246_11 = W*in
   wire signed [14:0] m246_11;
   assign m246_11 =15'b0;

   // m246_12 = W*in
   wire signed [14:0] m246_12;
   assign m246_12 ={ {3{in246[14]}} , in246[14:3] };

   // m246_13 = W*in
   wire signed [14:0] m246_13;
   assign m246_13 =15'b0;

   // m246_14 = W*in
   wire signed [14:0] m246_14;
   assign m246_14 =15'b0;

   // m246_15 = W*in
   wire signed [14:0] m246_15;
   assign m246_15 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_16 = W*in
   wire signed [14:0] m246_16;
   assign m246_16 =15'b0;

   // m246_17 = W*in
   wire signed [14:0] m246_17;
   assign m246_17 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_18 = W*in
   wire signed [14:0] m246_18;
   assign m246_18 =15'b0;

   // m246_19 = W*in
   wire signed [14:0] m246_19;
   assign m246_19 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_20 = W*in
   wire signed [14:0] m246_20;
   assign m246_20 =15'b0;

   // m246_21 = W*in
   wire signed [14:0] m246_21;
   assign m246_21 ={ {4{neg246[14]}} , neg246[14:4] };

   // m246_22 = W*in
   wire signed [14:0] m246_22;
   assign m246_22 ={ {3{in246[14]}} , in246[14:3] };

   // m246_23 = W*in
   wire signed [14:0] m246_23;
   assign m246_23 ={ {3{in246[14]}} , in246[14:3] };

   // m246_24 = W*in
   wire signed [14:0] m246_24;
   assign m246_24 ={ {3{in246[14]}} , in246[14:3] };

   // m246_25 = W*in
   wire signed [14:0] m246_25;
   assign m246_25 =15'b0;

   // m246_26 = W*in
   wire signed [14:0] m246_26;
   assign m246_26 ={ {2{in246[14]}} , in246[14:2] };

   // m246_27 = W*in
   wire signed [14:0] m246_27;
   assign m246_27 =15'b0;

   // m246_28 = W*in
   wire signed [14:0] m246_28;
   assign m246_28 ={ {4{neg246[14]}} , neg246[14:4] };

   // m246_29 = W*in
   wire signed [14:0] m246_29;
   assign m246_29 ={ {2{in246[14]}} , in246[14:2] };

   // m246_30 = W*in
   wire signed [14:0] m246_30;
   assign m246_30 =15'b0;

   // m246_31 = W*in
   wire signed [14:0] m246_31;
   assign m246_31 ={ {3{in246[14]}} , in246[14:3] };

   // m246_32 = W*in
   wire signed [14:0] m246_32;
   assign m246_32 =15'b0;

   // m246_33 = W*in
   wire signed [14:0] m246_33;
   assign m246_33 =15'b0;

   // m246_34 = W*in
   wire signed [14:0] m246_34;
   assign m246_34 ={ {3{in246[14]}} , in246[14:3] };

   // m246_35 = W*in
   wire signed [14:0] m246_35;
   assign m246_35 =15'b0;

   // m246_36 = W*in
   wire signed [14:0] m246_36;
   assign m246_36 =15'b0;

   // m246_37 = W*in
   wire signed [14:0] m246_37;
   assign m246_37 =15'b0;

   // m246_38 = W*in
   wire signed [14:0] m246_38;
   assign m246_38 =15'b0;

   // m246_39 = W*in
   wire signed [14:0] m246_39;
   assign m246_39 =15'b0;

   // m246_40 = W*in
   wire signed [14:0] m246_40;
   assign m246_40 =15'b0;

   // m246_41 = W*in
   wire signed [14:0] m246_41;
   assign m246_41 =15'b0;

   // m246_42 = W*in
   wire signed [14:0] m246_42;
   assign m246_42 =15'b0;

   // m246_43 = W*in
   wire signed [14:0] m246_43;
   assign m246_43 =15'b0;

   // m246_44 = W*in
   wire signed [14:0] m246_44;
   assign m246_44 =15'b0;

   // m246_45 = W*in
   wire signed [14:0] m246_45;
   assign m246_45 ={ {3{in246[14]}} , in246[14:3] };

   // m246_46 = W*in
   wire signed [14:0] m246_46;
   assign m246_46 ={ {4{neg246[14]}} , neg246[14:4] };

   // m246_47 = W*in
   wire signed [14:0] m246_47;
   assign m246_47 ={ {3{in246[14]}} , in246[14:3] };

   // m246_48 = W*in
   wire signed [14:0] m246_48;
   assign m246_48 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_49 = W*in
   wire signed [14:0] m246_49;
   assign m246_49 =15'b0;

   // m246_50 = W*in
   wire signed [14:0] m246_50;
   assign m246_50 =15'b0;

   // m246_51 = W*in
   wire signed [14:0] m246_51;
   assign m246_51 =15'b0;

   // m246_52 = W*in
   wire signed [14:0] m246_52;
   assign m246_52 =15'b0;

   // m246_53 = W*in
   wire signed [14:0] m246_53;
   assign m246_53 =15'b0;

   // m246_54 = W*in
   wire signed [14:0] m246_54;
   assign m246_54 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_55 = W*in
   wire signed [14:0] m246_55;
   assign m246_55 =15'b0;

   // m246_56 = W*in
   wire signed [14:0] m246_56;
   assign m246_56 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_57 = W*in
   wire signed [14:0] m246_57;
   assign m246_57 =15'b0;

   // m246_58 = W*in
   wire signed [14:0] m246_58;
   assign m246_58 =15'b0;

   // m246_59 = W*in
   wire signed [14:0] m246_59;
   assign m246_59 =15'b0;

   // m246_60 = W*in
   wire signed [14:0] m246_60;
   assign m246_60 =15'b0;

   // m246_61 = W*in
   wire signed [14:0] m246_61;
   assign m246_61 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_62 = W*in
   wire signed [14:0] m246_62;
   assign m246_62 =15'b0;

   // m246_63 = W*in
   wire signed [14:0] m246_63;
   assign m246_63 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_64 = W*in
   wire signed [14:0] m246_64;
   assign m246_64 =15'b0;

   // m246_65 = W*in
   wire signed [14:0] m246_65;
   assign m246_65 =15'b0;

   // m246_66 = W*in
   wire signed [14:0] m246_66;
   assign m246_66 ={ {4{neg246[14]}} , neg246[14:4] };

   // m246_67 = W*in
   wire signed [14:0] m246_67;
   assign m246_67 =15'b0;

   // m246_68 = W*in
   wire signed [14:0] m246_68;
   assign m246_68 =15'b0;

   // m246_69 = W*in
   wire signed [14:0] m246_69;
   assign m246_69 ={ {4{neg246[14]}} , neg246[14:4] };

   // m246_70 = W*in
   wire signed [14:0] m246_70;
   assign m246_70 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_71 = W*in
   wire signed [14:0] m246_71;
   assign m246_71 =15'b0;

   // m246_72 = W*in
   wire signed [14:0] m246_72;
   assign m246_72 =15'b0;

   // m246_73 = W*in
   wire signed [14:0] m246_73;
   assign m246_73 ={ {3{in246[14]}} , in246[14:3] };

   // m246_74 = W*in
   wire signed [14:0] m246_74;
   assign m246_74 ={ {3{in246[14]}} , in246[14:3] };

   // m246_75 = W*in
   wire signed [14:0] m246_75;
   assign m246_75 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_76 = W*in
   wire signed [14:0] m246_76;
   assign m246_76 ={ {4{in246[14]}} , in246[14:4] };

   // m246_77 = W*in
   wire signed [14:0] m246_77;
   assign m246_77 =15'b0;

   // m246_78 = W*in
   wire signed [14:0] m246_78;
   assign m246_78 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_79 = W*in
   wire signed [14:0] m246_79;
   assign m246_79 =15'b0;

   // m246_80 = W*in
   wire signed [14:0] m246_80;
   assign m246_80 =15'b0;

   // m246_81 = W*in
   wire signed [14:0] m246_81;
   assign m246_81 =15'b0;

   // m246_82 = W*in
   wire signed [14:0] m246_82;
   assign m246_82 =15'b0;

   // m246_83 = W*in
   wire signed [14:0] m246_83;
   assign m246_83 =15'b0;

   // m246_84 = W*in
   wire signed [14:0] m246_84;
   assign m246_84 =15'b0;

   // m246_85 = W*in
   wire signed [14:0] m246_85;
   assign m246_85 ={ {3{in246[14]}} , in246[14:3] };

   // m246_86 = W*in
   wire signed [14:0] m246_86;
   assign m246_86 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_87 = W*in
   wire signed [14:0] m246_87;
   assign m246_87 =15'b0;

   // m246_88 = W*in
   wire signed [14:0] m246_88;
   assign m246_88 ={ {3{in246[14]}} , in246[14:3] };

   // m246_89 = W*in
   wire signed [14:0] m246_89;
   assign m246_89 =15'b0;

   // m246_90 = W*in
   wire signed [14:0] m246_90;
   assign m246_90 =15'b0;

   // m246_91 = W*in
   wire signed [14:0] m246_91;
   assign m246_91 =15'b0;

   // m246_92 = W*in
   wire signed [14:0] m246_92;
   assign m246_92 =15'b0;

   // m246_93 = W*in
   wire signed [14:0] m246_93;
   assign m246_93 =15'b0;

   // m246_94 = W*in
   wire signed [14:0] m246_94;
   assign m246_94 =15'b0;

   // m246_95 = W*in
   wire signed [14:0] m246_95;
   assign m246_95 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_96 = W*in
   wire signed [14:0] m246_96;
   assign m246_96 =15'b0;

   // m246_97 = W*in
   wire signed [14:0] m246_97;
   assign m246_97 ={ {3{neg246[14]}} , neg246[14:3] };

   // m246_98 = W*in
   wire signed [14:0] m246_98;
   assign m246_98 =15'b0;

   // m246_99 = W*in
   wire signed [14:0] m246_99;
   assign m246_99 =15'b0;

   // m246_100 = W*in
   wire signed [14:0] m246_100;
   assign m246_100 =15'b0;

   // m247_1 = W*in
   wire signed [14:0] m247_1;
   assign m247_1 ={ {3{neg247[14]}} , neg247[14:3] };

   // m247_2 = W*in
   wire signed [14:0] m247_2;
   assign m247_2 =15'b0;

   // m247_3 = W*in
   wire signed [14:0] m247_3;
   assign m247_3 =15'b0;

   // m247_4 = W*in
   wire signed [14:0] m247_4;
   assign m247_4 =15'b0;

   // m247_5 = W*in
   wire signed [14:0] m247_5;
   assign m247_5 =15'b0;

   // m247_6 = W*in
   wire signed [14:0] m247_6;
   assign m247_6 =15'b0;

   // m247_7 = W*in
   wire signed [14:0] m247_7;
   assign m247_7 =15'b0;

   // m247_8 = W*in
   wire signed [14:0] m247_8;
   assign m247_8 =15'b0;

   // m247_9 = W*in
   wire signed [14:0] m247_9;
   assign m247_9 ={ {3{neg247[14]}} , neg247[14:3] };

   // m247_10 = W*in
   wire signed [14:0] m247_10;
   assign m247_10 =15'b0;

   // m247_11 = W*in
   wire signed [14:0] m247_11;
   assign m247_11 =15'b0;

   // m247_12 = W*in
   wire signed [14:0] m247_12;
   assign m247_12 =15'b0;

   // m247_13 = W*in
   wire signed [14:0] m247_13;
   assign m247_13 =15'b0;

   // m247_14 = W*in
   wire signed [14:0] m247_14;
   assign m247_14 =15'b0;

   // m247_15 = W*in
   wire signed [14:0] m247_15;
   assign m247_15 ={ {3{in247[14]}} , in247[14:3] };

   // m247_16 = W*in
   wire signed [14:0] m247_16;
   assign m247_16 =15'b0;

   // m247_17 = W*in
   wire signed [14:0] m247_17;
   assign m247_17 =15'b0;

   // m247_18 = W*in
   wire signed [14:0] m247_18;
   assign m247_18 =15'b0;

   // m247_19 = W*in
   wire signed [14:0] m247_19;
   assign m247_19 =15'b0;

   // m247_20 = W*in
   wire signed [14:0] m247_20;
   assign m247_20 =15'b0;

   // m247_21 = W*in
   wire signed [14:0] m247_21;
   assign m247_21 =15'b0;

   // m247_22 = W*in
   wire signed [14:0] m247_22;
   assign m247_22 =15'b0;

   // m247_23 = W*in
   wire signed [14:0] m247_23;
   assign m247_23 =15'b0;

   // m247_24 = W*in
   wire signed [14:0] m247_24;
   assign m247_24 =15'b0;

   // m247_25 = W*in
   wire signed [14:0] m247_25;
   assign m247_25 =15'b0;

   // m247_26 = W*in
   wire signed [14:0] m247_26;
   assign m247_26 =15'b0;

   // m247_27 = W*in
   wire signed [14:0] m247_27;
   assign m247_27 =15'b0;

   // m247_28 = W*in
   wire signed [14:0] m247_28;
   assign m247_28 ={ {4{neg247[14]}} , neg247[14:4] };

   // m247_29 = W*in
   wire signed [14:0] m247_29;
   assign m247_29 ={ {4{neg247[14]}} , neg247[14:4] };

   // m247_30 = W*in
   wire signed [14:0] m247_30;
   assign m247_30 =15'b0;

   // m247_31 = W*in
   wire signed [14:0] m247_31;
   assign m247_31 =15'b0;

   // m247_32 = W*in
   wire signed [14:0] m247_32;
   assign m247_32 =15'b0;

   // m247_33 = W*in
   wire signed [14:0] m247_33;
   assign m247_33 =15'b0;

   // m247_34 = W*in
   wire signed [14:0] m247_34;
   assign m247_34 =15'b0;

   // m247_35 = W*in
   wire signed [14:0] m247_35;
   assign m247_35 =15'b0;

   // m247_36 = W*in
   wire signed [14:0] m247_36;
   assign m247_36 =15'b0;

   // m247_37 = W*in
   wire signed [14:0] m247_37;
   assign m247_37 =15'b0;

   // m247_38 = W*in
   wire signed [14:0] m247_38;
   assign m247_38 =15'b0;

   // m247_39 = W*in
   wire signed [14:0] m247_39;
   assign m247_39 ={ {4{neg247[14]}} , neg247[14:4] };

   // m247_40 = W*in
   wire signed [14:0] m247_40;
   assign m247_40 =15'b0;

   // m247_41 = W*in
   wire signed [14:0] m247_41;
   assign m247_41 =15'b0;

   // m247_42 = W*in
   wire signed [14:0] m247_42;
   assign m247_42 =15'b0;

   // m247_43 = W*in
   wire signed [14:0] m247_43;
   assign m247_43 =15'b0;

   // m247_44 = W*in
   wire signed [14:0] m247_44;
   assign m247_44 =15'b0;

   // m247_45 = W*in
   wire signed [14:0] m247_45;
   assign m247_45 =15'b0;

   // m247_46 = W*in
   wire signed [14:0] m247_46;
   assign m247_46 =15'b0;

   // m247_47 = W*in
   wire signed [14:0] m247_47;
   assign m247_47 =15'b0;

   // m247_48 = W*in
   wire signed [14:0] m247_48;
   assign m247_48 ={ {3{in247[14]}} , in247[14:3] };

   // m247_49 = W*in
   wire signed [14:0] m247_49;
   assign m247_49 =15'b0;

   // m247_50 = W*in
   wire signed [14:0] m247_50;
   assign m247_50 =15'b0;

   // m247_51 = W*in
   wire signed [14:0] m247_51;
   assign m247_51 =15'b0;

   // m247_52 = W*in
   wire signed [14:0] m247_52;
   assign m247_52 =15'b0;

   // m247_53 = W*in
   wire signed [14:0] m247_53;
   assign m247_53 =15'b0;

   // m247_54 = W*in
   wire signed [14:0] m247_54;
   assign m247_54 =15'b0;

   // m247_55 = W*in
   wire signed [14:0] m247_55;
   assign m247_55 =15'b0;

   // m247_56 = W*in
   wire signed [14:0] m247_56;
   assign m247_56 =15'b0;

   // m247_57 = W*in
   wire signed [14:0] m247_57;
   assign m247_57 =15'b0;

   // m247_58 = W*in
   wire signed [14:0] m247_58;
   assign m247_58 =15'b0;

   // m247_59 = W*in
   wire signed [14:0] m247_59;
   assign m247_59 =15'b0;

   // m247_60 = W*in
   wire signed [14:0] m247_60;
   assign m247_60 =15'b0;

   // m247_61 = W*in
   wire signed [14:0] m247_61;
   assign m247_61 =15'b0;

   // m247_62 = W*in
   wire signed [14:0] m247_62;
   assign m247_62 =15'b0;

   // m247_63 = W*in
   wire signed [14:0] m247_63;
   assign m247_63 =15'b0;

   // m247_64 = W*in
   wire signed [14:0] m247_64;
   assign m247_64 =15'b0;

   // m247_65 = W*in
   wire signed [14:0] m247_65;
   assign m247_65 =15'b0;

   // m247_66 = W*in
   wire signed [14:0] m247_66;
   assign m247_66 =15'b0;

   // m247_67 = W*in
   wire signed [14:0] m247_67;
   assign m247_67 ={ {3{in247[14]}} , in247[14:3] };

   // m247_68 = W*in
   wire signed [14:0] m247_68;
   assign m247_68 =15'b0;

   // m247_69 = W*in
   wire signed [14:0] m247_69;
   assign m247_69 =15'b0;

   // m247_70 = W*in
   wire signed [14:0] m247_70;
   assign m247_70 =15'b0;

   // m247_71 = W*in
   wire signed [14:0] m247_71;
   assign m247_71 =15'b0;

   // m247_72 = W*in
   wire signed [14:0] m247_72;
   assign m247_72 =15'b0;

   // m247_73 = W*in
   wire signed [14:0] m247_73;
   assign m247_73 =15'b0;

   // m247_74 = W*in
   wire signed [14:0] m247_74;
   assign m247_74 ={ {4{neg247[14]}} , neg247[14:4] };

   // m247_75 = W*in
   wire signed [14:0] m247_75;
   assign m247_75 =15'b0;

   // m247_76 = W*in
   wire signed [14:0] m247_76;
   assign m247_76 ={ {4{neg247[14]}} , neg247[14:4] };

   // m247_77 = W*in
   wire signed [14:0] m247_77;
   assign m247_77 =15'b0;

   // m247_78 = W*in
   wire signed [14:0] m247_78;
   assign m247_78 ={ {3{in247[14]}} , in247[14:3] };

   // m247_79 = W*in
   wire signed [14:0] m247_79;
   assign m247_79 =15'b0;

   // m247_80 = W*in
   wire signed [14:0] m247_80;
   assign m247_80 =15'b0;

   // m247_81 = W*in
   wire signed [14:0] m247_81;
   assign m247_81 =15'b0;

   // m247_82 = W*in
   wire signed [14:0] m247_82;
   assign m247_82 =15'b0;

   // m247_83 = W*in
   wire signed [14:0] m247_83;
   assign m247_83 =15'b0;

   // m247_84 = W*in
   wire signed [14:0] m247_84;
   assign m247_84 ={ {4{neg247[14]}} , neg247[14:4] };

   // m247_85 = W*in
   wire signed [14:0] m247_85;
   assign m247_85 =15'b0;

   // m247_86 = W*in
   wire signed [14:0] m247_86;
   assign m247_86 =15'b0;

   // m247_87 = W*in
   wire signed [14:0] m247_87;
   assign m247_87 =15'b0;

   // m247_88 = W*in
   wire signed [14:0] m247_88;
   assign m247_88 =15'b0;

   // m247_89 = W*in
   wire signed [14:0] m247_89;
   assign m247_89 =15'b0;

   // m247_90 = W*in
   wire signed [14:0] m247_90;
   assign m247_90 =15'b0;

   // m247_91 = W*in
   wire signed [14:0] m247_91;
   assign m247_91 =15'b0;

   // m247_92 = W*in
   wire signed [14:0] m247_92;
   assign m247_92 =15'b0;

   // m247_93 = W*in
   wire signed [14:0] m247_93;
   assign m247_93 =15'b0;

   // m247_94 = W*in
   wire signed [14:0] m247_94;
   assign m247_94 =15'b0;

   // m247_95 = W*in
   wire signed [14:0] m247_95;
   assign m247_95 =15'b0;

   // m247_96 = W*in
   wire signed [14:0] m247_96;
   assign m247_96 =15'b0;

   // m247_97 = W*in
   wire signed [14:0] m247_97;
   assign m247_97 =15'b0;

   // m247_98 = W*in
   wire signed [14:0] m247_98;
   assign m247_98 ={ {3{in247[14]}} , in247[14:3] };

   // m247_99 = W*in
   wire signed [14:0] m247_99;
   assign m247_99 =15'b0;

   // m247_100 = W*in
   wire signed [14:0] m247_100;
   assign m247_100 =15'b0;

   // m248_1 = W*in
   wire signed [14:0] m248_1;
   assign m248_1 =15'b0;

   // m248_2 = W*in
   wire signed [14:0] m248_2;
   assign m248_2 =15'b0;

   // m248_3 = W*in
   wire signed [14:0] m248_3;
   assign m248_3 =15'b0;

   // m248_4 = W*in
   wire signed [14:0] m248_4;
   assign m248_4 ={ {3{neg248[14]}} , neg248[14:3] };

   // m248_5 = W*in
   wire signed [14:0] m248_5;
   assign m248_5 =15'b0;

   // m248_6 = W*in
   wire signed [14:0] m248_6;
   assign m248_6 =15'b0;

   // m248_7 = W*in
   wire signed [14:0] m248_7;
   assign m248_7 =15'b0;

   // m248_8 = W*in
   wire signed [14:0] m248_8;
   assign m248_8 =15'b0;

   // m248_9 = W*in
   wire signed [14:0] m248_9;
   assign m248_9 =15'b0;

   // m248_10 = W*in
   wire signed [14:0] m248_10;
   assign m248_10 =15'b0;

   // m248_11 = W*in
   wire signed [14:0] m248_11;
   assign m248_11 =15'b0;

   // m248_12 = W*in
   wire signed [14:0] m248_12;
   assign m248_12 =15'b0;

   // m248_13 = W*in
   wire signed [14:0] m248_13;
   assign m248_13 =15'b0;

   // m248_14 = W*in
   wire signed [14:0] m248_14;
   assign m248_14 =15'b0;

   // m248_15 = W*in
   wire signed [14:0] m248_15;
   assign m248_15 =15'b0;

   // m248_16 = W*in
   wire signed [14:0] m248_16;
   assign m248_16 =15'b0;

   // m248_17 = W*in
   wire signed [14:0] m248_17;
   assign m248_17 =15'b0;

   // m248_18 = W*in
   wire signed [14:0] m248_18;
   assign m248_18 =15'b0;

   // m248_19 = W*in
   wire signed [14:0] m248_19;
   assign m248_19 ={ {2{in248[14]}} , in248[14:2] };

   // m248_20 = W*in
   wire signed [14:0] m248_20;
   assign m248_20 =15'b0;

   // m248_21 = W*in
   wire signed [14:0] m248_21;
   assign m248_21 =15'b0;

   // m248_22 = W*in
   wire signed [14:0] m248_22;
   assign m248_22 =15'b0;

   // m248_23 = W*in
   wire signed [14:0] m248_23;
   assign m248_23 =15'b0;

   // m248_24 = W*in
   wire signed [14:0] m248_24;
   assign m248_24 =15'b0;

   // m248_25 = W*in
   wire signed [14:0] m248_25;
   assign m248_25 =15'b0;

   // m248_26 = W*in
   wire signed [14:0] m248_26;
   assign m248_26 =15'b0;

   // m248_27 = W*in
   wire signed [14:0] m248_27;
   assign m248_27 =15'b0;

   // m248_28 = W*in
   wire signed [14:0] m248_28;
   assign m248_28 =15'b0;

   // m248_29 = W*in
   wire signed [14:0] m248_29;
   assign m248_29 =15'b0;

   // m248_30 = W*in
   wire signed [14:0] m248_30;
   assign m248_30 =15'b0;

   // m248_31 = W*in
   wire signed [14:0] m248_31;
   assign m248_31 =15'b0;

   // m248_32 = W*in
   wire signed [14:0] m248_32;
   assign m248_32 =15'b0;

   // m248_33 = W*in
   wire signed [14:0] m248_33;
   assign m248_33 ={ {4{in248[14]}} , in248[14:4] };

   // m248_34 = W*in
   wire signed [14:0] m248_34;
   assign m248_34 =15'b0;

   // m248_35 = W*in
   wire signed [14:0] m248_35;
   assign m248_35 ={ {4{in248[14]}} , in248[14:4] };

   // m248_36 = W*in
   wire signed [14:0] m248_36;
   assign m248_36 =15'b0;

   // m248_37 = W*in
   wire signed [14:0] m248_37;
   assign m248_37 =15'b0;

   // m248_38 = W*in
   wire signed [14:0] m248_38;
   assign m248_38 =15'b0;

   // m248_39 = W*in
   wire signed [14:0] m248_39;
   assign m248_39 =15'b0;

   // m248_40 = W*in
   wire signed [14:0] m248_40;
   assign m248_40 =15'b0;

   // m248_41 = W*in
   wire signed [14:0] m248_41;
   assign m248_41 =15'b0;

   // m248_42 = W*in
   wire signed [14:0] m248_42;
   assign m248_42 =15'b0;

   // m248_43 = W*in
   wire signed [14:0] m248_43;
   assign m248_43 =15'b0;

   // m248_44 = W*in
   wire signed [14:0] m248_44;
   assign m248_44 ={ {4{in248[14]}} , in248[14:4] };

   // m248_45 = W*in
   wire signed [14:0] m248_45;
   assign m248_45 =15'b0;

   // m248_46 = W*in
   wire signed [14:0] m248_46;
   assign m248_46 =15'b0;

   // m248_47 = W*in
   wire signed [14:0] m248_47;
   assign m248_47 =15'b0;

   // m248_48 = W*in
   wire signed [14:0] m248_48;
   assign m248_48 =15'b0;

   // m248_49 = W*in
   wire signed [14:0] m248_49;
   assign m248_49 =15'b0;

   // m248_50 = W*in
   wire signed [14:0] m248_50;
   assign m248_50 =15'b0;

   // m248_51 = W*in
   wire signed [14:0] m248_51;
   assign m248_51 =15'b0;

   // m248_52 = W*in
   wire signed [14:0] m248_52;
   assign m248_52 =15'b0;

   // m248_53 = W*in
   wire signed [14:0] m248_53;
   assign m248_53 =15'b0;

   // m248_54 = W*in
   wire signed [14:0] m248_54;
   assign m248_54 ={ {3{in248[14]}} , in248[14:3] };

   // m248_55 = W*in
   wire signed [14:0] m248_55;
   assign m248_55 =15'b0;

   // m248_56 = W*in
   wire signed [14:0] m248_56;
   assign m248_56 =15'b0;

   // m248_57 = W*in
   wire signed [14:0] m248_57;
   assign m248_57 =15'b0;

   // m248_58 = W*in
   wire signed [14:0] m248_58;
   assign m248_58 =15'b0;

   // m248_59 = W*in
   wire signed [14:0] m248_59;
   assign m248_59 =15'b0;

   // m248_60 = W*in
   wire signed [14:0] m248_60;
   assign m248_60 =15'b0;

   // m248_61 = W*in
   wire signed [14:0] m248_61;
   assign m248_61 =15'b0;

   // m248_62 = W*in
   wire signed [14:0] m248_62;
   assign m248_62 ={ {4{in248[14]}} , in248[14:4] };

   // m248_63 = W*in
   wire signed [14:0] m248_63;
   assign m248_63 =15'b0;

   // m248_64 = W*in
   wire signed [14:0] m248_64;
   assign m248_64 =15'b0;

   // m248_65 = W*in
   wire signed [14:0] m248_65;
   assign m248_65 =15'b0;

   // m248_66 = W*in
   wire signed [14:0] m248_66;
   assign m248_66 ={ {3{neg248[14]}} , neg248[14:3] };

   // m248_67 = W*in
   wire signed [14:0] m248_67;
   assign m248_67 =15'b0;

   // m248_68 = W*in
   wire signed [14:0] m248_68;
   assign m248_68 =15'b0;

   // m248_69 = W*in
   wire signed [14:0] m248_69;
   assign m248_69 =15'b0;

   // m248_70 = W*in
   wire signed [14:0] m248_70;
   assign m248_70 ={ {4{in248[14]}} , in248[14:4] };

   // m248_71 = W*in
   wire signed [14:0] m248_71;
   assign m248_71 =15'b0;

   // m248_72 = W*in
   wire signed [14:0] m248_72;
   assign m248_72 =15'b0;

   // m248_73 = W*in
   wire signed [14:0] m248_73;
   assign m248_73 =15'b0;

   // m248_74 = W*in
   wire signed [14:0] m248_74;
   assign m248_74 =15'b0;

   // m248_75 = W*in
   wire signed [14:0] m248_75;
   assign m248_75 =15'b0;

   // m248_76 = W*in
   wire signed [14:0] m248_76;
   assign m248_76 =15'b0;

   // m248_77 = W*in
   wire signed [14:0] m248_77;
   assign m248_77 =15'b0;

   // m248_78 = W*in
   wire signed [14:0] m248_78;
   assign m248_78 =15'b0;

   // m248_79 = W*in
   wire signed [14:0] m248_79;
   assign m248_79 ={ {4{neg248[14]}} , neg248[14:4] };

   // m248_80 = W*in
   wire signed [14:0] m248_80;
   assign m248_80 ={ {3{neg248[14]}} , neg248[14:3] };

   // m248_81 = W*in
   wire signed [14:0] m248_81;
   assign m248_81 =15'b0;

   // m248_82 = W*in
   wire signed [14:0] m248_82;
   assign m248_82 =15'b0;

   // m248_83 = W*in
   wire signed [14:0] m248_83;
   assign m248_83 =15'b0;

   // m248_84 = W*in
   wire signed [14:0] m248_84;
   assign m248_84 =15'b0;

   // m248_85 = W*in
   wire signed [14:0] m248_85;
   assign m248_85 ={ {2{neg248[14]}} , neg248[14:2] };

   // m248_86 = W*in
   wire signed [14:0] m248_86;
   assign m248_86 =15'b0;

   // m248_87 = W*in
   wire signed [14:0] m248_87;
   assign m248_87 ={ {4{in248[14]}} , in248[14:4] };

   // m248_88 = W*in
   wire signed [14:0] m248_88;
   assign m248_88 =15'b0;

   // m248_89 = W*in
   wire signed [14:0] m248_89;
   assign m248_89 =15'b0;

   // m248_90 = W*in
   wire signed [14:0] m248_90;
   assign m248_90 ={ {4{in248[14]}} , in248[14:4] };

   // m248_91 = W*in
   wire signed [14:0] m248_91;
   assign m248_91 =15'b0;

   // m248_92 = W*in
   wire signed [14:0] m248_92;
   assign m248_92 ={ {4{neg248[14]}} , neg248[14:4] };

   // m248_93 = W*in
   wire signed [14:0] m248_93;
   assign m248_93 =15'b0;

   // m248_94 = W*in
   wire signed [14:0] m248_94;
   assign m248_94 =15'b0;

   // m248_95 = W*in
   wire signed [14:0] m248_95;
   assign m248_95 =15'b0;

   // m248_96 = W*in
   wire signed [14:0] m248_96;
   assign m248_96 =15'b0;

   // m248_97 = W*in
   wire signed [14:0] m248_97;
   assign m248_97 =15'b0;

   // m248_98 = W*in
   wire signed [14:0] m248_98;
   assign m248_98 =15'b0;

   // m248_99 = W*in
   wire signed [14:0] m248_99;
   assign m248_99 =15'b0;

   // m248_100 = W*in
   wire signed [14:0] m248_100;
   assign m248_100 ={ {4{neg248[14]}} , neg248[14:4] };

   // m249_1 = W*in
   wire signed [14:0] m249_1;
   assign m249_1 =15'b0;

   // m249_2 = W*in
   wire signed [14:0] m249_2;
   assign m249_2 =15'b0;

   // m249_3 = W*in
   wire signed [14:0] m249_3;
   assign m249_3 =15'b0;

   // m249_4 = W*in
   wire signed [14:0] m249_4;
   assign m249_4 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_5 = W*in
   wire signed [14:0] m249_5;
   assign m249_5 =15'b0;

   // m249_6 = W*in
   wire signed [14:0] m249_6;
   assign m249_6 =15'b0;

   // m249_7 = W*in
   wire signed [14:0] m249_7;
   assign m249_7 =15'b0;

   // m249_8 = W*in
   wire signed [14:0] m249_8;
   assign m249_8 =15'b0;

   // m249_9 = W*in
   wire signed [14:0] m249_9;
   assign m249_9 =15'b0;

   // m249_10 = W*in
   wire signed [14:0] m249_10;
   assign m249_10 =15'b0;

   // m249_11 = W*in
   wire signed [14:0] m249_11;
   assign m249_11 =15'b0;

   // m249_12 = W*in
   wire signed [14:0] m249_12;
   assign m249_12 =15'b0;

   // m249_13 = W*in
   wire signed [14:0] m249_13;
   assign m249_13 =15'b0;

   // m249_14 = W*in
   wire signed [14:0] m249_14;
   assign m249_14 =15'b0;

   // m249_15 = W*in
   wire signed [14:0] m249_15;
   assign m249_15 =15'b0;

   // m249_16 = W*in
   wire signed [14:0] m249_16;
   assign m249_16 ={ {3{in249[14]}} , in249[14:3] };

   // m249_17 = W*in
   wire signed [14:0] m249_17;
   assign m249_17 =15'b0;

   // m249_18 = W*in
   wire signed [14:0] m249_18;
   assign m249_18 ={ {3{neg249[14]}} , neg249[14:3] };

   // m249_19 = W*in
   wire signed [14:0] m249_19;
   assign m249_19 ={ {4{in249[14]}} , in249[14:4] };

   // m249_20 = W*in
   wire signed [14:0] m249_20;
   assign m249_20 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_21 = W*in
   wire signed [14:0] m249_21;
   assign m249_21 =15'b0;

   // m249_22 = W*in
   wire signed [14:0] m249_22;
   assign m249_22 =15'b0;

   // m249_23 = W*in
   wire signed [14:0] m249_23;
   assign m249_23 =15'b0;

   // m249_24 = W*in
   wire signed [14:0] m249_24;
   assign m249_24 =15'b0;

   // m249_25 = W*in
   wire signed [14:0] m249_25;
   assign m249_25 ={ {3{in249[14]}} , in249[14:3] };

   // m249_26 = W*in
   wire signed [14:0] m249_26;
   assign m249_26 ={ {3{in249[14]}} , in249[14:3] };

   // m249_27 = W*in
   wire signed [14:0] m249_27;
   assign m249_27 =15'b0;

   // m249_28 = W*in
   wire signed [14:0] m249_28;
   assign m249_28 ={ {3{neg249[14]}} , neg249[14:3] };

   // m249_29 = W*in
   wire signed [14:0] m249_29;
   assign m249_29 =15'b0;

   // m249_30 = W*in
   wire signed [14:0] m249_30;
   assign m249_30 =15'b0;

   // m249_31 = W*in
   wire signed [14:0] m249_31;
   assign m249_31 =15'b0;

   // m249_32 = W*in
   wire signed [14:0] m249_32;
   assign m249_32 ={ {3{in249[14]}} , in249[14:3] };

   // m249_33 = W*in
   wire signed [14:0] m249_33;
   assign m249_33 ={ {3{neg249[14]}} , neg249[14:3] };

   // m249_34 = W*in
   wire signed [14:0] m249_34;
   assign m249_34 =15'b0;

   // m249_35 = W*in
   wire signed [14:0] m249_35;
   assign m249_35 =15'b0;

   // m249_36 = W*in
   wire signed [14:0] m249_36;
   assign m249_36 =15'b0;

   // m249_37 = W*in
   wire signed [14:0] m249_37;
   assign m249_37 =15'b0;

   // m249_38 = W*in
   wire signed [14:0] m249_38;
   assign m249_38 =15'b0;

   // m249_39 = W*in
   wire signed [14:0] m249_39;
   assign m249_39 =15'b0;

   // m249_40 = W*in
   wire signed [14:0] m249_40;
   assign m249_40 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_41 = W*in
   wire signed [14:0] m249_41;
   assign m249_41 =15'b0;

   // m249_42 = W*in
   wire signed [14:0] m249_42;
   assign m249_42 =15'b0;

   // m249_43 = W*in
   wire signed [14:0] m249_43;
   assign m249_43 ={ {3{in249[14]}} , in249[14:3] };

   // m249_44 = W*in
   wire signed [14:0] m249_44;
   assign m249_44 =15'b0;

   // m249_45 = W*in
   wire signed [14:0] m249_45;
   assign m249_45 =15'b0;

   // m249_46 = W*in
   wire signed [14:0] m249_46;
   assign m249_46 ={ {4{in249[14]}} , in249[14:4] };

   // m249_47 = W*in
   wire signed [14:0] m249_47;
   assign m249_47 =15'b0;

   // m249_48 = W*in
   wire signed [14:0] m249_48;
   assign m249_48 =15'b0;

   // m249_49 = W*in
   wire signed [14:0] m249_49;
   assign m249_49 =15'b0;

   // m249_50 = W*in
   wire signed [14:0] m249_50;
   assign m249_50 ={ {3{in249[14]}} , in249[14:3] };

   // m249_51 = W*in
   wire signed [14:0] m249_51;
   assign m249_51 =15'b0;

   // m249_52 = W*in
   wire signed [14:0] m249_52;
   assign m249_52 =15'b0;

   // m249_53 = W*in
   wire signed [14:0] m249_53;
   assign m249_53 =15'b0;

   // m249_54 = W*in
   wire signed [14:0] m249_54;
   assign m249_54 =15'b0;

   // m249_55 = W*in
   wire signed [14:0] m249_55;
   assign m249_55 ={ {3{neg249[14]}} , neg249[14:3] };

   // m249_56 = W*in
   wire signed [14:0] m249_56;
   assign m249_56 ={ {3{neg249[14]}} , neg249[14:3] };

   // m249_57 = W*in
   wire signed [14:0] m249_57;
   assign m249_57 =15'b0;

   // m249_58 = W*in
   wire signed [14:0] m249_58;
   assign m249_58 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_59 = W*in
   wire signed [14:0] m249_59;
   assign m249_59 =15'b0;

   // m249_60 = W*in
   wire signed [14:0] m249_60;
   assign m249_60 =15'b0;

   // m249_61 = W*in
   wire signed [14:0] m249_61;
   assign m249_61 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_62 = W*in
   wire signed [14:0] m249_62;
   assign m249_62 =15'b0;

   // m249_63 = W*in
   wire signed [14:0] m249_63;
   assign m249_63 =15'b0;

   // m249_64 = W*in
   wire signed [14:0] m249_64;
   assign m249_64 =15'b0;

   // m249_65 = W*in
   wire signed [14:0] m249_65;
   assign m249_65 ={ {3{in249[14]}} , in249[14:3] };

   // m249_66 = W*in
   wire signed [14:0] m249_66;
   assign m249_66 =15'b0;

   // m249_67 = W*in
   wire signed [14:0] m249_67;
   assign m249_67 =15'b0;

   // m249_68 = W*in
   wire signed [14:0] m249_68;
   assign m249_68 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_69 = W*in
   wire signed [14:0] m249_69;
   assign m249_69 ={ {3{in249[14]}} , in249[14:3] };

   // m249_70 = W*in
   wire signed [14:0] m249_70;
   assign m249_70 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_71 = W*in
   wire signed [14:0] m249_71;
   assign m249_71 =15'b0;

   // m249_72 = W*in
   wire signed [14:0] m249_72;
   assign m249_72 =15'b0;

   // m249_73 = W*in
   wire signed [14:0] m249_73;
   assign m249_73 =15'b0;

   // m249_74 = W*in
   wire signed [14:0] m249_74;
   assign m249_74 ={ {3{neg249[14]}} , neg249[14:3] };

   // m249_75 = W*in
   wire signed [14:0] m249_75;
   assign m249_75 =15'b0;

   // m249_76 = W*in
   wire signed [14:0] m249_76;
   assign m249_76 ={ {4{in249[14]}} , in249[14:4] };

   // m249_77 = W*in
   wire signed [14:0] m249_77;
   assign m249_77 =15'b0;

   // m249_78 = W*in
   wire signed [14:0] m249_78;
   assign m249_78 ={ {4{neg249[14]}} , neg249[14:4] };

   // m249_79 = W*in
   wire signed [14:0] m249_79;
   assign m249_79 =15'b0;

   // m249_80 = W*in
   wire signed [14:0] m249_80;
   assign m249_80 =15'b0;

   // m249_81 = W*in
   wire signed [14:0] m249_81;
   assign m249_81 =15'b0;

   // m249_82 = W*in
   wire signed [14:0] m249_82;
   assign m249_82 =15'b0;

   // m249_83 = W*in
   wire signed [14:0] m249_83;
   assign m249_83 =15'b0;

   // m249_84 = W*in
   wire signed [14:0] m249_84;
   assign m249_84 =15'b0;

   // m249_85 = W*in
   wire signed [14:0] m249_85;
   assign m249_85 =15'b0;

   // m249_86 = W*in
   wire signed [14:0] m249_86;
   assign m249_86 =15'b0;

   // m249_87 = W*in
   wire signed [14:0] m249_87;
   assign m249_87 =15'b0;

   // m249_88 = W*in
   wire signed [14:0] m249_88;
   assign m249_88 =15'b0;

   // m249_89 = W*in
   wire signed [14:0] m249_89;
   assign m249_89 =15'b0;

   // m249_90 = W*in
   wire signed [14:0] m249_90;
   assign m249_90 =15'b0;

   // m249_91 = W*in
   wire signed [14:0] m249_91;
   assign m249_91 =15'b0;

   // m249_92 = W*in
   wire signed [14:0] m249_92;
   assign m249_92 ={ {3{in249[14]}} , in249[14:3] };

   // m249_93 = W*in
   wire signed [14:0] m249_93;
   assign m249_93 =15'b0;

   // m249_94 = W*in
   wire signed [14:0] m249_94;
   assign m249_94 =15'b0;

   // m249_95 = W*in
   wire signed [14:0] m249_95;
   assign m249_95 =15'b0;

   // m249_96 = W*in
   wire signed [14:0] m249_96;
   assign m249_96 =15'b0;

   // m249_97 = W*in
   wire signed [14:0] m249_97;
   assign m249_97 =15'b0;

   // m249_98 = W*in
   wire signed [14:0] m249_98;
   assign m249_98 =15'b0;

   // m249_99 = W*in
   wire signed [14:0] m249_99;
   assign m249_99 =15'b0;

   // m249_100 = W*in
   wire signed [14:0] m249_100;
   assign m249_100 =15'b0;

   // m250_1 = W*in
   wire signed [14:0] m250_1;
   assign m250_1 =15'b0;

   // m250_2 = W*in
   wire signed [14:0] m250_2;
   assign m250_2 =15'b0;

   // m250_3 = W*in
   wire signed [14:0] m250_3;
   assign m250_3 =15'b0;

   // m250_4 = W*in
   wire signed [14:0] m250_4;
   assign m250_4 =15'b0;

   // m250_5 = W*in
   wire signed [14:0] m250_5;
   assign m250_5 ={ {4{in250[14]}} , in250[14:4] };

   // m250_6 = W*in
   wire signed [14:0] m250_6;
   assign m250_6 =15'b0;

   // m250_7 = W*in
   wire signed [14:0] m250_7;
   assign m250_7 =15'b0;

   // m250_8 = W*in
   wire signed [14:0] m250_8;
   assign m250_8 =15'b0;

   // m250_9 = W*in
   wire signed [14:0] m250_9;
   assign m250_9 =15'b0;

   // m250_10 = W*in
   wire signed [14:0] m250_10;
   assign m250_10 =15'b0;

   // m250_11 = W*in
   wire signed [14:0] m250_11;
   assign m250_11 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_12 = W*in
   wire signed [14:0] m250_12;
   assign m250_12 =15'b0;

   // m250_13 = W*in
   wire signed [14:0] m250_13;
   assign m250_13 =15'b0;

   // m250_14 = W*in
   wire signed [14:0] m250_14;
   assign m250_14 =15'b0;

   // m250_15 = W*in
   wire signed [14:0] m250_15;
   assign m250_15 =15'b0;

   // m250_16 = W*in
   wire signed [14:0] m250_16;
   assign m250_16 =15'b0;

   // m250_17 = W*in
   wire signed [14:0] m250_17;
   assign m250_17 =15'b0;

   // m250_18 = W*in
   wire signed [14:0] m250_18;
   assign m250_18 ={ {4{in250[14]}} , in250[14:4] };

   // m250_19 = W*in
   wire signed [14:0] m250_19;
   assign m250_19 =15'b0;

   // m250_20 = W*in
   wire signed [14:0] m250_20;
   assign m250_20 =15'b0;

   // m250_21 = W*in
   wire signed [14:0] m250_21;
   assign m250_21 ={ {4{neg250[14]}} , neg250[14:4] };

   // m250_22 = W*in
   wire signed [14:0] m250_22;
   assign m250_22 ={ {3{in250[14]}} , in250[14:3] };

   // m250_23 = W*in
   wire signed [14:0] m250_23;
   assign m250_23 =15'b0;

   // m250_24 = W*in
   wire signed [14:0] m250_24;
   assign m250_24 =15'b0;

   // m250_25 = W*in
   wire signed [14:0] m250_25;
   assign m250_25 =15'b0;

   // m250_26 = W*in
   wire signed [14:0] m250_26;
   assign m250_26 =15'b0;

   // m250_27 = W*in
   wire signed [14:0] m250_27;
   assign m250_27 ={ {4{neg250[14]}} , neg250[14:4] };

   // m250_28 = W*in
   wire signed [14:0] m250_28;
   assign m250_28 =15'b0;

   // m250_29 = W*in
   wire signed [14:0] m250_29;
   assign m250_29 =15'b0;

   // m250_30 = W*in
   wire signed [14:0] m250_30;
   assign m250_30 =15'b0;

   // m250_31 = W*in
   wire signed [14:0] m250_31;
   assign m250_31 =15'b0;

   // m250_32 = W*in
   wire signed [14:0] m250_32;
   assign m250_32 =15'b0;

   // m250_33 = W*in
   wire signed [14:0] m250_33;
   assign m250_33 =15'b0;

   // m250_34 = W*in
   wire signed [14:0] m250_34;
   assign m250_34 =15'b0;

   // m250_35 = W*in
   wire signed [14:0] m250_35;
   assign m250_35 =15'b0;

   // m250_36 = W*in
   wire signed [14:0] m250_36;
   assign m250_36 =15'b0;

   // m250_37 = W*in
   wire signed [14:0] m250_37;
   assign m250_37 =15'b0;

   // m250_38 = W*in
   wire signed [14:0] m250_38;
   assign m250_38 =15'b0;

   // m250_39 = W*in
   wire signed [14:0] m250_39;
   assign m250_39 =15'b0;

   // m250_40 = W*in
   wire signed [14:0] m250_40;
   assign m250_40 =15'b0;

   // m250_41 = W*in
   wire signed [14:0] m250_41;
   assign m250_41 ={ {4{neg250[14]}} , neg250[14:4] };

   // m250_42 = W*in
   wire signed [14:0] m250_42;
   assign m250_42 =15'b0;

   // m250_43 = W*in
   wire signed [14:0] m250_43;
   assign m250_43 =15'b0;

   // m250_44 = W*in
   wire signed [14:0] m250_44;
   assign m250_44 =15'b0;

   // m250_45 = W*in
   wire signed [14:0] m250_45;
   assign m250_45 =15'b0;

   // m250_46 = W*in
   wire signed [14:0] m250_46;
   assign m250_46 =15'b0;

   // m250_47 = W*in
   wire signed [14:0] m250_47;
   assign m250_47 =15'b0;

   // m250_48 = W*in
   wire signed [14:0] m250_48;
   assign m250_48 =15'b0;

   // m250_49 = W*in
   wire signed [14:0] m250_49;
   assign m250_49 =15'b0;

   // m250_50 = W*in
   wire signed [14:0] m250_50;
   assign m250_50 =15'b0;

   // m250_51 = W*in
   wire signed [14:0] m250_51;
   assign m250_51 =15'b0;

   // m250_52 = W*in
   wire signed [14:0] m250_52;
   assign m250_52 =15'b0;

   // m250_53 = W*in
   wire signed [14:0] m250_53;
   assign m250_53 =15'b0;

   // m250_54 = W*in
   wire signed [14:0] m250_54;
   assign m250_54 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_55 = W*in
   wire signed [14:0] m250_55;
   assign m250_55 =15'b0;

   // m250_56 = W*in
   wire signed [14:0] m250_56;
   assign m250_56 =15'b0;

   // m250_57 = W*in
   wire signed [14:0] m250_57;
   assign m250_57 ={ {3{in250[14]}} , in250[14:3] };

   // m250_58 = W*in
   wire signed [14:0] m250_58;
   assign m250_58 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_59 = W*in
   wire signed [14:0] m250_59;
   assign m250_59 =15'b0;

   // m250_60 = W*in
   wire signed [14:0] m250_60;
   assign m250_60 =15'b0;

   // m250_61 = W*in
   wire signed [14:0] m250_61;
   assign m250_61 =15'b0;

   // m250_62 = W*in
   wire signed [14:0] m250_62;
   assign m250_62 =15'b0;

   // m250_63 = W*in
   wire signed [14:0] m250_63;
   assign m250_63 =15'b0;

   // m250_64 = W*in
   wire signed [14:0] m250_64;
   assign m250_64 ={ {3{in250[14]}} , in250[14:3] };

   // m250_65 = W*in
   wire signed [14:0] m250_65;
   assign m250_65 =15'b0;

   // m250_66 = W*in
   wire signed [14:0] m250_66;
   assign m250_66 =15'b0;

   // m250_67 = W*in
   wire signed [14:0] m250_67;
   assign m250_67 =15'b0;

   // m250_68 = W*in
   wire signed [14:0] m250_68;
   assign m250_68 =15'b0;

   // m250_69 = W*in
   wire signed [14:0] m250_69;
   assign m250_69 =15'b0;

   // m250_70 = W*in
   wire signed [14:0] m250_70;
   assign m250_70 =15'b0;

   // m250_71 = W*in
   wire signed [14:0] m250_71;
   assign m250_71 =15'b0;

   // m250_72 = W*in
   wire signed [14:0] m250_72;
   assign m250_72 =15'b0;

   // m250_73 = W*in
   wire signed [14:0] m250_73;
   assign m250_73 =15'b0;

   // m250_74 = W*in
   wire signed [14:0] m250_74;
   assign m250_74 =15'b0;

   // m250_75 = W*in
   wire signed [14:0] m250_75;
   assign m250_75 =15'b0;

   // m250_76 = W*in
   wire signed [14:0] m250_76;
   assign m250_76 =15'b0;

   // m250_77 = W*in
   wire signed [14:0] m250_77;
   assign m250_77 =15'b0;

   // m250_78 = W*in
   wire signed [14:0] m250_78;
   assign m250_78 =15'b0;

   // m250_79 = W*in
   wire signed [14:0] m250_79;
   assign m250_79 =15'b0;

   // m250_80 = W*in
   wire signed [14:0] m250_80;
   assign m250_80 =15'b0;

   // m250_81 = W*in
   wire signed [14:0] m250_81;
   assign m250_81 =15'b0;

   // m250_82 = W*in
   wire signed [14:0] m250_82;
   assign m250_82 =15'b0;

   // m250_83 = W*in
   wire signed [14:0] m250_83;
   assign m250_83 =15'b0;

   // m250_84 = W*in
   wire signed [14:0] m250_84;
   assign m250_84 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_85 = W*in
   wire signed [14:0] m250_85;
   assign m250_85 ={ {3{in250[14]}} , in250[14:3] };

   // m250_86 = W*in
   wire signed [14:0] m250_86;
   assign m250_86 =15'b0;

   // m250_87 = W*in
   wire signed [14:0] m250_87;
   assign m250_87 ={ {2{in250[14]}} , in250[14:2] };

   // m250_88 = W*in
   wire signed [14:0] m250_88;
   assign m250_88 =15'b0;

   // m250_89 = W*in
   wire signed [14:0] m250_89;
   assign m250_89 =15'b0;

   // m250_90 = W*in
   wire signed [14:0] m250_90;
   assign m250_90 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_91 = W*in
   wire signed [14:0] m250_91;
   assign m250_91 ={ {4{in250[14]}} , in250[14:4] };

   // m250_92 = W*in
   wire signed [14:0] m250_92;
   assign m250_92 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_93 = W*in
   wire signed [14:0] m250_93;
   assign m250_93 ={ {3{neg250[14]}} , neg250[14:3] };

   // m250_94 = W*in
   wire signed [14:0] m250_94;
   assign m250_94 =15'b0;

   // m250_95 = W*in
   wire signed [14:0] m250_95;
   assign m250_95 =15'b0;

   // m250_96 = W*in
   wire signed [14:0] m250_96;
   assign m250_96 =15'b0;

   // m250_97 = W*in
   wire signed [14:0] m250_97;
   assign m250_97 ={ {4{neg250[14]}} , neg250[14:4] };

   // m250_98 = W*in
   wire signed [14:0] m250_98;
   assign m250_98 =15'b0;

   // m250_99 = W*in
   wire signed [14:0] m250_99;
   assign m250_99 =15'b0;

   // m250_100 = W*in
   wire signed [14:0] m250_100;
   assign m250_100 =15'b0;

   // m251_1 = W*in
   wire signed [14:0] m251_1;
   assign m251_1 =15'b0;

   // m251_2 = W*in
   wire signed [14:0] m251_2;
   assign m251_2 =15'b0;

   // m251_3 = W*in
   wire signed [14:0] m251_3;
   assign m251_3 =15'b0;

   // m251_4 = W*in
   wire signed [14:0] m251_4;
   assign m251_4 =15'b0;

   // m251_5 = W*in
   wire signed [14:0] m251_5;
   assign m251_5 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_6 = W*in
   wire signed [14:0] m251_6;
   assign m251_6 =15'b0;

   // m251_7 = W*in
   wire signed [14:0] m251_7;
   assign m251_7 =15'b0;

   // m251_8 = W*in
   wire signed [14:0] m251_8;
   assign m251_8 =15'b0;

   // m251_9 = W*in
   wire signed [14:0] m251_9;
   assign m251_9 =15'b0;

   // m251_10 = W*in
   wire signed [14:0] m251_10;
   assign m251_10 =15'b0;

   // m251_11 = W*in
   wire signed [14:0] m251_11;
   assign m251_11 ={ {2{in251[14]}} , in251[14:2] };

   // m251_12 = W*in
   wire signed [14:0] m251_12;
   assign m251_12 =15'b0;

   // m251_13 = W*in
   wire signed [14:0] m251_13;
   assign m251_13 =15'b0;

   // m251_14 = W*in
   wire signed [14:0] m251_14;
   assign m251_14 =15'b0;

   // m251_15 = W*in
   wire signed [14:0] m251_15;
   assign m251_15 =15'b0;

   // m251_16 = W*in
   wire signed [14:0] m251_16;
   assign m251_16 ={ {2{neg251[14]}} , neg251[14:2] };

   // m251_17 = W*in
   wire signed [14:0] m251_17;
   assign m251_17 =15'b0;

   // m251_18 = W*in
   wire signed [14:0] m251_18;
   assign m251_18 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_19 = W*in
   wire signed [14:0] m251_19;
   assign m251_19 ={ {3{in251[14]}} , in251[14:3] };

   // m251_20 = W*in
   wire signed [14:0] m251_20;
   assign m251_20 ={ {4{neg251[14]}} , neg251[14:4] };

   // m251_21 = W*in
   wire signed [14:0] m251_21;
   assign m251_21 =15'b0;

   // m251_22 = W*in
   wire signed [14:0] m251_22;
   assign m251_22 =15'b0;

   // m251_23 = W*in
   wire signed [14:0] m251_23;
   assign m251_23 =15'b0;

   // m251_24 = W*in
   wire signed [14:0] m251_24;
   assign m251_24 =15'b0;

   // m251_25 = W*in
   wire signed [14:0] m251_25;
   assign m251_25 =15'b0;

   // m251_26 = W*in
   wire signed [14:0] m251_26;
   assign m251_26 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_27 = W*in
   wire signed [14:0] m251_27;
   assign m251_27 =15'b0;

   // m251_28 = W*in
   wire signed [14:0] m251_28;
   assign m251_28 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_29 = W*in
   wire signed [14:0] m251_29;
   assign m251_29 =15'b0;

   // m251_30 = W*in
   wire signed [14:0] m251_30;
   assign m251_30 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_31 = W*in
   wire signed [14:0] m251_31;
   assign m251_31 =15'b0;

   // m251_32 = W*in
   wire signed [14:0] m251_32;
   assign m251_32 ={ {3{in251[14]}} , in251[14:3] };

   // m251_33 = W*in
   wire signed [14:0] m251_33;
   assign m251_33 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_34 = W*in
   wire signed [14:0] m251_34;
   assign m251_34 =15'b0;

   // m251_35 = W*in
   wire signed [14:0] m251_35;
   assign m251_35 =15'b0;

   // m251_36 = W*in
   wire signed [14:0] m251_36;
   assign m251_36 =15'b0;

   // m251_37 = W*in
   wire signed [14:0] m251_37;
   assign m251_37 ={ {3{in251[14]}} , in251[14:3] };

   // m251_38 = W*in
   wire signed [14:0] m251_38;
   assign m251_38 =15'b0;

   // m251_39 = W*in
   wire signed [14:0] m251_39;
   assign m251_39 =15'b0;

   // m251_40 = W*in
   wire signed [14:0] m251_40;
   assign m251_40 =15'b0;

   // m251_41 = W*in
   wire signed [14:0] m251_41;
   assign m251_41 =15'b0;

   // m251_42 = W*in
   wire signed [14:0] m251_42;
   assign m251_42 =15'b0;

   // m251_43 = W*in
   wire signed [14:0] m251_43;
   assign m251_43 =15'b0;

   // m251_44 = W*in
   wire signed [14:0] m251_44;
   assign m251_44 ={ {3{in251[14]}} , in251[14:3] };

   // m251_45 = W*in
   wire signed [14:0] m251_45;
   assign m251_45 =15'b0;

   // m251_46 = W*in
   wire signed [14:0] m251_46;
   assign m251_46 =15'b0;

   // m251_47 = W*in
   wire signed [14:0] m251_47;
   assign m251_47 =15'b0;

   // m251_48 = W*in
   wire signed [14:0] m251_48;
   assign m251_48 =15'b0;

   // m251_49 = W*in
   wire signed [14:0] m251_49;
   assign m251_49 =15'b0;

   // m251_50 = W*in
   wire signed [14:0] m251_50;
   assign m251_50 =15'b0;

   // m251_51 = W*in
   wire signed [14:0] m251_51;
   assign m251_51 =15'b0;

   // m251_52 = W*in
   wire signed [14:0] m251_52;
   assign m251_52 =15'b0;

   // m251_53 = W*in
   wire signed [14:0] m251_53;
   assign m251_53 =15'b0;

   // m251_54 = W*in
   wire signed [14:0] m251_54;
   assign m251_54 =15'b0;

   // m251_55 = W*in
   wire signed [14:0] m251_55;
   assign m251_55 =15'b0;

   // m251_56 = W*in
   wire signed [14:0] m251_56;
   assign m251_56 =15'b0;

   // m251_57 = W*in
   wire signed [14:0] m251_57;
   assign m251_57 =15'b0;

   // m251_58 = W*in
   wire signed [14:0] m251_58;
   assign m251_58 ={ {4{neg251[14]}} , neg251[14:4] };

   // m251_59 = W*in
   wire signed [14:0] m251_59;
   assign m251_59 =15'b0;

   // m251_60 = W*in
   wire signed [14:0] m251_60;
   assign m251_60 =15'b0;

   // m251_61 = W*in
   wire signed [14:0] m251_61;
   assign m251_61 =15'b0;

   // m251_62 = W*in
   wire signed [14:0] m251_62;
   assign m251_62 =15'b0;

   // m251_63 = W*in
   wire signed [14:0] m251_63;
   assign m251_63 =15'b0;

   // m251_64 = W*in
   wire signed [14:0] m251_64;
   assign m251_64 =15'b0;

   // m251_65 = W*in
   wire signed [14:0] m251_65;
   assign m251_65 =15'b0;

   // m251_66 = W*in
   wire signed [14:0] m251_66;
   assign m251_66 ={ {4{in251[14]}} , in251[14:4] };

   // m251_67 = W*in
   wire signed [14:0] m251_67;
   assign m251_67 =15'b0;

   // m251_68 = W*in
   wire signed [14:0] m251_68;
   assign m251_68 =15'b0;

   // m251_69 = W*in
   wire signed [14:0] m251_69;
   assign m251_69 =15'b0;

   // m251_70 = W*in
   wire signed [14:0] m251_70;
   assign m251_70 =15'b0;

   // m251_71 = W*in
   wire signed [14:0] m251_71;
   assign m251_71 =15'b0;

   // m251_72 = W*in
   wire signed [14:0] m251_72;
   assign m251_72 =15'b0;

   // m251_73 = W*in
   wire signed [14:0] m251_73;
   assign m251_73 =15'b0;

   // m251_74 = W*in
   wire signed [14:0] m251_74;
   assign m251_74 =15'b0;

   // m251_75 = W*in
   wire signed [14:0] m251_75;
   assign m251_75 =15'b0;

   // m251_76 = W*in
   wire signed [14:0] m251_76;
   assign m251_76 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_77 = W*in
   wire signed [14:0] m251_77;
   assign m251_77 =15'b0;

   // m251_78 = W*in
   wire signed [14:0] m251_78;
   assign m251_78 =15'b0;

   // m251_79 = W*in
   wire signed [14:0] m251_79;
   assign m251_79 =15'b0;

   // m251_80 = W*in
   wire signed [14:0] m251_80;
   assign m251_80 =15'b0;

   // m251_81 = W*in
   wire signed [14:0] m251_81;
   assign m251_81 =15'b0;

   // m251_82 = W*in
   wire signed [14:0] m251_82;
   assign m251_82 =15'b0;

   // m251_83 = W*in
   wire signed [14:0] m251_83;
   assign m251_83 =15'b0;

   // m251_84 = W*in
   wire signed [14:0] m251_84;
   assign m251_84 =15'b0;

   // m251_85 = W*in
   wire signed [14:0] m251_85;
   assign m251_85 =15'b0;

   // m251_86 = W*in
   wire signed [14:0] m251_86;
   assign m251_86 =15'b0;

   // m251_87 = W*in
   wire signed [14:0] m251_87;
   assign m251_87 =15'b0;

   // m251_88 = W*in
   wire signed [14:0] m251_88;
   assign m251_88 =15'b0;

   // m251_89 = W*in
   wire signed [14:0] m251_89;
   assign m251_89 =15'b0;

   // m251_90 = W*in
   wire signed [14:0] m251_90;
   assign m251_90 =15'b0;

   // m251_91 = W*in
   wire signed [14:0] m251_91;
   assign m251_91 =15'b0;

   // m251_92 = W*in
   wire signed [14:0] m251_92;
   assign m251_92 =15'b0;

   // m251_93 = W*in
   wire signed [14:0] m251_93;
   assign m251_93 ={ {3{neg251[14]}} , neg251[14:3] };

   // m251_94 = W*in
   wire signed [14:0] m251_94;
   assign m251_94 =15'b0;

   // m251_95 = W*in
   wire signed [14:0] m251_95;
   assign m251_95 ={ {4{in251[14]}} , in251[14:4] };

   // m251_96 = W*in
   wire signed [14:0] m251_96;
   assign m251_96 =15'b0;

   // m251_97 = W*in
   wire signed [14:0] m251_97;
   assign m251_97 =15'b0;

   // m251_98 = W*in
   wire signed [14:0] m251_98;
   assign m251_98 =15'b0;

   // m251_99 = W*in
   wire signed [14:0] m251_99;
   assign m251_99 =15'b0;

   // m251_100 = W*in
   wire signed [14:0] m251_100;
   assign m251_100 =15'b0;

   // m252_1 = W*in
   wire signed [14:0] m252_1;
   assign m252_1 =15'b0;

   // m252_2 = W*in
   wire signed [14:0] m252_2;
   assign m252_2 =15'b0;

   // m252_3 = W*in
   wire signed [14:0] m252_3;
   assign m252_3 =15'b0;

   // m252_4 = W*in
   wire signed [14:0] m252_4;
   assign m252_4 =15'b0;

   // m252_5 = W*in
   wire signed [14:0] m252_5;
   assign m252_5 =15'b0;

   // m252_6 = W*in
   wire signed [14:0] m252_6;
   assign m252_6 =15'b0;

   // m252_7 = W*in
   wire signed [14:0] m252_7;
   assign m252_7 =15'b0;

   // m252_8 = W*in
   wire signed [14:0] m252_8;
   assign m252_8 ={ {3{neg252[14]}} , neg252[14:3] };

   // m252_9 = W*in
   wire signed [14:0] m252_9;
   assign m252_9 =15'b0;

   // m252_10 = W*in
   wire signed [14:0] m252_10;
   assign m252_10 =15'b0;

   // m252_11 = W*in
   wire signed [14:0] m252_11;
   assign m252_11 ={ {3{in252[14]}} , in252[14:3] };

   // m252_12 = W*in
   wire signed [14:0] m252_12;
   assign m252_12 =15'b0;

   // m252_13 = W*in
   wire signed [14:0] m252_13;
   assign m252_13 =15'b0;

   // m252_14 = W*in
   wire signed [14:0] m252_14;
   assign m252_14 =15'b0;

   // m252_15 = W*in
   wire signed [14:0] m252_15;
   assign m252_15 ={ {3{in252[14]}} , in252[14:3] };

   // m252_16 = W*in
   wire signed [14:0] m252_16;
   assign m252_16 =15'b0;

   // m252_17 = W*in
   wire signed [14:0] m252_17;
   assign m252_17 =15'b0;

   // m252_18 = W*in
   wire signed [14:0] m252_18;
   assign m252_18 =15'b0;

   // m252_19 = W*in
   wire signed [14:0] m252_19;
   assign m252_19 =15'b0;

   // m252_20 = W*in
   wire signed [14:0] m252_20;
   assign m252_20 =15'b0;

   // m252_21 = W*in
   wire signed [14:0] m252_21;
   assign m252_21 =15'b0;

   // m252_22 = W*in
   wire signed [14:0] m252_22;
   assign m252_22 =15'b0;

   // m252_23 = W*in
   wire signed [14:0] m252_23;
   assign m252_23 ={ {3{neg252[14]}} , neg252[14:3] };

   // m252_24 = W*in
   wire signed [14:0] m252_24;
   assign m252_24 =15'b0;

   // m252_25 = W*in
   wire signed [14:0] m252_25;
   assign m252_25 =15'b0;

   // m252_26 = W*in
   wire signed [14:0] m252_26;
   assign m252_26 =15'b0;

   // m252_27 = W*in
   wire signed [14:0] m252_27;
   assign m252_27 =15'b0;

   // m252_28 = W*in
   wire signed [14:0] m252_28;
   assign m252_28 =15'b0;

   // m252_29 = W*in
   wire signed [14:0] m252_29;
   assign m252_29 ={ {4{neg252[14]}} , neg252[14:4] };

   // m252_30 = W*in
   wire signed [14:0] m252_30;
   assign m252_30 =15'b0;

   // m252_31 = W*in
   wire signed [14:0] m252_31;
   assign m252_31 =15'b0;

   // m252_32 = W*in
   wire signed [14:0] m252_32;
   assign m252_32 =15'b0;

   // m252_33 = W*in
   wire signed [14:0] m252_33;
   assign m252_33 =15'b0;

   // m252_34 = W*in
   wire signed [14:0] m252_34;
   assign m252_34 =15'b0;

   // m252_35 = W*in
   wire signed [14:0] m252_35;
   assign m252_35 =15'b0;

   // m252_36 = W*in
   wire signed [14:0] m252_36;
   assign m252_36 =15'b0;

   // m252_37 = W*in
   wire signed [14:0] m252_37;
   assign m252_37 =15'b0;

   // m252_38 = W*in
   wire signed [14:0] m252_38;
   assign m252_38 =15'b0;

   // m252_39 = W*in
   wire signed [14:0] m252_39;
   assign m252_39 =15'b0;

   // m252_40 = W*in
   wire signed [14:0] m252_40;
   assign m252_40 =15'b0;

   // m252_41 = W*in
   wire signed [14:0] m252_41;
   assign m252_41 =15'b0;

   // m252_42 = W*in
   wire signed [14:0] m252_42;
   assign m252_42 =15'b0;

   // m252_43 = W*in
   wire signed [14:0] m252_43;
   assign m252_43 =15'b0;

   // m252_44 = W*in
   wire signed [14:0] m252_44;
   assign m252_44 =15'b0;

   // m252_45 = W*in
   wire signed [14:0] m252_45;
   assign m252_45 =15'b0;

   // m252_46 = W*in
   wire signed [14:0] m252_46;
   assign m252_46 ={ {4{neg252[14]}} , neg252[14:4] };

   // m252_47 = W*in
   wire signed [14:0] m252_47;
   assign m252_47 =15'b0;

   // m252_48 = W*in
   wire signed [14:0] m252_48;
   assign m252_48 =15'b0;

   // m252_49 = W*in
   wire signed [14:0] m252_49;
   assign m252_49 =15'b0;

   // m252_50 = W*in
   wire signed [14:0] m252_50;
   assign m252_50 =15'b0;

   // m252_51 = W*in
   wire signed [14:0] m252_51;
   assign m252_51 =15'b0;

   // m252_52 = W*in
   wire signed [14:0] m252_52;
   assign m252_52 =15'b0;

   // m252_53 = W*in
   wire signed [14:0] m252_53;
   assign m252_53 =15'b0;

   // m252_54 = W*in
   wire signed [14:0] m252_54;
   assign m252_54 =15'b0;

   // m252_55 = W*in
   wire signed [14:0] m252_55;
   assign m252_55 =15'b0;

   // m252_56 = W*in
   wire signed [14:0] m252_56;
   assign m252_56 =15'b0;

   // m252_57 = W*in
   wire signed [14:0] m252_57;
   assign m252_57 ={ {4{neg252[14]}} , neg252[14:4] };

   // m252_58 = W*in
   wire signed [14:0] m252_58;
   assign m252_58 =15'b0;

   // m252_59 = W*in
   wire signed [14:0] m252_59;
   assign m252_59 =15'b0;

   // m252_60 = W*in
   wire signed [14:0] m252_60;
   assign m252_60 =15'b0;

   // m252_61 = W*in
   wire signed [14:0] m252_61;
   assign m252_61 ={ {3{in252[14]}} , in252[14:3] };

   // m252_62 = W*in
   wire signed [14:0] m252_62;
   assign m252_62 =15'b0;

   // m252_63 = W*in
   wire signed [14:0] m252_63;
   assign m252_63 ={ {4{neg252[14]}} , neg252[14:4] };

   // m252_64 = W*in
   wire signed [14:0] m252_64;
   assign m252_64 ={ {3{in252[14]}} , in252[14:3] };

   // m252_65 = W*in
   wire signed [14:0] m252_65;
   assign m252_65 =15'b0;

   // m252_66 = W*in
   wire signed [14:0] m252_66;
   assign m252_66 =15'b0;

   // m252_67 = W*in
   wire signed [14:0] m252_67;
   assign m252_67 ={ {3{in252[14]}} , in252[14:3] };

   // m252_68 = W*in
   wire signed [14:0] m252_68;
   assign m252_68 ={ {4{in252[14]}} , in252[14:4] };

   // m252_69 = W*in
   wire signed [14:0] m252_69;
   assign m252_69 ={ {3{in252[14]}} , in252[14:3] };

   // m252_70 = W*in
   wire signed [14:0] m252_70;
   assign m252_70 =15'b0;

   // m252_71 = W*in
   wire signed [14:0] m252_71;
   assign m252_71 =15'b0;

   // m252_72 = W*in
   wire signed [14:0] m252_72;
   assign m252_72 =15'b0;

   // m252_73 = W*in
   wire signed [14:0] m252_73;
   assign m252_73 ={ {3{in252[14]}} , in252[14:3] };

   // m252_74 = W*in
   wire signed [14:0] m252_74;
   assign m252_74 ={ {4{neg252[14]}} , neg252[14:4] };

   // m252_75 = W*in
   wire signed [14:0] m252_75;
   assign m252_75 =15'b0;

   // m252_76 = W*in
   wire signed [14:0] m252_76;
   assign m252_76 ={ {3{neg252[14]}} , neg252[14:3] };

   // m252_77 = W*in
   wire signed [14:0] m252_77;
   assign m252_77 =15'b0;

   // m252_78 = W*in
   wire signed [14:0] m252_78;
   assign m252_78 ={ {4{in252[14]}} , in252[14:4] };

   // m252_79 = W*in
   wire signed [14:0] m252_79;
   assign m252_79 =15'b0;

   // m252_80 = W*in
   wire signed [14:0] m252_80;
   assign m252_80 =15'b0;

   // m252_81 = W*in
   wire signed [14:0] m252_81;
   assign m252_81 =15'b0;

   // m252_82 = W*in
   wire signed [14:0] m252_82;
   assign m252_82 =15'b0;

   // m252_83 = W*in
   wire signed [14:0] m252_83;
   assign m252_83 =15'b0;

   // m252_84 = W*in
   wire signed [14:0] m252_84;
   assign m252_84 =15'b0;

   // m252_85 = W*in
   wire signed [14:0] m252_85;
   assign m252_85 =15'b0;

   // m252_86 = W*in
   wire signed [14:0] m252_86;
   assign m252_86 =15'b0;

   // m252_87 = W*in
   wire signed [14:0] m252_87;
   assign m252_87 =15'b0;

   // m252_88 = W*in
   wire signed [14:0] m252_88;
   assign m252_88 ={ {3{neg252[14]}} , neg252[14:3] };

   // m252_89 = W*in
   wire signed [14:0] m252_89;
   assign m252_89 =15'b0;

   // m252_90 = W*in
   wire signed [14:0] m252_90;
   assign m252_90 =15'b0;

   // m252_91 = W*in
   wire signed [14:0] m252_91;
   assign m252_91 =15'b0;

   // m252_92 = W*in
   wire signed [14:0] m252_92;
   assign m252_92 ={ {3{in252[14]}} , in252[14:3] };

   // m252_93 = W*in
   wire signed [14:0] m252_93;
   assign m252_93 ={ {4{neg252[14]}} , neg252[14:4] };

   // m252_94 = W*in
   wire signed [14:0] m252_94;
   assign m252_94 =15'b0;

   // m252_95 = W*in
   wire signed [14:0] m252_95;
   assign m252_95 =15'b0;

   // m252_96 = W*in
   wire signed [14:0] m252_96;
   assign m252_96 =15'b0;

   // m252_97 = W*in
   wire signed [14:0] m252_97;
   assign m252_97 =15'b0;

   // m252_98 = W*in
   wire signed [14:0] m252_98;
   assign m252_98 ={ {3{in252[14]}} , in252[14:3] };

   // m252_99 = W*in
   wire signed [14:0] m252_99;
   assign m252_99 =15'b0;

   // m252_100 = W*in
   wire signed [14:0] m252_100;
   assign m252_100 ={ {3{neg252[14]}} , neg252[14:3] };

   // m253_1 = W*in
   wire signed [14:0] m253_1;
   assign m253_1 =15'b0;

   // m253_2 = W*in
   wire signed [14:0] m253_2;
   assign m253_2 =15'b0;

   // m253_3 = W*in
   wire signed [14:0] m253_3;
   assign m253_3 =15'b0;

   // m253_4 = W*in
   wire signed [14:0] m253_4;
   assign m253_4 =15'b0;

   // m253_5 = W*in
   wire signed [14:0] m253_5;
   assign m253_5 ={ {3{in253[14]}} , in253[14:3] };

   // m253_6 = W*in
   wire signed [14:0] m253_6;
   assign m253_6 ={ {4{neg253[14]}} , neg253[14:4] };

   // m253_7 = W*in
   wire signed [14:0] m253_7;
   assign m253_7 =15'b0;

   // m253_8 = W*in
   wire signed [14:0] m253_8;
   assign m253_8 =15'b0;

   // m253_9 = W*in
   wire signed [14:0] m253_9;
   assign m253_9 =15'b0;

   // m253_10 = W*in
   wire signed [14:0] m253_10;
   assign m253_10 =15'b0;

   // m253_11 = W*in
   wire signed [14:0] m253_11;
   assign m253_11 =15'b0;

   // m253_12 = W*in
   wire signed [14:0] m253_12;
   assign m253_12 =15'b0;

   // m253_13 = W*in
   wire signed [14:0] m253_13;
   assign m253_13 ={ {4{in253[14]}} , in253[14:4] };

   // m253_14 = W*in
   wire signed [14:0] m253_14;
   assign m253_14 =15'b0;

   // m253_15 = W*in
   wire signed [14:0] m253_15;
   assign m253_15 =15'b0;

   // m253_16 = W*in
   wire signed [14:0] m253_16;
   assign m253_16 =15'b0;

   // m253_17 = W*in
   wire signed [14:0] m253_17;
   assign m253_17 =15'b0;

   // m253_18 = W*in
   wire signed [14:0] m253_18;
   assign m253_18 =15'b0;

   // m253_19 = W*in
   wire signed [14:0] m253_19;
   assign m253_19 =15'b0;

   // m253_20 = W*in
   wire signed [14:0] m253_20;
   assign m253_20 =15'b0;

   // m253_21 = W*in
   wire signed [14:0] m253_21;
   assign m253_21 =15'b0;

   // m253_22 = W*in
   wire signed [14:0] m253_22;
   assign m253_22 =15'b0;

   // m253_23 = W*in
   wire signed [14:0] m253_23;
   assign m253_23 =15'b0;

   // m253_24 = W*in
   wire signed [14:0] m253_24;
   assign m253_24 =15'b0;

   // m253_25 = W*in
   wire signed [14:0] m253_25;
   assign m253_25 =15'b0;

   // m253_26 = W*in
   wire signed [14:0] m253_26;
   assign m253_26 =15'b0;

   // m253_27 = W*in
   wire signed [14:0] m253_27;
   assign m253_27 =15'b0;

   // m253_28 = W*in
   wire signed [14:0] m253_28;
   assign m253_28 ={ {4{neg253[14]}} , neg253[14:4] };

   // m253_29 = W*in
   wire signed [14:0] m253_29;
   assign m253_29 =15'b0;

   // m253_30 = W*in
   wire signed [14:0] m253_30;
   assign m253_30 =15'b0;

   // m253_31 = W*in
   wire signed [14:0] m253_31;
   assign m253_31 =15'b0;

   // m253_32 = W*in
   wire signed [14:0] m253_32;
   assign m253_32 =15'b0;

   // m253_33 = W*in
   wire signed [14:0] m253_33;
   assign m253_33 =15'b0;

   // m253_34 = W*in
   wire signed [14:0] m253_34;
   assign m253_34 =15'b0;

   // m253_35 = W*in
   wire signed [14:0] m253_35;
   assign m253_35 =15'b0;

   // m253_36 = W*in
   wire signed [14:0] m253_36;
   assign m253_36 =15'b0;

   // m253_37 = W*in
   wire signed [14:0] m253_37;
   assign m253_37 =15'b0;

   // m253_38 = W*in
   wire signed [14:0] m253_38;
   assign m253_38 =15'b0;

   // m253_39 = W*in
   wire signed [14:0] m253_39;
   assign m253_39 =15'b0;

   // m253_40 = W*in
   wire signed [14:0] m253_40;
   assign m253_40 =15'b0;

   // m253_41 = W*in
   wire signed [14:0] m253_41;
   assign m253_41 =15'b0;

   // m253_42 = W*in
   wire signed [14:0] m253_42;
   assign m253_42 =15'b0;

   // m253_43 = W*in
   wire signed [14:0] m253_43;
   assign m253_43 =15'b0;

   // m253_44 = W*in
   wire signed [14:0] m253_44;
   assign m253_44 =15'b0;

   // m253_45 = W*in
   wire signed [14:0] m253_45;
   assign m253_45 =15'b0;

   // m253_46 = W*in
   wire signed [14:0] m253_46;
   assign m253_46 =15'b0;

   // m253_47 = W*in
   wire signed [14:0] m253_47;
   assign m253_47 =15'b0;

   // m253_48 = W*in
   wire signed [14:0] m253_48;
   assign m253_48 =15'b0;

   // m253_49 = W*in
   wire signed [14:0] m253_49;
   assign m253_49 =15'b0;

   // m253_50 = W*in
   wire signed [14:0] m253_50;
   assign m253_50 =15'b0;

   // m253_51 = W*in
   wire signed [14:0] m253_51;
   assign m253_51 =15'b0;

   // m253_52 = W*in
   wire signed [14:0] m253_52;
   assign m253_52 =15'b0;

   // m253_53 = W*in
   wire signed [14:0] m253_53;
   assign m253_53 =15'b0;

   // m253_54 = W*in
   wire signed [14:0] m253_54;
   assign m253_54 =15'b0;

   // m253_55 = W*in
   wire signed [14:0] m253_55;
   assign m253_55 =15'b0;

   // m253_56 = W*in
   wire signed [14:0] m253_56;
   assign m253_56 =15'b0;

   // m253_57 = W*in
   wire signed [14:0] m253_57;
   assign m253_57 =15'b0;

   // m253_58 = W*in
   wire signed [14:0] m253_58;
   assign m253_58 =15'b0;

   // m253_59 = W*in
   wire signed [14:0] m253_59;
   assign m253_59 =15'b0;

   // m253_60 = W*in
   wire signed [14:0] m253_60;
   assign m253_60 =15'b0;

   // m253_61 = W*in
   wire signed [14:0] m253_61;
   assign m253_61 =15'b0;

   // m253_62 = W*in
   wire signed [14:0] m253_62;
   assign m253_62 =15'b0;

   // m253_63 = W*in
   wire signed [14:0] m253_63;
   assign m253_63 =15'b0;

   // m253_64 = W*in
   wire signed [14:0] m253_64;
   assign m253_64 ={ {3{in253[14]}} , in253[14:3] };

   // m253_65 = W*in
   wire signed [14:0] m253_65;
   assign m253_65 =15'b0;

   // m253_66 = W*in
   wire signed [14:0] m253_66;
   assign m253_66 =15'b0;

   // m253_67 = W*in
   wire signed [14:0] m253_67;
   assign m253_67 =15'b0;

   // m253_68 = W*in
   wire signed [14:0] m253_68;
   assign m253_68 =15'b0;

   // m253_69 = W*in
   wire signed [14:0] m253_69;
   assign m253_69 =15'b0;

   // m253_70 = W*in
   wire signed [14:0] m253_70;
   assign m253_70 =15'b0;

   // m253_71 = W*in
   wire signed [14:0] m253_71;
   assign m253_71 =15'b0;

   // m253_72 = W*in
   wire signed [14:0] m253_72;
   assign m253_72 =15'b0;

   // m253_73 = W*in
   wire signed [14:0] m253_73;
   assign m253_73 =15'b0;

   // m253_74 = W*in
   wire signed [14:0] m253_74;
   assign m253_74 =15'b0;

   // m253_75 = W*in
   wire signed [14:0] m253_75;
   assign m253_75 =15'b0;

   // m253_76 = W*in
   wire signed [14:0] m253_76;
   assign m253_76 =15'b0;

   // m253_77 = W*in
   wire signed [14:0] m253_77;
   assign m253_77 ={ {4{neg253[14]}} , neg253[14:4] };

   // m253_78 = W*in
   wire signed [14:0] m253_78;
   assign m253_78 =15'b0;

   // m253_79 = W*in
   wire signed [14:0] m253_79;
   assign m253_79 =15'b0;

   // m253_80 = W*in
   wire signed [14:0] m253_80;
   assign m253_80 =15'b0;

   // m253_81 = W*in
   wire signed [14:0] m253_81;
   assign m253_81 =15'b0;

   // m253_82 = W*in
   wire signed [14:0] m253_82;
   assign m253_82 =15'b0;

   // m253_83 = W*in
   wire signed [14:0] m253_83;
   assign m253_83 =15'b0;

   // m253_84 = W*in
   wire signed [14:0] m253_84;
   assign m253_84 =15'b0;

   // m253_85 = W*in
   wire signed [14:0] m253_85;
   assign m253_85 =15'b0;

   // m253_86 = W*in
   wire signed [14:0] m253_86;
   assign m253_86 ={ {3{neg253[14]}} , neg253[14:3] };

   // m253_87 = W*in
   wire signed [14:0] m253_87;
   assign m253_87 ={ {3{in253[14]}} , in253[14:3] };

   // m253_88 = W*in
   wire signed [14:0] m253_88;
   assign m253_88 ={ {3{neg253[14]}} , neg253[14:3] };

   // m253_89 = W*in
   wire signed [14:0] m253_89;
   assign m253_89 =15'b0;

   // m253_90 = W*in
   wire signed [14:0] m253_90;
   assign m253_90 =15'b0;

   // m253_91 = W*in
   wire signed [14:0] m253_91;
   assign m253_91 =15'b0;

   // m253_92 = W*in
   wire signed [14:0] m253_92;
   assign m253_92 =15'b0;

   // m253_93 = W*in
   wire signed [14:0] m253_93;
   assign m253_93 =15'b0;

   // m253_94 = W*in
   wire signed [14:0] m253_94;
   assign m253_94 =15'b0;

   // m253_95 = W*in
   wire signed [14:0] m253_95;
   assign m253_95 =15'b0;

   // m253_96 = W*in
   wire signed [14:0] m253_96;
   assign m253_96 =15'b0;

   // m253_97 = W*in
   wire signed [14:0] m253_97;
   assign m253_97 =15'b0;

   // m253_98 = W*in
   wire signed [14:0] m253_98;
   assign m253_98 =15'b0;

   // m253_99 = W*in
   wire signed [14:0] m253_99;
   assign m253_99 =15'b0;

   // m253_100 = W*in
   wire signed [14:0] m253_100;
   assign m253_100 =15'b0;

   // m254_1 = W*in
   wire signed [14:0] m254_1;
   assign m254_1 =15'b0;

   // m254_2 = W*in
   wire signed [14:0] m254_2;
   assign m254_2 =15'b0;

   // m254_3 = W*in
   wire signed [14:0] m254_3;
   assign m254_3 =15'b0;

   // m254_4 = W*in
   wire signed [14:0] m254_4;
   assign m254_4 =15'b0;

   // m254_5 = W*in
   wire signed [14:0] m254_5;
   assign m254_5 =15'b0;

   // m254_6 = W*in
   wire signed [14:0] m254_6;
   assign m254_6 =15'b0;

   // m254_7 = W*in
   wire signed [14:0] m254_7;
   assign m254_7 =15'b0;

   // m254_8 = W*in
   wire signed [14:0] m254_8;
   assign m254_8 =15'b0;

   // m254_9 = W*in
   wire signed [14:0] m254_9;
   assign m254_9 =15'b0;

   // m254_10 = W*in
   wire signed [14:0] m254_10;
   assign m254_10 ={ {2{in254[14]}} , in254[14:2] };

   // m254_11 = W*in
   wire signed [14:0] m254_11;
   assign m254_11 =15'b0;

   // m254_12 = W*in
   wire signed [14:0] m254_12;
   assign m254_12 =15'b0;

   // m254_13 = W*in
   wire signed [14:0] m254_13;
   assign m254_13 =15'b0;

   // m254_14 = W*in
   wire signed [14:0] m254_14;
   assign m254_14 =15'b0;

   // m254_15 = W*in
   wire signed [14:0] m254_15;
   assign m254_15 =15'b0;

   // m254_16 = W*in
   wire signed [14:0] m254_16;
   assign m254_16 =15'b0;

   // m254_17 = W*in
   wire signed [14:0] m254_17;
   assign m254_17 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_18 = W*in
   wire signed [14:0] m254_18;
   assign m254_18 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_19 = W*in
   wire signed [14:0] m254_19;
   assign m254_19 ={ {4{in254[14]}} , in254[14:4] };

   // m254_20 = W*in
   wire signed [14:0] m254_20;
   assign m254_20 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_21 = W*in
   wire signed [14:0] m254_21;
   assign m254_21 =15'b0;

   // m254_22 = W*in
   wire signed [14:0] m254_22;
   assign m254_22 =15'b0;

   // m254_23 = W*in
   wire signed [14:0] m254_23;
   assign m254_23 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_24 = W*in
   wire signed [14:0] m254_24;
   assign m254_24 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_25 = W*in
   wire signed [14:0] m254_25;
   assign m254_25 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_26 = W*in
   wire signed [14:0] m254_26;
   assign m254_26 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_27 = W*in
   wire signed [14:0] m254_27;
   assign m254_27 =15'b0;

   // m254_28 = W*in
   wire signed [14:0] m254_28;
   assign m254_28 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_29 = W*in
   wire signed [14:0] m254_29;
   assign m254_29 =15'b0;

   // m254_30 = W*in
   wire signed [14:0] m254_30;
   assign m254_30 =15'b0;

   // m254_31 = W*in
   wire signed [14:0] m254_31;
   assign m254_31 =15'b0;

   // m254_32 = W*in
   wire signed [14:0] m254_32;
   assign m254_32 ={ {4{in254[14]}} , in254[14:4] };

   // m254_33 = W*in
   wire signed [14:0] m254_33;
   assign m254_33 =15'b0;

   // m254_34 = W*in
   wire signed [14:0] m254_34;
   assign m254_34 =15'b0;

   // m254_35 = W*in
   wire signed [14:0] m254_35;
   assign m254_35 =15'b0;

   // m254_36 = W*in
   wire signed [14:0] m254_36;
   assign m254_36 =15'b0;

   // m254_37 = W*in
   wire signed [14:0] m254_37;
   assign m254_37 =15'b0;

   // m254_38 = W*in
   wire signed [14:0] m254_38;
   assign m254_38 =15'b0;

   // m254_39 = W*in
   wire signed [14:0] m254_39;
   assign m254_39 =15'b0;

   // m254_40 = W*in
   wire signed [14:0] m254_40;
   assign m254_40 =15'b0;

   // m254_41 = W*in
   wire signed [14:0] m254_41;
   assign m254_41 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_42 = W*in
   wire signed [14:0] m254_42;
   assign m254_42 =15'b0;

   // m254_43 = W*in
   wire signed [14:0] m254_43;
   assign m254_43 ={ {3{in254[14]}} , in254[14:3] };

   // m254_44 = W*in
   wire signed [14:0] m254_44;
   assign m254_44 =15'b0;

   // m254_45 = W*in
   wire signed [14:0] m254_45;
   assign m254_45 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_46 = W*in
   wire signed [14:0] m254_46;
   assign m254_46 ={ {3{in254[14]}} , in254[14:3] };

   // m254_47 = W*in
   wire signed [14:0] m254_47;
   assign m254_47 =15'b0;

   // m254_48 = W*in
   wire signed [14:0] m254_48;
   assign m254_48 =15'b0;

   // m254_49 = W*in
   wire signed [14:0] m254_49;
   assign m254_49 =15'b0;

   // m254_50 = W*in
   wire signed [14:0] m254_50;
   assign m254_50 =15'b0;

   // m254_51 = W*in
   wire signed [14:0] m254_51;
   assign m254_51 =15'b0;

   // m254_52 = W*in
   wire signed [14:0] m254_52;
   assign m254_52 =15'b0;

   // m254_53 = W*in
   wire signed [14:0] m254_53;
   assign m254_53 =15'b0;

   // m254_54 = W*in
   wire signed [14:0] m254_54;
   assign m254_54 =15'b0;

   // m254_55 = W*in
   wire signed [14:0] m254_55;
   assign m254_55 =15'b0;

   // m254_56 = W*in
   wire signed [14:0] m254_56;
   assign m254_56 =15'b0;

   // m254_57 = W*in
   wire signed [14:0] m254_57;
   assign m254_57 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_58 = W*in
   wire signed [14:0] m254_58;
   assign m254_58 =15'b0;

   // m254_59 = W*in
   wire signed [14:0] m254_59;
   assign m254_59 =15'b0;

   // m254_60 = W*in
   wire signed [14:0] m254_60;
   assign m254_60 =15'b0;

   // m254_61 = W*in
   wire signed [14:0] m254_61;
   assign m254_61 =15'b0;

   // m254_62 = W*in
   wire signed [14:0] m254_62;
   assign m254_62 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_63 = W*in
   wire signed [14:0] m254_63;
   assign m254_63 ={ {3{in254[14]}} , in254[14:3] };

   // m254_64 = W*in
   wire signed [14:0] m254_64;
   assign m254_64 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_65 = W*in
   wire signed [14:0] m254_65;
   assign m254_65 =15'b0;

   // m254_66 = W*in
   wire signed [14:0] m254_66;
   assign m254_66 ={ {3{in254[14]}} , in254[14:3] };

   // m254_67 = W*in
   wire signed [14:0] m254_67;
   assign m254_67 =15'b0;

   // m254_68 = W*in
   wire signed [14:0] m254_68;
   assign m254_68 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_69 = W*in
   wire signed [14:0] m254_69;
   assign m254_69 ={ {4{in254[14]}} , in254[14:4] };

   // m254_70 = W*in
   wire signed [14:0] m254_70;
   assign m254_70 =15'b0;

   // m254_71 = W*in
   wire signed [14:0] m254_71;
   assign m254_71 =15'b0;

   // m254_72 = W*in
   wire signed [14:0] m254_72;
   assign m254_72 =15'b0;

   // m254_73 = W*in
   wire signed [14:0] m254_73;
   assign m254_73 =15'b0;

   // m254_74 = W*in
   wire signed [14:0] m254_74;
   assign m254_74 =15'b0;

   // m254_75 = W*in
   wire signed [14:0] m254_75;
   assign m254_75 =15'b0;

   // m254_76 = W*in
   wire signed [14:0] m254_76;
   assign m254_76 =15'b0;

   // m254_77 = W*in
   wire signed [14:0] m254_77;
   assign m254_77 =15'b0;

   // m254_78 = W*in
   wire signed [14:0] m254_78;
   assign m254_78 ={ {4{neg254[14]}} , neg254[14:4] };

   // m254_79 = W*in
   wire signed [14:0] m254_79;
   assign m254_79 ={ {3{in254[14]}} , in254[14:3] };

   // m254_80 = W*in
   wire signed [14:0] m254_80;
   assign m254_80 ={ {3{in254[14]}} , in254[14:3] };

   // m254_81 = W*in
   wire signed [14:0] m254_81;
   assign m254_81 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_82 = W*in
   wire signed [14:0] m254_82;
   assign m254_82 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_83 = W*in
   wire signed [14:0] m254_83;
   assign m254_83 ={ {3{in254[14]}} , in254[14:3] };

   // m254_84 = W*in
   wire signed [14:0] m254_84;
   assign m254_84 ={ {3{in254[14]}} , in254[14:3] };

   // m254_85 = W*in
   wire signed [14:0] m254_85;
   assign m254_85 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_86 = W*in
   wire signed [14:0] m254_86;
   assign m254_86 =15'b0;

   // m254_87 = W*in
   wire signed [14:0] m254_87;
   assign m254_87 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_88 = W*in
   wire signed [14:0] m254_88;
   assign m254_88 ={ {3{neg254[14]}} , neg254[14:3] };

   // m254_89 = W*in
   wire signed [14:0] m254_89;
   assign m254_89 =15'b0;

   // m254_90 = W*in
   wire signed [14:0] m254_90;
   assign m254_90 =15'b0;

   // m254_91 = W*in
   wire signed [14:0] m254_91;
   assign m254_91 =15'b0;

   // m254_92 = W*in
   wire signed [14:0] m254_92;
   assign m254_92 =15'b0;

   // m254_93 = W*in
   wire signed [14:0] m254_93;
   assign m254_93 ={ {3{in254[14]}} , in254[14:3] };

   // m254_94 = W*in
   wire signed [14:0] m254_94;
   assign m254_94 =15'b0;

   // m254_95 = W*in
   wire signed [14:0] m254_95;
   assign m254_95 =15'b0;

   // m254_96 = W*in
   wire signed [14:0] m254_96;
   assign m254_96 =15'b0;

   // m254_97 = W*in
   wire signed [14:0] m254_97;
   assign m254_97 =15'b0;

   // m254_98 = W*in
   wire signed [14:0] m254_98;
   assign m254_98 =15'b0;

   // m254_99 = W*in
   wire signed [14:0] m254_99;
   assign m254_99 =15'b0;

   // m254_100 = W*in
   wire signed [14:0] m254_100;
   assign m254_100 ={ {3{in254[14]}} , in254[14:3] };

   // m255_1 = W*in
   wire signed [14:0] m255_1;
   assign m255_1 =15'b0;

   // m255_2 = W*in
   wire signed [14:0] m255_2;
   assign m255_2 =15'b0;

   // m255_3 = W*in
   wire signed [14:0] m255_3;
   assign m255_3 =15'b0;

   // m255_4 = W*in
   wire signed [14:0] m255_4;
   assign m255_4 =15'b0;

   // m255_5 = W*in
   wire signed [14:0] m255_5;
   assign m255_5 =15'b0;

   // m255_6 = W*in
   wire signed [14:0] m255_6;
   assign m255_6 =15'b0;

   // m255_7 = W*in
   wire signed [14:0] m255_7;
   assign m255_7 =15'b0;

   // m255_8 = W*in
   wire signed [14:0] m255_8;
   assign m255_8 =15'b0;

   // m255_9 = W*in
   wire signed [14:0] m255_9;
   assign m255_9 =15'b0;

   // m255_10 = W*in
   wire signed [14:0] m255_10;
   assign m255_10 ={ {3{in255[14]}} , in255[14:3] };

   // m255_11 = W*in
   wire signed [14:0] m255_11;
   assign m255_11 =15'b0;

   // m255_12 = W*in
   wire signed [14:0] m255_12;
   assign m255_12 =15'b0;

   // m255_13 = W*in
   wire signed [14:0] m255_13;
   assign m255_13 =15'b0;

   // m255_14 = W*in
   wire signed [14:0] m255_14;
   assign m255_14 =15'b0;

   // m255_15 = W*in
   wire signed [14:0] m255_15;
   assign m255_15 =15'b0;

   // m255_16 = W*in
   wire signed [14:0] m255_16;
   assign m255_16 =15'b0;

   // m255_17 = W*in
   wire signed [14:0] m255_17;
   assign m255_17 =15'b0;

   // m255_18 = W*in
   wire signed [14:0] m255_18;
   assign m255_18 =15'b0;

   // m255_19 = W*in
   wire signed [14:0] m255_19;
   assign m255_19 ={ {4{in255[14]}} , in255[14:4] };

   // m255_20 = W*in
   wire signed [14:0] m255_20;
   assign m255_20 =15'b0;

   // m255_21 = W*in
   wire signed [14:0] m255_21;
   assign m255_21 =15'b0;

   // m255_22 = W*in
   wire signed [14:0] m255_22;
   assign m255_22 =15'b0;

   // m255_23 = W*in
   wire signed [14:0] m255_23;
   assign m255_23 =15'b0;

   // m255_24 = W*in
   wire signed [14:0] m255_24;
   assign m255_24 ={ {3{neg255[14]}} , neg255[14:3] };

   // m255_25 = W*in
   wire signed [14:0] m255_25;
   assign m255_25 =15'b0;

   // m255_26 = W*in
   wire signed [14:0] m255_26;
   assign m255_26 =15'b0;

   // m255_27 = W*in
   wire signed [14:0] m255_27;
   assign m255_27 =15'b0;

   // m255_28 = W*in
   wire signed [14:0] m255_28;
   assign m255_28 =15'b0;

   // m255_29 = W*in
   wire signed [14:0] m255_29;
   assign m255_29 =15'b0;

   // m255_30 = W*in
   wire signed [14:0] m255_30;
   assign m255_30 =15'b0;

   // m255_31 = W*in
   wire signed [14:0] m255_31;
   assign m255_31 =15'b0;

   // m255_32 = W*in
   wire signed [14:0] m255_32;
   assign m255_32 =15'b0;

   // m255_33 = W*in
   wire signed [14:0] m255_33;
   assign m255_33 =15'b0;

   // m255_34 = W*in
   wire signed [14:0] m255_34;
   assign m255_34 =15'b0;

   // m255_35 = W*in
   wire signed [14:0] m255_35;
   assign m255_35 =15'b0;

   // m255_36 = W*in
   wire signed [14:0] m255_36;
   assign m255_36 =15'b0;

   // m255_37 = W*in
   wire signed [14:0] m255_37;
   assign m255_37 =15'b0;

   // m255_38 = W*in
   wire signed [14:0] m255_38;
   assign m255_38 =15'b0;

   // m255_39 = W*in
   wire signed [14:0] m255_39;
   assign m255_39 =15'b0;

   // m255_40 = W*in
   wire signed [14:0] m255_40;
   assign m255_40 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_41 = W*in
   wire signed [14:0] m255_41;
   assign m255_41 =15'b0;

   // m255_42 = W*in
   wire signed [14:0] m255_42;
   assign m255_42 =15'b0;

   // m255_43 = W*in
   wire signed [14:0] m255_43;
   assign m255_43 =15'b0;

   // m255_44 = W*in
   wire signed [14:0] m255_44;
   assign m255_44 =15'b0;

   // m255_45 = W*in
   wire signed [14:0] m255_45;
   assign m255_45 =15'b0;

   // m255_46 = W*in
   wire signed [14:0] m255_46;
   assign m255_46 ={ {4{in255[14]}} , in255[14:4] };

   // m255_47 = W*in
   wire signed [14:0] m255_47;
   assign m255_47 =15'b0;

   // m255_48 = W*in
   wire signed [14:0] m255_48;
   assign m255_48 =15'b0;

   // m255_49 = W*in
   wire signed [14:0] m255_49;
   assign m255_49 =15'b0;

   // m255_50 = W*in
   wire signed [14:0] m255_50;
   assign m255_50 =15'b0;

   // m255_51 = W*in
   wire signed [14:0] m255_51;
   assign m255_51 =15'b0;

   // m255_52 = W*in
   wire signed [14:0] m255_52;
   assign m255_52 =15'b0;

   // m255_53 = W*in
   wire signed [14:0] m255_53;
   assign m255_53 =15'b0;

   // m255_54 = W*in
   wire signed [14:0] m255_54;
   assign m255_54 =15'b0;

   // m255_55 = W*in
   wire signed [14:0] m255_55;
   assign m255_55 =15'b0;

   // m255_56 = W*in
   wire signed [14:0] m255_56;
   assign m255_56 =15'b0;

   // m255_57 = W*in
   wire signed [14:0] m255_57;
   assign m255_57 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_58 = W*in
   wire signed [14:0] m255_58;
   assign m255_58 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_59 = W*in
   wire signed [14:0] m255_59;
   assign m255_59 =15'b0;

   // m255_60 = W*in
   wire signed [14:0] m255_60;
   assign m255_60 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_61 = W*in
   wire signed [14:0] m255_61;
   assign m255_61 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_62 = W*in
   wire signed [14:0] m255_62;
   assign m255_62 ={ {3{neg255[14]}} , neg255[14:3] };

   // m255_63 = W*in
   wire signed [14:0] m255_63;
   assign m255_63 =15'b0;

   // m255_64 = W*in
   wire signed [14:0] m255_64;
   assign m255_64 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_65 = W*in
   wire signed [14:0] m255_65;
   assign m255_65 =15'b0;

   // m255_66 = W*in
   wire signed [14:0] m255_66;
   assign m255_66 ={ {4{in255[14]}} , in255[14:4] };

   // m255_67 = W*in
   wire signed [14:0] m255_67;
   assign m255_67 =15'b0;

   // m255_68 = W*in
   wire signed [14:0] m255_68;
   assign m255_68 ={ {4{neg255[14]}} , neg255[14:4] };

   // m255_69 = W*in
   wire signed [14:0] m255_69;
   assign m255_69 =15'b0;

   // m255_70 = W*in
   wire signed [14:0] m255_70;
   assign m255_70 ={ {4{in255[14]}} , in255[14:4] };

   // m255_71 = W*in
   wire signed [14:0] m255_71;
   assign m255_71 =15'b0;

   // m255_72 = W*in
   wire signed [14:0] m255_72;
   assign m255_72 =15'b0;

   // m255_73 = W*in
   wire signed [14:0] m255_73;
   assign m255_73 =15'b0;

   // m255_74 = W*in
   wire signed [14:0] m255_74;
   assign m255_74 =15'b0;

   // m255_75 = W*in
   wire signed [14:0] m255_75;
   assign m255_75 =15'b0;

   // m255_76 = W*in
   wire signed [14:0] m255_76;
   assign m255_76 =15'b0;

   // m255_77 = W*in
   wire signed [14:0] m255_77;
   assign m255_77 =15'b0;

   // m255_78 = W*in
   wire signed [14:0] m255_78;
   assign m255_78 =15'b0;

   // m255_79 = W*in
   wire signed [14:0] m255_79;
   assign m255_79 =15'b0;

   // m255_80 = W*in
   wire signed [14:0] m255_80;
   assign m255_80 =15'b0;

   // m255_81 = W*in
   wire signed [14:0] m255_81;
   assign m255_81 ={ {3{neg255[14]}} , neg255[14:3] };

   // m255_82 = W*in
   wire signed [14:0] m255_82;
   assign m255_82 =15'b0;

   // m255_83 = W*in
   wire signed [14:0] m255_83;
   assign m255_83 =15'b0;

   // m255_84 = W*in
   wire signed [14:0] m255_84;
   assign m255_84 =15'b0;

   // m255_85 = W*in
   wire signed [14:0] m255_85;
   assign m255_85 ={ {3{neg255[14]}} , neg255[14:3] };

   // m255_86 = W*in
   wire signed [14:0] m255_86;
   assign m255_86 =15'b0;

   // m255_87 = W*in
   wire signed [14:0] m255_87;
   assign m255_87 ={ {3{neg255[14]}} , neg255[14:3] };

   // m255_88 = W*in
   wire signed [14:0] m255_88;
   assign m255_88 =15'b0;

   // m255_89 = W*in
   wire signed [14:0] m255_89;
   assign m255_89 =15'b0;

   // m255_90 = W*in
   wire signed [14:0] m255_90;
   assign m255_90 =15'b0;

   // m255_91 = W*in
   wire signed [14:0] m255_91;
   assign m255_91 =15'b0;

   // m255_92 = W*in
   wire signed [14:0] m255_92;
   assign m255_92 =15'b0;

   // m255_93 = W*in
   wire signed [14:0] m255_93;
   assign m255_93 =15'b0;

   // m255_94 = W*in
   wire signed [14:0] m255_94;
   assign m255_94 =15'b0;

   // m255_95 = W*in
   wire signed [14:0] m255_95;
   assign m255_95 =15'b0;

   // m255_96 = W*in
   wire signed [14:0] m255_96;
   assign m255_96 =15'b0;

   // m255_97 = W*in
   wire signed [14:0] m255_97;
   assign m255_97 =15'b0;

   // m255_98 = W*in
   wire signed [14:0] m255_98;
   assign m255_98 =15'b0;

   // m255_99 = W*in
   wire signed [14:0] m255_99;
   assign m255_99 =15'b0;

   // m255_100 = W*in
   wire signed [14:0] m255_100;
   assign m255_100 =15'b0;

   // m256_1 = W*in
   wire signed [14:0] m256_1;
   assign m256_1 =15'b0;

   // m256_2 = W*in
   wire signed [14:0] m256_2;
   assign m256_2 =15'b0;

   // m256_3 = W*in
   wire signed [14:0] m256_3;
   assign m256_3 =15'b0;

   // m256_4 = W*in
   wire signed [14:0] m256_4;
   assign m256_4 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_5 = W*in
   wire signed [14:0] m256_5;
   assign m256_5 =15'b0;

   // m256_6 = W*in
   wire signed [14:0] m256_6;
   assign m256_6 =15'b0;

   // m256_7 = W*in
   wire signed [14:0] m256_7;
   assign m256_7 =15'b0;

   // m256_8 = W*in
   wire signed [14:0] m256_8;
   assign m256_8 =15'b0;

   // m256_9 = W*in
   wire signed [14:0] m256_9;
   assign m256_9 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_10 = W*in
   wire signed [14:0] m256_10;
   assign m256_10 =15'b0;

   // m256_11 = W*in
   wire signed [14:0] m256_11;
   assign m256_11 ={ {3{in256[14]}} , in256[14:3] };

   // m256_12 = W*in
   wire signed [14:0] m256_12;
   assign m256_12 =15'b0;

   // m256_13 = W*in
   wire signed [14:0] m256_13;
   assign m256_13 =15'b0;

   // m256_14 = W*in
   wire signed [14:0] m256_14;
   assign m256_14 =15'b0;

   // m256_15 = W*in
   wire signed [14:0] m256_15;
   assign m256_15 =15'b0;

   // m256_16 = W*in
   wire signed [14:0] m256_16;
   assign m256_16 ={ {3{in256[14]}} , in256[14:3] };

   // m256_17 = W*in
   wire signed [14:0] m256_17;
   assign m256_17 =15'b0;

   // m256_18 = W*in
   wire signed [14:0] m256_18;
   assign m256_18 =15'b0;

   // m256_19 = W*in
   wire signed [14:0] m256_19;
   assign m256_19 =15'b0;

   // m256_20 = W*in
   wire signed [14:0] m256_20;
   assign m256_20 =15'b0;

   // m256_21 = W*in
   wire signed [14:0] m256_21;
   assign m256_21 =15'b0;

   // m256_22 = W*in
   wire signed [14:0] m256_22;
   assign m256_22 ={ {3{in256[14]}} , in256[14:3] };

   // m256_23 = W*in
   wire signed [14:0] m256_23;
   assign m256_23 =15'b0;

   // m256_24 = W*in
   wire signed [14:0] m256_24;
   assign m256_24 ={ {4{in256[14]}} , in256[14:4] };

   // m256_25 = W*in
   wire signed [14:0] m256_25;
   assign m256_25 =15'b0;

   // m256_26 = W*in
   wire signed [14:0] m256_26;
   assign m256_26 =15'b0;

   // m256_27 = W*in
   wire signed [14:0] m256_27;
   assign m256_27 =15'b0;

   // m256_28 = W*in
   wire signed [14:0] m256_28;
   assign m256_28 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_29 = W*in
   wire signed [14:0] m256_29;
   assign m256_29 ={ {4{in256[14]}} , in256[14:4] };

   // m256_30 = W*in
   wire signed [14:0] m256_30;
   assign m256_30 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_31 = W*in
   wire signed [14:0] m256_31;
   assign m256_31 =15'b0;

   // m256_32 = W*in
   wire signed [14:0] m256_32;
   assign m256_32 ={ {4{neg256[14]}} , neg256[14:4] };

   // m256_33 = W*in
   wire signed [14:0] m256_33;
   assign m256_33 =15'b0;

   // m256_34 = W*in
   wire signed [14:0] m256_34;
   assign m256_34 =15'b0;

   // m256_35 = W*in
   wire signed [14:0] m256_35;
   assign m256_35 =15'b0;

   // m256_36 = W*in
   wire signed [14:0] m256_36;
   assign m256_36 =15'b0;

   // m256_37 = W*in
   wire signed [14:0] m256_37;
   assign m256_37 =15'b0;

   // m256_38 = W*in
   wire signed [14:0] m256_38;
   assign m256_38 =15'b0;

   // m256_39 = W*in
   wire signed [14:0] m256_39;
   assign m256_39 =15'b0;

   // m256_40 = W*in
   wire signed [14:0] m256_40;
   assign m256_40 =15'b0;

   // m256_41 = W*in
   wire signed [14:0] m256_41;
   assign m256_41 =15'b0;

   // m256_42 = W*in
   wire signed [14:0] m256_42;
   assign m256_42 =15'b0;

   // m256_43 = W*in
   wire signed [14:0] m256_43;
   assign m256_43 =15'b0;

   // m256_44 = W*in
   wire signed [14:0] m256_44;
   assign m256_44 =15'b0;

   // m256_45 = W*in
   wire signed [14:0] m256_45;
   assign m256_45 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_46 = W*in
   wire signed [14:0] m256_46;
   assign m256_46 ={ {3{in256[14]}} , in256[14:3] };

   // m256_47 = W*in
   wire signed [14:0] m256_47;
   assign m256_47 =15'b0;

   // m256_48 = W*in
   wire signed [14:0] m256_48;
   assign m256_48 =15'b0;

   // m256_49 = W*in
   wire signed [14:0] m256_49;
   assign m256_49 =15'b0;

   // m256_50 = W*in
   wire signed [14:0] m256_50;
   assign m256_50 =15'b0;

   // m256_51 = W*in
   wire signed [14:0] m256_51;
   assign m256_51 ={ {3{in256[14]}} , in256[14:3] };

   // m256_52 = W*in
   wire signed [14:0] m256_52;
   assign m256_52 =15'b0;

   // m256_53 = W*in
   wire signed [14:0] m256_53;
   assign m256_53 =15'b0;

   // m256_54 = W*in
   wire signed [14:0] m256_54;
   assign m256_54 =15'b0;

   // m256_55 = W*in
   wire signed [14:0] m256_55;
   assign m256_55 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_56 = W*in
   wire signed [14:0] m256_56;
   assign m256_56 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_57 = W*in
   wire signed [14:0] m256_57;
   assign m256_57 =15'b0;

   // m256_58 = W*in
   wire signed [14:0] m256_58;
   assign m256_58 =15'b0;

   // m256_59 = W*in
   wire signed [14:0] m256_59;
   assign m256_59 =15'b0;

   // m256_60 = W*in
   wire signed [14:0] m256_60;
   assign m256_60 =15'b0;

   // m256_61 = W*in
   wire signed [14:0] m256_61;
   assign m256_61 =15'b0;

   // m256_62 = W*in
   wire signed [14:0] m256_62;
   assign m256_62 =15'b0;

   // m256_63 = W*in
   wire signed [14:0] m256_63;
   assign m256_63 ={ {4{in256[14]}} , in256[14:4] };

   // m256_64 = W*in
   wire signed [14:0] m256_64;
   assign m256_64 =15'b0;

   // m256_65 = W*in
   wire signed [14:0] m256_65;
   assign m256_65 ={ {3{in256[14]}} , in256[14:3] };

   // m256_66 = W*in
   wire signed [14:0] m256_66;
   assign m256_66 =15'b0;

   // m256_67 = W*in
   wire signed [14:0] m256_67;
   assign m256_67 =15'b0;

   // m256_68 = W*in
   wire signed [14:0] m256_68;
   assign m256_68 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_69 = W*in
   wire signed [14:0] m256_69;
   assign m256_69 =15'b0;

   // m256_70 = W*in
   wire signed [14:0] m256_70;
   assign m256_70 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_71 = W*in
   wire signed [14:0] m256_71;
   assign m256_71 =15'b0;

   // m256_72 = W*in
   wire signed [14:0] m256_72;
   assign m256_72 ={ {3{in256[14]}} , in256[14:3] };

   // m256_73 = W*in
   wire signed [14:0] m256_73;
   assign m256_73 =15'b0;

   // m256_74 = W*in
   wire signed [14:0] m256_74;
   assign m256_74 ={ {4{neg256[14]}} , neg256[14:4] };

   // m256_75 = W*in
   wire signed [14:0] m256_75;
   assign m256_75 =15'b0;

   // m256_76 = W*in
   wire signed [14:0] m256_76;
   assign m256_76 =15'b0;

   // m256_77 = W*in
   wire signed [14:0] m256_77;
   assign m256_77 =15'b0;

   // m256_78 = W*in
   wire signed [14:0] m256_78;
   assign m256_78 =15'b0;

   // m256_79 = W*in
   wire signed [14:0] m256_79;
   assign m256_79 ={ {3{in256[14]}} , in256[14:3] };

   // m256_80 = W*in
   wire signed [14:0] m256_80;
   assign m256_80 ={ {3{in256[14]}} , in256[14:3] };

   // m256_81 = W*in
   wire signed [14:0] m256_81;
   assign m256_81 ={ {3{in256[14]}} , in256[14:3] };

   // m256_82 = W*in
   wire signed [14:0] m256_82;
   assign m256_82 =15'b0;

   // m256_83 = W*in
   wire signed [14:0] m256_83;
   assign m256_83 =15'b0;

   // m256_84 = W*in
   wire signed [14:0] m256_84;
   assign m256_84 =15'b0;

   // m256_85 = W*in
   wire signed [14:0] m256_85;
   assign m256_85 =15'b0;

   // m256_86 = W*in
   wire signed [14:0] m256_86;
   assign m256_86 =15'b0;

   // m256_87 = W*in
   wire signed [14:0] m256_87;
   assign m256_87 =15'b0;

   // m256_88 = W*in
   wire signed [14:0] m256_88;
   assign m256_88 =15'b0;

   // m256_89 = W*in
   wire signed [14:0] m256_89;
   assign m256_89 =15'b0;

   // m256_90 = W*in
   wire signed [14:0] m256_90;
   assign m256_90 =15'b0;

   // m256_91 = W*in
   wire signed [14:0] m256_91;
   assign m256_91 =15'b0;

   // m256_92 = W*in
   wire signed [14:0] m256_92;
   assign m256_92 =15'b0;

   // m256_93 = W*in
   wire signed [14:0] m256_93;
   assign m256_93 =15'b0;

   // m256_94 = W*in
   wire signed [14:0] m256_94;
   assign m256_94 =15'b0;

   // m256_95 = W*in
   wire signed [14:0] m256_95;
   assign m256_95 =15'b0;

   // m256_96 = W*in
   wire signed [14:0] m256_96;
   assign m256_96 =15'b0;

   // m256_97 = W*in
   wire signed [14:0] m256_97;
   assign m256_97 =15'b0;

   // m256_98 = W*in
   wire signed [14:0] m256_98;
   assign m256_98 =15'b0;

   // m256_99 = W*in
   wire signed [14:0] m256_99;
   assign m256_99 ={ {3{neg256[14]}} , neg256[14:3] };

   // m256_100 = W*in
   wire signed [14:0] m256_100;
   assign m256_100 =15'b0;

   // m257_1 = W*in
   wire signed [14:0] m257_1;
   assign m257_1 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_2 = W*in
   wire signed [14:0] m257_2;
   assign m257_2 =15'b0;

   // m257_3 = W*in
   wire signed [14:0] m257_3;
   assign m257_3 =15'b0;

   // m257_4 = W*in
   wire signed [14:0] m257_4;
   assign m257_4 =15'b0;

   // m257_5 = W*in
   wire signed [14:0] m257_5;
   assign m257_5 =15'b0;

   // m257_6 = W*in
   wire signed [14:0] m257_6;
   assign m257_6 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_7 = W*in
   wire signed [14:0] m257_7;
   assign m257_7 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_8 = W*in
   wire signed [14:0] m257_8;
   assign m257_8 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_9 = W*in
   wire signed [14:0] m257_9;
   assign m257_9 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_10 = W*in
   wire signed [14:0] m257_10;
   assign m257_10 =15'b0;

   // m257_11 = W*in
   wire signed [14:0] m257_11;
   assign m257_11 =15'b0;

   // m257_12 = W*in
   wire signed [14:0] m257_12;
   assign m257_12 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_13 = W*in
   wire signed [14:0] m257_13;
   assign m257_13 =15'b0;

   // m257_14 = W*in
   wire signed [14:0] m257_14;
   assign m257_14 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_15 = W*in
   wire signed [14:0] m257_15;
   assign m257_15 ={ {3{in257[14]}} , in257[14:3] };

   // m257_16 = W*in
   wire signed [14:0] m257_16;
   assign m257_16 =15'b0;

   // m257_17 = W*in
   wire signed [14:0] m257_17;
   assign m257_17 ={ {3{in257[14]}} , in257[14:3] };

   // m257_18 = W*in
   wire signed [14:0] m257_18;
   assign m257_18 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_19 = W*in
   wire signed [14:0] m257_19;
   assign m257_19 ={ {4{in257[14]}} , in257[14:4] };

   // m257_20 = W*in
   wire signed [14:0] m257_20;
   assign m257_20 =15'b0;

   // m257_21 = W*in
   wire signed [14:0] m257_21;
   assign m257_21 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_22 = W*in
   wire signed [14:0] m257_22;
   assign m257_22 =15'b0;

   // m257_23 = W*in
   wire signed [14:0] m257_23;
   assign m257_23 =15'b0;

   // m257_24 = W*in
   wire signed [14:0] m257_24;
   assign m257_24 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_25 = W*in
   wire signed [14:0] m257_25;
   assign m257_25 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_26 = W*in
   wire signed [14:0] m257_26;
   assign m257_26 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_27 = W*in
   wire signed [14:0] m257_27;
   assign m257_27 ={ {4{in257[14]}} , in257[14:4] };

   // m257_28 = W*in
   wire signed [14:0] m257_28;
   assign m257_28 =15'b0;

   // m257_29 = W*in
   wire signed [14:0] m257_29;
   assign m257_29 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_30 = W*in
   wire signed [14:0] m257_30;
   assign m257_30 =15'b0;

   // m257_31 = W*in
   wire signed [14:0] m257_31;
   assign m257_31 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_32 = W*in
   wire signed [14:0] m257_32;
   assign m257_32 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_33 = W*in
   wire signed [14:0] m257_33;
   assign m257_33 =15'b0;

   // m257_34 = W*in
   wire signed [14:0] m257_34;
   assign m257_34 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_35 = W*in
   wire signed [14:0] m257_35;
   assign m257_35 =15'b0;

   // m257_36 = W*in
   wire signed [14:0] m257_36;
   assign m257_36 =15'b0;

   // m257_37 = W*in
   wire signed [14:0] m257_37;
   assign m257_37 =15'b0;

   // m257_38 = W*in
   wire signed [14:0] m257_38;
   assign m257_38 =15'b0;

   // m257_39 = W*in
   wire signed [14:0] m257_39;
   assign m257_39 =15'b0;

   // m257_40 = W*in
   wire signed [14:0] m257_40;
   assign m257_40 =15'b0;

   // m257_41 = W*in
   wire signed [14:0] m257_41;
   assign m257_41 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_42 = W*in
   wire signed [14:0] m257_42;
   assign m257_42 =15'b0;

   // m257_43 = W*in
   wire signed [14:0] m257_43;
   assign m257_43 =15'b0;

   // m257_44 = W*in
   wire signed [14:0] m257_44;
   assign m257_44 =15'b0;

   // m257_45 = W*in
   wire signed [14:0] m257_45;
   assign m257_45 =15'b0;

   // m257_46 = W*in
   wire signed [14:0] m257_46;
   assign m257_46 ={ {4{in257[14]}} , in257[14:4] };

   // m257_47 = W*in
   wire signed [14:0] m257_47;
   assign m257_47 =15'b0;

   // m257_48 = W*in
   wire signed [14:0] m257_48;
   assign m257_48 =15'b0;

   // m257_49 = W*in
   wire signed [14:0] m257_49;
   assign m257_49 ={ {3{in257[14]}} , in257[14:3] };

   // m257_50 = W*in
   wire signed [14:0] m257_50;
   assign m257_50 =15'b0;

   // m257_51 = W*in
   wire signed [14:0] m257_51;
   assign m257_51 =15'b0;

   // m257_52 = W*in
   wire signed [14:0] m257_52;
   assign m257_52 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_53 = W*in
   wire signed [14:0] m257_53;
   assign m257_53 =15'b0;

   // m257_54 = W*in
   wire signed [14:0] m257_54;
   assign m257_54 =15'b0;

   // m257_55 = W*in
   wire signed [14:0] m257_55;
   assign m257_55 =15'b0;

   // m257_56 = W*in
   wire signed [14:0] m257_56;
   assign m257_56 ={ {3{in257[14]}} , in257[14:3] };

   // m257_57 = W*in
   wire signed [14:0] m257_57;
   assign m257_57 =15'b0;

   // m257_58 = W*in
   wire signed [14:0] m257_58;
   assign m257_58 ={ {4{in257[14]}} , in257[14:4] };

   // m257_59 = W*in
   wire signed [14:0] m257_59;
   assign m257_59 ={ {4{in257[14]}} , in257[14:4] };

   // m257_60 = W*in
   wire signed [14:0] m257_60;
   assign m257_60 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_61 = W*in
   wire signed [14:0] m257_61;
   assign m257_61 ={ {4{in257[14]}} , in257[14:4] };

   // m257_62 = W*in
   wire signed [14:0] m257_62;
   assign m257_62 =15'b0;

   // m257_63 = W*in
   wire signed [14:0] m257_63;
   assign m257_63 =15'b0;

   // m257_64 = W*in
   wire signed [14:0] m257_64;
   assign m257_64 ={ {4{in257[14]}} , in257[14:4] };

   // m257_65 = W*in
   wire signed [14:0] m257_65;
   assign m257_65 =15'b0;

   // m257_66 = W*in
   wire signed [14:0] m257_66;
   assign m257_66 =15'b0;

   // m257_67 = W*in
   wire signed [14:0] m257_67;
   assign m257_67 ={ {3{in257[14]}} , in257[14:3] };

   // m257_68 = W*in
   wire signed [14:0] m257_68;
   assign m257_68 =15'b0;

   // m257_69 = W*in
   wire signed [14:0] m257_69;
   assign m257_69 ={ {3{in257[14]}} , in257[14:3] };

   // m257_70 = W*in
   wire signed [14:0] m257_70;
   assign m257_70 =15'b0;

   // m257_71 = W*in
   wire signed [14:0] m257_71;
   assign m257_71 =15'b0;

   // m257_72 = W*in
   wire signed [14:0] m257_72;
   assign m257_72 =15'b0;

   // m257_73 = W*in
   wire signed [14:0] m257_73;
   assign m257_73 =15'b0;

   // m257_74 = W*in
   wire signed [14:0] m257_74;
   assign m257_74 =15'b0;

   // m257_75 = W*in
   wire signed [14:0] m257_75;
   assign m257_75 =15'b0;

   // m257_76 = W*in
   wire signed [14:0] m257_76;
   assign m257_76 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_77 = W*in
   wire signed [14:0] m257_77;
   assign m257_77 =15'b0;

   // m257_78 = W*in
   wire signed [14:0] m257_78;
   assign m257_78 ={ {4{neg257[14]}} , neg257[14:4] };

   // m257_79 = W*in
   wire signed [14:0] m257_79;
   assign m257_79 =15'b0;

   // m257_80 = W*in
   wire signed [14:0] m257_80;
   assign m257_80 =15'b0;

   // m257_81 = W*in
   wire signed [14:0] m257_81;
   assign m257_81 =15'b0;

   // m257_82 = W*in
   wire signed [14:0] m257_82;
   assign m257_82 =15'b0;

   // m257_83 = W*in
   wire signed [14:0] m257_83;
   assign m257_83 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_84 = W*in
   wire signed [14:0] m257_84;
   assign m257_84 =15'b0;

   // m257_85 = W*in
   wire signed [14:0] m257_85;
   assign m257_85 =15'b0;

   // m257_86 = W*in
   wire signed [14:0] m257_86;
   assign m257_86 ={ {3{in257[14]}} , in257[14:3] };

   // m257_87 = W*in
   wire signed [14:0] m257_87;
   assign m257_87 =15'b0;

   // m257_88 = W*in
   wire signed [14:0] m257_88;
   assign m257_88 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_89 = W*in
   wire signed [14:0] m257_89;
   assign m257_89 =15'b0;

   // m257_90 = W*in
   wire signed [14:0] m257_90;
   assign m257_90 =15'b0;

   // m257_91 = W*in
   wire signed [14:0] m257_91;
   assign m257_91 =15'b0;

   // m257_92 = W*in
   wire signed [14:0] m257_92;
   assign m257_92 =15'b0;

   // m257_93 = W*in
   wire signed [14:0] m257_93;
   assign m257_93 =15'b0;

   // m257_94 = W*in
   wire signed [14:0] m257_94;
   assign m257_94 =15'b0;

   // m257_95 = W*in
   wire signed [14:0] m257_95;
   assign m257_95 =15'b0;

   // m257_96 = W*in
   wire signed [14:0] m257_96;
   assign m257_96 ={ {3{neg257[14]}} , neg257[14:3] };

   // m257_97 = W*in
   wire signed [14:0] m257_97;
   assign m257_97 =15'b0;

   // m257_98 = W*in
   wire signed [14:0] m257_98;
   assign m257_98 =15'b0;

   // m257_99 = W*in
   wire signed [14:0] m257_99;
   assign m257_99 =15'b0;

   // m257_100 = W*in
   wire signed [14:0] m257_100;
   assign m257_100 =15'b0;

   // m258_1 = W*in
   wire signed [14:0] m258_1;
   assign m258_1 =15'b0;

   // m258_2 = W*in
   wire signed [14:0] m258_2;
   assign m258_2 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_3 = W*in
   wire signed [14:0] m258_3;
   assign m258_3 =15'b0;

   // m258_4 = W*in
   wire signed [14:0] m258_4;
   assign m258_4 =15'b0;

   // m258_5 = W*in
   wire signed [14:0] m258_5;
   assign m258_5 ={ {2{neg258[14]}} , neg258[14:2] };

   // m258_6 = W*in
   wire signed [14:0] m258_6;
   assign m258_6 =15'b0;

   // m258_7 = W*in
   wire signed [14:0] m258_7;
   assign m258_7 =15'b0;

   // m258_8 = W*in
   wire signed [14:0] m258_8;
   assign m258_8 =15'b0;

   // m258_9 = W*in
   wire signed [14:0] m258_9;
   assign m258_9 =15'b0;

   // m258_10 = W*in
   wire signed [14:0] m258_10;
   assign m258_10 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_11 = W*in
   wire signed [14:0] m258_11;
   assign m258_11 =15'b0;

   // m258_12 = W*in
   wire signed [14:0] m258_12;
   assign m258_12 =15'b0;

   // m258_13 = W*in
   wire signed [14:0] m258_13;
   assign m258_13 =15'b0;

   // m258_14 = W*in
   wire signed [14:0] m258_14;
   assign m258_14 =15'b0;

   // m258_15 = W*in
   wire signed [14:0] m258_15;
   assign m258_15 =15'b0;

   // m258_16 = W*in
   wire signed [14:0] m258_16;
   assign m258_16 ={ {2{neg258[14]}} , neg258[14:2] };

   // m258_17 = W*in
   wire signed [14:0] m258_17;
   assign m258_17 ={ {3{in258[14]}} , in258[14:3] };

   // m258_18 = W*in
   wire signed [14:0] m258_18;
   assign m258_18 =15'b0;

   // m258_19 = W*in
   wire signed [14:0] m258_19;
   assign m258_19 =15'b0;

   // m258_20 = W*in
   wire signed [14:0] m258_20;
   assign m258_20 =15'b0;

   // m258_21 = W*in
   wire signed [14:0] m258_21;
   assign m258_21 =15'b0;

   // m258_22 = W*in
   wire signed [14:0] m258_22;
   assign m258_22 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_23 = W*in
   wire signed [14:0] m258_23;
   assign m258_23 ={ {3{in258[14]}} , in258[14:3] };

   // m258_24 = W*in
   wire signed [14:0] m258_24;
   assign m258_24 =15'b0;

   // m258_25 = W*in
   wire signed [14:0] m258_25;
   assign m258_25 =15'b0;

   // m258_26 = W*in
   wire signed [14:0] m258_26;
   assign m258_26 =15'b0;

   // m258_27 = W*in
   wire signed [14:0] m258_27;
   assign m258_27 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_28 = W*in
   wire signed [14:0] m258_28;
   assign m258_28 =15'b0;

   // m258_29 = W*in
   wire signed [14:0] m258_29;
   assign m258_29 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_30 = W*in
   wire signed [14:0] m258_30;
   assign m258_30 =15'b0;

   // m258_31 = W*in
   wire signed [14:0] m258_31;
   assign m258_31 ={ {4{neg258[14]}} , neg258[14:4] };

   // m258_32 = W*in
   wire signed [14:0] m258_32;
   assign m258_32 =15'b0;

   // m258_33 = W*in
   wire signed [14:0] m258_33;
   assign m258_33 =15'b0;

   // m258_34 = W*in
   wire signed [14:0] m258_34;
   assign m258_34 =15'b0;

   // m258_35 = W*in
   wire signed [14:0] m258_35;
   assign m258_35 =15'b0;

   // m258_36 = W*in
   wire signed [14:0] m258_36;
   assign m258_36 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_37 = W*in
   wire signed [14:0] m258_37;
   assign m258_37 =15'b0;

   // m258_38 = W*in
   wire signed [14:0] m258_38;
   assign m258_38 =15'b0;

   // m258_39 = W*in
   wire signed [14:0] m258_39;
   assign m258_39 =15'b0;

   // m258_40 = W*in
   wire signed [14:0] m258_40;
   assign m258_40 =15'b0;

   // m258_41 = W*in
   wire signed [14:0] m258_41;
   assign m258_41 ={ {3{in258[14]}} , in258[14:3] };

   // m258_42 = W*in
   wire signed [14:0] m258_42;
   assign m258_42 =15'b0;

   // m258_43 = W*in
   wire signed [14:0] m258_43;
   assign m258_43 =15'b0;

   // m258_44 = W*in
   wire signed [14:0] m258_44;
   assign m258_44 =15'b0;

   // m258_45 = W*in
   wire signed [14:0] m258_45;
   assign m258_45 =15'b0;

   // m258_46 = W*in
   wire signed [14:0] m258_46;
   assign m258_46 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_47 = W*in
   wire signed [14:0] m258_47;
   assign m258_47 =15'b0;

   // m258_48 = W*in
   wire signed [14:0] m258_48;
   assign m258_48 =15'b0;

   // m258_49 = W*in
   wire signed [14:0] m258_49;
   assign m258_49 ={ {3{in258[14]}} , in258[14:3] };

   // m258_50 = W*in
   wire signed [14:0] m258_50;
   assign m258_50 =15'b0;

   // m258_51 = W*in
   wire signed [14:0] m258_51;
   assign m258_51 =15'b0;

   // m258_52 = W*in
   wire signed [14:0] m258_52;
   assign m258_52 ={ {3{in258[14]}} , in258[14:3] };

   // m258_53 = W*in
   wire signed [14:0] m258_53;
   assign m258_53 =15'b0;

   // m258_54 = W*in
   wire signed [14:0] m258_54;
   assign m258_54 =15'b0;

   // m258_55 = W*in
   wire signed [14:0] m258_55;
   assign m258_55 =15'b0;

   // m258_56 = W*in
   wire signed [14:0] m258_56;
   assign m258_56 =15'b0;

   // m258_57 = W*in
   wire signed [14:0] m258_57;
   assign m258_57 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_58 = W*in
   wire signed [14:0] m258_58;
   assign m258_58 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_59 = W*in
   wire signed [14:0] m258_59;
   assign m258_59 =15'b0;

   // m258_60 = W*in
   wire signed [14:0] m258_60;
   assign m258_60 =15'b0;

   // m258_61 = W*in
   wire signed [14:0] m258_61;
   assign m258_61 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_62 = W*in
   wire signed [14:0] m258_62;
   assign m258_62 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_63 = W*in
   wire signed [14:0] m258_63;
   assign m258_63 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_64 = W*in
   wire signed [14:0] m258_64;
   assign m258_64 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_65 = W*in
   wire signed [14:0] m258_65;
   assign m258_65 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_66 = W*in
   wire signed [14:0] m258_66;
   assign m258_66 =15'b0;

   // m258_67 = W*in
   wire signed [14:0] m258_67;
   assign m258_67 =15'b0;

   // m258_68 = W*in
   wire signed [14:0] m258_68;
   assign m258_68 ={ {4{neg258[14]}} , neg258[14:4] };

   // m258_69 = W*in
   wire signed [14:0] m258_69;
   assign m258_69 =15'b0;

   // m258_70 = W*in
   wire signed [14:0] m258_70;
   assign m258_70 ={ {2{in258[14]}} , in258[14:2] };

   // m258_71 = W*in
   wire signed [14:0] m258_71;
   assign m258_71 ={ {3{in258[14]}} , in258[14:3] };

   // m258_72 = W*in
   wire signed [14:0] m258_72;
   assign m258_72 =15'b0;

   // m258_73 = W*in
   wire signed [14:0] m258_73;
   assign m258_73 =15'b0;

   // m258_74 = W*in
   wire signed [14:0] m258_74;
   assign m258_74 =15'b0;

   // m258_75 = W*in
   wire signed [14:0] m258_75;
   assign m258_75 =15'b0;

   // m258_76 = W*in
   wire signed [14:0] m258_76;
   assign m258_76 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_77 = W*in
   wire signed [14:0] m258_77;
   assign m258_77 =15'b0;

   // m258_78 = W*in
   wire signed [14:0] m258_78;
   assign m258_78 =15'b0;

   // m258_79 = W*in
   wire signed [14:0] m258_79;
   assign m258_79 =15'b0;

   // m258_80 = W*in
   wire signed [14:0] m258_80;
   assign m258_80 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_81 = W*in
   wire signed [14:0] m258_81;
   assign m258_81 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_82 = W*in
   wire signed [14:0] m258_82;
   assign m258_82 ={ {2{neg258[14]}} , neg258[14:2] };

   // m258_83 = W*in
   wire signed [14:0] m258_83;
   assign m258_83 =15'b0;

   // m258_84 = W*in
   wire signed [14:0] m258_84;
   assign m258_84 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_85 = W*in
   wire signed [14:0] m258_85;
   assign m258_85 =15'b0;

   // m258_86 = W*in
   wire signed [14:0] m258_86;
   assign m258_86 =15'b0;

   // m258_87 = W*in
   wire signed [14:0] m258_87;
   assign m258_87 =15'b0;

   // m258_88 = W*in
   wire signed [14:0] m258_88;
   assign m258_88 =15'b0;

   // m258_89 = W*in
   wire signed [14:0] m258_89;
   assign m258_89 ={ {3{in258[14]}} , in258[14:3] };

   // m258_90 = W*in
   wire signed [14:0] m258_90;
   assign m258_90 =15'b0;

   // m258_91 = W*in
   wire signed [14:0] m258_91;
   assign m258_91 =15'b0;

   // m258_92 = W*in
   wire signed [14:0] m258_92;
   assign m258_92 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_93 = W*in
   wire signed [14:0] m258_93;
   assign m258_93 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_94 = W*in
   wire signed [14:0] m258_94;
   assign m258_94 =15'b0;

   // m258_95 = W*in
   wire signed [14:0] m258_95;
   assign m258_95 ={ {3{in258[14]}} , in258[14:3] };

   // m258_96 = W*in
   wire signed [14:0] m258_96;
   assign m258_96 ={ {3{in258[14]}} , in258[14:3] };

   // m258_97 = W*in
   wire signed [14:0] m258_97;
   assign m258_97 ={ {3{neg258[14]}} , neg258[14:3] };

   // m258_98 = W*in
   wire signed [14:0] m258_98;
   assign m258_98 ={ {3{in258[14]}} , in258[14:3] };

   // m258_99 = W*in
   wire signed [14:0] m258_99;
   assign m258_99 =15'b0;

   // m258_100 = W*in
   wire signed [14:0] m258_100;
   assign m258_100 =15'b0;

   // m259_1 = W*in
   wire signed [14:0] m259_1;
   assign m259_1 =15'b0;

   // m259_2 = W*in
   wire signed [14:0] m259_2;
   assign m259_2 =15'b0;

   // m259_3 = W*in
   wire signed [14:0] m259_3;
   assign m259_3 =15'b0;

   // m259_4 = W*in
   wire signed [14:0] m259_4;
   assign m259_4 =15'b0;

   // m259_5 = W*in
   wire signed [14:0] m259_5;
   assign m259_5 =15'b0;

   // m259_6 = W*in
   wire signed [14:0] m259_6;
   assign m259_6 =15'b0;

   // m259_7 = W*in
   wire signed [14:0] m259_7;
   assign m259_7 =15'b0;

   // m259_8 = W*in
   wire signed [14:0] m259_8;
   assign m259_8 =15'b0;

   // m259_9 = W*in
   wire signed [14:0] m259_9;
   assign m259_9 =15'b0;

   // m259_10 = W*in
   wire signed [14:0] m259_10;
   assign m259_10 ={ {3{in259[14]}} , in259[14:3] };

   // m259_11 = W*in
   wire signed [14:0] m259_11;
   assign m259_11 =15'b0;

   // m259_12 = W*in
   wire signed [14:0] m259_12;
   assign m259_12 =15'b0;

   // m259_13 = W*in
   wire signed [14:0] m259_13;
   assign m259_13 =15'b0;

   // m259_14 = W*in
   wire signed [14:0] m259_14;
   assign m259_14 =15'b0;

   // m259_15 = W*in
   wire signed [14:0] m259_15;
   assign m259_15 =15'b0;

   // m259_16 = W*in
   wire signed [14:0] m259_16;
   assign m259_16 =15'b0;

   // m259_17 = W*in
   wire signed [14:0] m259_17;
   assign m259_17 ={ {3{neg259[14]}} , neg259[14:3] };

   // m259_18 = W*in
   wire signed [14:0] m259_18;
   assign m259_18 =15'b0;

   // m259_19 = W*in
   wire signed [14:0] m259_19;
   assign m259_19 =15'b0;

   // m259_20 = W*in
   wire signed [14:0] m259_20;
   assign m259_20 =15'b0;

   // m259_21 = W*in
   wire signed [14:0] m259_21;
   assign m259_21 =15'b0;

   // m259_22 = W*in
   wire signed [14:0] m259_22;
   assign m259_22 =15'b0;

   // m259_23 = W*in
   wire signed [14:0] m259_23;
   assign m259_23 =15'b0;

   // m259_24 = W*in
   wire signed [14:0] m259_24;
   assign m259_24 =15'b0;

   // m259_25 = W*in
   wire signed [14:0] m259_25;
   assign m259_25 =15'b0;

   // m259_26 = W*in
   wire signed [14:0] m259_26;
   assign m259_26 =15'b0;

   // m259_27 = W*in
   wire signed [14:0] m259_27;
   assign m259_27 ={ {4{neg259[14]}} , neg259[14:4] };

   // m259_28 = W*in
   wire signed [14:0] m259_28;
   assign m259_28 =15'b0;

   // m259_29 = W*in
   wire signed [14:0] m259_29;
   assign m259_29 =15'b0;

   // m259_30 = W*in
   wire signed [14:0] m259_30;
   assign m259_30 =15'b0;

   // m259_31 = W*in
   wire signed [14:0] m259_31;
   assign m259_31 =15'b0;

   // m259_32 = W*in
   wire signed [14:0] m259_32;
   assign m259_32 =15'b0;

   // m259_33 = W*in
   wire signed [14:0] m259_33;
   assign m259_33 =15'b0;

   // m259_34 = W*in
   wire signed [14:0] m259_34;
   assign m259_34 =15'b0;

   // m259_35 = W*in
   wire signed [14:0] m259_35;
   assign m259_35 =15'b0;

   // m259_36 = W*in
   wire signed [14:0] m259_36;
   assign m259_36 =15'b0;

   // m259_37 = W*in
   wire signed [14:0] m259_37;
   assign m259_37 ={ {2{in259[14]}} , in259[14:2] };

   // m259_38 = W*in
   wire signed [14:0] m259_38;
   assign m259_38 =15'b0;

   // m259_39 = W*in
   wire signed [14:0] m259_39;
   assign m259_39 =15'b0;

   // m259_40 = W*in
   wire signed [14:0] m259_40;
   assign m259_40 =15'b0;

   // m259_41 = W*in
   wire signed [14:0] m259_41;
   assign m259_41 =15'b0;

   // m259_42 = W*in
   wire signed [14:0] m259_42;
   assign m259_42 =15'b0;

   // m259_43 = W*in
   wire signed [14:0] m259_43;
   assign m259_43 =15'b0;

   // m259_44 = W*in
   wire signed [14:0] m259_44;
   assign m259_44 =15'b0;

   // m259_45 = W*in
   wire signed [14:0] m259_45;
   assign m259_45 =15'b0;

   // m259_46 = W*in
   wire signed [14:0] m259_46;
   assign m259_46 =15'b0;

   // m259_47 = W*in
   wire signed [14:0] m259_47;
   assign m259_47 =15'b0;

   // m259_48 = W*in
   wire signed [14:0] m259_48;
   assign m259_48 =15'b0;

   // m259_49 = W*in
   wire signed [14:0] m259_49;
   assign m259_49 =15'b0;

   // m259_50 = W*in
   wire signed [14:0] m259_50;
   assign m259_50 =15'b0;

   // m259_51 = W*in
   wire signed [14:0] m259_51;
   assign m259_51 =15'b0;

   // m259_52 = W*in
   wire signed [14:0] m259_52;
   assign m259_52 =15'b0;

   // m259_53 = W*in
   wire signed [14:0] m259_53;
   assign m259_53 =15'b0;

   // m259_54 = W*in
   wire signed [14:0] m259_54;
   assign m259_54 =15'b0;

   // m259_55 = W*in
   wire signed [14:0] m259_55;
   assign m259_55 =15'b0;

   // m259_56 = W*in
   wire signed [14:0] m259_56;
   assign m259_56 =15'b0;

   // m259_57 = W*in
   wire signed [14:0] m259_57;
   assign m259_57 =15'b0;

   // m259_58 = W*in
   wire signed [14:0] m259_58;
   assign m259_58 =15'b0;

   // m259_59 = W*in
   wire signed [14:0] m259_59;
   assign m259_59 =15'b0;

   // m259_60 = W*in
   wire signed [14:0] m259_60;
   assign m259_60 =15'b0;

   // m259_61 = W*in
   wire signed [14:0] m259_61;
   assign m259_61 =15'b0;

   // m259_62 = W*in
   wire signed [14:0] m259_62;
   assign m259_62 =15'b0;

   // m259_63 = W*in
   wire signed [14:0] m259_63;
   assign m259_63 ={ {3{in259[14]}} , in259[14:3] };

   // m259_64 = W*in
   wire signed [14:0] m259_64;
   assign m259_64 =15'b0;

   // m259_65 = W*in
   wire signed [14:0] m259_65;
   assign m259_65 =15'b0;

   // m259_66 = W*in
   wire signed [14:0] m259_66;
   assign m259_66 =15'b0;

   // m259_67 = W*in
   wire signed [14:0] m259_67;
   assign m259_67 =15'b0;

   // m259_68 = W*in
   wire signed [14:0] m259_68;
   assign m259_68 =15'b0;

   // m259_69 = W*in
   wire signed [14:0] m259_69;
   assign m259_69 =15'b0;

   // m259_70 = W*in
   wire signed [14:0] m259_70;
   assign m259_70 =15'b0;

   // m259_71 = W*in
   wire signed [14:0] m259_71;
   assign m259_71 =15'b0;

   // m259_72 = W*in
   wire signed [14:0] m259_72;
   assign m259_72 =15'b0;

   // m259_73 = W*in
   wire signed [14:0] m259_73;
   assign m259_73 =15'b0;

   // m259_74 = W*in
   wire signed [14:0] m259_74;
   assign m259_74 =15'b0;

   // m259_75 = W*in
   wire signed [14:0] m259_75;
   assign m259_75 ={ {3{neg259[14]}} , neg259[14:3] };

   // m259_76 = W*in
   wire signed [14:0] m259_76;
   assign m259_76 =15'b0;

   // m259_77 = W*in
   wire signed [14:0] m259_77;
   assign m259_77 =15'b0;

   // m259_78 = W*in
   wire signed [14:0] m259_78;
   assign m259_78 =15'b0;

   // m259_79 = W*in
   wire signed [14:0] m259_79;
   assign m259_79 =15'b0;

   // m259_80 = W*in
   wire signed [14:0] m259_80;
   assign m259_80 =15'b0;

   // m259_81 = W*in
   wire signed [14:0] m259_81;
   assign m259_81 =15'b0;

   // m259_82 = W*in
   wire signed [14:0] m259_82;
   assign m259_82 =15'b0;

   // m259_83 = W*in
   wire signed [14:0] m259_83;
   assign m259_83 =15'b0;

   // m259_84 = W*in
   wire signed [14:0] m259_84;
   assign m259_84 =15'b0;

   // m259_85 = W*in
   wire signed [14:0] m259_85;
   assign m259_85 =15'b0;

   // m259_86 = W*in
   wire signed [14:0] m259_86;
   assign m259_86 =15'b0;

   // m259_87 = W*in
   wire signed [14:0] m259_87;
   assign m259_87 =15'b0;

   // m259_88 = W*in
   wire signed [14:0] m259_88;
   assign m259_88 =15'b0;

   // m259_89 = W*in
   wire signed [14:0] m259_89;
   assign m259_89 =15'b0;

   // m259_90 = W*in
   wire signed [14:0] m259_90;
   assign m259_90 =15'b0;

   // m259_91 = W*in
   wire signed [14:0] m259_91;
   assign m259_91 ={ {3{in259[14]}} , in259[14:3] };

   // m259_92 = W*in
   wire signed [14:0] m259_92;
   assign m259_92 =15'b0;

   // m259_93 = W*in
   wire signed [14:0] m259_93;
   assign m259_93 =15'b0;

   // m259_94 = W*in
   wire signed [14:0] m259_94;
   assign m259_94 =15'b0;

   // m259_95 = W*in
   wire signed [14:0] m259_95;
   assign m259_95 =15'b0;

   // m259_96 = W*in
   wire signed [14:0] m259_96;
   assign m259_96 =15'b0;

   // m259_97 = W*in
   wire signed [14:0] m259_97;
   assign m259_97 =15'b0;

   // m259_98 = W*in
   wire signed [14:0] m259_98;
   assign m259_98 =15'b0;

   // m259_99 = W*in
   wire signed [14:0] m259_99;
   assign m259_99 =15'b0;

   // m259_100 = W*in
   wire signed [14:0] m259_100;
   assign m259_100 =15'b0;

   // m260_1 = W*in
   wire signed [14:0] m260_1;
   assign m260_1 ={ {4{neg260[14]}} , neg260[14:4] };

   // m260_2 = W*in
   wire signed [14:0] m260_2;
   assign m260_2 =15'b0;

   // m260_3 = W*in
   wire signed [14:0] m260_3;
   assign m260_3 =15'b0;

   // m260_4 = W*in
   wire signed [14:0] m260_4;
   assign m260_4 ={ {4{in260[14]}} , in260[14:4] };

   // m260_5 = W*in
   wire signed [14:0] m260_5;
   assign m260_5 =15'b0;

   // m260_6 = W*in
   wire signed [14:0] m260_6;
   assign m260_6 =15'b0;

   // m260_7 = W*in
   wire signed [14:0] m260_7;
   assign m260_7 =15'b0;

   // m260_8 = W*in
   wire signed [14:0] m260_8;
   assign m260_8 =15'b0;

   // m260_9 = W*in
   wire signed [14:0] m260_9;
   assign m260_9 =15'b0;

   // m260_10 = W*in
   wire signed [14:0] m260_10;
   assign m260_10 ={ {3{neg260[14]}} , neg260[14:3] };

   // m260_11 = W*in
   wire signed [14:0] m260_11;
   assign m260_11 =15'b0;

   // m260_12 = W*in
   wire signed [14:0] m260_12;
   assign m260_12 =15'b0;

   // m260_13 = W*in
   wire signed [14:0] m260_13;
   assign m260_13 =15'b0;

   // m260_14 = W*in
   wire signed [14:0] m260_14;
   assign m260_14 =15'b0;

   // m260_15 = W*in
   wire signed [14:0] m260_15;
   assign m260_15 =15'b0;

   // m260_16 = W*in
   wire signed [14:0] m260_16;
   assign m260_16 =15'b0;

   // m260_17 = W*in
   wire signed [14:0] m260_17;
   assign m260_17 =15'b0;

   // m260_18 = W*in
   wire signed [14:0] m260_18;
   assign m260_18 =15'b0;

   // m260_19 = W*in
   wire signed [14:0] m260_19;
   assign m260_19 =15'b0;

   // m260_20 = W*in
   wire signed [14:0] m260_20;
   assign m260_20 =15'b0;

   // m260_21 = W*in
   wire signed [14:0] m260_21;
   assign m260_21 =15'b0;

   // m260_22 = W*in
   wire signed [14:0] m260_22;
   assign m260_22 =15'b0;

   // m260_23 = W*in
   wire signed [14:0] m260_23;
   assign m260_23 =15'b0;

   // m260_24 = W*in
   wire signed [14:0] m260_24;
   assign m260_24 =15'b0;

   // m260_25 = W*in
   wire signed [14:0] m260_25;
   assign m260_25 =15'b0;

   // m260_26 = W*in
   wire signed [14:0] m260_26;
   assign m260_26 =15'b0;

   // m260_27 = W*in
   wire signed [14:0] m260_27;
   assign m260_27 =15'b0;

   // m260_28 = W*in
   wire signed [14:0] m260_28;
   assign m260_28 =15'b0;

   // m260_29 = W*in
   wire signed [14:0] m260_29;
   assign m260_29 =15'b0;

   // m260_30 = W*in
   wire signed [14:0] m260_30;
   assign m260_30 =15'b0;

   // m260_31 = W*in
   wire signed [14:0] m260_31;
   assign m260_31 =15'b0;

   // m260_32 = W*in
   wire signed [14:0] m260_32;
   assign m260_32 ={ {4{neg260[14]}} , neg260[14:4] };

   // m260_33 = W*in
   wire signed [14:0] m260_33;
   assign m260_33 =15'b0;

   // m260_34 = W*in
   wire signed [14:0] m260_34;
   assign m260_34 =15'b0;

   // m260_35 = W*in
   wire signed [14:0] m260_35;
   assign m260_35 =15'b0;

   // m260_36 = W*in
   wire signed [14:0] m260_36;
   assign m260_36 =15'b0;

   // m260_37 = W*in
   wire signed [14:0] m260_37;
   assign m260_37 =15'b0;

   // m260_38 = W*in
   wire signed [14:0] m260_38;
   assign m260_38 =15'b0;

   // m260_39 = W*in
   wire signed [14:0] m260_39;
   assign m260_39 =15'b0;

   // m260_40 = W*in
   wire signed [14:0] m260_40;
   assign m260_40 =15'b0;

   // m260_41 = W*in
   wire signed [14:0] m260_41;
   assign m260_41 =15'b0;

   // m260_42 = W*in
   wire signed [14:0] m260_42;
   assign m260_42 =15'b0;

   // m260_43 = W*in
   wire signed [14:0] m260_43;
   assign m260_43 =15'b0;

   // m260_44 = W*in
   wire signed [14:0] m260_44;
   assign m260_44 ={ {2{in260[14]}} , in260[14:2] };

   // m260_45 = W*in
   wire signed [14:0] m260_45;
   assign m260_45 =15'b0;

   // m260_46 = W*in
   wire signed [14:0] m260_46;
   assign m260_46 =15'b0;

   // m260_47 = W*in
   wire signed [14:0] m260_47;
   assign m260_47 =15'b0;

   // m260_48 = W*in
   wire signed [14:0] m260_48;
   assign m260_48 =15'b0;

   // m260_49 = W*in
   wire signed [14:0] m260_49;
   assign m260_49 =15'b0;

   // m260_50 = W*in
   wire signed [14:0] m260_50;
   assign m260_50 =15'b0;

   // m260_51 = W*in
   wire signed [14:0] m260_51;
   assign m260_51 =15'b0;

   // m260_52 = W*in
   wire signed [14:0] m260_52;
   assign m260_52 =15'b0;

   // m260_53 = W*in
   wire signed [14:0] m260_53;
   assign m260_53 =15'b0;

   // m260_54 = W*in
   wire signed [14:0] m260_54;
   assign m260_54 =15'b0;

   // m260_55 = W*in
   wire signed [14:0] m260_55;
   assign m260_55 =15'b0;

   // m260_56 = W*in
   wire signed [14:0] m260_56;
   assign m260_56 ={ {4{neg260[14]}} , neg260[14:4] };

   // m260_57 = W*in
   wire signed [14:0] m260_57;
   assign m260_57 =15'b0;

   // m260_58 = W*in
   wire signed [14:0] m260_58;
   assign m260_58 =15'b0;

   // m260_59 = W*in
   wire signed [14:0] m260_59;
   assign m260_59 =15'b0;

   // m260_60 = W*in
   wire signed [14:0] m260_60;
   assign m260_60 =15'b0;

   // m260_61 = W*in
   wire signed [14:0] m260_61;
   assign m260_61 =15'b0;

   // m260_62 = W*in
   wire signed [14:0] m260_62;
   assign m260_62 =15'b0;

   // m260_63 = W*in
   wire signed [14:0] m260_63;
   assign m260_63 =15'b0;

   // m260_64 = W*in
   wire signed [14:0] m260_64;
   assign m260_64 =15'b0;

   // m260_65 = W*in
   wire signed [14:0] m260_65;
   assign m260_65 =15'b0;

   // m260_66 = W*in
   wire signed [14:0] m260_66;
   assign m260_66 =15'b0;

   // m260_67 = W*in
   wire signed [14:0] m260_67;
   assign m260_67 =15'b0;

   // m260_68 = W*in
   wire signed [14:0] m260_68;
   assign m260_68 =15'b0;

   // m260_69 = W*in
   wire signed [14:0] m260_69;
   assign m260_69 ={ {4{in260[14]}} , in260[14:4] };

   // m260_70 = W*in
   wire signed [14:0] m260_70;
   assign m260_70 =15'b0;

   // m260_71 = W*in
   wire signed [14:0] m260_71;
   assign m260_71 =15'b0;

   // m260_72 = W*in
   wire signed [14:0] m260_72;
   assign m260_72 =15'b0;

   // m260_73 = W*in
   wire signed [14:0] m260_73;
   assign m260_73 =15'b0;

   // m260_74 = W*in
   wire signed [14:0] m260_74;
   assign m260_74 ={ {4{neg260[14]}} , neg260[14:4] };

   // m260_75 = W*in
   wire signed [14:0] m260_75;
   assign m260_75 =15'b0;

   // m260_76 = W*in
   wire signed [14:0] m260_76;
   assign m260_76 =15'b0;

   // m260_77 = W*in
   wire signed [14:0] m260_77;
   assign m260_77 =15'b0;

   // m260_78 = W*in
   wire signed [14:0] m260_78;
   assign m260_78 =15'b0;

   // m260_79 = W*in
   wire signed [14:0] m260_79;
   assign m260_79 =15'b0;

   // m260_80 = W*in
   wire signed [14:0] m260_80;
   assign m260_80 =15'b0;

   // m260_81 = W*in
   wire signed [14:0] m260_81;
   assign m260_81 =15'b0;

   // m260_82 = W*in
   wire signed [14:0] m260_82;
   assign m260_82 ={ {3{neg260[14]}} , neg260[14:3] };

   // m260_83 = W*in
   wire signed [14:0] m260_83;
   assign m260_83 =15'b0;

   // m260_84 = W*in
   wire signed [14:0] m260_84;
   assign m260_84 =15'b0;

   // m260_85 = W*in
   wire signed [14:0] m260_85;
   assign m260_85 =15'b0;

   // m260_86 = W*in
   wire signed [14:0] m260_86;
   assign m260_86 =15'b0;

   // m260_87 = W*in
   wire signed [14:0] m260_87;
   assign m260_87 =15'b0;

   // m260_88 = W*in
   wire signed [14:0] m260_88;
   assign m260_88 =15'b0;

   // m260_89 = W*in
   wire signed [14:0] m260_89;
   assign m260_89 =15'b0;

   // m260_90 = W*in
   wire signed [14:0] m260_90;
   assign m260_90 =15'b0;

   // m260_91 = W*in
   wire signed [14:0] m260_91;
   assign m260_91 =15'b0;

   // m260_92 = W*in
   wire signed [14:0] m260_92;
   assign m260_92 =15'b0;

   // m260_93 = W*in
   wire signed [14:0] m260_93;
   assign m260_93 =15'b0;

   // m260_94 = W*in
   wire signed [14:0] m260_94;
   assign m260_94 =15'b0;

   // m260_95 = W*in
   wire signed [14:0] m260_95;
   assign m260_95 =15'b0;

   // m260_96 = W*in
   wire signed [14:0] m260_96;
   assign m260_96 =15'b0;

   // m260_97 = W*in
   wire signed [14:0] m260_97;
   assign m260_97 =15'b0;

   // m260_98 = W*in
   wire signed [14:0] m260_98;
   assign m260_98 =15'b0;

   // m260_99 = W*in
   wire signed [14:0] m260_99;
   assign m260_99 =15'b0;

   // m260_100 = W*in
   wire signed [14:0] m260_100;
   assign m260_100 =15'b0;

   // m261_1 = W*in
   wire signed [14:0] m261_1;
   assign m261_1 =15'b0;

   // m261_2 = W*in
   wire signed [14:0] m261_2;
   assign m261_2 =15'b0;

   // m261_3 = W*in
   wire signed [14:0] m261_3;
   assign m261_3 =15'b0;

   // m261_4 = W*in
   wire signed [14:0] m261_4;
   assign m261_4 =15'b0;

   // m261_5 = W*in
   wire signed [14:0] m261_5;
   assign m261_5 =15'b0;

   // m261_6 = W*in
   wire signed [14:0] m261_6;
   assign m261_6 =15'b0;

   // m261_7 = W*in
   wire signed [14:0] m261_7;
   assign m261_7 =15'b0;

   // m261_8 = W*in
   wire signed [14:0] m261_8;
   assign m261_8 =15'b0;

   // m261_9 = W*in
   wire signed [14:0] m261_9;
   assign m261_9 =15'b0;

   // m261_10 = W*in
   wire signed [14:0] m261_10;
   assign m261_10 =15'b0;

   // m261_11 = W*in
   wire signed [14:0] m261_11;
   assign m261_11 =15'b0;

   // m261_12 = W*in
   wire signed [14:0] m261_12;
   assign m261_12 =15'b0;

   // m261_13 = W*in
   wire signed [14:0] m261_13;
   assign m261_13 ={ {3{neg261[14]}} , neg261[14:3] };

   // m261_14 = W*in
   wire signed [14:0] m261_14;
   assign m261_14 =15'b0;

   // m261_15 = W*in
   wire signed [14:0] m261_15;
   assign m261_15 =15'b0;

   // m261_16 = W*in
   wire signed [14:0] m261_16;
   assign m261_16 =15'b0;

   // m261_17 = W*in
   wire signed [14:0] m261_17;
   assign m261_17 =15'b0;

   // m261_18 = W*in
   wire signed [14:0] m261_18;
   assign m261_18 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_19 = W*in
   wire signed [14:0] m261_19;
   assign m261_19 =15'b0;

   // m261_20 = W*in
   wire signed [14:0] m261_20;
   assign m261_20 =15'b0;

   // m261_21 = W*in
   wire signed [14:0] m261_21;
   assign m261_21 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_22 = W*in
   wire signed [14:0] m261_22;
   assign m261_22 =15'b0;

   // m261_23 = W*in
   wire signed [14:0] m261_23;
   assign m261_23 =15'b0;

   // m261_24 = W*in
   wire signed [14:0] m261_24;
   assign m261_24 ={ {4{in261[14]}} , in261[14:4] };

   // m261_25 = W*in
   wire signed [14:0] m261_25;
   assign m261_25 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_26 = W*in
   wire signed [14:0] m261_26;
   assign m261_26 =15'b0;

   // m261_27 = W*in
   wire signed [14:0] m261_27;
   assign m261_27 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_28 = W*in
   wire signed [14:0] m261_28;
   assign m261_28 =15'b0;

   // m261_29 = W*in
   wire signed [14:0] m261_29;
   assign m261_29 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_30 = W*in
   wire signed [14:0] m261_30;
   assign m261_30 =15'b0;

   // m261_31 = W*in
   wire signed [14:0] m261_31;
   assign m261_31 =15'b0;

   // m261_32 = W*in
   wire signed [14:0] m261_32;
   assign m261_32 =15'b0;

   // m261_33 = W*in
   wire signed [14:0] m261_33;
   assign m261_33 =15'b0;

   // m261_34 = W*in
   wire signed [14:0] m261_34;
   assign m261_34 =15'b0;

   // m261_35 = W*in
   wire signed [14:0] m261_35;
   assign m261_35 =15'b0;

   // m261_36 = W*in
   wire signed [14:0] m261_36;
   assign m261_36 =15'b0;

   // m261_37 = W*in
   wire signed [14:0] m261_37;
   assign m261_37 =15'b0;

   // m261_38 = W*in
   wire signed [14:0] m261_38;
   assign m261_38 =15'b0;

   // m261_39 = W*in
   wire signed [14:0] m261_39;
   assign m261_39 =15'b0;

   // m261_40 = W*in
   wire signed [14:0] m261_40;
   assign m261_40 ={ {4{in261[14]}} , in261[14:4] };

   // m261_41 = W*in
   wire signed [14:0] m261_41;
   assign m261_41 =15'b0;

   // m261_42 = W*in
   wire signed [14:0] m261_42;
   assign m261_42 =15'b0;

   // m261_43 = W*in
   wire signed [14:0] m261_43;
   assign m261_43 =15'b0;

   // m261_44 = W*in
   wire signed [14:0] m261_44;
   assign m261_44 =15'b0;

   // m261_45 = W*in
   wire signed [14:0] m261_45;
   assign m261_45 =15'b0;

   // m261_46 = W*in
   wire signed [14:0] m261_46;
   assign m261_46 =15'b0;

   // m261_47 = W*in
   wire signed [14:0] m261_47;
   assign m261_47 =15'b0;

   // m261_48 = W*in
   wire signed [14:0] m261_48;
   assign m261_48 =15'b0;

   // m261_49 = W*in
   wire signed [14:0] m261_49;
   assign m261_49 =15'b0;

   // m261_50 = W*in
   wire signed [14:0] m261_50;
   assign m261_50 =15'b0;

   // m261_51 = W*in
   wire signed [14:0] m261_51;
   assign m261_51 =15'b0;

   // m261_52 = W*in
   wire signed [14:0] m261_52;
   assign m261_52 =15'b0;

   // m261_53 = W*in
   wire signed [14:0] m261_53;
   assign m261_53 =15'b0;

   // m261_54 = W*in
   wire signed [14:0] m261_54;
   assign m261_54 =15'b0;

   // m261_55 = W*in
   wire signed [14:0] m261_55;
   assign m261_55 =15'b0;

   // m261_56 = W*in
   wire signed [14:0] m261_56;
   assign m261_56 =15'b0;

   // m261_57 = W*in
   wire signed [14:0] m261_57;
   assign m261_57 =15'b0;

   // m261_58 = W*in
   wire signed [14:0] m261_58;
   assign m261_58 =15'b0;

   // m261_59 = W*in
   wire signed [14:0] m261_59;
   assign m261_59 ={ {4{in261[14]}} , in261[14:4] };

   // m261_60 = W*in
   wire signed [14:0] m261_60;
   assign m261_60 =15'b0;

   // m261_61 = W*in
   wire signed [14:0] m261_61;
   assign m261_61 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_62 = W*in
   wire signed [14:0] m261_62;
   assign m261_62 =15'b0;

   // m261_63 = W*in
   wire signed [14:0] m261_63;
   assign m261_63 =15'b0;

   // m261_64 = W*in
   wire signed [14:0] m261_64;
   assign m261_64 =15'b0;

   // m261_65 = W*in
   wire signed [14:0] m261_65;
   assign m261_65 =15'b0;

   // m261_66 = W*in
   wire signed [14:0] m261_66;
   assign m261_66 =15'b0;

   // m261_67 = W*in
   wire signed [14:0] m261_67;
   assign m261_67 =15'b0;

   // m261_68 = W*in
   wire signed [14:0] m261_68;
   assign m261_68 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_69 = W*in
   wire signed [14:0] m261_69;
   assign m261_69 =15'b0;

   // m261_70 = W*in
   wire signed [14:0] m261_70;
   assign m261_70 ={ {4{in261[14]}} , in261[14:4] };

   // m261_71 = W*in
   wire signed [14:0] m261_71;
   assign m261_71 =15'b0;

   // m261_72 = W*in
   wire signed [14:0] m261_72;
   assign m261_72 =15'b0;

   // m261_73 = W*in
   wire signed [14:0] m261_73;
   assign m261_73 =15'b0;

   // m261_74 = W*in
   wire signed [14:0] m261_74;
   assign m261_74 =15'b0;

   // m261_75 = W*in
   wire signed [14:0] m261_75;
   assign m261_75 =15'b0;

   // m261_76 = W*in
   wire signed [14:0] m261_76;
   assign m261_76 =15'b0;

   // m261_77 = W*in
   wire signed [14:0] m261_77;
   assign m261_77 =15'b0;

   // m261_78 = W*in
   wire signed [14:0] m261_78;
   assign m261_78 ={ {4{neg261[14]}} , neg261[14:4] };

   // m261_79 = W*in
   wire signed [14:0] m261_79;
   assign m261_79 =15'b0;

   // m261_80 = W*in
   wire signed [14:0] m261_80;
   assign m261_80 =15'b0;

   // m261_81 = W*in
   wire signed [14:0] m261_81;
   assign m261_81 =15'b0;

   // m261_82 = W*in
   wire signed [14:0] m261_82;
   assign m261_82 =15'b0;

   // m261_83 = W*in
   wire signed [14:0] m261_83;
   assign m261_83 =15'b0;

   // m261_84 = W*in
   wire signed [14:0] m261_84;
   assign m261_84 =15'b0;

   // m261_85 = W*in
   wire signed [14:0] m261_85;
   assign m261_85 =15'b0;

   // m261_86 = W*in
   wire signed [14:0] m261_86;
   assign m261_86 =15'b0;

   // m261_87 = W*in
   wire signed [14:0] m261_87;
   assign m261_87 =15'b0;

   // m261_88 = W*in
   wire signed [14:0] m261_88;
   assign m261_88 =15'b0;

   // m261_89 = W*in
   wire signed [14:0] m261_89;
   assign m261_89 =15'b0;

   // m261_90 = W*in
   wire signed [14:0] m261_90;
   assign m261_90 =15'b0;

   // m261_91 = W*in
   wire signed [14:0] m261_91;
   assign m261_91 =15'b0;

   // m261_92 = W*in
   wire signed [14:0] m261_92;
   assign m261_92 =15'b0;

   // m261_93 = W*in
   wire signed [14:0] m261_93;
   assign m261_93 =15'b0;

   // m261_94 = W*in
   wire signed [14:0] m261_94;
   assign m261_94 =15'b0;

   // m261_95 = W*in
   wire signed [14:0] m261_95;
   assign m261_95 =15'b0;

   // m261_96 = W*in
   wire signed [14:0] m261_96;
   assign m261_96 =15'b0;

   // m261_97 = W*in
   wire signed [14:0] m261_97;
   assign m261_97 =15'b0;

   // m261_98 = W*in
   wire signed [14:0] m261_98;
   assign m261_98 =15'b0;

   // m261_99 = W*in
   wire signed [14:0] m261_99;
   assign m261_99 =15'b0;

   // m261_100 = W*in
   wire signed [14:0] m261_100;
   assign m261_100 =15'b0;

   // m262_1 = W*in
   wire signed [14:0] m262_1;
   assign m262_1 =15'b0;

   // m262_2 = W*in
   wire signed [14:0] m262_2;
   assign m262_2 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_3 = W*in
   wire signed [14:0] m262_3;
   assign m262_3 =15'b0;

   // m262_4 = W*in
   wire signed [14:0] m262_4;
   assign m262_4 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_5 = W*in
   wire signed [14:0] m262_5;
   assign m262_5 =15'b0;

   // m262_6 = W*in
   wire signed [14:0] m262_6;
   assign m262_6 ={ {3{in262[14]}} , in262[14:3] };

   // m262_7 = W*in
   wire signed [14:0] m262_7;
   assign m262_7 ={ {3{in262[14]}} , in262[14:3] };

   // m262_8 = W*in
   wire signed [14:0] m262_8;
   assign m262_8 ={ {3{in262[14]}} , in262[14:3] };

   // m262_9 = W*in
   wire signed [14:0] m262_9;
   assign m262_9 =15'b0;

   // m262_10 = W*in
   wire signed [14:0] m262_10;
   assign m262_10 ={ {3{in262[14]}} , in262[14:3] };

   // m262_11 = W*in
   wire signed [14:0] m262_11;
   assign m262_11 =15'b0;

   // m262_12 = W*in
   wire signed [14:0] m262_12;
   assign m262_12 =15'b0;

   // m262_13 = W*in
   wire signed [14:0] m262_13;
   assign m262_13 =15'b0;

   // m262_14 = W*in
   wire signed [14:0] m262_14;
   assign m262_14 ={ {3{in262[14]}} , in262[14:3] };

   // m262_15 = W*in
   wire signed [14:0] m262_15;
   assign m262_15 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_16 = W*in
   wire signed [14:0] m262_16;
   assign m262_16 =15'b0;

   // m262_17 = W*in
   wire signed [14:0] m262_17;
   assign m262_17 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_18 = W*in
   wire signed [14:0] m262_18;
   assign m262_18 ={ {4{in262[14]}} , in262[14:4] };

   // m262_19 = W*in
   wire signed [14:0] m262_19;
   assign m262_19 =15'b0;

   // m262_20 = W*in
   wire signed [14:0] m262_20;
   assign m262_20 =15'b0;

   // m262_21 = W*in
   wire signed [14:0] m262_21;
   assign m262_21 =15'b0;

   // m262_22 = W*in
   wire signed [14:0] m262_22;
   assign m262_22 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_23 = W*in
   wire signed [14:0] m262_23;
   assign m262_23 =15'b0;

   // m262_24 = W*in
   wire signed [14:0] m262_24;
   assign m262_24 ={ {3{in262[14]}} , in262[14:3] };

   // m262_25 = W*in
   wire signed [14:0] m262_25;
   assign m262_25 =15'b0;

   // m262_26 = W*in
   wire signed [14:0] m262_26;
   assign m262_26 =15'b0;

   // m262_27 = W*in
   wire signed [14:0] m262_27;
   assign m262_27 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_28 = W*in
   wire signed [14:0] m262_28;
   assign m262_28 =15'b0;

   // m262_29 = W*in
   wire signed [14:0] m262_29;
   assign m262_29 =15'b0;

   // m262_30 = W*in
   wire signed [14:0] m262_30;
   assign m262_30 =15'b0;

   // m262_31 = W*in
   wire signed [14:0] m262_31;
   assign m262_31 ={ {3{in262[14]}} , in262[14:3] };

   // m262_32 = W*in
   wire signed [14:0] m262_32;
   assign m262_32 =15'b0;

   // m262_33 = W*in
   wire signed [14:0] m262_33;
   assign m262_33 =15'b0;

   // m262_34 = W*in
   wire signed [14:0] m262_34;
   assign m262_34 =15'b0;

   // m262_35 = W*in
   wire signed [14:0] m262_35;
   assign m262_35 =15'b0;

   // m262_36 = W*in
   wire signed [14:0] m262_36;
   assign m262_36 =15'b0;

   // m262_37 = W*in
   wire signed [14:0] m262_37;
   assign m262_37 =15'b0;

   // m262_38 = W*in
   wire signed [14:0] m262_38;
   assign m262_38 =15'b0;

   // m262_39 = W*in
   wire signed [14:0] m262_39;
   assign m262_39 =15'b0;

   // m262_40 = W*in
   wire signed [14:0] m262_40;
   assign m262_40 ={ {4{neg262[14]}} , neg262[14:4] };

   // m262_41 = W*in
   wire signed [14:0] m262_41;
   assign m262_41 =15'b0;

   // m262_42 = W*in
   wire signed [14:0] m262_42;
   assign m262_42 =15'b0;

   // m262_43 = W*in
   wire signed [14:0] m262_43;
   assign m262_43 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_44 = W*in
   wire signed [14:0] m262_44;
   assign m262_44 =15'b0;

   // m262_45 = W*in
   wire signed [14:0] m262_45;
   assign m262_45 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_46 = W*in
   wire signed [14:0] m262_46;
   assign m262_46 =15'b0;

   // m262_47 = W*in
   wire signed [14:0] m262_47;
   assign m262_47 ={ {3{in262[14]}} , in262[14:3] };

   // m262_48 = W*in
   wire signed [14:0] m262_48;
   assign m262_48 =15'b0;

   // m262_49 = W*in
   wire signed [14:0] m262_49;
   assign m262_49 =15'b0;

   // m262_50 = W*in
   wire signed [14:0] m262_50;
   assign m262_50 =15'b0;

   // m262_51 = W*in
   wire signed [14:0] m262_51;
   assign m262_51 ={ {3{in262[14]}} , in262[14:3] };

   // m262_52 = W*in
   wire signed [14:0] m262_52;
   assign m262_52 =15'b0;

   // m262_53 = W*in
   wire signed [14:0] m262_53;
   assign m262_53 =15'b0;

   // m262_54 = W*in
   wire signed [14:0] m262_54;
   assign m262_54 =15'b0;

   // m262_55 = W*in
   wire signed [14:0] m262_55;
   assign m262_55 =15'b0;

   // m262_56 = W*in
   wire signed [14:0] m262_56;
   assign m262_56 =15'b0;

   // m262_57 = W*in
   wire signed [14:0] m262_57;
   assign m262_57 ={ {4{in262[14]}} , in262[14:4] };

   // m262_58 = W*in
   wire signed [14:0] m262_58;
   assign m262_58 ={ {4{neg262[14]}} , neg262[14:4] };

   // m262_59 = W*in
   wire signed [14:0] m262_59;
   assign m262_59 ={ {4{neg262[14]}} , neg262[14:4] };

   // m262_60 = W*in
   wire signed [14:0] m262_60;
   assign m262_60 =15'b0;

   // m262_61 = W*in
   wire signed [14:0] m262_61;
   assign m262_61 =15'b0;

   // m262_62 = W*in
   wire signed [14:0] m262_62;
   assign m262_62 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_63 = W*in
   wire signed [14:0] m262_63;
   assign m262_63 ={ {2{in262[14]}} , in262[14:2] };

   // m262_64 = W*in
   wire signed [14:0] m262_64;
   assign m262_64 ={ {4{neg262[14]}} , neg262[14:4] };

   // m262_65 = W*in
   wire signed [14:0] m262_65;
   assign m262_65 =15'b0;

   // m262_66 = W*in
   wire signed [14:0] m262_66;
   assign m262_66 ={ {4{in262[14]}} , in262[14:4] };

   // m262_67 = W*in
   wire signed [14:0] m262_67;
   assign m262_67 =15'b0;

   // m262_68 = W*in
   wire signed [14:0] m262_68;
   assign m262_68 =15'b0;

   // m262_69 = W*in
   wire signed [14:0] m262_69;
   assign m262_69 =15'b0;

   // m262_70 = W*in
   wire signed [14:0] m262_70;
   assign m262_70 =15'b0;

   // m262_71 = W*in
   wire signed [14:0] m262_71;
   assign m262_71 ={ {3{in262[14]}} , in262[14:3] };

   // m262_72 = W*in
   wire signed [14:0] m262_72;
   assign m262_72 =15'b0;

   // m262_73 = W*in
   wire signed [14:0] m262_73;
   assign m262_73 ={ {3{in262[14]}} , in262[14:3] };

   // m262_74 = W*in
   wire signed [14:0] m262_74;
   assign m262_74 ={ {4{neg262[14]}} , neg262[14:4] };

   // m262_75 = W*in
   wire signed [14:0] m262_75;
   assign m262_75 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_76 = W*in
   wire signed [14:0] m262_76;
   assign m262_76 ={ {4{neg262[14]}} , neg262[14:4] };

   // m262_77 = W*in
   wire signed [14:0] m262_77;
   assign m262_77 ={ {3{in262[14]}} , in262[14:3] };

   // m262_78 = W*in
   wire signed [14:0] m262_78;
   assign m262_78 =15'b0;

   // m262_79 = W*in
   wire signed [14:0] m262_79;
   assign m262_79 =15'b0;

   // m262_80 = W*in
   wire signed [14:0] m262_80;
   assign m262_80 =15'b0;

   // m262_81 = W*in
   wire signed [14:0] m262_81;
   assign m262_81 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_82 = W*in
   wire signed [14:0] m262_82;
   assign m262_82 =15'b0;

   // m262_83 = W*in
   wire signed [14:0] m262_83;
   assign m262_83 =15'b0;

   // m262_84 = W*in
   wire signed [14:0] m262_84;
   assign m262_84 =15'b0;

   // m262_85 = W*in
   wire signed [14:0] m262_85;
   assign m262_85 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_86 = W*in
   wire signed [14:0] m262_86;
   assign m262_86 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_87 = W*in
   wire signed [14:0] m262_87;
   assign m262_87 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_88 = W*in
   wire signed [14:0] m262_88;
   assign m262_88 =15'b0;

   // m262_89 = W*in
   wire signed [14:0] m262_89;
   assign m262_89 ={ {3{in262[14]}} , in262[14:3] };

   // m262_90 = W*in
   wire signed [14:0] m262_90;
   assign m262_90 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_91 = W*in
   wire signed [14:0] m262_91;
   assign m262_91 ={ {3{in262[14]}} , in262[14:3] };

   // m262_92 = W*in
   wire signed [14:0] m262_92;
   assign m262_92 =15'b0;

   // m262_93 = W*in
   wire signed [14:0] m262_93;
   assign m262_93 =15'b0;

   // m262_94 = W*in
   wire signed [14:0] m262_94;
   assign m262_94 =15'b0;

   // m262_95 = W*in
   wire signed [14:0] m262_95;
   assign m262_95 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_96 = W*in
   wire signed [14:0] m262_96;
   assign m262_96 ={ {3{in262[14]}} , in262[14:3] };

   // m262_97 = W*in
   wire signed [14:0] m262_97;
   assign m262_97 ={ {3{neg262[14]}} , neg262[14:3] };

   // m262_98 = W*in
   wire signed [14:0] m262_98;
   assign m262_98 =15'b0;

   // m262_99 = W*in
   wire signed [14:0] m262_99;
   assign m262_99 =15'b0;

   // m262_100 = W*in
   wire signed [14:0] m262_100;
   assign m262_100 =15'b0;

   // m263_1 = W*in
   wire signed [14:0] m263_1;
   assign m263_1 =15'b0;

   // m263_2 = W*in
   wire signed [14:0] m263_2;
   assign m263_2 =15'b0;

   // m263_3 = W*in
   wire signed [14:0] m263_3;
   assign m263_3 =15'b0;

   // m263_4 = W*in
   wire signed [14:0] m263_4;
   assign m263_4 =15'b0;

   // m263_5 = W*in
   wire signed [14:0] m263_5;
   assign m263_5 =15'b0;

   // m263_6 = W*in
   wire signed [14:0] m263_6;
   assign m263_6 =15'b0;

   // m263_7 = W*in
   wire signed [14:0] m263_7;
   assign m263_7 =15'b0;

   // m263_8 = W*in
   wire signed [14:0] m263_8;
   assign m263_8 =15'b0;

   // m263_9 = W*in
   wire signed [14:0] m263_9;
   assign m263_9 =15'b0;

   // m263_10 = W*in
   wire signed [14:0] m263_10;
   assign m263_10 =15'b0;

   // m263_11 = W*in
   wire signed [14:0] m263_11;
   assign m263_11 ={ {3{neg263[14]}} , neg263[14:3] };

   // m263_12 = W*in
   wire signed [14:0] m263_12;
   assign m263_12 =15'b0;

   // m263_13 = W*in
   wire signed [14:0] m263_13;
   assign m263_13 =15'b0;

   // m263_14 = W*in
   wire signed [14:0] m263_14;
   assign m263_14 =15'b0;

   // m263_15 = W*in
   wire signed [14:0] m263_15;
   assign m263_15 ={ {4{in263[14]}} , in263[14:4] };

   // m263_16 = W*in
   wire signed [14:0] m263_16;
   assign m263_16 =15'b0;

   // m263_17 = W*in
   wire signed [14:0] m263_17;
   assign m263_17 =15'b0;

   // m263_18 = W*in
   wire signed [14:0] m263_18;
   assign m263_18 =15'b0;

   // m263_19 = W*in
   wire signed [14:0] m263_19;
   assign m263_19 =15'b0;

   // m263_20 = W*in
   wire signed [14:0] m263_20;
   assign m263_20 ={ {3{in263[14]}} , in263[14:3] };

   // m263_21 = W*in
   wire signed [14:0] m263_21;
   assign m263_21 =15'b0;

   // m263_22 = W*in
   wire signed [14:0] m263_22;
   assign m263_22 =15'b0;

   // m263_23 = W*in
   wire signed [14:0] m263_23;
   assign m263_23 =15'b0;

   // m263_24 = W*in
   wire signed [14:0] m263_24;
   assign m263_24 =15'b0;

   // m263_25 = W*in
   wire signed [14:0] m263_25;
   assign m263_25 =15'b0;

   // m263_26 = W*in
   wire signed [14:0] m263_26;
   assign m263_26 ={ {4{neg263[14]}} , neg263[14:4] };

   // m263_27 = W*in
   wire signed [14:0] m263_27;
   assign m263_27 =15'b0;

   // m263_28 = W*in
   wire signed [14:0] m263_28;
   assign m263_28 =15'b0;

   // m263_29 = W*in
   wire signed [14:0] m263_29;
   assign m263_29 =15'b0;

   // m263_30 = W*in
   wire signed [14:0] m263_30;
   assign m263_30 =15'b0;

   // m263_31 = W*in
   wire signed [14:0] m263_31;
   assign m263_31 =15'b0;

   // m263_32 = W*in
   wire signed [14:0] m263_32;
   assign m263_32 =15'b0;

   // m263_33 = W*in
   wire signed [14:0] m263_33;
   assign m263_33 =15'b0;

   // m263_34 = W*in
   wire signed [14:0] m263_34;
   assign m263_34 =15'b0;

   // m263_35 = W*in
   wire signed [14:0] m263_35;
   assign m263_35 =15'b0;

   // m263_36 = W*in
   wire signed [14:0] m263_36;
   assign m263_36 =15'b0;

   // m263_37 = W*in
   wire signed [14:0] m263_37;
   assign m263_37 =15'b0;

   // m263_38 = W*in
   wire signed [14:0] m263_38;
   assign m263_38 =15'b0;

   // m263_39 = W*in
   wire signed [14:0] m263_39;
   assign m263_39 ={ {3{neg263[14]}} , neg263[14:3] };

   // m263_40 = W*in
   wire signed [14:0] m263_40;
   assign m263_40 =15'b0;

   // m263_41 = W*in
   wire signed [14:0] m263_41;
   assign m263_41 =15'b0;

   // m263_42 = W*in
   wire signed [14:0] m263_42;
   assign m263_42 =15'b0;

   // m263_43 = W*in
   wire signed [14:0] m263_43;
   assign m263_43 =15'b0;

   // m263_44 = W*in
   wire signed [14:0] m263_44;
   assign m263_44 =15'b0;

   // m263_45 = W*in
   wire signed [14:0] m263_45;
   assign m263_45 ={ {3{neg263[14]}} , neg263[14:3] };

   // m263_46 = W*in
   wire signed [14:0] m263_46;
   assign m263_46 =15'b0;

   // m263_47 = W*in
   wire signed [14:0] m263_47;
   assign m263_47 =15'b0;

   // m263_48 = W*in
   wire signed [14:0] m263_48;
   assign m263_48 =15'b0;

   // m263_49 = W*in
   wire signed [14:0] m263_49;
   assign m263_49 =15'b0;

   // m263_50 = W*in
   wire signed [14:0] m263_50;
   assign m263_50 =15'b0;

   // m263_51 = W*in
   wire signed [14:0] m263_51;
   assign m263_51 =15'b0;

   // m263_52 = W*in
   wire signed [14:0] m263_52;
   assign m263_52 =15'b0;

   // m263_53 = W*in
   wire signed [14:0] m263_53;
   assign m263_53 =15'b0;

   // m263_54 = W*in
   wire signed [14:0] m263_54;
   assign m263_54 =15'b0;

   // m263_55 = W*in
   wire signed [14:0] m263_55;
   assign m263_55 =15'b0;

   // m263_56 = W*in
   wire signed [14:0] m263_56;
   assign m263_56 =15'b0;

   // m263_57 = W*in
   wire signed [14:0] m263_57;
   assign m263_57 =15'b0;

   // m263_58 = W*in
   wire signed [14:0] m263_58;
   assign m263_58 =15'b0;

   // m263_59 = W*in
   wire signed [14:0] m263_59;
   assign m263_59 =15'b0;

   // m263_60 = W*in
   wire signed [14:0] m263_60;
   assign m263_60 =15'b0;

   // m263_61 = W*in
   wire signed [14:0] m263_61;
   assign m263_61 =15'b0;

   // m263_62 = W*in
   wire signed [14:0] m263_62;
   assign m263_62 =15'b0;

   // m263_63 = W*in
   wire signed [14:0] m263_63;
   assign m263_63 =15'b0;

   // m263_64 = W*in
   wire signed [14:0] m263_64;
   assign m263_64 =15'b0;

   // m263_65 = W*in
   wire signed [14:0] m263_65;
   assign m263_65 =15'b0;

   // m263_66 = W*in
   wire signed [14:0] m263_66;
   assign m263_66 =15'b0;

   // m263_67 = W*in
   wire signed [14:0] m263_67;
   assign m263_67 ={ {3{in263[14]}} , in263[14:3] };

   // m263_68 = W*in
   wire signed [14:0] m263_68;
   assign m263_68 ={ {4{in263[14]}} , in263[14:4] };

   // m263_69 = W*in
   wire signed [14:0] m263_69;
   assign m263_69 =15'b0;

   // m263_70 = W*in
   wire signed [14:0] m263_70;
   assign m263_70 ={ {3{neg263[14]}} , neg263[14:3] };

   // m263_71 = W*in
   wire signed [14:0] m263_71;
   assign m263_71 =15'b0;

   // m263_72 = W*in
   wire signed [14:0] m263_72;
   assign m263_72 =15'b0;

   // m263_73 = W*in
   wire signed [14:0] m263_73;
   assign m263_73 =15'b0;

   // m263_74 = W*in
   wire signed [14:0] m263_74;
   assign m263_74 =15'b0;

   // m263_75 = W*in
   wire signed [14:0] m263_75;
   assign m263_75 =15'b0;

   // m263_76 = W*in
   wire signed [14:0] m263_76;
   assign m263_76 ={ {4{neg263[14]}} , neg263[14:4] };

   // m263_77 = W*in
   wire signed [14:0] m263_77;
   assign m263_77 =15'b0;

   // m263_78 = W*in
   wire signed [14:0] m263_78;
   assign m263_78 =15'b0;

   // m263_79 = W*in
   wire signed [14:0] m263_79;
   assign m263_79 =15'b0;

   // m263_80 = W*in
   wire signed [14:0] m263_80;
   assign m263_80 ={ {4{neg263[14]}} , neg263[14:4] };

   // m263_81 = W*in
   wire signed [14:0] m263_81;
   assign m263_81 =15'b0;

   // m263_82 = W*in
   wire signed [14:0] m263_82;
   assign m263_82 =15'b0;

   // m263_83 = W*in
   wire signed [14:0] m263_83;
   assign m263_83 =15'b0;

   // m263_84 = W*in
   wire signed [14:0] m263_84;
   assign m263_84 =15'b0;

   // m263_85 = W*in
   wire signed [14:0] m263_85;
   assign m263_85 =15'b0;

   // m263_86 = W*in
   wire signed [14:0] m263_86;
   assign m263_86 =15'b0;

   // m263_87 = W*in
   wire signed [14:0] m263_87;
   assign m263_87 =15'b0;

   // m263_88 = W*in
   wire signed [14:0] m263_88;
   assign m263_88 ={ {3{in263[14]}} , in263[14:3] };

   // m263_89 = W*in
   wire signed [14:0] m263_89;
   assign m263_89 =15'b0;

   // m263_90 = W*in
   wire signed [14:0] m263_90;
   assign m263_90 =15'b0;

   // m263_91 = W*in
   wire signed [14:0] m263_91;
   assign m263_91 =15'b0;

   // m263_92 = W*in
   wire signed [14:0] m263_92;
   assign m263_92 =15'b0;

   // m263_93 = W*in
   wire signed [14:0] m263_93;
   assign m263_93 ={ {3{neg263[14]}} , neg263[14:3] };

   // m263_94 = W*in
   wire signed [14:0] m263_94;
   assign m263_94 =15'b0;

   // m263_95 = W*in
   wire signed [14:0] m263_95;
   assign m263_95 ={ {4{in263[14]}} , in263[14:4] };

   // m263_96 = W*in
   wire signed [14:0] m263_96;
   assign m263_96 =15'b0;

   // m263_97 = W*in
   wire signed [14:0] m263_97;
   assign m263_97 =15'b0;

   // m263_98 = W*in
   wire signed [14:0] m263_98;
   assign m263_98 =15'b0;

   // m263_99 = W*in
   wire signed [14:0] m263_99;
   assign m263_99 =15'b0;

   // m263_100 = W*in
   wire signed [14:0] m263_100;
   assign m263_100 ={ {4{neg263[14]}} , neg263[14:4] };

   //Perceptron Adders
   assign out1 = m1_1+m2_1+m3_1+m4_1+m5_1+m6_1+m7_1+m8_1+m9_1+m10_1+m11_1+m12_1+m13_1+m14_1+m15_1+m16_1+m17_1+m18_1+m19_1+m20_1+m21_1+m22_1+m23_1+m24_1+m25_1+m26_1+m27_1+m28_1+m29_1+m30_1+m31_1+m32_1+m33_1+m34_1+m35_1+m36_1+m37_1+m38_1+m39_1+m40_1+m41_1+m42_1+m43_1+m44_1+m45_1+m46_1+m47_1+m48_1+m49_1+m50_1+m51_1+m52_1+m53_1+m54_1+m55_1+m56_1+m57_1+m58_1+m59_1+m60_1+m61_1+m62_1+m63_1+m64_1+m65_1+m66_1+m67_1+m68_1+m69_1+m70_1+m71_1+m72_1+m73_1+m74_1+m75_1+m76_1+m77_1+m78_1+m79_1+m80_1+m81_1+m82_1+m83_1+m84_1+m85_1+m86_1+m87_1+m88_1+m89_1+m90_1+m91_1+m92_1+m93_1+m94_1+m95_1+m96_1+m97_1+m98_1+m99_1+m100_1+m101_1+m102_1+m103_1+m104_1+m105_1+m106_1+m107_1+m108_1+m109_1+m110_1+m111_1+m112_1+m113_1+m114_1+m115_1+m116_1+m117_1+m118_1+m119_1+m120_1+m121_1+m122_1+m123_1+m124_1+m125_1+m126_1+m127_1+m128_1+m129_1+m130_1+m131_1+m132_1+m133_1+m134_1+m135_1+m136_1+m137_1+m138_1+m139_1+m140_1+m141_1+m142_1+m143_1+m144_1+m145_1+m146_1+m147_1+m148_1+m149_1+m150_1+m151_1+m152_1+m153_1+m154_1+m155_1+m156_1+m157_1+m158_1+m159_1+m160_1+m161_1+m162_1+m163_1+m164_1+m165_1+m166_1+m167_1+m168_1+m169_1+m170_1+m171_1+m172_1+m173_1+m174_1+m175_1+m176_1+m177_1+m178_1+m179_1+m180_1+m181_1+m182_1+m183_1+m184_1+m185_1+m186_1+m187_1+m188_1+m189_1+m190_1+m191_1+m192_1+m193_1+m194_1+m195_1+m196_1+m197_1+m198_1+m199_1+m200_1+m201_1+m202_1+m203_1+m204_1+m205_1+m206_1+m207_1+m208_1+m209_1+m210_1+m211_1+m212_1+m213_1+m214_1+m215_1+m216_1+m217_1+m218_1+m219_1+m220_1+m221_1+m222_1+m223_1+m224_1+m225_1+m226_1+m227_1+m228_1+m229_1+m230_1+m231_1+m232_1+m233_1+m234_1+m235_1+m236_1+m237_1+m238_1+m239_1+m240_1+m241_1+m242_1+m243_1+m244_1+m245_1+m246_1+m247_1+m248_1+m249_1+m250_1+m251_1+m252_1+m253_1+m254_1+m255_1+m256_1+m257_1+m258_1+m259_1+m260_1+m261_1+m262_1+m263_1+b1;
   assign out2 = m1_2+m2_2+m3_2+m4_2+m5_2+m6_2+m7_2+m8_2+m9_2+m10_2+m11_2+m12_2+m13_2+m14_2+m15_2+m16_2+m17_2+m18_2+m19_2+m20_2+m21_2+m22_2+m23_2+m24_2+m25_2+m26_2+m27_2+m28_2+m29_2+m30_2+m31_2+m32_2+m33_2+m34_2+m35_2+m36_2+m37_2+m38_2+m39_2+m40_2+m41_2+m42_2+m43_2+m44_2+m45_2+m46_2+m47_2+m48_2+m49_2+m50_2+m51_2+m52_2+m53_2+m54_2+m55_2+m56_2+m57_2+m58_2+m59_2+m60_2+m61_2+m62_2+m63_2+m64_2+m65_2+m66_2+m67_2+m68_2+m69_2+m70_2+m71_2+m72_2+m73_2+m74_2+m75_2+m76_2+m77_2+m78_2+m79_2+m80_2+m81_2+m82_2+m83_2+m84_2+m85_2+m86_2+m87_2+m88_2+m89_2+m90_2+m91_2+m92_2+m93_2+m94_2+m95_2+m96_2+m97_2+m98_2+m99_2+m100_2+m101_2+m102_2+m103_2+m104_2+m105_2+m106_2+m107_2+m108_2+m109_2+m110_2+m111_2+m112_2+m113_2+m114_2+m115_2+m116_2+m117_2+m118_2+m119_2+m120_2+m121_2+m122_2+m123_2+m124_2+m125_2+m126_2+m127_2+m128_2+m129_2+m130_2+m131_2+m132_2+m133_2+m134_2+m135_2+m136_2+m137_2+m138_2+m139_2+m140_2+m141_2+m142_2+m143_2+m144_2+m145_2+m146_2+m147_2+m148_2+m149_2+m150_2+m151_2+m152_2+m153_2+m154_2+m155_2+m156_2+m157_2+m158_2+m159_2+m160_2+m161_2+m162_2+m163_2+m164_2+m165_2+m166_2+m167_2+m168_2+m169_2+m170_2+m171_2+m172_2+m173_2+m174_2+m175_2+m176_2+m177_2+m178_2+m179_2+m180_2+m181_2+m182_2+m183_2+m184_2+m185_2+m186_2+m187_2+m188_2+m189_2+m190_2+m191_2+m192_2+m193_2+m194_2+m195_2+m196_2+m197_2+m198_2+m199_2+m200_2+m201_2+m202_2+m203_2+m204_2+m205_2+m206_2+m207_2+m208_2+m209_2+m210_2+m211_2+m212_2+m213_2+m214_2+m215_2+m216_2+m217_2+m218_2+m219_2+m220_2+m221_2+m222_2+m223_2+m224_2+m225_2+m226_2+m227_2+m228_2+m229_2+m230_2+m231_2+m232_2+m233_2+m234_2+m235_2+m236_2+m237_2+m238_2+m239_2+m240_2+m241_2+m242_2+m243_2+m244_2+m245_2+m246_2+m247_2+m248_2+m249_2+m250_2+m251_2+m252_2+m253_2+m254_2+m255_2+m256_2+m257_2+m258_2+m259_2+m260_2+m261_2+m262_2+m263_2+b2;
   assign out3 = m1_3+m2_3+m3_3+m4_3+m5_3+m6_3+m7_3+m8_3+m9_3+m10_3+m11_3+m12_3+m13_3+m14_3+m15_3+m16_3+m17_3+m18_3+m19_3+m20_3+m21_3+m22_3+m23_3+m24_3+m25_3+m26_3+m27_3+m28_3+m29_3+m30_3+m31_3+m32_3+m33_3+m34_3+m35_3+m36_3+m37_3+m38_3+m39_3+m40_3+m41_3+m42_3+m43_3+m44_3+m45_3+m46_3+m47_3+m48_3+m49_3+m50_3+m51_3+m52_3+m53_3+m54_3+m55_3+m56_3+m57_3+m58_3+m59_3+m60_3+m61_3+m62_3+m63_3+m64_3+m65_3+m66_3+m67_3+m68_3+m69_3+m70_3+m71_3+m72_3+m73_3+m74_3+m75_3+m76_3+m77_3+m78_3+m79_3+m80_3+m81_3+m82_3+m83_3+m84_3+m85_3+m86_3+m87_3+m88_3+m89_3+m90_3+m91_3+m92_3+m93_3+m94_3+m95_3+m96_3+m97_3+m98_3+m99_3+m100_3+m101_3+m102_3+m103_3+m104_3+m105_3+m106_3+m107_3+m108_3+m109_3+m110_3+m111_3+m112_3+m113_3+m114_3+m115_3+m116_3+m117_3+m118_3+m119_3+m120_3+m121_3+m122_3+m123_3+m124_3+m125_3+m126_3+m127_3+m128_3+m129_3+m130_3+m131_3+m132_3+m133_3+m134_3+m135_3+m136_3+m137_3+m138_3+m139_3+m140_3+m141_3+m142_3+m143_3+m144_3+m145_3+m146_3+m147_3+m148_3+m149_3+m150_3+m151_3+m152_3+m153_3+m154_3+m155_3+m156_3+m157_3+m158_3+m159_3+m160_3+m161_3+m162_3+m163_3+m164_3+m165_3+m166_3+m167_3+m168_3+m169_3+m170_3+m171_3+m172_3+m173_3+m174_3+m175_3+m176_3+m177_3+m178_3+m179_3+m180_3+m181_3+m182_3+m183_3+m184_3+m185_3+m186_3+m187_3+m188_3+m189_3+m190_3+m191_3+m192_3+m193_3+m194_3+m195_3+m196_3+m197_3+m198_3+m199_3+m200_3+m201_3+m202_3+m203_3+m204_3+m205_3+m206_3+m207_3+m208_3+m209_3+m210_3+m211_3+m212_3+m213_3+m214_3+m215_3+m216_3+m217_3+m218_3+m219_3+m220_3+m221_3+m222_3+m223_3+m224_3+m225_3+m226_3+m227_3+m228_3+m229_3+m230_3+m231_3+m232_3+m233_3+m234_3+m235_3+m236_3+m237_3+m238_3+m239_3+m240_3+m241_3+m242_3+m243_3+m244_3+m245_3+m246_3+m247_3+m248_3+m249_3+m250_3+m251_3+m252_3+m253_3+m254_3+m255_3+m256_3+m257_3+m258_3+m259_3+m260_3+m261_3+m262_3+m263_3+b3;
   assign out4 = m1_4+m2_4+m3_4+m4_4+m5_4+m6_4+m7_4+m8_4+m9_4+m10_4+m11_4+m12_4+m13_4+m14_4+m15_4+m16_4+m17_4+m18_4+m19_4+m20_4+m21_4+m22_4+m23_4+m24_4+m25_4+m26_4+m27_4+m28_4+m29_4+m30_4+m31_4+m32_4+m33_4+m34_4+m35_4+m36_4+m37_4+m38_4+m39_4+m40_4+m41_4+m42_4+m43_4+m44_4+m45_4+m46_4+m47_4+m48_4+m49_4+m50_4+m51_4+m52_4+m53_4+m54_4+m55_4+m56_4+m57_4+m58_4+m59_4+m60_4+m61_4+m62_4+m63_4+m64_4+m65_4+m66_4+m67_4+m68_4+m69_4+m70_4+m71_4+m72_4+m73_4+m74_4+m75_4+m76_4+m77_4+m78_4+m79_4+m80_4+m81_4+m82_4+m83_4+m84_4+m85_4+m86_4+m87_4+m88_4+m89_4+m90_4+m91_4+m92_4+m93_4+m94_4+m95_4+m96_4+m97_4+m98_4+m99_4+m100_4+m101_4+m102_4+m103_4+m104_4+m105_4+m106_4+m107_4+m108_4+m109_4+m110_4+m111_4+m112_4+m113_4+m114_4+m115_4+m116_4+m117_4+m118_4+m119_4+m120_4+m121_4+m122_4+m123_4+m124_4+m125_4+m126_4+m127_4+m128_4+m129_4+m130_4+m131_4+m132_4+m133_4+m134_4+m135_4+m136_4+m137_4+m138_4+m139_4+m140_4+m141_4+m142_4+m143_4+m144_4+m145_4+m146_4+m147_4+m148_4+m149_4+m150_4+m151_4+m152_4+m153_4+m154_4+m155_4+m156_4+m157_4+m158_4+m159_4+m160_4+m161_4+m162_4+m163_4+m164_4+m165_4+m166_4+m167_4+m168_4+m169_4+m170_4+m171_4+m172_4+m173_4+m174_4+m175_4+m176_4+m177_4+m178_4+m179_4+m180_4+m181_4+m182_4+m183_4+m184_4+m185_4+m186_4+m187_4+m188_4+m189_4+m190_4+m191_4+m192_4+m193_4+m194_4+m195_4+m196_4+m197_4+m198_4+m199_4+m200_4+m201_4+m202_4+m203_4+m204_4+m205_4+m206_4+m207_4+m208_4+m209_4+m210_4+m211_4+m212_4+m213_4+m214_4+m215_4+m216_4+m217_4+m218_4+m219_4+m220_4+m221_4+m222_4+m223_4+m224_4+m225_4+m226_4+m227_4+m228_4+m229_4+m230_4+m231_4+m232_4+m233_4+m234_4+m235_4+m236_4+m237_4+m238_4+m239_4+m240_4+m241_4+m242_4+m243_4+m244_4+m245_4+m246_4+m247_4+m248_4+m249_4+m250_4+m251_4+m252_4+m253_4+m254_4+m255_4+m256_4+m257_4+m258_4+m259_4+m260_4+m261_4+m262_4+m263_4+b4;
   assign out5 = m1_5+m2_5+m3_5+m4_5+m5_5+m6_5+m7_5+m8_5+m9_5+m10_5+m11_5+m12_5+m13_5+m14_5+m15_5+m16_5+m17_5+m18_5+m19_5+m20_5+m21_5+m22_5+m23_5+m24_5+m25_5+m26_5+m27_5+m28_5+m29_5+m30_5+m31_5+m32_5+m33_5+m34_5+m35_5+m36_5+m37_5+m38_5+m39_5+m40_5+m41_5+m42_5+m43_5+m44_5+m45_5+m46_5+m47_5+m48_5+m49_5+m50_5+m51_5+m52_5+m53_5+m54_5+m55_5+m56_5+m57_5+m58_5+m59_5+m60_5+m61_5+m62_5+m63_5+m64_5+m65_5+m66_5+m67_5+m68_5+m69_5+m70_5+m71_5+m72_5+m73_5+m74_5+m75_5+m76_5+m77_5+m78_5+m79_5+m80_5+m81_5+m82_5+m83_5+m84_5+m85_5+m86_5+m87_5+m88_5+m89_5+m90_5+m91_5+m92_5+m93_5+m94_5+m95_5+m96_5+m97_5+m98_5+m99_5+m100_5+m101_5+m102_5+m103_5+m104_5+m105_5+m106_5+m107_5+m108_5+m109_5+m110_5+m111_5+m112_5+m113_5+m114_5+m115_5+m116_5+m117_5+m118_5+m119_5+m120_5+m121_5+m122_5+m123_5+m124_5+m125_5+m126_5+m127_5+m128_5+m129_5+m130_5+m131_5+m132_5+m133_5+m134_5+m135_5+m136_5+m137_5+m138_5+m139_5+m140_5+m141_5+m142_5+m143_5+m144_5+m145_5+m146_5+m147_5+m148_5+m149_5+m150_5+m151_5+m152_5+m153_5+m154_5+m155_5+m156_5+m157_5+m158_5+m159_5+m160_5+m161_5+m162_5+m163_5+m164_5+m165_5+m166_5+m167_5+m168_5+m169_5+m170_5+m171_5+m172_5+m173_5+m174_5+m175_5+m176_5+m177_5+m178_5+m179_5+m180_5+m181_5+m182_5+m183_5+m184_5+m185_5+m186_5+m187_5+m188_5+m189_5+m190_5+m191_5+m192_5+m193_5+m194_5+m195_5+m196_5+m197_5+m198_5+m199_5+m200_5+m201_5+m202_5+m203_5+m204_5+m205_5+m206_5+m207_5+m208_5+m209_5+m210_5+m211_5+m212_5+m213_5+m214_5+m215_5+m216_5+m217_5+m218_5+m219_5+m220_5+m221_5+m222_5+m223_5+m224_5+m225_5+m226_5+m227_5+m228_5+m229_5+m230_5+m231_5+m232_5+m233_5+m234_5+m235_5+m236_5+m237_5+m238_5+m239_5+m240_5+m241_5+m242_5+m243_5+m244_5+m245_5+m246_5+m247_5+m248_5+m249_5+m250_5+m251_5+m252_5+m253_5+m254_5+m255_5+m256_5+m257_5+m258_5+m259_5+m260_5+m261_5+m262_5+m263_5+b5;
   assign out6 = m1_6+m2_6+m3_6+m4_6+m5_6+m6_6+m7_6+m8_6+m9_6+m10_6+m11_6+m12_6+m13_6+m14_6+m15_6+m16_6+m17_6+m18_6+m19_6+m20_6+m21_6+m22_6+m23_6+m24_6+m25_6+m26_6+m27_6+m28_6+m29_6+m30_6+m31_6+m32_6+m33_6+m34_6+m35_6+m36_6+m37_6+m38_6+m39_6+m40_6+m41_6+m42_6+m43_6+m44_6+m45_6+m46_6+m47_6+m48_6+m49_6+m50_6+m51_6+m52_6+m53_6+m54_6+m55_6+m56_6+m57_6+m58_6+m59_6+m60_6+m61_6+m62_6+m63_6+m64_6+m65_6+m66_6+m67_6+m68_6+m69_6+m70_6+m71_6+m72_6+m73_6+m74_6+m75_6+m76_6+m77_6+m78_6+m79_6+m80_6+m81_6+m82_6+m83_6+m84_6+m85_6+m86_6+m87_6+m88_6+m89_6+m90_6+m91_6+m92_6+m93_6+m94_6+m95_6+m96_6+m97_6+m98_6+m99_6+m100_6+m101_6+m102_6+m103_6+m104_6+m105_6+m106_6+m107_6+m108_6+m109_6+m110_6+m111_6+m112_6+m113_6+m114_6+m115_6+m116_6+m117_6+m118_6+m119_6+m120_6+m121_6+m122_6+m123_6+m124_6+m125_6+m126_6+m127_6+m128_6+m129_6+m130_6+m131_6+m132_6+m133_6+m134_6+m135_6+m136_6+m137_6+m138_6+m139_6+m140_6+m141_6+m142_6+m143_6+m144_6+m145_6+m146_6+m147_6+m148_6+m149_6+m150_6+m151_6+m152_6+m153_6+m154_6+m155_6+m156_6+m157_6+m158_6+m159_6+m160_6+m161_6+m162_6+m163_6+m164_6+m165_6+m166_6+m167_6+m168_6+m169_6+m170_6+m171_6+m172_6+m173_6+m174_6+m175_6+m176_6+m177_6+m178_6+m179_6+m180_6+m181_6+m182_6+m183_6+m184_6+m185_6+m186_6+m187_6+m188_6+m189_6+m190_6+m191_6+m192_6+m193_6+m194_6+m195_6+m196_6+m197_6+m198_6+m199_6+m200_6+m201_6+m202_6+m203_6+m204_6+m205_6+m206_6+m207_6+m208_6+m209_6+m210_6+m211_6+m212_6+m213_6+m214_6+m215_6+m216_6+m217_6+m218_6+m219_6+m220_6+m221_6+m222_6+m223_6+m224_6+m225_6+m226_6+m227_6+m228_6+m229_6+m230_6+m231_6+m232_6+m233_6+m234_6+m235_6+m236_6+m237_6+m238_6+m239_6+m240_6+m241_6+m242_6+m243_6+m244_6+m245_6+m246_6+m247_6+m248_6+m249_6+m250_6+m251_6+m252_6+m253_6+m254_6+m255_6+m256_6+m257_6+m258_6+m259_6+m260_6+m261_6+m262_6+m263_6+b6;
   assign out7 = m1_7+m2_7+m3_7+m4_7+m5_7+m6_7+m7_7+m8_7+m9_7+m10_7+m11_7+m12_7+m13_7+m14_7+m15_7+m16_7+m17_7+m18_7+m19_7+m20_7+m21_7+m22_7+m23_7+m24_7+m25_7+m26_7+m27_7+m28_7+m29_7+m30_7+m31_7+m32_7+m33_7+m34_7+m35_7+m36_7+m37_7+m38_7+m39_7+m40_7+m41_7+m42_7+m43_7+m44_7+m45_7+m46_7+m47_7+m48_7+m49_7+m50_7+m51_7+m52_7+m53_7+m54_7+m55_7+m56_7+m57_7+m58_7+m59_7+m60_7+m61_7+m62_7+m63_7+m64_7+m65_7+m66_7+m67_7+m68_7+m69_7+m70_7+m71_7+m72_7+m73_7+m74_7+m75_7+m76_7+m77_7+m78_7+m79_7+m80_7+m81_7+m82_7+m83_7+m84_7+m85_7+m86_7+m87_7+m88_7+m89_7+m90_7+m91_7+m92_7+m93_7+m94_7+m95_7+m96_7+m97_7+m98_7+m99_7+m100_7+m101_7+m102_7+m103_7+m104_7+m105_7+m106_7+m107_7+m108_7+m109_7+m110_7+m111_7+m112_7+m113_7+m114_7+m115_7+m116_7+m117_7+m118_7+m119_7+m120_7+m121_7+m122_7+m123_7+m124_7+m125_7+m126_7+m127_7+m128_7+m129_7+m130_7+m131_7+m132_7+m133_7+m134_7+m135_7+m136_7+m137_7+m138_7+m139_7+m140_7+m141_7+m142_7+m143_7+m144_7+m145_7+m146_7+m147_7+m148_7+m149_7+m150_7+m151_7+m152_7+m153_7+m154_7+m155_7+m156_7+m157_7+m158_7+m159_7+m160_7+m161_7+m162_7+m163_7+m164_7+m165_7+m166_7+m167_7+m168_7+m169_7+m170_7+m171_7+m172_7+m173_7+m174_7+m175_7+m176_7+m177_7+m178_7+m179_7+m180_7+m181_7+m182_7+m183_7+m184_7+m185_7+m186_7+m187_7+m188_7+m189_7+m190_7+m191_7+m192_7+m193_7+m194_7+m195_7+m196_7+m197_7+m198_7+m199_7+m200_7+m201_7+m202_7+m203_7+m204_7+m205_7+m206_7+m207_7+m208_7+m209_7+m210_7+m211_7+m212_7+m213_7+m214_7+m215_7+m216_7+m217_7+m218_7+m219_7+m220_7+m221_7+m222_7+m223_7+m224_7+m225_7+m226_7+m227_7+m228_7+m229_7+m230_7+m231_7+m232_7+m233_7+m234_7+m235_7+m236_7+m237_7+m238_7+m239_7+m240_7+m241_7+m242_7+m243_7+m244_7+m245_7+m246_7+m247_7+m248_7+m249_7+m250_7+m251_7+m252_7+m253_7+m254_7+m255_7+m256_7+m257_7+m258_7+m259_7+m260_7+m261_7+m262_7+m263_7+b7;
   assign out8 = m1_8+m2_8+m3_8+m4_8+m5_8+m6_8+m7_8+m8_8+m9_8+m10_8+m11_8+m12_8+m13_8+m14_8+m15_8+m16_8+m17_8+m18_8+m19_8+m20_8+m21_8+m22_8+m23_8+m24_8+m25_8+m26_8+m27_8+m28_8+m29_8+m30_8+m31_8+m32_8+m33_8+m34_8+m35_8+m36_8+m37_8+m38_8+m39_8+m40_8+m41_8+m42_8+m43_8+m44_8+m45_8+m46_8+m47_8+m48_8+m49_8+m50_8+m51_8+m52_8+m53_8+m54_8+m55_8+m56_8+m57_8+m58_8+m59_8+m60_8+m61_8+m62_8+m63_8+m64_8+m65_8+m66_8+m67_8+m68_8+m69_8+m70_8+m71_8+m72_8+m73_8+m74_8+m75_8+m76_8+m77_8+m78_8+m79_8+m80_8+m81_8+m82_8+m83_8+m84_8+m85_8+m86_8+m87_8+m88_8+m89_8+m90_8+m91_8+m92_8+m93_8+m94_8+m95_8+m96_8+m97_8+m98_8+m99_8+m100_8+m101_8+m102_8+m103_8+m104_8+m105_8+m106_8+m107_8+m108_8+m109_8+m110_8+m111_8+m112_8+m113_8+m114_8+m115_8+m116_8+m117_8+m118_8+m119_8+m120_8+m121_8+m122_8+m123_8+m124_8+m125_8+m126_8+m127_8+m128_8+m129_8+m130_8+m131_8+m132_8+m133_8+m134_8+m135_8+m136_8+m137_8+m138_8+m139_8+m140_8+m141_8+m142_8+m143_8+m144_8+m145_8+m146_8+m147_8+m148_8+m149_8+m150_8+m151_8+m152_8+m153_8+m154_8+m155_8+m156_8+m157_8+m158_8+m159_8+m160_8+m161_8+m162_8+m163_8+m164_8+m165_8+m166_8+m167_8+m168_8+m169_8+m170_8+m171_8+m172_8+m173_8+m174_8+m175_8+m176_8+m177_8+m178_8+m179_8+m180_8+m181_8+m182_8+m183_8+m184_8+m185_8+m186_8+m187_8+m188_8+m189_8+m190_8+m191_8+m192_8+m193_8+m194_8+m195_8+m196_8+m197_8+m198_8+m199_8+m200_8+m201_8+m202_8+m203_8+m204_8+m205_8+m206_8+m207_8+m208_8+m209_8+m210_8+m211_8+m212_8+m213_8+m214_8+m215_8+m216_8+m217_8+m218_8+m219_8+m220_8+m221_8+m222_8+m223_8+m224_8+m225_8+m226_8+m227_8+m228_8+m229_8+m230_8+m231_8+m232_8+m233_8+m234_8+m235_8+m236_8+m237_8+m238_8+m239_8+m240_8+m241_8+m242_8+m243_8+m244_8+m245_8+m246_8+m247_8+m248_8+m249_8+m250_8+m251_8+m252_8+m253_8+m254_8+m255_8+m256_8+m257_8+m258_8+m259_8+m260_8+m261_8+m262_8+m263_8+b8;
   assign out9 = m1_9+m2_9+m3_9+m4_9+m5_9+m6_9+m7_9+m8_9+m9_9+m10_9+m11_9+m12_9+m13_9+m14_9+m15_9+m16_9+m17_9+m18_9+m19_9+m20_9+m21_9+m22_9+m23_9+m24_9+m25_9+m26_9+m27_9+m28_9+m29_9+m30_9+m31_9+m32_9+m33_9+m34_9+m35_9+m36_9+m37_9+m38_9+m39_9+m40_9+m41_9+m42_9+m43_9+m44_9+m45_9+m46_9+m47_9+m48_9+m49_9+m50_9+m51_9+m52_9+m53_9+m54_9+m55_9+m56_9+m57_9+m58_9+m59_9+m60_9+m61_9+m62_9+m63_9+m64_9+m65_9+m66_9+m67_9+m68_9+m69_9+m70_9+m71_9+m72_9+m73_9+m74_9+m75_9+m76_9+m77_9+m78_9+m79_9+m80_9+m81_9+m82_9+m83_9+m84_9+m85_9+m86_9+m87_9+m88_9+m89_9+m90_9+m91_9+m92_9+m93_9+m94_9+m95_9+m96_9+m97_9+m98_9+m99_9+m100_9+m101_9+m102_9+m103_9+m104_9+m105_9+m106_9+m107_9+m108_9+m109_9+m110_9+m111_9+m112_9+m113_9+m114_9+m115_9+m116_9+m117_9+m118_9+m119_9+m120_9+m121_9+m122_9+m123_9+m124_9+m125_9+m126_9+m127_9+m128_9+m129_9+m130_9+m131_9+m132_9+m133_9+m134_9+m135_9+m136_9+m137_9+m138_9+m139_9+m140_9+m141_9+m142_9+m143_9+m144_9+m145_9+m146_9+m147_9+m148_9+m149_9+m150_9+m151_9+m152_9+m153_9+m154_9+m155_9+m156_9+m157_9+m158_9+m159_9+m160_9+m161_9+m162_9+m163_9+m164_9+m165_9+m166_9+m167_9+m168_9+m169_9+m170_9+m171_9+m172_9+m173_9+m174_9+m175_9+m176_9+m177_9+m178_9+m179_9+m180_9+m181_9+m182_9+m183_9+m184_9+m185_9+m186_9+m187_9+m188_9+m189_9+m190_9+m191_9+m192_9+m193_9+m194_9+m195_9+m196_9+m197_9+m198_9+m199_9+m200_9+m201_9+m202_9+m203_9+m204_9+m205_9+m206_9+m207_9+m208_9+m209_9+m210_9+m211_9+m212_9+m213_9+m214_9+m215_9+m216_9+m217_9+m218_9+m219_9+m220_9+m221_9+m222_9+m223_9+m224_9+m225_9+m226_9+m227_9+m228_9+m229_9+m230_9+m231_9+m232_9+m233_9+m234_9+m235_9+m236_9+m237_9+m238_9+m239_9+m240_9+m241_9+m242_9+m243_9+m244_9+m245_9+m246_9+m247_9+m248_9+m249_9+m250_9+m251_9+m252_9+m253_9+m254_9+m255_9+m256_9+m257_9+m258_9+m259_9+m260_9+m261_9+m262_9+m263_9+b9;
   assign out10 = m1_10+m2_10+m3_10+m4_10+m5_10+m6_10+m7_10+m8_10+m9_10+m10_10+m11_10+m12_10+m13_10+m14_10+m15_10+m16_10+m17_10+m18_10+m19_10+m20_10+m21_10+m22_10+m23_10+m24_10+m25_10+m26_10+m27_10+m28_10+m29_10+m30_10+m31_10+m32_10+m33_10+m34_10+m35_10+m36_10+m37_10+m38_10+m39_10+m40_10+m41_10+m42_10+m43_10+m44_10+m45_10+m46_10+m47_10+m48_10+m49_10+m50_10+m51_10+m52_10+m53_10+m54_10+m55_10+m56_10+m57_10+m58_10+m59_10+m60_10+m61_10+m62_10+m63_10+m64_10+m65_10+m66_10+m67_10+m68_10+m69_10+m70_10+m71_10+m72_10+m73_10+m74_10+m75_10+m76_10+m77_10+m78_10+m79_10+m80_10+m81_10+m82_10+m83_10+m84_10+m85_10+m86_10+m87_10+m88_10+m89_10+m90_10+m91_10+m92_10+m93_10+m94_10+m95_10+m96_10+m97_10+m98_10+m99_10+m100_10+m101_10+m102_10+m103_10+m104_10+m105_10+m106_10+m107_10+m108_10+m109_10+m110_10+m111_10+m112_10+m113_10+m114_10+m115_10+m116_10+m117_10+m118_10+m119_10+m120_10+m121_10+m122_10+m123_10+m124_10+m125_10+m126_10+m127_10+m128_10+m129_10+m130_10+m131_10+m132_10+m133_10+m134_10+m135_10+m136_10+m137_10+m138_10+m139_10+m140_10+m141_10+m142_10+m143_10+m144_10+m145_10+m146_10+m147_10+m148_10+m149_10+m150_10+m151_10+m152_10+m153_10+m154_10+m155_10+m156_10+m157_10+m158_10+m159_10+m160_10+m161_10+m162_10+m163_10+m164_10+m165_10+m166_10+m167_10+m168_10+m169_10+m170_10+m171_10+m172_10+m173_10+m174_10+m175_10+m176_10+m177_10+m178_10+m179_10+m180_10+m181_10+m182_10+m183_10+m184_10+m185_10+m186_10+m187_10+m188_10+m189_10+m190_10+m191_10+m192_10+m193_10+m194_10+m195_10+m196_10+m197_10+m198_10+m199_10+m200_10+m201_10+m202_10+m203_10+m204_10+m205_10+m206_10+m207_10+m208_10+m209_10+m210_10+m211_10+m212_10+m213_10+m214_10+m215_10+m216_10+m217_10+m218_10+m219_10+m220_10+m221_10+m222_10+m223_10+m224_10+m225_10+m226_10+m227_10+m228_10+m229_10+m230_10+m231_10+m232_10+m233_10+m234_10+m235_10+m236_10+m237_10+m238_10+m239_10+m240_10+m241_10+m242_10+m243_10+m244_10+m245_10+m246_10+m247_10+m248_10+m249_10+m250_10+m251_10+m252_10+m253_10+m254_10+m255_10+m256_10+m257_10+m258_10+m259_10+m260_10+m261_10+m262_10+m263_10+b10;
   assign out11 = m1_11+m2_11+m3_11+m4_11+m5_11+m6_11+m7_11+m8_11+m9_11+m10_11+m11_11+m12_11+m13_11+m14_11+m15_11+m16_11+m17_11+m18_11+m19_11+m20_11+m21_11+m22_11+m23_11+m24_11+m25_11+m26_11+m27_11+m28_11+m29_11+m30_11+m31_11+m32_11+m33_11+m34_11+m35_11+m36_11+m37_11+m38_11+m39_11+m40_11+m41_11+m42_11+m43_11+m44_11+m45_11+m46_11+m47_11+m48_11+m49_11+m50_11+m51_11+m52_11+m53_11+m54_11+m55_11+m56_11+m57_11+m58_11+m59_11+m60_11+m61_11+m62_11+m63_11+m64_11+m65_11+m66_11+m67_11+m68_11+m69_11+m70_11+m71_11+m72_11+m73_11+m74_11+m75_11+m76_11+m77_11+m78_11+m79_11+m80_11+m81_11+m82_11+m83_11+m84_11+m85_11+m86_11+m87_11+m88_11+m89_11+m90_11+m91_11+m92_11+m93_11+m94_11+m95_11+m96_11+m97_11+m98_11+m99_11+m100_11+m101_11+m102_11+m103_11+m104_11+m105_11+m106_11+m107_11+m108_11+m109_11+m110_11+m111_11+m112_11+m113_11+m114_11+m115_11+m116_11+m117_11+m118_11+m119_11+m120_11+m121_11+m122_11+m123_11+m124_11+m125_11+m126_11+m127_11+m128_11+m129_11+m130_11+m131_11+m132_11+m133_11+m134_11+m135_11+m136_11+m137_11+m138_11+m139_11+m140_11+m141_11+m142_11+m143_11+m144_11+m145_11+m146_11+m147_11+m148_11+m149_11+m150_11+m151_11+m152_11+m153_11+m154_11+m155_11+m156_11+m157_11+m158_11+m159_11+m160_11+m161_11+m162_11+m163_11+m164_11+m165_11+m166_11+m167_11+m168_11+m169_11+m170_11+m171_11+m172_11+m173_11+m174_11+m175_11+m176_11+m177_11+m178_11+m179_11+m180_11+m181_11+m182_11+m183_11+m184_11+m185_11+m186_11+m187_11+m188_11+m189_11+m190_11+m191_11+m192_11+m193_11+m194_11+m195_11+m196_11+m197_11+m198_11+m199_11+m200_11+m201_11+m202_11+m203_11+m204_11+m205_11+m206_11+m207_11+m208_11+m209_11+m210_11+m211_11+m212_11+m213_11+m214_11+m215_11+m216_11+m217_11+m218_11+m219_11+m220_11+m221_11+m222_11+m223_11+m224_11+m225_11+m226_11+m227_11+m228_11+m229_11+m230_11+m231_11+m232_11+m233_11+m234_11+m235_11+m236_11+m237_11+m238_11+m239_11+m240_11+m241_11+m242_11+m243_11+m244_11+m245_11+m246_11+m247_11+m248_11+m249_11+m250_11+m251_11+m252_11+m253_11+m254_11+m255_11+m256_11+m257_11+m258_11+m259_11+m260_11+m261_11+m262_11+m263_11+b11;
   assign out12 = m1_12+m2_12+m3_12+m4_12+m5_12+m6_12+m7_12+m8_12+m9_12+m10_12+m11_12+m12_12+m13_12+m14_12+m15_12+m16_12+m17_12+m18_12+m19_12+m20_12+m21_12+m22_12+m23_12+m24_12+m25_12+m26_12+m27_12+m28_12+m29_12+m30_12+m31_12+m32_12+m33_12+m34_12+m35_12+m36_12+m37_12+m38_12+m39_12+m40_12+m41_12+m42_12+m43_12+m44_12+m45_12+m46_12+m47_12+m48_12+m49_12+m50_12+m51_12+m52_12+m53_12+m54_12+m55_12+m56_12+m57_12+m58_12+m59_12+m60_12+m61_12+m62_12+m63_12+m64_12+m65_12+m66_12+m67_12+m68_12+m69_12+m70_12+m71_12+m72_12+m73_12+m74_12+m75_12+m76_12+m77_12+m78_12+m79_12+m80_12+m81_12+m82_12+m83_12+m84_12+m85_12+m86_12+m87_12+m88_12+m89_12+m90_12+m91_12+m92_12+m93_12+m94_12+m95_12+m96_12+m97_12+m98_12+m99_12+m100_12+m101_12+m102_12+m103_12+m104_12+m105_12+m106_12+m107_12+m108_12+m109_12+m110_12+m111_12+m112_12+m113_12+m114_12+m115_12+m116_12+m117_12+m118_12+m119_12+m120_12+m121_12+m122_12+m123_12+m124_12+m125_12+m126_12+m127_12+m128_12+m129_12+m130_12+m131_12+m132_12+m133_12+m134_12+m135_12+m136_12+m137_12+m138_12+m139_12+m140_12+m141_12+m142_12+m143_12+m144_12+m145_12+m146_12+m147_12+m148_12+m149_12+m150_12+m151_12+m152_12+m153_12+m154_12+m155_12+m156_12+m157_12+m158_12+m159_12+m160_12+m161_12+m162_12+m163_12+m164_12+m165_12+m166_12+m167_12+m168_12+m169_12+m170_12+m171_12+m172_12+m173_12+m174_12+m175_12+m176_12+m177_12+m178_12+m179_12+m180_12+m181_12+m182_12+m183_12+m184_12+m185_12+m186_12+m187_12+m188_12+m189_12+m190_12+m191_12+m192_12+m193_12+m194_12+m195_12+m196_12+m197_12+m198_12+m199_12+m200_12+m201_12+m202_12+m203_12+m204_12+m205_12+m206_12+m207_12+m208_12+m209_12+m210_12+m211_12+m212_12+m213_12+m214_12+m215_12+m216_12+m217_12+m218_12+m219_12+m220_12+m221_12+m222_12+m223_12+m224_12+m225_12+m226_12+m227_12+m228_12+m229_12+m230_12+m231_12+m232_12+m233_12+m234_12+m235_12+m236_12+m237_12+m238_12+m239_12+m240_12+m241_12+m242_12+m243_12+m244_12+m245_12+m246_12+m247_12+m248_12+m249_12+m250_12+m251_12+m252_12+m253_12+m254_12+m255_12+m256_12+m257_12+m258_12+m259_12+m260_12+m261_12+m262_12+m263_12+b12;
   assign out13 = m1_13+m2_13+m3_13+m4_13+m5_13+m6_13+m7_13+m8_13+m9_13+m10_13+m11_13+m12_13+m13_13+m14_13+m15_13+m16_13+m17_13+m18_13+m19_13+m20_13+m21_13+m22_13+m23_13+m24_13+m25_13+m26_13+m27_13+m28_13+m29_13+m30_13+m31_13+m32_13+m33_13+m34_13+m35_13+m36_13+m37_13+m38_13+m39_13+m40_13+m41_13+m42_13+m43_13+m44_13+m45_13+m46_13+m47_13+m48_13+m49_13+m50_13+m51_13+m52_13+m53_13+m54_13+m55_13+m56_13+m57_13+m58_13+m59_13+m60_13+m61_13+m62_13+m63_13+m64_13+m65_13+m66_13+m67_13+m68_13+m69_13+m70_13+m71_13+m72_13+m73_13+m74_13+m75_13+m76_13+m77_13+m78_13+m79_13+m80_13+m81_13+m82_13+m83_13+m84_13+m85_13+m86_13+m87_13+m88_13+m89_13+m90_13+m91_13+m92_13+m93_13+m94_13+m95_13+m96_13+m97_13+m98_13+m99_13+m100_13+m101_13+m102_13+m103_13+m104_13+m105_13+m106_13+m107_13+m108_13+m109_13+m110_13+m111_13+m112_13+m113_13+m114_13+m115_13+m116_13+m117_13+m118_13+m119_13+m120_13+m121_13+m122_13+m123_13+m124_13+m125_13+m126_13+m127_13+m128_13+m129_13+m130_13+m131_13+m132_13+m133_13+m134_13+m135_13+m136_13+m137_13+m138_13+m139_13+m140_13+m141_13+m142_13+m143_13+m144_13+m145_13+m146_13+m147_13+m148_13+m149_13+m150_13+m151_13+m152_13+m153_13+m154_13+m155_13+m156_13+m157_13+m158_13+m159_13+m160_13+m161_13+m162_13+m163_13+m164_13+m165_13+m166_13+m167_13+m168_13+m169_13+m170_13+m171_13+m172_13+m173_13+m174_13+m175_13+m176_13+m177_13+m178_13+m179_13+m180_13+m181_13+m182_13+m183_13+m184_13+m185_13+m186_13+m187_13+m188_13+m189_13+m190_13+m191_13+m192_13+m193_13+m194_13+m195_13+m196_13+m197_13+m198_13+m199_13+m200_13+m201_13+m202_13+m203_13+m204_13+m205_13+m206_13+m207_13+m208_13+m209_13+m210_13+m211_13+m212_13+m213_13+m214_13+m215_13+m216_13+m217_13+m218_13+m219_13+m220_13+m221_13+m222_13+m223_13+m224_13+m225_13+m226_13+m227_13+m228_13+m229_13+m230_13+m231_13+m232_13+m233_13+m234_13+m235_13+m236_13+m237_13+m238_13+m239_13+m240_13+m241_13+m242_13+m243_13+m244_13+m245_13+m246_13+m247_13+m248_13+m249_13+m250_13+m251_13+m252_13+m253_13+m254_13+m255_13+m256_13+m257_13+m258_13+m259_13+m260_13+m261_13+m262_13+m263_13+b13;
   assign out14 = m1_14+m2_14+m3_14+m4_14+m5_14+m6_14+m7_14+m8_14+m9_14+m10_14+m11_14+m12_14+m13_14+m14_14+m15_14+m16_14+m17_14+m18_14+m19_14+m20_14+m21_14+m22_14+m23_14+m24_14+m25_14+m26_14+m27_14+m28_14+m29_14+m30_14+m31_14+m32_14+m33_14+m34_14+m35_14+m36_14+m37_14+m38_14+m39_14+m40_14+m41_14+m42_14+m43_14+m44_14+m45_14+m46_14+m47_14+m48_14+m49_14+m50_14+m51_14+m52_14+m53_14+m54_14+m55_14+m56_14+m57_14+m58_14+m59_14+m60_14+m61_14+m62_14+m63_14+m64_14+m65_14+m66_14+m67_14+m68_14+m69_14+m70_14+m71_14+m72_14+m73_14+m74_14+m75_14+m76_14+m77_14+m78_14+m79_14+m80_14+m81_14+m82_14+m83_14+m84_14+m85_14+m86_14+m87_14+m88_14+m89_14+m90_14+m91_14+m92_14+m93_14+m94_14+m95_14+m96_14+m97_14+m98_14+m99_14+m100_14+m101_14+m102_14+m103_14+m104_14+m105_14+m106_14+m107_14+m108_14+m109_14+m110_14+m111_14+m112_14+m113_14+m114_14+m115_14+m116_14+m117_14+m118_14+m119_14+m120_14+m121_14+m122_14+m123_14+m124_14+m125_14+m126_14+m127_14+m128_14+m129_14+m130_14+m131_14+m132_14+m133_14+m134_14+m135_14+m136_14+m137_14+m138_14+m139_14+m140_14+m141_14+m142_14+m143_14+m144_14+m145_14+m146_14+m147_14+m148_14+m149_14+m150_14+m151_14+m152_14+m153_14+m154_14+m155_14+m156_14+m157_14+m158_14+m159_14+m160_14+m161_14+m162_14+m163_14+m164_14+m165_14+m166_14+m167_14+m168_14+m169_14+m170_14+m171_14+m172_14+m173_14+m174_14+m175_14+m176_14+m177_14+m178_14+m179_14+m180_14+m181_14+m182_14+m183_14+m184_14+m185_14+m186_14+m187_14+m188_14+m189_14+m190_14+m191_14+m192_14+m193_14+m194_14+m195_14+m196_14+m197_14+m198_14+m199_14+m200_14+m201_14+m202_14+m203_14+m204_14+m205_14+m206_14+m207_14+m208_14+m209_14+m210_14+m211_14+m212_14+m213_14+m214_14+m215_14+m216_14+m217_14+m218_14+m219_14+m220_14+m221_14+m222_14+m223_14+m224_14+m225_14+m226_14+m227_14+m228_14+m229_14+m230_14+m231_14+m232_14+m233_14+m234_14+m235_14+m236_14+m237_14+m238_14+m239_14+m240_14+m241_14+m242_14+m243_14+m244_14+m245_14+m246_14+m247_14+m248_14+m249_14+m250_14+m251_14+m252_14+m253_14+m254_14+m255_14+m256_14+m257_14+m258_14+m259_14+m260_14+m261_14+m262_14+m263_14+b14;
   assign out15 = m1_15+m2_15+m3_15+m4_15+m5_15+m6_15+m7_15+m8_15+m9_15+m10_15+m11_15+m12_15+m13_15+m14_15+m15_15+m16_15+m17_15+m18_15+m19_15+m20_15+m21_15+m22_15+m23_15+m24_15+m25_15+m26_15+m27_15+m28_15+m29_15+m30_15+m31_15+m32_15+m33_15+m34_15+m35_15+m36_15+m37_15+m38_15+m39_15+m40_15+m41_15+m42_15+m43_15+m44_15+m45_15+m46_15+m47_15+m48_15+m49_15+m50_15+m51_15+m52_15+m53_15+m54_15+m55_15+m56_15+m57_15+m58_15+m59_15+m60_15+m61_15+m62_15+m63_15+m64_15+m65_15+m66_15+m67_15+m68_15+m69_15+m70_15+m71_15+m72_15+m73_15+m74_15+m75_15+m76_15+m77_15+m78_15+m79_15+m80_15+m81_15+m82_15+m83_15+m84_15+m85_15+m86_15+m87_15+m88_15+m89_15+m90_15+m91_15+m92_15+m93_15+m94_15+m95_15+m96_15+m97_15+m98_15+m99_15+m100_15+m101_15+m102_15+m103_15+m104_15+m105_15+m106_15+m107_15+m108_15+m109_15+m110_15+m111_15+m112_15+m113_15+m114_15+m115_15+m116_15+m117_15+m118_15+m119_15+m120_15+m121_15+m122_15+m123_15+m124_15+m125_15+m126_15+m127_15+m128_15+m129_15+m130_15+m131_15+m132_15+m133_15+m134_15+m135_15+m136_15+m137_15+m138_15+m139_15+m140_15+m141_15+m142_15+m143_15+m144_15+m145_15+m146_15+m147_15+m148_15+m149_15+m150_15+m151_15+m152_15+m153_15+m154_15+m155_15+m156_15+m157_15+m158_15+m159_15+m160_15+m161_15+m162_15+m163_15+m164_15+m165_15+m166_15+m167_15+m168_15+m169_15+m170_15+m171_15+m172_15+m173_15+m174_15+m175_15+m176_15+m177_15+m178_15+m179_15+m180_15+m181_15+m182_15+m183_15+m184_15+m185_15+m186_15+m187_15+m188_15+m189_15+m190_15+m191_15+m192_15+m193_15+m194_15+m195_15+m196_15+m197_15+m198_15+m199_15+m200_15+m201_15+m202_15+m203_15+m204_15+m205_15+m206_15+m207_15+m208_15+m209_15+m210_15+m211_15+m212_15+m213_15+m214_15+m215_15+m216_15+m217_15+m218_15+m219_15+m220_15+m221_15+m222_15+m223_15+m224_15+m225_15+m226_15+m227_15+m228_15+m229_15+m230_15+m231_15+m232_15+m233_15+m234_15+m235_15+m236_15+m237_15+m238_15+m239_15+m240_15+m241_15+m242_15+m243_15+m244_15+m245_15+m246_15+m247_15+m248_15+m249_15+m250_15+m251_15+m252_15+m253_15+m254_15+m255_15+m256_15+m257_15+m258_15+m259_15+m260_15+m261_15+m262_15+m263_15+b15;
   assign out16 = m1_16+m2_16+m3_16+m4_16+m5_16+m6_16+m7_16+m8_16+m9_16+m10_16+m11_16+m12_16+m13_16+m14_16+m15_16+m16_16+m17_16+m18_16+m19_16+m20_16+m21_16+m22_16+m23_16+m24_16+m25_16+m26_16+m27_16+m28_16+m29_16+m30_16+m31_16+m32_16+m33_16+m34_16+m35_16+m36_16+m37_16+m38_16+m39_16+m40_16+m41_16+m42_16+m43_16+m44_16+m45_16+m46_16+m47_16+m48_16+m49_16+m50_16+m51_16+m52_16+m53_16+m54_16+m55_16+m56_16+m57_16+m58_16+m59_16+m60_16+m61_16+m62_16+m63_16+m64_16+m65_16+m66_16+m67_16+m68_16+m69_16+m70_16+m71_16+m72_16+m73_16+m74_16+m75_16+m76_16+m77_16+m78_16+m79_16+m80_16+m81_16+m82_16+m83_16+m84_16+m85_16+m86_16+m87_16+m88_16+m89_16+m90_16+m91_16+m92_16+m93_16+m94_16+m95_16+m96_16+m97_16+m98_16+m99_16+m100_16+m101_16+m102_16+m103_16+m104_16+m105_16+m106_16+m107_16+m108_16+m109_16+m110_16+m111_16+m112_16+m113_16+m114_16+m115_16+m116_16+m117_16+m118_16+m119_16+m120_16+m121_16+m122_16+m123_16+m124_16+m125_16+m126_16+m127_16+m128_16+m129_16+m130_16+m131_16+m132_16+m133_16+m134_16+m135_16+m136_16+m137_16+m138_16+m139_16+m140_16+m141_16+m142_16+m143_16+m144_16+m145_16+m146_16+m147_16+m148_16+m149_16+m150_16+m151_16+m152_16+m153_16+m154_16+m155_16+m156_16+m157_16+m158_16+m159_16+m160_16+m161_16+m162_16+m163_16+m164_16+m165_16+m166_16+m167_16+m168_16+m169_16+m170_16+m171_16+m172_16+m173_16+m174_16+m175_16+m176_16+m177_16+m178_16+m179_16+m180_16+m181_16+m182_16+m183_16+m184_16+m185_16+m186_16+m187_16+m188_16+m189_16+m190_16+m191_16+m192_16+m193_16+m194_16+m195_16+m196_16+m197_16+m198_16+m199_16+m200_16+m201_16+m202_16+m203_16+m204_16+m205_16+m206_16+m207_16+m208_16+m209_16+m210_16+m211_16+m212_16+m213_16+m214_16+m215_16+m216_16+m217_16+m218_16+m219_16+m220_16+m221_16+m222_16+m223_16+m224_16+m225_16+m226_16+m227_16+m228_16+m229_16+m230_16+m231_16+m232_16+m233_16+m234_16+m235_16+m236_16+m237_16+m238_16+m239_16+m240_16+m241_16+m242_16+m243_16+m244_16+m245_16+m246_16+m247_16+m248_16+m249_16+m250_16+m251_16+m252_16+m253_16+m254_16+m255_16+m256_16+m257_16+m258_16+m259_16+m260_16+m261_16+m262_16+m263_16+b16;
   assign out17 = m1_17+m2_17+m3_17+m4_17+m5_17+m6_17+m7_17+m8_17+m9_17+m10_17+m11_17+m12_17+m13_17+m14_17+m15_17+m16_17+m17_17+m18_17+m19_17+m20_17+m21_17+m22_17+m23_17+m24_17+m25_17+m26_17+m27_17+m28_17+m29_17+m30_17+m31_17+m32_17+m33_17+m34_17+m35_17+m36_17+m37_17+m38_17+m39_17+m40_17+m41_17+m42_17+m43_17+m44_17+m45_17+m46_17+m47_17+m48_17+m49_17+m50_17+m51_17+m52_17+m53_17+m54_17+m55_17+m56_17+m57_17+m58_17+m59_17+m60_17+m61_17+m62_17+m63_17+m64_17+m65_17+m66_17+m67_17+m68_17+m69_17+m70_17+m71_17+m72_17+m73_17+m74_17+m75_17+m76_17+m77_17+m78_17+m79_17+m80_17+m81_17+m82_17+m83_17+m84_17+m85_17+m86_17+m87_17+m88_17+m89_17+m90_17+m91_17+m92_17+m93_17+m94_17+m95_17+m96_17+m97_17+m98_17+m99_17+m100_17+m101_17+m102_17+m103_17+m104_17+m105_17+m106_17+m107_17+m108_17+m109_17+m110_17+m111_17+m112_17+m113_17+m114_17+m115_17+m116_17+m117_17+m118_17+m119_17+m120_17+m121_17+m122_17+m123_17+m124_17+m125_17+m126_17+m127_17+m128_17+m129_17+m130_17+m131_17+m132_17+m133_17+m134_17+m135_17+m136_17+m137_17+m138_17+m139_17+m140_17+m141_17+m142_17+m143_17+m144_17+m145_17+m146_17+m147_17+m148_17+m149_17+m150_17+m151_17+m152_17+m153_17+m154_17+m155_17+m156_17+m157_17+m158_17+m159_17+m160_17+m161_17+m162_17+m163_17+m164_17+m165_17+m166_17+m167_17+m168_17+m169_17+m170_17+m171_17+m172_17+m173_17+m174_17+m175_17+m176_17+m177_17+m178_17+m179_17+m180_17+m181_17+m182_17+m183_17+m184_17+m185_17+m186_17+m187_17+m188_17+m189_17+m190_17+m191_17+m192_17+m193_17+m194_17+m195_17+m196_17+m197_17+m198_17+m199_17+m200_17+m201_17+m202_17+m203_17+m204_17+m205_17+m206_17+m207_17+m208_17+m209_17+m210_17+m211_17+m212_17+m213_17+m214_17+m215_17+m216_17+m217_17+m218_17+m219_17+m220_17+m221_17+m222_17+m223_17+m224_17+m225_17+m226_17+m227_17+m228_17+m229_17+m230_17+m231_17+m232_17+m233_17+m234_17+m235_17+m236_17+m237_17+m238_17+m239_17+m240_17+m241_17+m242_17+m243_17+m244_17+m245_17+m246_17+m247_17+m248_17+m249_17+m250_17+m251_17+m252_17+m253_17+m254_17+m255_17+m256_17+m257_17+m258_17+m259_17+m260_17+m261_17+m262_17+m263_17+b17;
   assign out18 = m1_18+m2_18+m3_18+m4_18+m5_18+m6_18+m7_18+m8_18+m9_18+m10_18+m11_18+m12_18+m13_18+m14_18+m15_18+m16_18+m17_18+m18_18+m19_18+m20_18+m21_18+m22_18+m23_18+m24_18+m25_18+m26_18+m27_18+m28_18+m29_18+m30_18+m31_18+m32_18+m33_18+m34_18+m35_18+m36_18+m37_18+m38_18+m39_18+m40_18+m41_18+m42_18+m43_18+m44_18+m45_18+m46_18+m47_18+m48_18+m49_18+m50_18+m51_18+m52_18+m53_18+m54_18+m55_18+m56_18+m57_18+m58_18+m59_18+m60_18+m61_18+m62_18+m63_18+m64_18+m65_18+m66_18+m67_18+m68_18+m69_18+m70_18+m71_18+m72_18+m73_18+m74_18+m75_18+m76_18+m77_18+m78_18+m79_18+m80_18+m81_18+m82_18+m83_18+m84_18+m85_18+m86_18+m87_18+m88_18+m89_18+m90_18+m91_18+m92_18+m93_18+m94_18+m95_18+m96_18+m97_18+m98_18+m99_18+m100_18+m101_18+m102_18+m103_18+m104_18+m105_18+m106_18+m107_18+m108_18+m109_18+m110_18+m111_18+m112_18+m113_18+m114_18+m115_18+m116_18+m117_18+m118_18+m119_18+m120_18+m121_18+m122_18+m123_18+m124_18+m125_18+m126_18+m127_18+m128_18+m129_18+m130_18+m131_18+m132_18+m133_18+m134_18+m135_18+m136_18+m137_18+m138_18+m139_18+m140_18+m141_18+m142_18+m143_18+m144_18+m145_18+m146_18+m147_18+m148_18+m149_18+m150_18+m151_18+m152_18+m153_18+m154_18+m155_18+m156_18+m157_18+m158_18+m159_18+m160_18+m161_18+m162_18+m163_18+m164_18+m165_18+m166_18+m167_18+m168_18+m169_18+m170_18+m171_18+m172_18+m173_18+m174_18+m175_18+m176_18+m177_18+m178_18+m179_18+m180_18+m181_18+m182_18+m183_18+m184_18+m185_18+m186_18+m187_18+m188_18+m189_18+m190_18+m191_18+m192_18+m193_18+m194_18+m195_18+m196_18+m197_18+m198_18+m199_18+m200_18+m201_18+m202_18+m203_18+m204_18+m205_18+m206_18+m207_18+m208_18+m209_18+m210_18+m211_18+m212_18+m213_18+m214_18+m215_18+m216_18+m217_18+m218_18+m219_18+m220_18+m221_18+m222_18+m223_18+m224_18+m225_18+m226_18+m227_18+m228_18+m229_18+m230_18+m231_18+m232_18+m233_18+m234_18+m235_18+m236_18+m237_18+m238_18+m239_18+m240_18+m241_18+m242_18+m243_18+m244_18+m245_18+m246_18+m247_18+m248_18+m249_18+m250_18+m251_18+m252_18+m253_18+m254_18+m255_18+m256_18+m257_18+m258_18+m259_18+m260_18+m261_18+m262_18+m263_18+b18;
   assign out19 = m1_19+m2_19+m3_19+m4_19+m5_19+m6_19+m7_19+m8_19+m9_19+m10_19+m11_19+m12_19+m13_19+m14_19+m15_19+m16_19+m17_19+m18_19+m19_19+m20_19+m21_19+m22_19+m23_19+m24_19+m25_19+m26_19+m27_19+m28_19+m29_19+m30_19+m31_19+m32_19+m33_19+m34_19+m35_19+m36_19+m37_19+m38_19+m39_19+m40_19+m41_19+m42_19+m43_19+m44_19+m45_19+m46_19+m47_19+m48_19+m49_19+m50_19+m51_19+m52_19+m53_19+m54_19+m55_19+m56_19+m57_19+m58_19+m59_19+m60_19+m61_19+m62_19+m63_19+m64_19+m65_19+m66_19+m67_19+m68_19+m69_19+m70_19+m71_19+m72_19+m73_19+m74_19+m75_19+m76_19+m77_19+m78_19+m79_19+m80_19+m81_19+m82_19+m83_19+m84_19+m85_19+m86_19+m87_19+m88_19+m89_19+m90_19+m91_19+m92_19+m93_19+m94_19+m95_19+m96_19+m97_19+m98_19+m99_19+m100_19+m101_19+m102_19+m103_19+m104_19+m105_19+m106_19+m107_19+m108_19+m109_19+m110_19+m111_19+m112_19+m113_19+m114_19+m115_19+m116_19+m117_19+m118_19+m119_19+m120_19+m121_19+m122_19+m123_19+m124_19+m125_19+m126_19+m127_19+m128_19+m129_19+m130_19+m131_19+m132_19+m133_19+m134_19+m135_19+m136_19+m137_19+m138_19+m139_19+m140_19+m141_19+m142_19+m143_19+m144_19+m145_19+m146_19+m147_19+m148_19+m149_19+m150_19+m151_19+m152_19+m153_19+m154_19+m155_19+m156_19+m157_19+m158_19+m159_19+m160_19+m161_19+m162_19+m163_19+m164_19+m165_19+m166_19+m167_19+m168_19+m169_19+m170_19+m171_19+m172_19+m173_19+m174_19+m175_19+m176_19+m177_19+m178_19+m179_19+m180_19+m181_19+m182_19+m183_19+m184_19+m185_19+m186_19+m187_19+m188_19+m189_19+m190_19+m191_19+m192_19+m193_19+m194_19+m195_19+m196_19+m197_19+m198_19+m199_19+m200_19+m201_19+m202_19+m203_19+m204_19+m205_19+m206_19+m207_19+m208_19+m209_19+m210_19+m211_19+m212_19+m213_19+m214_19+m215_19+m216_19+m217_19+m218_19+m219_19+m220_19+m221_19+m222_19+m223_19+m224_19+m225_19+m226_19+m227_19+m228_19+m229_19+m230_19+m231_19+m232_19+m233_19+m234_19+m235_19+m236_19+m237_19+m238_19+m239_19+m240_19+m241_19+m242_19+m243_19+m244_19+m245_19+m246_19+m247_19+m248_19+m249_19+m250_19+m251_19+m252_19+m253_19+m254_19+m255_19+m256_19+m257_19+m258_19+m259_19+m260_19+m261_19+m262_19+m263_19+b19;
   assign out20 = m1_20+m2_20+m3_20+m4_20+m5_20+m6_20+m7_20+m8_20+m9_20+m10_20+m11_20+m12_20+m13_20+m14_20+m15_20+m16_20+m17_20+m18_20+m19_20+m20_20+m21_20+m22_20+m23_20+m24_20+m25_20+m26_20+m27_20+m28_20+m29_20+m30_20+m31_20+m32_20+m33_20+m34_20+m35_20+m36_20+m37_20+m38_20+m39_20+m40_20+m41_20+m42_20+m43_20+m44_20+m45_20+m46_20+m47_20+m48_20+m49_20+m50_20+m51_20+m52_20+m53_20+m54_20+m55_20+m56_20+m57_20+m58_20+m59_20+m60_20+m61_20+m62_20+m63_20+m64_20+m65_20+m66_20+m67_20+m68_20+m69_20+m70_20+m71_20+m72_20+m73_20+m74_20+m75_20+m76_20+m77_20+m78_20+m79_20+m80_20+m81_20+m82_20+m83_20+m84_20+m85_20+m86_20+m87_20+m88_20+m89_20+m90_20+m91_20+m92_20+m93_20+m94_20+m95_20+m96_20+m97_20+m98_20+m99_20+m100_20+m101_20+m102_20+m103_20+m104_20+m105_20+m106_20+m107_20+m108_20+m109_20+m110_20+m111_20+m112_20+m113_20+m114_20+m115_20+m116_20+m117_20+m118_20+m119_20+m120_20+m121_20+m122_20+m123_20+m124_20+m125_20+m126_20+m127_20+m128_20+m129_20+m130_20+m131_20+m132_20+m133_20+m134_20+m135_20+m136_20+m137_20+m138_20+m139_20+m140_20+m141_20+m142_20+m143_20+m144_20+m145_20+m146_20+m147_20+m148_20+m149_20+m150_20+m151_20+m152_20+m153_20+m154_20+m155_20+m156_20+m157_20+m158_20+m159_20+m160_20+m161_20+m162_20+m163_20+m164_20+m165_20+m166_20+m167_20+m168_20+m169_20+m170_20+m171_20+m172_20+m173_20+m174_20+m175_20+m176_20+m177_20+m178_20+m179_20+m180_20+m181_20+m182_20+m183_20+m184_20+m185_20+m186_20+m187_20+m188_20+m189_20+m190_20+m191_20+m192_20+m193_20+m194_20+m195_20+m196_20+m197_20+m198_20+m199_20+m200_20+m201_20+m202_20+m203_20+m204_20+m205_20+m206_20+m207_20+m208_20+m209_20+m210_20+m211_20+m212_20+m213_20+m214_20+m215_20+m216_20+m217_20+m218_20+m219_20+m220_20+m221_20+m222_20+m223_20+m224_20+m225_20+m226_20+m227_20+m228_20+m229_20+m230_20+m231_20+m232_20+m233_20+m234_20+m235_20+m236_20+m237_20+m238_20+m239_20+m240_20+m241_20+m242_20+m243_20+m244_20+m245_20+m246_20+m247_20+m248_20+m249_20+m250_20+m251_20+m252_20+m253_20+m254_20+m255_20+m256_20+m257_20+m258_20+m259_20+m260_20+m261_20+m262_20+m263_20+b20;
   assign out21 = m1_21+m2_21+m3_21+m4_21+m5_21+m6_21+m7_21+m8_21+m9_21+m10_21+m11_21+m12_21+m13_21+m14_21+m15_21+m16_21+m17_21+m18_21+m19_21+m20_21+m21_21+m22_21+m23_21+m24_21+m25_21+m26_21+m27_21+m28_21+m29_21+m30_21+m31_21+m32_21+m33_21+m34_21+m35_21+m36_21+m37_21+m38_21+m39_21+m40_21+m41_21+m42_21+m43_21+m44_21+m45_21+m46_21+m47_21+m48_21+m49_21+m50_21+m51_21+m52_21+m53_21+m54_21+m55_21+m56_21+m57_21+m58_21+m59_21+m60_21+m61_21+m62_21+m63_21+m64_21+m65_21+m66_21+m67_21+m68_21+m69_21+m70_21+m71_21+m72_21+m73_21+m74_21+m75_21+m76_21+m77_21+m78_21+m79_21+m80_21+m81_21+m82_21+m83_21+m84_21+m85_21+m86_21+m87_21+m88_21+m89_21+m90_21+m91_21+m92_21+m93_21+m94_21+m95_21+m96_21+m97_21+m98_21+m99_21+m100_21+m101_21+m102_21+m103_21+m104_21+m105_21+m106_21+m107_21+m108_21+m109_21+m110_21+m111_21+m112_21+m113_21+m114_21+m115_21+m116_21+m117_21+m118_21+m119_21+m120_21+m121_21+m122_21+m123_21+m124_21+m125_21+m126_21+m127_21+m128_21+m129_21+m130_21+m131_21+m132_21+m133_21+m134_21+m135_21+m136_21+m137_21+m138_21+m139_21+m140_21+m141_21+m142_21+m143_21+m144_21+m145_21+m146_21+m147_21+m148_21+m149_21+m150_21+m151_21+m152_21+m153_21+m154_21+m155_21+m156_21+m157_21+m158_21+m159_21+m160_21+m161_21+m162_21+m163_21+m164_21+m165_21+m166_21+m167_21+m168_21+m169_21+m170_21+m171_21+m172_21+m173_21+m174_21+m175_21+m176_21+m177_21+m178_21+m179_21+m180_21+m181_21+m182_21+m183_21+m184_21+m185_21+m186_21+m187_21+m188_21+m189_21+m190_21+m191_21+m192_21+m193_21+m194_21+m195_21+m196_21+m197_21+m198_21+m199_21+m200_21+m201_21+m202_21+m203_21+m204_21+m205_21+m206_21+m207_21+m208_21+m209_21+m210_21+m211_21+m212_21+m213_21+m214_21+m215_21+m216_21+m217_21+m218_21+m219_21+m220_21+m221_21+m222_21+m223_21+m224_21+m225_21+m226_21+m227_21+m228_21+m229_21+m230_21+m231_21+m232_21+m233_21+m234_21+m235_21+m236_21+m237_21+m238_21+m239_21+m240_21+m241_21+m242_21+m243_21+m244_21+m245_21+m246_21+m247_21+m248_21+m249_21+m250_21+m251_21+m252_21+m253_21+m254_21+m255_21+m256_21+m257_21+m258_21+m259_21+m260_21+m261_21+m262_21+m263_21+b21;
   assign out22 = m1_22+m2_22+m3_22+m4_22+m5_22+m6_22+m7_22+m8_22+m9_22+m10_22+m11_22+m12_22+m13_22+m14_22+m15_22+m16_22+m17_22+m18_22+m19_22+m20_22+m21_22+m22_22+m23_22+m24_22+m25_22+m26_22+m27_22+m28_22+m29_22+m30_22+m31_22+m32_22+m33_22+m34_22+m35_22+m36_22+m37_22+m38_22+m39_22+m40_22+m41_22+m42_22+m43_22+m44_22+m45_22+m46_22+m47_22+m48_22+m49_22+m50_22+m51_22+m52_22+m53_22+m54_22+m55_22+m56_22+m57_22+m58_22+m59_22+m60_22+m61_22+m62_22+m63_22+m64_22+m65_22+m66_22+m67_22+m68_22+m69_22+m70_22+m71_22+m72_22+m73_22+m74_22+m75_22+m76_22+m77_22+m78_22+m79_22+m80_22+m81_22+m82_22+m83_22+m84_22+m85_22+m86_22+m87_22+m88_22+m89_22+m90_22+m91_22+m92_22+m93_22+m94_22+m95_22+m96_22+m97_22+m98_22+m99_22+m100_22+m101_22+m102_22+m103_22+m104_22+m105_22+m106_22+m107_22+m108_22+m109_22+m110_22+m111_22+m112_22+m113_22+m114_22+m115_22+m116_22+m117_22+m118_22+m119_22+m120_22+m121_22+m122_22+m123_22+m124_22+m125_22+m126_22+m127_22+m128_22+m129_22+m130_22+m131_22+m132_22+m133_22+m134_22+m135_22+m136_22+m137_22+m138_22+m139_22+m140_22+m141_22+m142_22+m143_22+m144_22+m145_22+m146_22+m147_22+m148_22+m149_22+m150_22+m151_22+m152_22+m153_22+m154_22+m155_22+m156_22+m157_22+m158_22+m159_22+m160_22+m161_22+m162_22+m163_22+m164_22+m165_22+m166_22+m167_22+m168_22+m169_22+m170_22+m171_22+m172_22+m173_22+m174_22+m175_22+m176_22+m177_22+m178_22+m179_22+m180_22+m181_22+m182_22+m183_22+m184_22+m185_22+m186_22+m187_22+m188_22+m189_22+m190_22+m191_22+m192_22+m193_22+m194_22+m195_22+m196_22+m197_22+m198_22+m199_22+m200_22+m201_22+m202_22+m203_22+m204_22+m205_22+m206_22+m207_22+m208_22+m209_22+m210_22+m211_22+m212_22+m213_22+m214_22+m215_22+m216_22+m217_22+m218_22+m219_22+m220_22+m221_22+m222_22+m223_22+m224_22+m225_22+m226_22+m227_22+m228_22+m229_22+m230_22+m231_22+m232_22+m233_22+m234_22+m235_22+m236_22+m237_22+m238_22+m239_22+m240_22+m241_22+m242_22+m243_22+m244_22+m245_22+m246_22+m247_22+m248_22+m249_22+m250_22+m251_22+m252_22+m253_22+m254_22+m255_22+m256_22+m257_22+m258_22+m259_22+m260_22+m261_22+m262_22+m263_22+b22;
   assign out23 = m1_23+m2_23+m3_23+m4_23+m5_23+m6_23+m7_23+m8_23+m9_23+m10_23+m11_23+m12_23+m13_23+m14_23+m15_23+m16_23+m17_23+m18_23+m19_23+m20_23+m21_23+m22_23+m23_23+m24_23+m25_23+m26_23+m27_23+m28_23+m29_23+m30_23+m31_23+m32_23+m33_23+m34_23+m35_23+m36_23+m37_23+m38_23+m39_23+m40_23+m41_23+m42_23+m43_23+m44_23+m45_23+m46_23+m47_23+m48_23+m49_23+m50_23+m51_23+m52_23+m53_23+m54_23+m55_23+m56_23+m57_23+m58_23+m59_23+m60_23+m61_23+m62_23+m63_23+m64_23+m65_23+m66_23+m67_23+m68_23+m69_23+m70_23+m71_23+m72_23+m73_23+m74_23+m75_23+m76_23+m77_23+m78_23+m79_23+m80_23+m81_23+m82_23+m83_23+m84_23+m85_23+m86_23+m87_23+m88_23+m89_23+m90_23+m91_23+m92_23+m93_23+m94_23+m95_23+m96_23+m97_23+m98_23+m99_23+m100_23+m101_23+m102_23+m103_23+m104_23+m105_23+m106_23+m107_23+m108_23+m109_23+m110_23+m111_23+m112_23+m113_23+m114_23+m115_23+m116_23+m117_23+m118_23+m119_23+m120_23+m121_23+m122_23+m123_23+m124_23+m125_23+m126_23+m127_23+m128_23+m129_23+m130_23+m131_23+m132_23+m133_23+m134_23+m135_23+m136_23+m137_23+m138_23+m139_23+m140_23+m141_23+m142_23+m143_23+m144_23+m145_23+m146_23+m147_23+m148_23+m149_23+m150_23+m151_23+m152_23+m153_23+m154_23+m155_23+m156_23+m157_23+m158_23+m159_23+m160_23+m161_23+m162_23+m163_23+m164_23+m165_23+m166_23+m167_23+m168_23+m169_23+m170_23+m171_23+m172_23+m173_23+m174_23+m175_23+m176_23+m177_23+m178_23+m179_23+m180_23+m181_23+m182_23+m183_23+m184_23+m185_23+m186_23+m187_23+m188_23+m189_23+m190_23+m191_23+m192_23+m193_23+m194_23+m195_23+m196_23+m197_23+m198_23+m199_23+m200_23+m201_23+m202_23+m203_23+m204_23+m205_23+m206_23+m207_23+m208_23+m209_23+m210_23+m211_23+m212_23+m213_23+m214_23+m215_23+m216_23+m217_23+m218_23+m219_23+m220_23+m221_23+m222_23+m223_23+m224_23+m225_23+m226_23+m227_23+m228_23+m229_23+m230_23+m231_23+m232_23+m233_23+m234_23+m235_23+m236_23+m237_23+m238_23+m239_23+m240_23+m241_23+m242_23+m243_23+m244_23+m245_23+m246_23+m247_23+m248_23+m249_23+m250_23+m251_23+m252_23+m253_23+m254_23+m255_23+m256_23+m257_23+m258_23+m259_23+m260_23+m261_23+m262_23+m263_23+b23;
   assign out24 = m1_24+m2_24+m3_24+m4_24+m5_24+m6_24+m7_24+m8_24+m9_24+m10_24+m11_24+m12_24+m13_24+m14_24+m15_24+m16_24+m17_24+m18_24+m19_24+m20_24+m21_24+m22_24+m23_24+m24_24+m25_24+m26_24+m27_24+m28_24+m29_24+m30_24+m31_24+m32_24+m33_24+m34_24+m35_24+m36_24+m37_24+m38_24+m39_24+m40_24+m41_24+m42_24+m43_24+m44_24+m45_24+m46_24+m47_24+m48_24+m49_24+m50_24+m51_24+m52_24+m53_24+m54_24+m55_24+m56_24+m57_24+m58_24+m59_24+m60_24+m61_24+m62_24+m63_24+m64_24+m65_24+m66_24+m67_24+m68_24+m69_24+m70_24+m71_24+m72_24+m73_24+m74_24+m75_24+m76_24+m77_24+m78_24+m79_24+m80_24+m81_24+m82_24+m83_24+m84_24+m85_24+m86_24+m87_24+m88_24+m89_24+m90_24+m91_24+m92_24+m93_24+m94_24+m95_24+m96_24+m97_24+m98_24+m99_24+m100_24+m101_24+m102_24+m103_24+m104_24+m105_24+m106_24+m107_24+m108_24+m109_24+m110_24+m111_24+m112_24+m113_24+m114_24+m115_24+m116_24+m117_24+m118_24+m119_24+m120_24+m121_24+m122_24+m123_24+m124_24+m125_24+m126_24+m127_24+m128_24+m129_24+m130_24+m131_24+m132_24+m133_24+m134_24+m135_24+m136_24+m137_24+m138_24+m139_24+m140_24+m141_24+m142_24+m143_24+m144_24+m145_24+m146_24+m147_24+m148_24+m149_24+m150_24+m151_24+m152_24+m153_24+m154_24+m155_24+m156_24+m157_24+m158_24+m159_24+m160_24+m161_24+m162_24+m163_24+m164_24+m165_24+m166_24+m167_24+m168_24+m169_24+m170_24+m171_24+m172_24+m173_24+m174_24+m175_24+m176_24+m177_24+m178_24+m179_24+m180_24+m181_24+m182_24+m183_24+m184_24+m185_24+m186_24+m187_24+m188_24+m189_24+m190_24+m191_24+m192_24+m193_24+m194_24+m195_24+m196_24+m197_24+m198_24+m199_24+m200_24+m201_24+m202_24+m203_24+m204_24+m205_24+m206_24+m207_24+m208_24+m209_24+m210_24+m211_24+m212_24+m213_24+m214_24+m215_24+m216_24+m217_24+m218_24+m219_24+m220_24+m221_24+m222_24+m223_24+m224_24+m225_24+m226_24+m227_24+m228_24+m229_24+m230_24+m231_24+m232_24+m233_24+m234_24+m235_24+m236_24+m237_24+m238_24+m239_24+m240_24+m241_24+m242_24+m243_24+m244_24+m245_24+m246_24+m247_24+m248_24+m249_24+m250_24+m251_24+m252_24+m253_24+m254_24+m255_24+m256_24+m257_24+m258_24+m259_24+m260_24+m261_24+m262_24+m263_24+b24;
   assign out25 = m1_25+m2_25+m3_25+m4_25+m5_25+m6_25+m7_25+m8_25+m9_25+m10_25+m11_25+m12_25+m13_25+m14_25+m15_25+m16_25+m17_25+m18_25+m19_25+m20_25+m21_25+m22_25+m23_25+m24_25+m25_25+m26_25+m27_25+m28_25+m29_25+m30_25+m31_25+m32_25+m33_25+m34_25+m35_25+m36_25+m37_25+m38_25+m39_25+m40_25+m41_25+m42_25+m43_25+m44_25+m45_25+m46_25+m47_25+m48_25+m49_25+m50_25+m51_25+m52_25+m53_25+m54_25+m55_25+m56_25+m57_25+m58_25+m59_25+m60_25+m61_25+m62_25+m63_25+m64_25+m65_25+m66_25+m67_25+m68_25+m69_25+m70_25+m71_25+m72_25+m73_25+m74_25+m75_25+m76_25+m77_25+m78_25+m79_25+m80_25+m81_25+m82_25+m83_25+m84_25+m85_25+m86_25+m87_25+m88_25+m89_25+m90_25+m91_25+m92_25+m93_25+m94_25+m95_25+m96_25+m97_25+m98_25+m99_25+m100_25+m101_25+m102_25+m103_25+m104_25+m105_25+m106_25+m107_25+m108_25+m109_25+m110_25+m111_25+m112_25+m113_25+m114_25+m115_25+m116_25+m117_25+m118_25+m119_25+m120_25+m121_25+m122_25+m123_25+m124_25+m125_25+m126_25+m127_25+m128_25+m129_25+m130_25+m131_25+m132_25+m133_25+m134_25+m135_25+m136_25+m137_25+m138_25+m139_25+m140_25+m141_25+m142_25+m143_25+m144_25+m145_25+m146_25+m147_25+m148_25+m149_25+m150_25+m151_25+m152_25+m153_25+m154_25+m155_25+m156_25+m157_25+m158_25+m159_25+m160_25+m161_25+m162_25+m163_25+m164_25+m165_25+m166_25+m167_25+m168_25+m169_25+m170_25+m171_25+m172_25+m173_25+m174_25+m175_25+m176_25+m177_25+m178_25+m179_25+m180_25+m181_25+m182_25+m183_25+m184_25+m185_25+m186_25+m187_25+m188_25+m189_25+m190_25+m191_25+m192_25+m193_25+m194_25+m195_25+m196_25+m197_25+m198_25+m199_25+m200_25+m201_25+m202_25+m203_25+m204_25+m205_25+m206_25+m207_25+m208_25+m209_25+m210_25+m211_25+m212_25+m213_25+m214_25+m215_25+m216_25+m217_25+m218_25+m219_25+m220_25+m221_25+m222_25+m223_25+m224_25+m225_25+m226_25+m227_25+m228_25+m229_25+m230_25+m231_25+m232_25+m233_25+m234_25+m235_25+m236_25+m237_25+m238_25+m239_25+m240_25+m241_25+m242_25+m243_25+m244_25+m245_25+m246_25+m247_25+m248_25+m249_25+m250_25+m251_25+m252_25+m253_25+m254_25+m255_25+m256_25+m257_25+m258_25+m259_25+m260_25+m261_25+m262_25+m263_25+b25;
   assign out26 = m1_26+m2_26+m3_26+m4_26+m5_26+m6_26+m7_26+m8_26+m9_26+m10_26+m11_26+m12_26+m13_26+m14_26+m15_26+m16_26+m17_26+m18_26+m19_26+m20_26+m21_26+m22_26+m23_26+m24_26+m25_26+m26_26+m27_26+m28_26+m29_26+m30_26+m31_26+m32_26+m33_26+m34_26+m35_26+m36_26+m37_26+m38_26+m39_26+m40_26+m41_26+m42_26+m43_26+m44_26+m45_26+m46_26+m47_26+m48_26+m49_26+m50_26+m51_26+m52_26+m53_26+m54_26+m55_26+m56_26+m57_26+m58_26+m59_26+m60_26+m61_26+m62_26+m63_26+m64_26+m65_26+m66_26+m67_26+m68_26+m69_26+m70_26+m71_26+m72_26+m73_26+m74_26+m75_26+m76_26+m77_26+m78_26+m79_26+m80_26+m81_26+m82_26+m83_26+m84_26+m85_26+m86_26+m87_26+m88_26+m89_26+m90_26+m91_26+m92_26+m93_26+m94_26+m95_26+m96_26+m97_26+m98_26+m99_26+m100_26+m101_26+m102_26+m103_26+m104_26+m105_26+m106_26+m107_26+m108_26+m109_26+m110_26+m111_26+m112_26+m113_26+m114_26+m115_26+m116_26+m117_26+m118_26+m119_26+m120_26+m121_26+m122_26+m123_26+m124_26+m125_26+m126_26+m127_26+m128_26+m129_26+m130_26+m131_26+m132_26+m133_26+m134_26+m135_26+m136_26+m137_26+m138_26+m139_26+m140_26+m141_26+m142_26+m143_26+m144_26+m145_26+m146_26+m147_26+m148_26+m149_26+m150_26+m151_26+m152_26+m153_26+m154_26+m155_26+m156_26+m157_26+m158_26+m159_26+m160_26+m161_26+m162_26+m163_26+m164_26+m165_26+m166_26+m167_26+m168_26+m169_26+m170_26+m171_26+m172_26+m173_26+m174_26+m175_26+m176_26+m177_26+m178_26+m179_26+m180_26+m181_26+m182_26+m183_26+m184_26+m185_26+m186_26+m187_26+m188_26+m189_26+m190_26+m191_26+m192_26+m193_26+m194_26+m195_26+m196_26+m197_26+m198_26+m199_26+m200_26+m201_26+m202_26+m203_26+m204_26+m205_26+m206_26+m207_26+m208_26+m209_26+m210_26+m211_26+m212_26+m213_26+m214_26+m215_26+m216_26+m217_26+m218_26+m219_26+m220_26+m221_26+m222_26+m223_26+m224_26+m225_26+m226_26+m227_26+m228_26+m229_26+m230_26+m231_26+m232_26+m233_26+m234_26+m235_26+m236_26+m237_26+m238_26+m239_26+m240_26+m241_26+m242_26+m243_26+m244_26+m245_26+m246_26+m247_26+m248_26+m249_26+m250_26+m251_26+m252_26+m253_26+m254_26+m255_26+m256_26+m257_26+m258_26+m259_26+m260_26+m261_26+m262_26+m263_26+b26;
   assign out27 = m1_27+m2_27+m3_27+m4_27+m5_27+m6_27+m7_27+m8_27+m9_27+m10_27+m11_27+m12_27+m13_27+m14_27+m15_27+m16_27+m17_27+m18_27+m19_27+m20_27+m21_27+m22_27+m23_27+m24_27+m25_27+m26_27+m27_27+m28_27+m29_27+m30_27+m31_27+m32_27+m33_27+m34_27+m35_27+m36_27+m37_27+m38_27+m39_27+m40_27+m41_27+m42_27+m43_27+m44_27+m45_27+m46_27+m47_27+m48_27+m49_27+m50_27+m51_27+m52_27+m53_27+m54_27+m55_27+m56_27+m57_27+m58_27+m59_27+m60_27+m61_27+m62_27+m63_27+m64_27+m65_27+m66_27+m67_27+m68_27+m69_27+m70_27+m71_27+m72_27+m73_27+m74_27+m75_27+m76_27+m77_27+m78_27+m79_27+m80_27+m81_27+m82_27+m83_27+m84_27+m85_27+m86_27+m87_27+m88_27+m89_27+m90_27+m91_27+m92_27+m93_27+m94_27+m95_27+m96_27+m97_27+m98_27+m99_27+m100_27+m101_27+m102_27+m103_27+m104_27+m105_27+m106_27+m107_27+m108_27+m109_27+m110_27+m111_27+m112_27+m113_27+m114_27+m115_27+m116_27+m117_27+m118_27+m119_27+m120_27+m121_27+m122_27+m123_27+m124_27+m125_27+m126_27+m127_27+m128_27+m129_27+m130_27+m131_27+m132_27+m133_27+m134_27+m135_27+m136_27+m137_27+m138_27+m139_27+m140_27+m141_27+m142_27+m143_27+m144_27+m145_27+m146_27+m147_27+m148_27+m149_27+m150_27+m151_27+m152_27+m153_27+m154_27+m155_27+m156_27+m157_27+m158_27+m159_27+m160_27+m161_27+m162_27+m163_27+m164_27+m165_27+m166_27+m167_27+m168_27+m169_27+m170_27+m171_27+m172_27+m173_27+m174_27+m175_27+m176_27+m177_27+m178_27+m179_27+m180_27+m181_27+m182_27+m183_27+m184_27+m185_27+m186_27+m187_27+m188_27+m189_27+m190_27+m191_27+m192_27+m193_27+m194_27+m195_27+m196_27+m197_27+m198_27+m199_27+m200_27+m201_27+m202_27+m203_27+m204_27+m205_27+m206_27+m207_27+m208_27+m209_27+m210_27+m211_27+m212_27+m213_27+m214_27+m215_27+m216_27+m217_27+m218_27+m219_27+m220_27+m221_27+m222_27+m223_27+m224_27+m225_27+m226_27+m227_27+m228_27+m229_27+m230_27+m231_27+m232_27+m233_27+m234_27+m235_27+m236_27+m237_27+m238_27+m239_27+m240_27+m241_27+m242_27+m243_27+m244_27+m245_27+m246_27+m247_27+m248_27+m249_27+m250_27+m251_27+m252_27+m253_27+m254_27+m255_27+m256_27+m257_27+m258_27+m259_27+m260_27+m261_27+m262_27+m263_27+b27;
   assign out28 = m1_28+m2_28+m3_28+m4_28+m5_28+m6_28+m7_28+m8_28+m9_28+m10_28+m11_28+m12_28+m13_28+m14_28+m15_28+m16_28+m17_28+m18_28+m19_28+m20_28+m21_28+m22_28+m23_28+m24_28+m25_28+m26_28+m27_28+m28_28+m29_28+m30_28+m31_28+m32_28+m33_28+m34_28+m35_28+m36_28+m37_28+m38_28+m39_28+m40_28+m41_28+m42_28+m43_28+m44_28+m45_28+m46_28+m47_28+m48_28+m49_28+m50_28+m51_28+m52_28+m53_28+m54_28+m55_28+m56_28+m57_28+m58_28+m59_28+m60_28+m61_28+m62_28+m63_28+m64_28+m65_28+m66_28+m67_28+m68_28+m69_28+m70_28+m71_28+m72_28+m73_28+m74_28+m75_28+m76_28+m77_28+m78_28+m79_28+m80_28+m81_28+m82_28+m83_28+m84_28+m85_28+m86_28+m87_28+m88_28+m89_28+m90_28+m91_28+m92_28+m93_28+m94_28+m95_28+m96_28+m97_28+m98_28+m99_28+m100_28+m101_28+m102_28+m103_28+m104_28+m105_28+m106_28+m107_28+m108_28+m109_28+m110_28+m111_28+m112_28+m113_28+m114_28+m115_28+m116_28+m117_28+m118_28+m119_28+m120_28+m121_28+m122_28+m123_28+m124_28+m125_28+m126_28+m127_28+m128_28+m129_28+m130_28+m131_28+m132_28+m133_28+m134_28+m135_28+m136_28+m137_28+m138_28+m139_28+m140_28+m141_28+m142_28+m143_28+m144_28+m145_28+m146_28+m147_28+m148_28+m149_28+m150_28+m151_28+m152_28+m153_28+m154_28+m155_28+m156_28+m157_28+m158_28+m159_28+m160_28+m161_28+m162_28+m163_28+m164_28+m165_28+m166_28+m167_28+m168_28+m169_28+m170_28+m171_28+m172_28+m173_28+m174_28+m175_28+m176_28+m177_28+m178_28+m179_28+m180_28+m181_28+m182_28+m183_28+m184_28+m185_28+m186_28+m187_28+m188_28+m189_28+m190_28+m191_28+m192_28+m193_28+m194_28+m195_28+m196_28+m197_28+m198_28+m199_28+m200_28+m201_28+m202_28+m203_28+m204_28+m205_28+m206_28+m207_28+m208_28+m209_28+m210_28+m211_28+m212_28+m213_28+m214_28+m215_28+m216_28+m217_28+m218_28+m219_28+m220_28+m221_28+m222_28+m223_28+m224_28+m225_28+m226_28+m227_28+m228_28+m229_28+m230_28+m231_28+m232_28+m233_28+m234_28+m235_28+m236_28+m237_28+m238_28+m239_28+m240_28+m241_28+m242_28+m243_28+m244_28+m245_28+m246_28+m247_28+m248_28+m249_28+m250_28+m251_28+m252_28+m253_28+m254_28+m255_28+m256_28+m257_28+m258_28+m259_28+m260_28+m261_28+m262_28+m263_28+b28;
   assign out29 = m1_29+m2_29+m3_29+m4_29+m5_29+m6_29+m7_29+m8_29+m9_29+m10_29+m11_29+m12_29+m13_29+m14_29+m15_29+m16_29+m17_29+m18_29+m19_29+m20_29+m21_29+m22_29+m23_29+m24_29+m25_29+m26_29+m27_29+m28_29+m29_29+m30_29+m31_29+m32_29+m33_29+m34_29+m35_29+m36_29+m37_29+m38_29+m39_29+m40_29+m41_29+m42_29+m43_29+m44_29+m45_29+m46_29+m47_29+m48_29+m49_29+m50_29+m51_29+m52_29+m53_29+m54_29+m55_29+m56_29+m57_29+m58_29+m59_29+m60_29+m61_29+m62_29+m63_29+m64_29+m65_29+m66_29+m67_29+m68_29+m69_29+m70_29+m71_29+m72_29+m73_29+m74_29+m75_29+m76_29+m77_29+m78_29+m79_29+m80_29+m81_29+m82_29+m83_29+m84_29+m85_29+m86_29+m87_29+m88_29+m89_29+m90_29+m91_29+m92_29+m93_29+m94_29+m95_29+m96_29+m97_29+m98_29+m99_29+m100_29+m101_29+m102_29+m103_29+m104_29+m105_29+m106_29+m107_29+m108_29+m109_29+m110_29+m111_29+m112_29+m113_29+m114_29+m115_29+m116_29+m117_29+m118_29+m119_29+m120_29+m121_29+m122_29+m123_29+m124_29+m125_29+m126_29+m127_29+m128_29+m129_29+m130_29+m131_29+m132_29+m133_29+m134_29+m135_29+m136_29+m137_29+m138_29+m139_29+m140_29+m141_29+m142_29+m143_29+m144_29+m145_29+m146_29+m147_29+m148_29+m149_29+m150_29+m151_29+m152_29+m153_29+m154_29+m155_29+m156_29+m157_29+m158_29+m159_29+m160_29+m161_29+m162_29+m163_29+m164_29+m165_29+m166_29+m167_29+m168_29+m169_29+m170_29+m171_29+m172_29+m173_29+m174_29+m175_29+m176_29+m177_29+m178_29+m179_29+m180_29+m181_29+m182_29+m183_29+m184_29+m185_29+m186_29+m187_29+m188_29+m189_29+m190_29+m191_29+m192_29+m193_29+m194_29+m195_29+m196_29+m197_29+m198_29+m199_29+m200_29+m201_29+m202_29+m203_29+m204_29+m205_29+m206_29+m207_29+m208_29+m209_29+m210_29+m211_29+m212_29+m213_29+m214_29+m215_29+m216_29+m217_29+m218_29+m219_29+m220_29+m221_29+m222_29+m223_29+m224_29+m225_29+m226_29+m227_29+m228_29+m229_29+m230_29+m231_29+m232_29+m233_29+m234_29+m235_29+m236_29+m237_29+m238_29+m239_29+m240_29+m241_29+m242_29+m243_29+m244_29+m245_29+m246_29+m247_29+m248_29+m249_29+m250_29+m251_29+m252_29+m253_29+m254_29+m255_29+m256_29+m257_29+m258_29+m259_29+m260_29+m261_29+m262_29+m263_29+b29;
   assign out30 = m1_30+m2_30+m3_30+m4_30+m5_30+m6_30+m7_30+m8_30+m9_30+m10_30+m11_30+m12_30+m13_30+m14_30+m15_30+m16_30+m17_30+m18_30+m19_30+m20_30+m21_30+m22_30+m23_30+m24_30+m25_30+m26_30+m27_30+m28_30+m29_30+m30_30+m31_30+m32_30+m33_30+m34_30+m35_30+m36_30+m37_30+m38_30+m39_30+m40_30+m41_30+m42_30+m43_30+m44_30+m45_30+m46_30+m47_30+m48_30+m49_30+m50_30+m51_30+m52_30+m53_30+m54_30+m55_30+m56_30+m57_30+m58_30+m59_30+m60_30+m61_30+m62_30+m63_30+m64_30+m65_30+m66_30+m67_30+m68_30+m69_30+m70_30+m71_30+m72_30+m73_30+m74_30+m75_30+m76_30+m77_30+m78_30+m79_30+m80_30+m81_30+m82_30+m83_30+m84_30+m85_30+m86_30+m87_30+m88_30+m89_30+m90_30+m91_30+m92_30+m93_30+m94_30+m95_30+m96_30+m97_30+m98_30+m99_30+m100_30+m101_30+m102_30+m103_30+m104_30+m105_30+m106_30+m107_30+m108_30+m109_30+m110_30+m111_30+m112_30+m113_30+m114_30+m115_30+m116_30+m117_30+m118_30+m119_30+m120_30+m121_30+m122_30+m123_30+m124_30+m125_30+m126_30+m127_30+m128_30+m129_30+m130_30+m131_30+m132_30+m133_30+m134_30+m135_30+m136_30+m137_30+m138_30+m139_30+m140_30+m141_30+m142_30+m143_30+m144_30+m145_30+m146_30+m147_30+m148_30+m149_30+m150_30+m151_30+m152_30+m153_30+m154_30+m155_30+m156_30+m157_30+m158_30+m159_30+m160_30+m161_30+m162_30+m163_30+m164_30+m165_30+m166_30+m167_30+m168_30+m169_30+m170_30+m171_30+m172_30+m173_30+m174_30+m175_30+m176_30+m177_30+m178_30+m179_30+m180_30+m181_30+m182_30+m183_30+m184_30+m185_30+m186_30+m187_30+m188_30+m189_30+m190_30+m191_30+m192_30+m193_30+m194_30+m195_30+m196_30+m197_30+m198_30+m199_30+m200_30+m201_30+m202_30+m203_30+m204_30+m205_30+m206_30+m207_30+m208_30+m209_30+m210_30+m211_30+m212_30+m213_30+m214_30+m215_30+m216_30+m217_30+m218_30+m219_30+m220_30+m221_30+m222_30+m223_30+m224_30+m225_30+m226_30+m227_30+m228_30+m229_30+m230_30+m231_30+m232_30+m233_30+m234_30+m235_30+m236_30+m237_30+m238_30+m239_30+m240_30+m241_30+m242_30+m243_30+m244_30+m245_30+m246_30+m247_30+m248_30+m249_30+m250_30+m251_30+m252_30+m253_30+m254_30+m255_30+m256_30+m257_30+m258_30+m259_30+m260_30+m261_30+m262_30+m263_30+b30;
   assign out31 = m1_31+m2_31+m3_31+m4_31+m5_31+m6_31+m7_31+m8_31+m9_31+m10_31+m11_31+m12_31+m13_31+m14_31+m15_31+m16_31+m17_31+m18_31+m19_31+m20_31+m21_31+m22_31+m23_31+m24_31+m25_31+m26_31+m27_31+m28_31+m29_31+m30_31+m31_31+m32_31+m33_31+m34_31+m35_31+m36_31+m37_31+m38_31+m39_31+m40_31+m41_31+m42_31+m43_31+m44_31+m45_31+m46_31+m47_31+m48_31+m49_31+m50_31+m51_31+m52_31+m53_31+m54_31+m55_31+m56_31+m57_31+m58_31+m59_31+m60_31+m61_31+m62_31+m63_31+m64_31+m65_31+m66_31+m67_31+m68_31+m69_31+m70_31+m71_31+m72_31+m73_31+m74_31+m75_31+m76_31+m77_31+m78_31+m79_31+m80_31+m81_31+m82_31+m83_31+m84_31+m85_31+m86_31+m87_31+m88_31+m89_31+m90_31+m91_31+m92_31+m93_31+m94_31+m95_31+m96_31+m97_31+m98_31+m99_31+m100_31+m101_31+m102_31+m103_31+m104_31+m105_31+m106_31+m107_31+m108_31+m109_31+m110_31+m111_31+m112_31+m113_31+m114_31+m115_31+m116_31+m117_31+m118_31+m119_31+m120_31+m121_31+m122_31+m123_31+m124_31+m125_31+m126_31+m127_31+m128_31+m129_31+m130_31+m131_31+m132_31+m133_31+m134_31+m135_31+m136_31+m137_31+m138_31+m139_31+m140_31+m141_31+m142_31+m143_31+m144_31+m145_31+m146_31+m147_31+m148_31+m149_31+m150_31+m151_31+m152_31+m153_31+m154_31+m155_31+m156_31+m157_31+m158_31+m159_31+m160_31+m161_31+m162_31+m163_31+m164_31+m165_31+m166_31+m167_31+m168_31+m169_31+m170_31+m171_31+m172_31+m173_31+m174_31+m175_31+m176_31+m177_31+m178_31+m179_31+m180_31+m181_31+m182_31+m183_31+m184_31+m185_31+m186_31+m187_31+m188_31+m189_31+m190_31+m191_31+m192_31+m193_31+m194_31+m195_31+m196_31+m197_31+m198_31+m199_31+m200_31+m201_31+m202_31+m203_31+m204_31+m205_31+m206_31+m207_31+m208_31+m209_31+m210_31+m211_31+m212_31+m213_31+m214_31+m215_31+m216_31+m217_31+m218_31+m219_31+m220_31+m221_31+m222_31+m223_31+m224_31+m225_31+m226_31+m227_31+m228_31+m229_31+m230_31+m231_31+m232_31+m233_31+m234_31+m235_31+m236_31+m237_31+m238_31+m239_31+m240_31+m241_31+m242_31+m243_31+m244_31+m245_31+m246_31+m247_31+m248_31+m249_31+m250_31+m251_31+m252_31+m253_31+m254_31+m255_31+m256_31+m257_31+m258_31+m259_31+m260_31+m261_31+m262_31+m263_31+b31;
   assign out32 = m1_32+m2_32+m3_32+m4_32+m5_32+m6_32+m7_32+m8_32+m9_32+m10_32+m11_32+m12_32+m13_32+m14_32+m15_32+m16_32+m17_32+m18_32+m19_32+m20_32+m21_32+m22_32+m23_32+m24_32+m25_32+m26_32+m27_32+m28_32+m29_32+m30_32+m31_32+m32_32+m33_32+m34_32+m35_32+m36_32+m37_32+m38_32+m39_32+m40_32+m41_32+m42_32+m43_32+m44_32+m45_32+m46_32+m47_32+m48_32+m49_32+m50_32+m51_32+m52_32+m53_32+m54_32+m55_32+m56_32+m57_32+m58_32+m59_32+m60_32+m61_32+m62_32+m63_32+m64_32+m65_32+m66_32+m67_32+m68_32+m69_32+m70_32+m71_32+m72_32+m73_32+m74_32+m75_32+m76_32+m77_32+m78_32+m79_32+m80_32+m81_32+m82_32+m83_32+m84_32+m85_32+m86_32+m87_32+m88_32+m89_32+m90_32+m91_32+m92_32+m93_32+m94_32+m95_32+m96_32+m97_32+m98_32+m99_32+m100_32+m101_32+m102_32+m103_32+m104_32+m105_32+m106_32+m107_32+m108_32+m109_32+m110_32+m111_32+m112_32+m113_32+m114_32+m115_32+m116_32+m117_32+m118_32+m119_32+m120_32+m121_32+m122_32+m123_32+m124_32+m125_32+m126_32+m127_32+m128_32+m129_32+m130_32+m131_32+m132_32+m133_32+m134_32+m135_32+m136_32+m137_32+m138_32+m139_32+m140_32+m141_32+m142_32+m143_32+m144_32+m145_32+m146_32+m147_32+m148_32+m149_32+m150_32+m151_32+m152_32+m153_32+m154_32+m155_32+m156_32+m157_32+m158_32+m159_32+m160_32+m161_32+m162_32+m163_32+m164_32+m165_32+m166_32+m167_32+m168_32+m169_32+m170_32+m171_32+m172_32+m173_32+m174_32+m175_32+m176_32+m177_32+m178_32+m179_32+m180_32+m181_32+m182_32+m183_32+m184_32+m185_32+m186_32+m187_32+m188_32+m189_32+m190_32+m191_32+m192_32+m193_32+m194_32+m195_32+m196_32+m197_32+m198_32+m199_32+m200_32+m201_32+m202_32+m203_32+m204_32+m205_32+m206_32+m207_32+m208_32+m209_32+m210_32+m211_32+m212_32+m213_32+m214_32+m215_32+m216_32+m217_32+m218_32+m219_32+m220_32+m221_32+m222_32+m223_32+m224_32+m225_32+m226_32+m227_32+m228_32+m229_32+m230_32+m231_32+m232_32+m233_32+m234_32+m235_32+m236_32+m237_32+m238_32+m239_32+m240_32+m241_32+m242_32+m243_32+m244_32+m245_32+m246_32+m247_32+m248_32+m249_32+m250_32+m251_32+m252_32+m253_32+m254_32+m255_32+m256_32+m257_32+m258_32+m259_32+m260_32+m261_32+m262_32+m263_32+b32;
   assign out33 = m1_33+m2_33+m3_33+m4_33+m5_33+m6_33+m7_33+m8_33+m9_33+m10_33+m11_33+m12_33+m13_33+m14_33+m15_33+m16_33+m17_33+m18_33+m19_33+m20_33+m21_33+m22_33+m23_33+m24_33+m25_33+m26_33+m27_33+m28_33+m29_33+m30_33+m31_33+m32_33+m33_33+m34_33+m35_33+m36_33+m37_33+m38_33+m39_33+m40_33+m41_33+m42_33+m43_33+m44_33+m45_33+m46_33+m47_33+m48_33+m49_33+m50_33+m51_33+m52_33+m53_33+m54_33+m55_33+m56_33+m57_33+m58_33+m59_33+m60_33+m61_33+m62_33+m63_33+m64_33+m65_33+m66_33+m67_33+m68_33+m69_33+m70_33+m71_33+m72_33+m73_33+m74_33+m75_33+m76_33+m77_33+m78_33+m79_33+m80_33+m81_33+m82_33+m83_33+m84_33+m85_33+m86_33+m87_33+m88_33+m89_33+m90_33+m91_33+m92_33+m93_33+m94_33+m95_33+m96_33+m97_33+m98_33+m99_33+m100_33+m101_33+m102_33+m103_33+m104_33+m105_33+m106_33+m107_33+m108_33+m109_33+m110_33+m111_33+m112_33+m113_33+m114_33+m115_33+m116_33+m117_33+m118_33+m119_33+m120_33+m121_33+m122_33+m123_33+m124_33+m125_33+m126_33+m127_33+m128_33+m129_33+m130_33+m131_33+m132_33+m133_33+m134_33+m135_33+m136_33+m137_33+m138_33+m139_33+m140_33+m141_33+m142_33+m143_33+m144_33+m145_33+m146_33+m147_33+m148_33+m149_33+m150_33+m151_33+m152_33+m153_33+m154_33+m155_33+m156_33+m157_33+m158_33+m159_33+m160_33+m161_33+m162_33+m163_33+m164_33+m165_33+m166_33+m167_33+m168_33+m169_33+m170_33+m171_33+m172_33+m173_33+m174_33+m175_33+m176_33+m177_33+m178_33+m179_33+m180_33+m181_33+m182_33+m183_33+m184_33+m185_33+m186_33+m187_33+m188_33+m189_33+m190_33+m191_33+m192_33+m193_33+m194_33+m195_33+m196_33+m197_33+m198_33+m199_33+m200_33+m201_33+m202_33+m203_33+m204_33+m205_33+m206_33+m207_33+m208_33+m209_33+m210_33+m211_33+m212_33+m213_33+m214_33+m215_33+m216_33+m217_33+m218_33+m219_33+m220_33+m221_33+m222_33+m223_33+m224_33+m225_33+m226_33+m227_33+m228_33+m229_33+m230_33+m231_33+m232_33+m233_33+m234_33+m235_33+m236_33+m237_33+m238_33+m239_33+m240_33+m241_33+m242_33+m243_33+m244_33+m245_33+m246_33+m247_33+m248_33+m249_33+m250_33+m251_33+m252_33+m253_33+m254_33+m255_33+m256_33+m257_33+m258_33+m259_33+m260_33+m261_33+m262_33+m263_33+b33;
   assign out34 = m1_34+m2_34+m3_34+m4_34+m5_34+m6_34+m7_34+m8_34+m9_34+m10_34+m11_34+m12_34+m13_34+m14_34+m15_34+m16_34+m17_34+m18_34+m19_34+m20_34+m21_34+m22_34+m23_34+m24_34+m25_34+m26_34+m27_34+m28_34+m29_34+m30_34+m31_34+m32_34+m33_34+m34_34+m35_34+m36_34+m37_34+m38_34+m39_34+m40_34+m41_34+m42_34+m43_34+m44_34+m45_34+m46_34+m47_34+m48_34+m49_34+m50_34+m51_34+m52_34+m53_34+m54_34+m55_34+m56_34+m57_34+m58_34+m59_34+m60_34+m61_34+m62_34+m63_34+m64_34+m65_34+m66_34+m67_34+m68_34+m69_34+m70_34+m71_34+m72_34+m73_34+m74_34+m75_34+m76_34+m77_34+m78_34+m79_34+m80_34+m81_34+m82_34+m83_34+m84_34+m85_34+m86_34+m87_34+m88_34+m89_34+m90_34+m91_34+m92_34+m93_34+m94_34+m95_34+m96_34+m97_34+m98_34+m99_34+m100_34+m101_34+m102_34+m103_34+m104_34+m105_34+m106_34+m107_34+m108_34+m109_34+m110_34+m111_34+m112_34+m113_34+m114_34+m115_34+m116_34+m117_34+m118_34+m119_34+m120_34+m121_34+m122_34+m123_34+m124_34+m125_34+m126_34+m127_34+m128_34+m129_34+m130_34+m131_34+m132_34+m133_34+m134_34+m135_34+m136_34+m137_34+m138_34+m139_34+m140_34+m141_34+m142_34+m143_34+m144_34+m145_34+m146_34+m147_34+m148_34+m149_34+m150_34+m151_34+m152_34+m153_34+m154_34+m155_34+m156_34+m157_34+m158_34+m159_34+m160_34+m161_34+m162_34+m163_34+m164_34+m165_34+m166_34+m167_34+m168_34+m169_34+m170_34+m171_34+m172_34+m173_34+m174_34+m175_34+m176_34+m177_34+m178_34+m179_34+m180_34+m181_34+m182_34+m183_34+m184_34+m185_34+m186_34+m187_34+m188_34+m189_34+m190_34+m191_34+m192_34+m193_34+m194_34+m195_34+m196_34+m197_34+m198_34+m199_34+m200_34+m201_34+m202_34+m203_34+m204_34+m205_34+m206_34+m207_34+m208_34+m209_34+m210_34+m211_34+m212_34+m213_34+m214_34+m215_34+m216_34+m217_34+m218_34+m219_34+m220_34+m221_34+m222_34+m223_34+m224_34+m225_34+m226_34+m227_34+m228_34+m229_34+m230_34+m231_34+m232_34+m233_34+m234_34+m235_34+m236_34+m237_34+m238_34+m239_34+m240_34+m241_34+m242_34+m243_34+m244_34+m245_34+m246_34+m247_34+m248_34+m249_34+m250_34+m251_34+m252_34+m253_34+m254_34+m255_34+m256_34+m257_34+m258_34+m259_34+m260_34+m261_34+m262_34+m263_34+b34;
   assign out35 = m1_35+m2_35+m3_35+m4_35+m5_35+m6_35+m7_35+m8_35+m9_35+m10_35+m11_35+m12_35+m13_35+m14_35+m15_35+m16_35+m17_35+m18_35+m19_35+m20_35+m21_35+m22_35+m23_35+m24_35+m25_35+m26_35+m27_35+m28_35+m29_35+m30_35+m31_35+m32_35+m33_35+m34_35+m35_35+m36_35+m37_35+m38_35+m39_35+m40_35+m41_35+m42_35+m43_35+m44_35+m45_35+m46_35+m47_35+m48_35+m49_35+m50_35+m51_35+m52_35+m53_35+m54_35+m55_35+m56_35+m57_35+m58_35+m59_35+m60_35+m61_35+m62_35+m63_35+m64_35+m65_35+m66_35+m67_35+m68_35+m69_35+m70_35+m71_35+m72_35+m73_35+m74_35+m75_35+m76_35+m77_35+m78_35+m79_35+m80_35+m81_35+m82_35+m83_35+m84_35+m85_35+m86_35+m87_35+m88_35+m89_35+m90_35+m91_35+m92_35+m93_35+m94_35+m95_35+m96_35+m97_35+m98_35+m99_35+m100_35+m101_35+m102_35+m103_35+m104_35+m105_35+m106_35+m107_35+m108_35+m109_35+m110_35+m111_35+m112_35+m113_35+m114_35+m115_35+m116_35+m117_35+m118_35+m119_35+m120_35+m121_35+m122_35+m123_35+m124_35+m125_35+m126_35+m127_35+m128_35+m129_35+m130_35+m131_35+m132_35+m133_35+m134_35+m135_35+m136_35+m137_35+m138_35+m139_35+m140_35+m141_35+m142_35+m143_35+m144_35+m145_35+m146_35+m147_35+m148_35+m149_35+m150_35+m151_35+m152_35+m153_35+m154_35+m155_35+m156_35+m157_35+m158_35+m159_35+m160_35+m161_35+m162_35+m163_35+m164_35+m165_35+m166_35+m167_35+m168_35+m169_35+m170_35+m171_35+m172_35+m173_35+m174_35+m175_35+m176_35+m177_35+m178_35+m179_35+m180_35+m181_35+m182_35+m183_35+m184_35+m185_35+m186_35+m187_35+m188_35+m189_35+m190_35+m191_35+m192_35+m193_35+m194_35+m195_35+m196_35+m197_35+m198_35+m199_35+m200_35+m201_35+m202_35+m203_35+m204_35+m205_35+m206_35+m207_35+m208_35+m209_35+m210_35+m211_35+m212_35+m213_35+m214_35+m215_35+m216_35+m217_35+m218_35+m219_35+m220_35+m221_35+m222_35+m223_35+m224_35+m225_35+m226_35+m227_35+m228_35+m229_35+m230_35+m231_35+m232_35+m233_35+m234_35+m235_35+m236_35+m237_35+m238_35+m239_35+m240_35+m241_35+m242_35+m243_35+m244_35+m245_35+m246_35+m247_35+m248_35+m249_35+m250_35+m251_35+m252_35+m253_35+m254_35+m255_35+m256_35+m257_35+m258_35+m259_35+m260_35+m261_35+m262_35+m263_35+b35;
   assign out36 = m1_36+m2_36+m3_36+m4_36+m5_36+m6_36+m7_36+m8_36+m9_36+m10_36+m11_36+m12_36+m13_36+m14_36+m15_36+m16_36+m17_36+m18_36+m19_36+m20_36+m21_36+m22_36+m23_36+m24_36+m25_36+m26_36+m27_36+m28_36+m29_36+m30_36+m31_36+m32_36+m33_36+m34_36+m35_36+m36_36+m37_36+m38_36+m39_36+m40_36+m41_36+m42_36+m43_36+m44_36+m45_36+m46_36+m47_36+m48_36+m49_36+m50_36+m51_36+m52_36+m53_36+m54_36+m55_36+m56_36+m57_36+m58_36+m59_36+m60_36+m61_36+m62_36+m63_36+m64_36+m65_36+m66_36+m67_36+m68_36+m69_36+m70_36+m71_36+m72_36+m73_36+m74_36+m75_36+m76_36+m77_36+m78_36+m79_36+m80_36+m81_36+m82_36+m83_36+m84_36+m85_36+m86_36+m87_36+m88_36+m89_36+m90_36+m91_36+m92_36+m93_36+m94_36+m95_36+m96_36+m97_36+m98_36+m99_36+m100_36+m101_36+m102_36+m103_36+m104_36+m105_36+m106_36+m107_36+m108_36+m109_36+m110_36+m111_36+m112_36+m113_36+m114_36+m115_36+m116_36+m117_36+m118_36+m119_36+m120_36+m121_36+m122_36+m123_36+m124_36+m125_36+m126_36+m127_36+m128_36+m129_36+m130_36+m131_36+m132_36+m133_36+m134_36+m135_36+m136_36+m137_36+m138_36+m139_36+m140_36+m141_36+m142_36+m143_36+m144_36+m145_36+m146_36+m147_36+m148_36+m149_36+m150_36+m151_36+m152_36+m153_36+m154_36+m155_36+m156_36+m157_36+m158_36+m159_36+m160_36+m161_36+m162_36+m163_36+m164_36+m165_36+m166_36+m167_36+m168_36+m169_36+m170_36+m171_36+m172_36+m173_36+m174_36+m175_36+m176_36+m177_36+m178_36+m179_36+m180_36+m181_36+m182_36+m183_36+m184_36+m185_36+m186_36+m187_36+m188_36+m189_36+m190_36+m191_36+m192_36+m193_36+m194_36+m195_36+m196_36+m197_36+m198_36+m199_36+m200_36+m201_36+m202_36+m203_36+m204_36+m205_36+m206_36+m207_36+m208_36+m209_36+m210_36+m211_36+m212_36+m213_36+m214_36+m215_36+m216_36+m217_36+m218_36+m219_36+m220_36+m221_36+m222_36+m223_36+m224_36+m225_36+m226_36+m227_36+m228_36+m229_36+m230_36+m231_36+m232_36+m233_36+m234_36+m235_36+m236_36+m237_36+m238_36+m239_36+m240_36+m241_36+m242_36+m243_36+m244_36+m245_36+m246_36+m247_36+m248_36+m249_36+m250_36+m251_36+m252_36+m253_36+m254_36+m255_36+m256_36+m257_36+m258_36+m259_36+m260_36+m261_36+m262_36+m263_36+b36;
   assign out37 = m1_37+m2_37+m3_37+m4_37+m5_37+m6_37+m7_37+m8_37+m9_37+m10_37+m11_37+m12_37+m13_37+m14_37+m15_37+m16_37+m17_37+m18_37+m19_37+m20_37+m21_37+m22_37+m23_37+m24_37+m25_37+m26_37+m27_37+m28_37+m29_37+m30_37+m31_37+m32_37+m33_37+m34_37+m35_37+m36_37+m37_37+m38_37+m39_37+m40_37+m41_37+m42_37+m43_37+m44_37+m45_37+m46_37+m47_37+m48_37+m49_37+m50_37+m51_37+m52_37+m53_37+m54_37+m55_37+m56_37+m57_37+m58_37+m59_37+m60_37+m61_37+m62_37+m63_37+m64_37+m65_37+m66_37+m67_37+m68_37+m69_37+m70_37+m71_37+m72_37+m73_37+m74_37+m75_37+m76_37+m77_37+m78_37+m79_37+m80_37+m81_37+m82_37+m83_37+m84_37+m85_37+m86_37+m87_37+m88_37+m89_37+m90_37+m91_37+m92_37+m93_37+m94_37+m95_37+m96_37+m97_37+m98_37+m99_37+m100_37+m101_37+m102_37+m103_37+m104_37+m105_37+m106_37+m107_37+m108_37+m109_37+m110_37+m111_37+m112_37+m113_37+m114_37+m115_37+m116_37+m117_37+m118_37+m119_37+m120_37+m121_37+m122_37+m123_37+m124_37+m125_37+m126_37+m127_37+m128_37+m129_37+m130_37+m131_37+m132_37+m133_37+m134_37+m135_37+m136_37+m137_37+m138_37+m139_37+m140_37+m141_37+m142_37+m143_37+m144_37+m145_37+m146_37+m147_37+m148_37+m149_37+m150_37+m151_37+m152_37+m153_37+m154_37+m155_37+m156_37+m157_37+m158_37+m159_37+m160_37+m161_37+m162_37+m163_37+m164_37+m165_37+m166_37+m167_37+m168_37+m169_37+m170_37+m171_37+m172_37+m173_37+m174_37+m175_37+m176_37+m177_37+m178_37+m179_37+m180_37+m181_37+m182_37+m183_37+m184_37+m185_37+m186_37+m187_37+m188_37+m189_37+m190_37+m191_37+m192_37+m193_37+m194_37+m195_37+m196_37+m197_37+m198_37+m199_37+m200_37+m201_37+m202_37+m203_37+m204_37+m205_37+m206_37+m207_37+m208_37+m209_37+m210_37+m211_37+m212_37+m213_37+m214_37+m215_37+m216_37+m217_37+m218_37+m219_37+m220_37+m221_37+m222_37+m223_37+m224_37+m225_37+m226_37+m227_37+m228_37+m229_37+m230_37+m231_37+m232_37+m233_37+m234_37+m235_37+m236_37+m237_37+m238_37+m239_37+m240_37+m241_37+m242_37+m243_37+m244_37+m245_37+m246_37+m247_37+m248_37+m249_37+m250_37+m251_37+m252_37+m253_37+m254_37+m255_37+m256_37+m257_37+m258_37+m259_37+m260_37+m261_37+m262_37+m263_37+b37;
   assign out38 = m1_38+m2_38+m3_38+m4_38+m5_38+m6_38+m7_38+m8_38+m9_38+m10_38+m11_38+m12_38+m13_38+m14_38+m15_38+m16_38+m17_38+m18_38+m19_38+m20_38+m21_38+m22_38+m23_38+m24_38+m25_38+m26_38+m27_38+m28_38+m29_38+m30_38+m31_38+m32_38+m33_38+m34_38+m35_38+m36_38+m37_38+m38_38+m39_38+m40_38+m41_38+m42_38+m43_38+m44_38+m45_38+m46_38+m47_38+m48_38+m49_38+m50_38+m51_38+m52_38+m53_38+m54_38+m55_38+m56_38+m57_38+m58_38+m59_38+m60_38+m61_38+m62_38+m63_38+m64_38+m65_38+m66_38+m67_38+m68_38+m69_38+m70_38+m71_38+m72_38+m73_38+m74_38+m75_38+m76_38+m77_38+m78_38+m79_38+m80_38+m81_38+m82_38+m83_38+m84_38+m85_38+m86_38+m87_38+m88_38+m89_38+m90_38+m91_38+m92_38+m93_38+m94_38+m95_38+m96_38+m97_38+m98_38+m99_38+m100_38+m101_38+m102_38+m103_38+m104_38+m105_38+m106_38+m107_38+m108_38+m109_38+m110_38+m111_38+m112_38+m113_38+m114_38+m115_38+m116_38+m117_38+m118_38+m119_38+m120_38+m121_38+m122_38+m123_38+m124_38+m125_38+m126_38+m127_38+m128_38+m129_38+m130_38+m131_38+m132_38+m133_38+m134_38+m135_38+m136_38+m137_38+m138_38+m139_38+m140_38+m141_38+m142_38+m143_38+m144_38+m145_38+m146_38+m147_38+m148_38+m149_38+m150_38+m151_38+m152_38+m153_38+m154_38+m155_38+m156_38+m157_38+m158_38+m159_38+m160_38+m161_38+m162_38+m163_38+m164_38+m165_38+m166_38+m167_38+m168_38+m169_38+m170_38+m171_38+m172_38+m173_38+m174_38+m175_38+m176_38+m177_38+m178_38+m179_38+m180_38+m181_38+m182_38+m183_38+m184_38+m185_38+m186_38+m187_38+m188_38+m189_38+m190_38+m191_38+m192_38+m193_38+m194_38+m195_38+m196_38+m197_38+m198_38+m199_38+m200_38+m201_38+m202_38+m203_38+m204_38+m205_38+m206_38+m207_38+m208_38+m209_38+m210_38+m211_38+m212_38+m213_38+m214_38+m215_38+m216_38+m217_38+m218_38+m219_38+m220_38+m221_38+m222_38+m223_38+m224_38+m225_38+m226_38+m227_38+m228_38+m229_38+m230_38+m231_38+m232_38+m233_38+m234_38+m235_38+m236_38+m237_38+m238_38+m239_38+m240_38+m241_38+m242_38+m243_38+m244_38+m245_38+m246_38+m247_38+m248_38+m249_38+m250_38+m251_38+m252_38+m253_38+m254_38+m255_38+m256_38+m257_38+m258_38+m259_38+m260_38+m261_38+m262_38+m263_38+b38;
   assign out39 = m1_39+m2_39+m3_39+m4_39+m5_39+m6_39+m7_39+m8_39+m9_39+m10_39+m11_39+m12_39+m13_39+m14_39+m15_39+m16_39+m17_39+m18_39+m19_39+m20_39+m21_39+m22_39+m23_39+m24_39+m25_39+m26_39+m27_39+m28_39+m29_39+m30_39+m31_39+m32_39+m33_39+m34_39+m35_39+m36_39+m37_39+m38_39+m39_39+m40_39+m41_39+m42_39+m43_39+m44_39+m45_39+m46_39+m47_39+m48_39+m49_39+m50_39+m51_39+m52_39+m53_39+m54_39+m55_39+m56_39+m57_39+m58_39+m59_39+m60_39+m61_39+m62_39+m63_39+m64_39+m65_39+m66_39+m67_39+m68_39+m69_39+m70_39+m71_39+m72_39+m73_39+m74_39+m75_39+m76_39+m77_39+m78_39+m79_39+m80_39+m81_39+m82_39+m83_39+m84_39+m85_39+m86_39+m87_39+m88_39+m89_39+m90_39+m91_39+m92_39+m93_39+m94_39+m95_39+m96_39+m97_39+m98_39+m99_39+m100_39+m101_39+m102_39+m103_39+m104_39+m105_39+m106_39+m107_39+m108_39+m109_39+m110_39+m111_39+m112_39+m113_39+m114_39+m115_39+m116_39+m117_39+m118_39+m119_39+m120_39+m121_39+m122_39+m123_39+m124_39+m125_39+m126_39+m127_39+m128_39+m129_39+m130_39+m131_39+m132_39+m133_39+m134_39+m135_39+m136_39+m137_39+m138_39+m139_39+m140_39+m141_39+m142_39+m143_39+m144_39+m145_39+m146_39+m147_39+m148_39+m149_39+m150_39+m151_39+m152_39+m153_39+m154_39+m155_39+m156_39+m157_39+m158_39+m159_39+m160_39+m161_39+m162_39+m163_39+m164_39+m165_39+m166_39+m167_39+m168_39+m169_39+m170_39+m171_39+m172_39+m173_39+m174_39+m175_39+m176_39+m177_39+m178_39+m179_39+m180_39+m181_39+m182_39+m183_39+m184_39+m185_39+m186_39+m187_39+m188_39+m189_39+m190_39+m191_39+m192_39+m193_39+m194_39+m195_39+m196_39+m197_39+m198_39+m199_39+m200_39+m201_39+m202_39+m203_39+m204_39+m205_39+m206_39+m207_39+m208_39+m209_39+m210_39+m211_39+m212_39+m213_39+m214_39+m215_39+m216_39+m217_39+m218_39+m219_39+m220_39+m221_39+m222_39+m223_39+m224_39+m225_39+m226_39+m227_39+m228_39+m229_39+m230_39+m231_39+m232_39+m233_39+m234_39+m235_39+m236_39+m237_39+m238_39+m239_39+m240_39+m241_39+m242_39+m243_39+m244_39+m245_39+m246_39+m247_39+m248_39+m249_39+m250_39+m251_39+m252_39+m253_39+m254_39+m255_39+m256_39+m257_39+m258_39+m259_39+m260_39+m261_39+m262_39+m263_39+b39;
   assign out40 = m1_40+m2_40+m3_40+m4_40+m5_40+m6_40+m7_40+m8_40+m9_40+m10_40+m11_40+m12_40+m13_40+m14_40+m15_40+m16_40+m17_40+m18_40+m19_40+m20_40+m21_40+m22_40+m23_40+m24_40+m25_40+m26_40+m27_40+m28_40+m29_40+m30_40+m31_40+m32_40+m33_40+m34_40+m35_40+m36_40+m37_40+m38_40+m39_40+m40_40+m41_40+m42_40+m43_40+m44_40+m45_40+m46_40+m47_40+m48_40+m49_40+m50_40+m51_40+m52_40+m53_40+m54_40+m55_40+m56_40+m57_40+m58_40+m59_40+m60_40+m61_40+m62_40+m63_40+m64_40+m65_40+m66_40+m67_40+m68_40+m69_40+m70_40+m71_40+m72_40+m73_40+m74_40+m75_40+m76_40+m77_40+m78_40+m79_40+m80_40+m81_40+m82_40+m83_40+m84_40+m85_40+m86_40+m87_40+m88_40+m89_40+m90_40+m91_40+m92_40+m93_40+m94_40+m95_40+m96_40+m97_40+m98_40+m99_40+m100_40+m101_40+m102_40+m103_40+m104_40+m105_40+m106_40+m107_40+m108_40+m109_40+m110_40+m111_40+m112_40+m113_40+m114_40+m115_40+m116_40+m117_40+m118_40+m119_40+m120_40+m121_40+m122_40+m123_40+m124_40+m125_40+m126_40+m127_40+m128_40+m129_40+m130_40+m131_40+m132_40+m133_40+m134_40+m135_40+m136_40+m137_40+m138_40+m139_40+m140_40+m141_40+m142_40+m143_40+m144_40+m145_40+m146_40+m147_40+m148_40+m149_40+m150_40+m151_40+m152_40+m153_40+m154_40+m155_40+m156_40+m157_40+m158_40+m159_40+m160_40+m161_40+m162_40+m163_40+m164_40+m165_40+m166_40+m167_40+m168_40+m169_40+m170_40+m171_40+m172_40+m173_40+m174_40+m175_40+m176_40+m177_40+m178_40+m179_40+m180_40+m181_40+m182_40+m183_40+m184_40+m185_40+m186_40+m187_40+m188_40+m189_40+m190_40+m191_40+m192_40+m193_40+m194_40+m195_40+m196_40+m197_40+m198_40+m199_40+m200_40+m201_40+m202_40+m203_40+m204_40+m205_40+m206_40+m207_40+m208_40+m209_40+m210_40+m211_40+m212_40+m213_40+m214_40+m215_40+m216_40+m217_40+m218_40+m219_40+m220_40+m221_40+m222_40+m223_40+m224_40+m225_40+m226_40+m227_40+m228_40+m229_40+m230_40+m231_40+m232_40+m233_40+m234_40+m235_40+m236_40+m237_40+m238_40+m239_40+m240_40+m241_40+m242_40+m243_40+m244_40+m245_40+m246_40+m247_40+m248_40+m249_40+m250_40+m251_40+m252_40+m253_40+m254_40+m255_40+m256_40+m257_40+m258_40+m259_40+m260_40+m261_40+m262_40+m263_40+b40;
   assign out41 = m1_41+m2_41+m3_41+m4_41+m5_41+m6_41+m7_41+m8_41+m9_41+m10_41+m11_41+m12_41+m13_41+m14_41+m15_41+m16_41+m17_41+m18_41+m19_41+m20_41+m21_41+m22_41+m23_41+m24_41+m25_41+m26_41+m27_41+m28_41+m29_41+m30_41+m31_41+m32_41+m33_41+m34_41+m35_41+m36_41+m37_41+m38_41+m39_41+m40_41+m41_41+m42_41+m43_41+m44_41+m45_41+m46_41+m47_41+m48_41+m49_41+m50_41+m51_41+m52_41+m53_41+m54_41+m55_41+m56_41+m57_41+m58_41+m59_41+m60_41+m61_41+m62_41+m63_41+m64_41+m65_41+m66_41+m67_41+m68_41+m69_41+m70_41+m71_41+m72_41+m73_41+m74_41+m75_41+m76_41+m77_41+m78_41+m79_41+m80_41+m81_41+m82_41+m83_41+m84_41+m85_41+m86_41+m87_41+m88_41+m89_41+m90_41+m91_41+m92_41+m93_41+m94_41+m95_41+m96_41+m97_41+m98_41+m99_41+m100_41+m101_41+m102_41+m103_41+m104_41+m105_41+m106_41+m107_41+m108_41+m109_41+m110_41+m111_41+m112_41+m113_41+m114_41+m115_41+m116_41+m117_41+m118_41+m119_41+m120_41+m121_41+m122_41+m123_41+m124_41+m125_41+m126_41+m127_41+m128_41+m129_41+m130_41+m131_41+m132_41+m133_41+m134_41+m135_41+m136_41+m137_41+m138_41+m139_41+m140_41+m141_41+m142_41+m143_41+m144_41+m145_41+m146_41+m147_41+m148_41+m149_41+m150_41+m151_41+m152_41+m153_41+m154_41+m155_41+m156_41+m157_41+m158_41+m159_41+m160_41+m161_41+m162_41+m163_41+m164_41+m165_41+m166_41+m167_41+m168_41+m169_41+m170_41+m171_41+m172_41+m173_41+m174_41+m175_41+m176_41+m177_41+m178_41+m179_41+m180_41+m181_41+m182_41+m183_41+m184_41+m185_41+m186_41+m187_41+m188_41+m189_41+m190_41+m191_41+m192_41+m193_41+m194_41+m195_41+m196_41+m197_41+m198_41+m199_41+m200_41+m201_41+m202_41+m203_41+m204_41+m205_41+m206_41+m207_41+m208_41+m209_41+m210_41+m211_41+m212_41+m213_41+m214_41+m215_41+m216_41+m217_41+m218_41+m219_41+m220_41+m221_41+m222_41+m223_41+m224_41+m225_41+m226_41+m227_41+m228_41+m229_41+m230_41+m231_41+m232_41+m233_41+m234_41+m235_41+m236_41+m237_41+m238_41+m239_41+m240_41+m241_41+m242_41+m243_41+m244_41+m245_41+m246_41+m247_41+m248_41+m249_41+m250_41+m251_41+m252_41+m253_41+m254_41+m255_41+m256_41+m257_41+m258_41+m259_41+m260_41+m261_41+m262_41+m263_41+b41;
   assign out42 = m1_42+m2_42+m3_42+m4_42+m5_42+m6_42+m7_42+m8_42+m9_42+m10_42+m11_42+m12_42+m13_42+m14_42+m15_42+m16_42+m17_42+m18_42+m19_42+m20_42+m21_42+m22_42+m23_42+m24_42+m25_42+m26_42+m27_42+m28_42+m29_42+m30_42+m31_42+m32_42+m33_42+m34_42+m35_42+m36_42+m37_42+m38_42+m39_42+m40_42+m41_42+m42_42+m43_42+m44_42+m45_42+m46_42+m47_42+m48_42+m49_42+m50_42+m51_42+m52_42+m53_42+m54_42+m55_42+m56_42+m57_42+m58_42+m59_42+m60_42+m61_42+m62_42+m63_42+m64_42+m65_42+m66_42+m67_42+m68_42+m69_42+m70_42+m71_42+m72_42+m73_42+m74_42+m75_42+m76_42+m77_42+m78_42+m79_42+m80_42+m81_42+m82_42+m83_42+m84_42+m85_42+m86_42+m87_42+m88_42+m89_42+m90_42+m91_42+m92_42+m93_42+m94_42+m95_42+m96_42+m97_42+m98_42+m99_42+m100_42+m101_42+m102_42+m103_42+m104_42+m105_42+m106_42+m107_42+m108_42+m109_42+m110_42+m111_42+m112_42+m113_42+m114_42+m115_42+m116_42+m117_42+m118_42+m119_42+m120_42+m121_42+m122_42+m123_42+m124_42+m125_42+m126_42+m127_42+m128_42+m129_42+m130_42+m131_42+m132_42+m133_42+m134_42+m135_42+m136_42+m137_42+m138_42+m139_42+m140_42+m141_42+m142_42+m143_42+m144_42+m145_42+m146_42+m147_42+m148_42+m149_42+m150_42+m151_42+m152_42+m153_42+m154_42+m155_42+m156_42+m157_42+m158_42+m159_42+m160_42+m161_42+m162_42+m163_42+m164_42+m165_42+m166_42+m167_42+m168_42+m169_42+m170_42+m171_42+m172_42+m173_42+m174_42+m175_42+m176_42+m177_42+m178_42+m179_42+m180_42+m181_42+m182_42+m183_42+m184_42+m185_42+m186_42+m187_42+m188_42+m189_42+m190_42+m191_42+m192_42+m193_42+m194_42+m195_42+m196_42+m197_42+m198_42+m199_42+m200_42+m201_42+m202_42+m203_42+m204_42+m205_42+m206_42+m207_42+m208_42+m209_42+m210_42+m211_42+m212_42+m213_42+m214_42+m215_42+m216_42+m217_42+m218_42+m219_42+m220_42+m221_42+m222_42+m223_42+m224_42+m225_42+m226_42+m227_42+m228_42+m229_42+m230_42+m231_42+m232_42+m233_42+m234_42+m235_42+m236_42+m237_42+m238_42+m239_42+m240_42+m241_42+m242_42+m243_42+m244_42+m245_42+m246_42+m247_42+m248_42+m249_42+m250_42+m251_42+m252_42+m253_42+m254_42+m255_42+m256_42+m257_42+m258_42+m259_42+m260_42+m261_42+m262_42+m263_42+b42;
   assign out43 = m1_43+m2_43+m3_43+m4_43+m5_43+m6_43+m7_43+m8_43+m9_43+m10_43+m11_43+m12_43+m13_43+m14_43+m15_43+m16_43+m17_43+m18_43+m19_43+m20_43+m21_43+m22_43+m23_43+m24_43+m25_43+m26_43+m27_43+m28_43+m29_43+m30_43+m31_43+m32_43+m33_43+m34_43+m35_43+m36_43+m37_43+m38_43+m39_43+m40_43+m41_43+m42_43+m43_43+m44_43+m45_43+m46_43+m47_43+m48_43+m49_43+m50_43+m51_43+m52_43+m53_43+m54_43+m55_43+m56_43+m57_43+m58_43+m59_43+m60_43+m61_43+m62_43+m63_43+m64_43+m65_43+m66_43+m67_43+m68_43+m69_43+m70_43+m71_43+m72_43+m73_43+m74_43+m75_43+m76_43+m77_43+m78_43+m79_43+m80_43+m81_43+m82_43+m83_43+m84_43+m85_43+m86_43+m87_43+m88_43+m89_43+m90_43+m91_43+m92_43+m93_43+m94_43+m95_43+m96_43+m97_43+m98_43+m99_43+m100_43+m101_43+m102_43+m103_43+m104_43+m105_43+m106_43+m107_43+m108_43+m109_43+m110_43+m111_43+m112_43+m113_43+m114_43+m115_43+m116_43+m117_43+m118_43+m119_43+m120_43+m121_43+m122_43+m123_43+m124_43+m125_43+m126_43+m127_43+m128_43+m129_43+m130_43+m131_43+m132_43+m133_43+m134_43+m135_43+m136_43+m137_43+m138_43+m139_43+m140_43+m141_43+m142_43+m143_43+m144_43+m145_43+m146_43+m147_43+m148_43+m149_43+m150_43+m151_43+m152_43+m153_43+m154_43+m155_43+m156_43+m157_43+m158_43+m159_43+m160_43+m161_43+m162_43+m163_43+m164_43+m165_43+m166_43+m167_43+m168_43+m169_43+m170_43+m171_43+m172_43+m173_43+m174_43+m175_43+m176_43+m177_43+m178_43+m179_43+m180_43+m181_43+m182_43+m183_43+m184_43+m185_43+m186_43+m187_43+m188_43+m189_43+m190_43+m191_43+m192_43+m193_43+m194_43+m195_43+m196_43+m197_43+m198_43+m199_43+m200_43+m201_43+m202_43+m203_43+m204_43+m205_43+m206_43+m207_43+m208_43+m209_43+m210_43+m211_43+m212_43+m213_43+m214_43+m215_43+m216_43+m217_43+m218_43+m219_43+m220_43+m221_43+m222_43+m223_43+m224_43+m225_43+m226_43+m227_43+m228_43+m229_43+m230_43+m231_43+m232_43+m233_43+m234_43+m235_43+m236_43+m237_43+m238_43+m239_43+m240_43+m241_43+m242_43+m243_43+m244_43+m245_43+m246_43+m247_43+m248_43+m249_43+m250_43+m251_43+m252_43+m253_43+m254_43+m255_43+m256_43+m257_43+m258_43+m259_43+m260_43+m261_43+m262_43+m263_43+b43;
   assign out44 = m1_44+m2_44+m3_44+m4_44+m5_44+m6_44+m7_44+m8_44+m9_44+m10_44+m11_44+m12_44+m13_44+m14_44+m15_44+m16_44+m17_44+m18_44+m19_44+m20_44+m21_44+m22_44+m23_44+m24_44+m25_44+m26_44+m27_44+m28_44+m29_44+m30_44+m31_44+m32_44+m33_44+m34_44+m35_44+m36_44+m37_44+m38_44+m39_44+m40_44+m41_44+m42_44+m43_44+m44_44+m45_44+m46_44+m47_44+m48_44+m49_44+m50_44+m51_44+m52_44+m53_44+m54_44+m55_44+m56_44+m57_44+m58_44+m59_44+m60_44+m61_44+m62_44+m63_44+m64_44+m65_44+m66_44+m67_44+m68_44+m69_44+m70_44+m71_44+m72_44+m73_44+m74_44+m75_44+m76_44+m77_44+m78_44+m79_44+m80_44+m81_44+m82_44+m83_44+m84_44+m85_44+m86_44+m87_44+m88_44+m89_44+m90_44+m91_44+m92_44+m93_44+m94_44+m95_44+m96_44+m97_44+m98_44+m99_44+m100_44+m101_44+m102_44+m103_44+m104_44+m105_44+m106_44+m107_44+m108_44+m109_44+m110_44+m111_44+m112_44+m113_44+m114_44+m115_44+m116_44+m117_44+m118_44+m119_44+m120_44+m121_44+m122_44+m123_44+m124_44+m125_44+m126_44+m127_44+m128_44+m129_44+m130_44+m131_44+m132_44+m133_44+m134_44+m135_44+m136_44+m137_44+m138_44+m139_44+m140_44+m141_44+m142_44+m143_44+m144_44+m145_44+m146_44+m147_44+m148_44+m149_44+m150_44+m151_44+m152_44+m153_44+m154_44+m155_44+m156_44+m157_44+m158_44+m159_44+m160_44+m161_44+m162_44+m163_44+m164_44+m165_44+m166_44+m167_44+m168_44+m169_44+m170_44+m171_44+m172_44+m173_44+m174_44+m175_44+m176_44+m177_44+m178_44+m179_44+m180_44+m181_44+m182_44+m183_44+m184_44+m185_44+m186_44+m187_44+m188_44+m189_44+m190_44+m191_44+m192_44+m193_44+m194_44+m195_44+m196_44+m197_44+m198_44+m199_44+m200_44+m201_44+m202_44+m203_44+m204_44+m205_44+m206_44+m207_44+m208_44+m209_44+m210_44+m211_44+m212_44+m213_44+m214_44+m215_44+m216_44+m217_44+m218_44+m219_44+m220_44+m221_44+m222_44+m223_44+m224_44+m225_44+m226_44+m227_44+m228_44+m229_44+m230_44+m231_44+m232_44+m233_44+m234_44+m235_44+m236_44+m237_44+m238_44+m239_44+m240_44+m241_44+m242_44+m243_44+m244_44+m245_44+m246_44+m247_44+m248_44+m249_44+m250_44+m251_44+m252_44+m253_44+m254_44+m255_44+m256_44+m257_44+m258_44+m259_44+m260_44+m261_44+m262_44+m263_44+b44;
   assign out45 = m1_45+m2_45+m3_45+m4_45+m5_45+m6_45+m7_45+m8_45+m9_45+m10_45+m11_45+m12_45+m13_45+m14_45+m15_45+m16_45+m17_45+m18_45+m19_45+m20_45+m21_45+m22_45+m23_45+m24_45+m25_45+m26_45+m27_45+m28_45+m29_45+m30_45+m31_45+m32_45+m33_45+m34_45+m35_45+m36_45+m37_45+m38_45+m39_45+m40_45+m41_45+m42_45+m43_45+m44_45+m45_45+m46_45+m47_45+m48_45+m49_45+m50_45+m51_45+m52_45+m53_45+m54_45+m55_45+m56_45+m57_45+m58_45+m59_45+m60_45+m61_45+m62_45+m63_45+m64_45+m65_45+m66_45+m67_45+m68_45+m69_45+m70_45+m71_45+m72_45+m73_45+m74_45+m75_45+m76_45+m77_45+m78_45+m79_45+m80_45+m81_45+m82_45+m83_45+m84_45+m85_45+m86_45+m87_45+m88_45+m89_45+m90_45+m91_45+m92_45+m93_45+m94_45+m95_45+m96_45+m97_45+m98_45+m99_45+m100_45+m101_45+m102_45+m103_45+m104_45+m105_45+m106_45+m107_45+m108_45+m109_45+m110_45+m111_45+m112_45+m113_45+m114_45+m115_45+m116_45+m117_45+m118_45+m119_45+m120_45+m121_45+m122_45+m123_45+m124_45+m125_45+m126_45+m127_45+m128_45+m129_45+m130_45+m131_45+m132_45+m133_45+m134_45+m135_45+m136_45+m137_45+m138_45+m139_45+m140_45+m141_45+m142_45+m143_45+m144_45+m145_45+m146_45+m147_45+m148_45+m149_45+m150_45+m151_45+m152_45+m153_45+m154_45+m155_45+m156_45+m157_45+m158_45+m159_45+m160_45+m161_45+m162_45+m163_45+m164_45+m165_45+m166_45+m167_45+m168_45+m169_45+m170_45+m171_45+m172_45+m173_45+m174_45+m175_45+m176_45+m177_45+m178_45+m179_45+m180_45+m181_45+m182_45+m183_45+m184_45+m185_45+m186_45+m187_45+m188_45+m189_45+m190_45+m191_45+m192_45+m193_45+m194_45+m195_45+m196_45+m197_45+m198_45+m199_45+m200_45+m201_45+m202_45+m203_45+m204_45+m205_45+m206_45+m207_45+m208_45+m209_45+m210_45+m211_45+m212_45+m213_45+m214_45+m215_45+m216_45+m217_45+m218_45+m219_45+m220_45+m221_45+m222_45+m223_45+m224_45+m225_45+m226_45+m227_45+m228_45+m229_45+m230_45+m231_45+m232_45+m233_45+m234_45+m235_45+m236_45+m237_45+m238_45+m239_45+m240_45+m241_45+m242_45+m243_45+m244_45+m245_45+m246_45+m247_45+m248_45+m249_45+m250_45+m251_45+m252_45+m253_45+m254_45+m255_45+m256_45+m257_45+m258_45+m259_45+m260_45+m261_45+m262_45+m263_45+b45;
   assign out46 = m1_46+m2_46+m3_46+m4_46+m5_46+m6_46+m7_46+m8_46+m9_46+m10_46+m11_46+m12_46+m13_46+m14_46+m15_46+m16_46+m17_46+m18_46+m19_46+m20_46+m21_46+m22_46+m23_46+m24_46+m25_46+m26_46+m27_46+m28_46+m29_46+m30_46+m31_46+m32_46+m33_46+m34_46+m35_46+m36_46+m37_46+m38_46+m39_46+m40_46+m41_46+m42_46+m43_46+m44_46+m45_46+m46_46+m47_46+m48_46+m49_46+m50_46+m51_46+m52_46+m53_46+m54_46+m55_46+m56_46+m57_46+m58_46+m59_46+m60_46+m61_46+m62_46+m63_46+m64_46+m65_46+m66_46+m67_46+m68_46+m69_46+m70_46+m71_46+m72_46+m73_46+m74_46+m75_46+m76_46+m77_46+m78_46+m79_46+m80_46+m81_46+m82_46+m83_46+m84_46+m85_46+m86_46+m87_46+m88_46+m89_46+m90_46+m91_46+m92_46+m93_46+m94_46+m95_46+m96_46+m97_46+m98_46+m99_46+m100_46+m101_46+m102_46+m103_46+m104_46+m105_46+m106_46+m107_46+m108_46+m109_46+m110_46+m111_46+m112_46+m113_46+m114_46+m115_46+m116_46+m117_46+m118_46+m119_46+m120_46+m121_46+m122_46+m123_46+m124_46+m125_46+m126_46+m127_46+m128_46+m129_46+m130_46+m131_46+m132_46+m133_46+m134_46+m135_46+m136_46+m137_46+m138_46+m139_46+m140_46+m141_46+m142_46+m143_46+m144_46+m145_46+m146_46+m147_46+m148_46+m149_46+m150_46+m151_46+m152_46+m153_46+m154_46+m155_46+m156_46+m157_46+m158_46+m159_46+m160_46+m161_46+m162_46+m163_46+m164_46+m165_46+m166_46+m167_46+m168_46+m169_46+m170_46+m171_46+m172_46+m173_46+m174_46+m175_46+m176_46+m177_46+m178_46+m179_46+m180_46+m181_46+m182_46+m183_46+m184_46+m185_46+m186_46+m187_46+m188_46+m189_46+m190_46+m191_46+m192_46+m193_46+m194_46+m195_46+m196_46+m197_46+m198_46+m199_46+m200_46+m201_46+m202_46+m203_46+m204_46+m205_46+m206_46+m207_46+m208_46+m209_46+m210_46+m211_46+m212_46+m213_46+m214_46+m215_46+m216_46+m217_46+m218_46+m219_46+m220_46+m221_46+m222_46+m223_46+m224_46+m225_46+m226_46+m227_46+m228_46+m229_46+m230_46+m231_46+m232_46+m233_46+m234_46+m235_46+m236_46+m237_46+m238_46+m239_46+m240_46+m241_46+m242_46+m243_46+m244_46+m245_46+m246_46+m247_46+m248_46+m249_46+m250_46+m251_46+m252_46+m253_46+m254_46+m255_46+m256_46+m257_46+m258_46+m259_46+m260_46+m261_46+m262_46+m263_46+b46;
   assign out47 = m1_47+m2_47+m3_47+m4_47+m5_47+m6_47+m7_47+m8_47+m9_47+m10_47+m11_47+m12_47+m13_47+m14_47+m15_47+m16_47+m17_47+m18_47+m19_47+m20_47+m21_47+m22_47+m23_47+m24_47+m25_47+m26_47+m27_47+m28_47+m29_47+m30_47+m31_47+m32_47+m33_47+m34_47+m35_47+m36_47+m37_47+m38_47+m39_47+m40_47+m41_47+m42_47+m43_47+m44_47+m45_47+m46_47+m47_47+m48_47+m49_47+m50_47+m51_47+m52_47+m53_47+m54_47+m55_47+m56_47+m57_47+m58_47+m59_47+m60_47+m61_47+m62_47+m63_47+m64_47+m65_47+m66_47+m67_47+m68_47+m69_47+m70_47+m71_47+m72_47+m73_47+m74_47+m75_47+m76_47+m77_47+m78_47+m79_47+m80_47+m81_47+m82_47+m83_47+m84_47+m85_47+m86_47+m87_47+m88_47+m89_47+m90_47+m91_47+m92_47+m93_47+m94_47+m95_47+m96_47+m97_47+m98_47+m99_47+m100_47+m101_47+m102_47+m103_47+m104_47+m105_47+m106_47+m107_47+m108_47+m109_47+m110_47+m111_47+m112_47+m113_47+m114_47+m115_47+m116_47+m117_47+m118_47+m119_47+m120_47+m121_47+m122_47+m123_47+m124_47+m125_47+m126_47+m127_47+m128_47+m129_47+m130_47+m131_47+m132_47+m133_47+m134_47+m135_47+m136_47+m137_47+m138_47+m139_47+m140_47+m141_47+m142_47+m143_47+m144_47+m145_47+m146_47+m147_47+m148_47+m149_47+m150_47+m151_47+m152_47+m153_47+m154_47+m155_47+m156_47+m157_47+m158_47+m159_47+m160_47+m161_47+m162_47+m163_47+m164_47+m165_47+m166_47+m167_47+m168_47+m169_47+m170_47+m171_47+m172_47+m173_47+m174_47+m175_47+m176_47+m177_47+m178_47+m179_47+m180_47+m181_47+m182_47+m183_47+m184_47+m185_47+m186_47+m187_47+m188_47+m189_47+m190_47+m191_47+m192_47+m193_47+m194_47+m195_47+m196_47+m197_47+m198_47+m199_47+m200_47+m201_47+m202_47+m203_47+m204_47+m205_47+m206_47+m207_47+m208_47+m209_47+m210_47+m211_47+m212_47+m213_47+m214_47+m215_47+m216_47+m217_47+m218_47+m219_47+m220_47+m221_47+m222_47+m223_47+m224_47+m225_47+m226_47+m227_47+m228_47+m229_47+m230_47+m231_47+m232_47+m233_47+m234_47+m235_47+m236_47+m237_47+m238_47+m239_47+m240_47+m241_47+m242_47+m243_47+m244_47+m245_47+m246_47+m247_47+m248_47+m249_47+m250_47+m251_47+m252_47+m253_47+m254_47+m255_47+m256_47+m257_47+m258_47+m259_47+m260_47+m261_47+m262_47+m263_47+b47;
   assign out48 = m1_48+m2_48+m3_48+m4_48+m5_48+m6_48+m7_48+m8_48+m9_48+m10_48+m11_48+m12_48+m13_48+m14_48+m15_48+m16_48+m17_48+m18_48+m19_48+m20_48+m21_48+m22_48+m23_48+m24_48+m25_48+m26_48+m27_48+m28_48+m29_48+m30_48+m31_48+m32_48+m33_48+m34_48+m35_48+m36_48+m37_48+m38_48+m39_48+m40_48+m41_48+m42_48+m43_48+m44_48+m45_48+m46_48+m47_48+m48_48+m49_48+m50_48+m51_48+m52_48+m53_48+m54_48+m55_48+m56_48+m57_48+m58_48+m59_48+m60_48+m61_48+m62_48+m63_48+m64_48+m65_48+m66_48+m67_48+m68_48+m69_48+m70_48+m71_48+m72_48+m73_48+m74_48+m75_48+m76_48+m77_48+m78_48+m79_48+m80_48+m81_48+m82_48+m83_48+m84_48+m85_48+m86_48+m87_48+m88_48+m89_48+m90_48+m91_48+m92_48+m93_48+m94_48+m95_48+m96_48+m97_48+m98_48+m99_48+m100_48+m101_48+m102_48+m103_48+m104_48+m105_48+m106_48+m107_48+m108_48+m109_48+m110_48+m111_48+m112_48+m113_48+m114_48+m115_48+m116_48+m117_48+m118_48+m119_48+m120_48+m121_48+m122_48+m123_48+m124_48+m125_48+m126_48+m127_48+m128_48+m129_48+m130_48+m131_48+m132_48+m133_48+m134_48+m135_48+m136_48+m137_48+m138_48+m139_48+m140_48+m141_48+m142_48+m143_48+m144_48+m145_48+m146_48+m147_48+m148_48+m149_48+m150_48+m151_48+m152_48+m153_48+m154_48+m155_48+m156_48+m157_48+m158_48+m159_48+m160_48+m161_48+m162_48+m163_48+m164_48+m165_48+m166_48+m167_48+m168_48+m169_48+m170_48+m171_48+m172_48+m173_48+m174_48+m175_48+m176_48+m177_48+m178_48+m179_48+m180_48+m181_48+m182_48+m183_48+m184_48+m185_48+m186_48+m187_48+m188_48+m189_48+m190_48+m191_48+m192_48+m193_48+m194_48+m195_48+m196_48+m197_48+m198_48+m199_48+m200_48+m201_48+m202_48+m203_48+m204_48+m205_48+m206_48+m207_48+m208_48+m209_48+m210_48+m211_48+m212_48+m213_48+m214_48+m215_48+m216_48+m217_48+m218_48+m219_48+m220_48+m221_48+m222_48+m223_48+m224_48+m225_48+m226_48+m227_48+m228_48+m229_48+m230_48+m231_48+m232_48+m233_48+m234_48+m235_48+m236_48+m237_48+m238_48+m239_48+m240_48+m241_48+m242_48+m243_48+m244_48+m245_48+m246_48+m247_48+m248_48+m249_48+m250_48+m251_48+m252_48+m253_48+m254_48+m255_48+m256_48+m257_48+m258_48+m259_48+m260_48+m261_48+m262_48+m263_48+b48;
   assign out49 = m1_49+m2_49+m3_49+m4_49+m5_49+m6_49+m7_49+m8_49+m9_49+m10_49+m11_49+m12_49+m13_49+m14_49+m15_49+m16_49+m17_49+m18_49+m19_49+m20_49+m21_49+m22_49+m23_49+m24_49+m25_49+m26_49+m27_49+m28_49+m29_49+m30_49+m31_49+m32_49+m33_49+m34_49+m35_49+m36_49+m37_49+m38_49+m39_49+m40_49+m41_49+m42_49+m43_49+m44_49+m45_49+m46_49+m47_49+m48_49+m49_49+m50_49+m51_49+m52_49+m53_49+m54_49+m55_49+m56_49+m57_49+m58_49+m59_49+m60_49+m61_49+m62_49+m63_49+m64_49+m65_49+m66_49+m67_49+m68_49+m69_49+m70_49+m71_49+m72_49+m73_49+m74_49+m75_49+m76_49+m77_49+m78_49+m79_49+m80_49+m81_49+m82_49+m83_49+m84_49+m85_49+m86_49+m87_49+m88_49+m89_49+m90_49+m91_49+m92_49+m93_49+m94_49+m95_49+m96_49+m97_49+m98_49+m99_49+m100_49+m101_49+m102_49+m103_49+m104_49+m105_49+m106_49+m107_49+m108_49+m109_49+m110_49+m111_49+m112_49+m113_49+m114_49+m115_49+m116_49+m117_49+m118_49+m119_49+m120_49+m121_49+m122_49+m123_49+m124_49+m125_49+m126_49+m127_49+m128_49+m129_49+m130_49+m131_49+m132_49+m133_49+m134_49+m135_49+m136_49+m137_49+m138_49+m139_49+m140_49+m141_49+m142_49+m143_49+m144_49+m145_49+m146_49+m147_49+m148_49+m149_49+m150_49+m151_49+m152_49+m153_49+m154_49+m155_49+m156_49+m157_49+m158_49+m159_49+m160_49+m161_49+m162_49+m163_49+m164_49+m165_49+m166_49+m167_49+m168_49+m169_49+m170_49+m171_49+m172_49+m173_49+m174_49+m175_49+m176_49+m177_49+m178_49+m179_49+m180_49+m181_49+m182_49+m183_49+m184_49+m185_49+m186_49+m187_49+m188_49+m189_49+m190_49+m191_49+m192_49+m193_49+m194_49+m195_49+m196_49+m197_49+m198_49+m199_49+m200_49+m201_49+m202_49+m203_49+m204_49+m205_49+m206_49+m207_49+m208_49+m209_49+m210_49+m211_49+m212_49+m213_49+m214_49+m215_49+m216_49+m217_49+m218_49+m219_49+m220_49+m221_49+m222_49+m223_49+m224_49+m225_49+m226_49+m227_49+m228_49+m229_49+m230_49+m231_49+m232_49+m233_49+m234_49+m235_49+m236_49+m237_49+m238_49+m239_49+m240_49+m241_49+m242_49+m243_49+m244_49+m245_49+m246_49+m247_49+m248_49+m249_49+m250_49+m251_49+m252_49+m253_49+m254_49+m255_49+m256_49+m257_49+m258_49+m259_49+m260_49+m261_49+m262_49+m263_49+b49;
   assign out50 = m1_50+m2_50+m3_50+m4_50+m5_50+m6_50+m7_50+m8_50+m9_50+m10_50+m11_50+m12_50+m13_50+m14_50+m15_50+m16_50+m17_50+m18_50+m19_50+m20_50+m21_50+m22_50+m23_50+m24_50+m25_50+m26_50+m27_50+m28_50+m29_50+m30_50+m31_50+m32_50+m33_50+m34_50+m35_50+m36_50+m37_50+m38_50+m39_50+m40_50+m41_50+m42_50+m43_50+m44_50+m45_50+m46_50+m47_50+m48_50+m49_50+m50_50+m51_50+m52_50+m53_50+m54_50+m55_50+m56_50+m57_50+m58_50+m59_50+m60_50+m61_50+m62_50+m63_50+m64_50+m65_50+m66_50+m67_50+m68_50+m69_50+m70_50+m71_50+m72_50+m73_50+m74_50+m75_50+m76_50+m77_50+m78_50+m79_50+m80_50+m81_50+m82_50+m83_50+m84_50+m85_50+m86_50+m87_50+m88_50+m89_50+m90_50+m91_50+m92_50+m93_50+m94_50+m95_50+m96_50+m97_50+m98_50+m99_50+m100_50+m101_50+m102_50+m103_50+m104_50+m105_50+m106_50+m107_50+m108_50+m109_50+m110_50+m111_50+m112_50+m113_50+m114_50+m115_50+m116_50+m117_50+m118_50+m119_50+m120_50+m121_50+m122_50+m123_50+m124_50+m125_50+m126_50+m127_50+m128_50+m129_50+m130_50+m131_50+m132_50+m133_50+m134_50+m135_50+m136_50+m137_50+m138_50+m139_50+m140_50+m141_50+m142_50+m143_50+m144_50+m145_50+m146_50+m147_50+m148_50+m149_50+m150_50+m151_50+m152_50+m153_50+m154_50+m155_50+m156_50+m157_50+m158_50+m159_50+m160_50+m161_50+m162_50+m163_50+m164_50+m165_50+m166_50+m167_50+m168_50+m169_50+m170_50+m171_50+m172_50+m173_50+m174_50+m175_50+m176_50+m177_50+m178_50+m179_50+m180_50+m181_50+m182_50+m183_50+m184_50+m185_50+m186_50+m187_50+m188_50+m189_50+m190_50+m191_50+m192_50+m193_50+m194_50+m195_50+m196_50+m197_50+m198_50+m199_50+m200_50+m201_50+m202_50+m203_50+m204_50+m205_50+m206_50+m207_50+m208_50+m209_50+m210_50+m211_50+m212_50+m213_50+m214_50+m215_50+m216_50+m217_50+m218_50+m219_50+m220_50+m221_50+m222_50+m223_50+m224_50+m225_50+m226_50+m227_50+m228_50+m229_50+m230_50+m231_50+m232_50+m233_50+m234_50+m235_50+m236_50+m237_50+m238_50+m239_50+m240_50+m241_50+m242_50+m243_50+m244_50+m245_50+m246_50+m247_50+m248_50+m249_50+m250_50+m251_50+m252_50+m253_50+m254_50+m255_50+m256_50+m257_50+m258_50+m259_50+m260_50+m261_50+m262_50+m263_50+b50;
   assign out51 = m1_51+m2_51+m3_51+m4_51+m5_51+m6_51+m7_51+m8_51+m9_51+m10_51+m11_51+m12_51+m13_51+m14_51+m15_51+m16_51+m17_51+m18_51+m19_51+m20_51+m21_51+m22_51+m23_51+m24_51+m25_51+m26_51+m27_51+m28_51+m29_51+m30_51+m31_51+m32_51+m33_51+m34_51+m35_51+m36_51+m37_51+m38_51+m39_51+m40_51+m41_51+m42_51+m43_51+m44_51+m45_51+m46_51+m47_51+m48_51+m49_51+m50_51+m51_51+m52_51+m53_51+m54_51+m55_51+m56_51+m57_51+m58_51+m59_51+m60_51+m61_51+m62_51+m63_51+m64_51+m65_51+m66_51+m67_51+m68_51+m69_51+m70_51+m71_51+m72_51+m73_51+m74_51+m75_51+m76_51+m77_51+m78_51+m79_51+m80_51+m81_51+m82_51+m83_51+m84_51+m85_51+m86_51+m87_51+m88_51+m89_51+m90_51+m91_51+m92_51+m93_51+m94_51+m95_51+m96_51+m97_51+m98_51+m99_51+m100_51+m101_51+m102_51+m103_51+m104_51+m105_51+m106_51+m107_51+m108_51+m109_51+m110_51+m111_51+m112_51+m113_51+m114_51+m115_51+m116_51+m117_51+m118_51+m119_51+m120_51+m121_51+m122_51+m123_51+m124_51+m125_51+m126_51+m127_51+m128_51+m129_51+m130_51+m131_51+m132_51+m133_51+m134_51+m135_51+m136_51+m137_51+m138_51+m139_51+m140_51+m141_51+m142_51+m143_51+m144_51+m145_51+m146_51+m147_51+m148_51+m149_51+m150_51+m151_51+m152_51+m153_51+m154_51+m155_51+m156_51+m157_51+m158_51+m159_51+m160_51+m161_51+m162_51+m163_51+m164_51+m165_51+m166_51+m167_51+m168_51+m169_51+m170_51+m171_51+m172_51+m173_51+m174_51+m175_51+m176_51+m177_51+m178_51+m179_51+m180_51+m181_51+m182_51+m183_51+m184_51+m185_51+m186_51+m187_51+m188_51+m189_51+m190_51+m191_51+m192_51+m193_51+m194_51+m195_51+m196_51+m197_51+m198_51+m199_51+m200_51+m201_51+m202_51+m203_51+m204_51+m205_51+m206_51+m207_51+m208_51+m209_51+m210_51+m211_51+m212_51+m213_51+m214_51+m215_51+m216_51+m217_51+m218_51+m219_51+m220_51+m221_51+m222_51+m223_51+m224_51+m225_51+m226_51+m227_51+m228_51+m229_51+m230_51+m231_51+m232_51+m233_51+m234_51+m235_51+m236_51+m237_51+m238_51+m239_51+m240_51+m241_51+m242_51+m243_51+m244_51+m245_51+m246_51+m247_51+m248_51+m249_51+m250_51+m251_51+m252_51+m253_51+m254_51+m255_51+m256_51+m257_51+m258_51+m259_51+m260_51+m261_51+m262_51+m263_51+b51;
   assign out52 = m1_52+m2_52+m3_52+m4_52+m5_52+m6_52+m7_52+m8_52+m9_52+m10_52+m11_52+m12_52+m13_52+m14_52+m15_52+m16_52+m17_52+m18_52+m19_52+m20_52+m21_52+m22_52+m23_52+m24_52+m25_52+m26_52+m27_52+m28_52+m29_52+m30_52+m31_52+m32_52+m33_52+m34_52+m35_52+m36_52+m37_52+m38_52+m39_52+m40_52+m41_52+m42_52+m43_52+m44_52+m45_52+m46_52+m47_52+m48_52+m49_52+m50_52+m51_52+m52_52+m53_52+m54_52+m55_52+m56_52+m57_52+m58_52+m59_52+m60_52+m61_52+m62_52+m63_52+m64_52+m65_52+m66_52+m67_52+m68_52+m69_52+m70_52+m71_52+m72_52+m73_52+m74_52+m75_52+m76_52+m77_52+m78_52+m79_52+m80_52+m81_52+m82_52+m83_52+m84_52+m85_52+m86_52+m87_52+m88_52+m89_52+m90_52+m91_52+m92_52+m93_52+m94_52+m95_52+m96_52+m97_52+m98_52+m99_52+m100_52+m101_52+m102_52+m103_52+m104_52+m105_52+m106_52+m107_52+m108_52+m109_52+m110_52+m111_52+m112_52+m113_52+m114_52+m115_52+m116_52+m117_52+m118_52+m119_52+m120_52+m121_52+m122_52+m123_52+m124_52+m125_52+m126_52+m127_52+m128_52+m129_52+m130_52+m131_52+m132_52+m133_52+m134_52+m135_52+m136_52+m137_52+m138_52+m139_52+m140_52+m141_52+m142_52+m143_52+m144_52+m145_52+m146_52+m147_52+m148_52+m149_52+m150_52+m151_52+m152_52+m153_52+m154_52+m155_52+m156_52+m157_52+m158_52+m159_52+m160_52+m161_52+m162_52+m163_52+m164_52+m165_52+m166_52+m167_52+m168_52+m169_52+m170_52+m171_52+m172_52+m173_52+m174_52+m175_52+m176_52+m177_52+m178_52+m179_52+m180_52+m181_52+m182_52+m183_52+m184_52+m185_52+m186_52+m187_52+m188_52+m189_52+m190_52+m191_52+m192_52+m193_52+m194_52+m195_52+m196_52+m197_52+m198_52+m199_52+m200_52+m201_52+m202_52+m203_52+m204_52+m205_52+m206_52+m207_52+m208_52+m209_52+m210_52+m211_52+m212_52+m213_52+m214_52+m215_52+m216_52+m217_52+m218_52+m219_52+m220_52+m221_52+m222_52+m223_52+m224_52+m225_52+m226_52+m227_52+m228_52+m229_52+m230_52+m231_52+m232_52+m233_52+m234_52+m235_52+m236_52+m237_52+m238_52+m239_52+m240_52+m241_52+m242_52+m243_52+m244_52+m245_52+m246_52+m247_52+m248_52+m249_52+m250_52+m251_52+m252_52+m253_52+m254_52+m255_52+m256_52+m257_52+m258_52+m259_52+m260_52+m261_52+m262_52+m263_52+b52;
   assign out53 = m1_53+m2_53+m3_53+m4_53+m5_53+m6_53+m7_53+m8_53+m9_53+m10_53+m11_53+m12_53+m13_53+m14_53+m15_53+m16_53+m17_53+m18_53+m19_53+m20_53+m21_53+m22_53+m23_53+m24_53+m25_53+m26_53+m27_53+m28_53+m29_53+m30_53+m31_53+m32_53+m33_53+m34_53+m35_53+m36_53+m37_53+m38_53+m39_53+m40_53+m41_53+m42_53+m43_53+m44_53+m45_53+m46_53+m47_53+m48_53+m49_53+m50_53+m51_53+m52_53+m53_53+m54_53+m55_53+m56_53+m57_53+m58_53+m59_53+m60_53+m61_53+m62_53+m63_53+m64_53+m65_53+m66_53+m67_53+m68_53+m69_53+m70_53+m71_53+m72_53+m73_53+m74_53+m75_53+m76_53+m77_53+m78_53+m79_53+m80_53+m81_53+m82_53+m83_53+m84_53+m85_53+m86_53+m87_53+m88_53+m89_53+m90_53+m91_53+m92_53+m93_53+m94_53+m95_53+m96_53+m97_53+m98_53+m99_53+m100_53+m101_53+m102_53+m103_53+m104_53+m105_53+m106_53+m107_53+m108_53+m109_53+m110_53+m111_53+m112_53+m113_53+m114_53+m115_53+m116_53+m117_53+m118_53+m119_53+m120_53+m121_53+m122_53+m123_53+m124_53+m125_53+m126_53+m127_53+m128_53+m129_53+m130_53+m131_53+m132_53+m133_53+m134_53+m135_53+m136_53+m137_53+m138_53+m139_53+m140_53+m141_53+m142_53+m143_53+m144_53+m145_53+m146_53+m147_53+m148_53+m149_53+m150_53+m151_53+m152_53+m153_53+m154_53+m155_53+m156_53+m157_53+m158_53+m159_53+m160_53+m161_53+m162_53+m163_53+m164_53+m165_53+m166_53+m167_53+m168_53+m169_53+m170_53+m171_53+m172_53+m173_53+m174_53+m175_53+m176_53+m177_53+m178_53+m179_53+m180_53+m181_53+m182_53+m183_53+m184_53+m185_53+m186_53+m187_53+m188_53+m189_53+m190_53+m191_53+m192_53+m193_53+m194_53+m195_53+m196_53+m197_53+m198_53+m199_53+m200_53+m201_53+m202_53+m203_53+m204_53+m205_53+m206_53+m207_53+m208_53+m209_53+m210_53+m211_53+m212_53+m213_53+m214_53+m215_53+m216_53+m217_53+m218_53+m219_53+m220_53+m221_53+m222_53+m223_53+m224_53+m225_53+m226_53+m227_53+m228_53+m229_53+m230_53+m231_53+m232_53+m233_53+m234_53+m235_53+m236_53+m237_53+m238_53+m239_53+m240_53+m241_53+m242_53+m243_53+m244_53+m245_53+m246_53+m247_53+m248_53+m249_53+m250_53+m251_53+m252_53+m253_53+m254_53+m255_53+m256_53+m257_53+m258_53+m259_53+m260_53+m261_53+m262_53+m263_53+b53;
   assign out54 = m1_54+m2_54+m3_54+m4_54+m5_54+m6_54+m7_54+m8_54+m9_54+m10_54+m11_54+m12_54+m13_54+m14_54+m15_54+m16_54+m17_54+m18_54+m19_54+m20_54+m21_54+m22_54+m23_54+m24_54+m25_54+m26_54+m27_54+m28_54+m29_54+m30_54+m31_54+m32_54+m33_54+m34_54+m35_54+m36_54+m37_54+m38_54+m39_54+m40_54+m41_54+m42_54+m43_54+m44_54+m45_54+m46_54+m47_54+m48_54+m49_54+m50_54+m51_54+m52_54+m53_54+m54_54+m55_54+m56_54+m57_54+m58_54+m59_54+m60_54+m61_54+m62_54+m63_54+m64_54+m65_54+m66_54+m67_54+m68_54+m69_54+m70_54+m71_54+m72_54+m73_54+m74_54+m75_54+m76_54+m77_54+m78_54+m79_54+m80_54+m81_54+m82_54+m83_54+m84_54+m85_54+m86_54+m87_54+m88_54+m89_54+m90_54+m91_54+m92_54+m93_54+m94_54+m95_54+m96_54+m97_54+m98_54+m99_54+m100_54+m101_54+m102_54+m103_54+m104_54+m105_54+m106_54+m107_54+m108_54+m109_54+m110_54+m111_54+m112_54+m113_54+m114_54+m115_54+m116_54+m117_54+m118_54+m119_54+m120_54+m121_54+m122_54+m123_54+m124_54+m125_54+m126_54+m127_54+m128_54+m129_54+m130_54+m131_54+m132_54+m133_54+m134_54+m135_54+m136_54+m137_54+m138_54+m139_54+m140_54+m141_54+m142_54+m143_54+m144_54+m145_54+m146_54+m147_54+m148_54+m149_54+m150_54+m151_54+m152_54+m153_54+m154_54+m155_54+m156_54+m157_54+m158_54+m159_54+m160_54+m161_54+m162_54+m163_54+m164_54+m165_54+m166_54+m167_54+m168_54+m169_54+m170_54+m171_54+m172_54+m173_54+m174_54+m175_54+m176_54+m177_54+m178_54+m179_54+m180_54+m181_54+m182_54+m183_54+m184_54+m185_54+m186_54+m187_54+m188_54+m189_54+m190_54+m191_54+m192_54+m193_54+m194_54+m195_54+m196_54+m197_54+m198_54+m199_54+m200_54+m201_54+m202_54+m203_54+m204_54+m205_54+m206_54+m207_54+m208_54+m209_54+m210_54+m211_54+m212_54+m213_54+m214_54+m215_54+m216_54+m217_54+m218_54+m219_54+m220_54+m221_54+m222_54+m223_54+m224_54+m225_54+m226_54+m227_54+m228_54+m229_54+m230_54+m231_54+m232_54+m233_54+m234_54+m235_54+m236_54+m237_54+m238_54+m239_54+m240_54+m241_54+m242_54+m243_54+m244_54+m245_54+m246_54+m247_54+m248_54+m249_54+m250_54+m251_54+m252_54+m253_54+m254_54+m255_54+m256_54+m257_54+m258_54+m259_54+m260_54+m261_54+m262_54+m263_54+b54;
   assign out55 = m1_55+m2_55+m3_55+m4_55+m5_55+m6_55+m7_55+m8_55+m9_55+m10_55+m11_55+m12_55+m13_55+m14_55+m15_55+m16_55+m17_55+m18_55+m19_55+m20_55+m21_55+m22_55+m23_55+m24_55+m25_55+m26_55+m27_55+m28_55+m29_55+m30_55+m31_55+m32_55+m33_55+m34_55+m35_55+m36_55+m37_55+m38_55+m39_55+m40_55+m41_55+m42_55+m43_55+m44_55+m45_55+m46_55+m47_55+m48_55+m49_55+m50_55+m51_55+m52_55+m53_55+m54_55+m55_55+m56_55+m57_55+m58_55+m59_55+m60_55+m61_55+m62_55+m63_55+m64_55+m65_55+m66_55+m67_55+m68_55+m69_55+m70_55+m71_55+m72_55+m73_55+m74_55+m75_55+m76_55+m77_55+m78_55+m79_55+m80_55+m81_55+m82_55+m83_55+m84_55+m85_55+m86_55+m87_55+m88_55+m89_55+m90_55+m91_55+m92_55+m93_55+m94_55+m95_55+m96_55+m97_55+m98_55+m99_55+m100_55+m101_55+m102_55+m103_55+m104_55+m105_55+m106_55+m107_55+m108_55+m109_55+m110_55+m111_55+m112_55+m113_55+m114_55+m115_55+m116_55+m117_55+m118_55+m119_55+m120_55+m121_55+m122_55+m123_55+m124_55+m125_55+m126_55+m127_55+m128_55+m129_55+m130_55+m131_55+m132_55+m133_55+m134_55+m135_55+m136_55+m137_55+m138_55+m139_55+m140_55+m141_55+m142_55+m143_55+m144_55+m145_55+m146_55+m147_55+m148_55+m149_55+m150_55+m151_55+m152_55+m153_55+m154_55+m155_55+m156_55+m157_55+m158_55+m159_55+m160_55+m161_55+m162_55+m163_55+m164_55+m165_55+m166_55+m167_55+m168_55+m169_55+m170_55+m171_55+m172_55+m173_55+m174_55+m175_55+m176_55+m177_55+m178_55+m179_55+m180_55+m181_55+m182_55+m183_55+m184_55+m185_55+m186_55+m187_55+m188_55+m189_55+m190_55+m191_55+m192_55+m193_55+m194_55+m195_55+m196_55+m197_55+m198_55+m199_55+m200_55+m201_55+m202_55+m203_55+m204_55+m205_55+m206_55+m207_55+m208_55+m209_55+m210_55+m211_55+m212_55+m213_55+m214_55+m215_55+m216_55+m217_55+m218_55+m219_55+m220_55+m221_55+m222_55+m223_55+m224_55+m225_55+m226_55+m227_55+m228_55+m229_55+m230_55+m231_55+m232_55+m233_55+m234_55+m235_55+m236_55+m237_55+m238_55+m239_55+m240_55+m241_55+m242_55+m243_55+m244_55+m245_55+m246_55+m247_55+m248_55+m249_55+m250_55+m251_55+m252_55+m253_55+m254_55+m255_55+m256_55+m257_55+m258_55+m259_55+m260_55+m261_55+m262_55+m263_55+b55;
   assign out56 = m1_56+m2_56+m3_56+m4_56+m5_56+m6_56+m7_56+m8_56+m9_56+m10_56+m11_56+m12_56+m13_56+m14_56+m15_56+m16_56+m17_56+m18_56+m19_56+m20_56+m21_56+m22_56+m23_56+m24_56+m25_56+m26_56+m27_56+m28_56+m29_56+m30_56+m31_56+m32_56+m33_56+m34_56+m35_56+m36_56+m37_56+m38_56+m39_56+m40_56+m41_56+m42_56+m43_56+m44_56+m45_56+m46_56+m47_56+m48_56+m49_56+m50_56+m51_56+m52_56+m53_56+m54_56+m55_56+m56_56+m57_56+m58_56+m59_56+m60_56+m61_56+m62_56+m63_56+m64_56+m65_56+m66_56+m67_56+m68_56+m69_56+m70_56+m71_56+m72_56+m73_56+m74_56+m75_56+m76_56+m77_56+m78_56+m79_56+m80_56+m81_56+m82_56+m83_56+m84_56+m85_56+m86_56+m87_56+m88_56+m89_56+m90_56+m91_56+m92_56+m93_56+m94_56+m95_56+m96_56+m97_56+m98_56+m99_56+m100_56+m101_56+m102_56+m103_56+m104_56+m105_56+m106_56+m107_56+m108_56+m109_56+m110_56+m111_56+m112_56+m113_56+m114_56+m115_56+m116_56+m117_56+m118_56+m119_56+m120_56+m121_56+m122_56+m123_56+m124_56+m125_56+m126_56+m127_56+m128_56+m129_56+m130_56+m131_56+m132_56+m133_56+m134_56+m135_56+m136_56+m137_56+m138_56+m139_56+m140_56+m141_56+m142_56+m143_56+m144_56+m145_56+m146_56+m147_56+m148_56+m149_56+m150_56+m151_56+m152_56+m153_56+m154_56+m155_56+m156_56+m157_56+m158_56+m159_56+m160_56+m161_56+m162_56+m163_56+m164_56+m165_56+m166_56+m167_56+m168_56+m169_56+m170_56+m171_56+m172_56+m173_56+m174_56+m175_56+m176_56+m177_56+m178_56+m179_56+m180_56+m181_56+m182_56+m183_56+m184_56+m185_56+m186_56+m187_56+m188_56+m189_56+m190_56+m191_56+m192_56+m193_56+m194_56+m195_56+m196_56+m197_56+m198_56+m199_56+m200_56+m201_56+m202_56+m203_56+m204_56+m205_56+m206_56+m207_56+m208_56+m209_56+m210_56+m211_56+m212_56+m213_56+m214_56+m215_56+m216_56+m217_56+m218_56+m219_56+m220_56+m221_56+m222_56+m223_56+m224_56+m225_56+m226_56+m227_56+m228_56+m229_56+m230_56+m231_56+m232_56+m233_56+m234_56+m235_56+m236_56+m237_56+m238_56+m239_56+m240_56+m241_56+m242_56+m243_56+m244_56+m245_56+m246_56+m247_56+m248_56+m249_56+m250_56+m251_56+m252_56+m253_56+m254_56+m255_56+m256_56+m257_56+m258_56+m259_56+m260_56+m261_56+m262_56+m263_56+b56;
   assign out57 = m1_57+m2_57+m3_57+m4_57+m5_57+m6_57+m7_57+m8_57+m9_57+m10_57+m11_57+m12_57+m13_57+m14_57+m15_57+m16_57+m17_57+m18_57+m19_57+m20_57+m21_57+m22_57+m23_57+m24_57+m25_57+m26_57+m27_57+m28_57+m29_57+m30_57+m31_57+m32_57+m33_57+m34_57+m35_57+m36_57+m37_57+m38_57+m39_57+m40_57+m41_57+m42_57+m43_57+m44_57+m45_57+m46_57+m47_57+m48_57+m49_57+m50_57+m51_57+m52_57+m53_57+m54_57+m55_57+m56_57+m57_57+m58_57+m59_57+m60_57+m61_57+m62_57+m63_57+m64_57+m65_57+m66_57+m67_57+m68_57+m69_57+m70_57+m71_57+m72_57+m73_57+m74_57+m75_57+m76_57+m77_57+m78_57+m79_57+m80_57+m81_57+m82_57+m83_57+m84_57+m85_57+m86_57+m87_57+m88_57+m89_57+m90_57+m91_57+m92_57+m93_57+m94_57+m95_57+m96_57+m97_57+m98_57+m99_57+m100_57+m101_57+m102_57+m103_57+m104_57+m105_57+m106_57+m107_57+m108_57+m109_57+m110_57+m111_57+m112_57+m113_57+m114_57+m115_57+m116_57+m117_57+m118_57+m119_57+m120_57+m121_57+m122_57+m123_57+m124_57+m125_57+m126_57+m127_57+m128_57+m129_57+m130_57+m131_57+m132_57+m133_57+m134_57+m135_57+m136_57+m137_57+m138_57+m139_57+m140_57+m141_57+m142_57+m143_57+m144_57+m145_57+m146_57+m147_57+m148_57+m149_57+m150_57+m151_57+m152_57+m153_57+m154_57+m155_57+m156_57+m157_57+m158_57+m159_57+m160_57+m161_57+m162_57+m163_57+m164_57+m165_57+m166_57+m167_57+m168_57+m169_57+m170_57+m171_57+m172_57+m173_57+m174_57+m175_57+m176_57+m177_57+m178_57+m179_57+m180_57+m181_57+m182_57+m183_57+m184_57+m185_57+m186_57+m187_57+m188_57+m189_57+m190_57+m191_57+m192_57+m193_57+m194_57+m195_57+m196_57+m197_57+m198_57+m199_57+m200_57+m201_57+m202_57+m203_57+m204_57+m205_57+m206_57+m207_57+m208_57+m209_57+m210_57+m211_57+m212_57+m213_57+m214_57+m215_57+m216_57+m217_57+m218_57+m219_57+m220_57+m221_57+m222_57+m223_57+m224_57+m225_57+m226_57+m227_57+m228_57+m229_57+m230_57+m231_57+m232_57+m233_57+m234_57+m235_57+m236_57+m237_57+m238_57+m239_57+m240_57+m241_57+m242_57+m243_57+m244_57+m245_57+m246_57+m247_57+m248_57+m249_57+m250_57+m251_57+m252_57+m253_57+m254_57+m255_57+m256_57+m257_57+m258_57+m259_57+m260_57+m261_57+m262_57+m263_57+b57;
   assign out58 = m1_58+m2_58+m3_58+m4_58+m5_58+m6_58+m7_58+m8_58+m9_58+m10_58+m11_58+m12_58+m13_58+m14_58+m15_58+m16_58+m17_58+m18_58+m19_58+m20_58+m21_58+m22_58+m23_58+m24_58+m25_58+m26_58+m27_58+m28_58+m29_58+m30_58+m31_58+m32_58+m33_58+m34_58+m35_58+m36_58+m37_58+m38_58+m39_58+m40_58+m41_58+m42_58+m43_58+m44_58+m45_58+m46_58+m47_58+m48_58+m49_58+m50_58+m51_58+m52_58+m53_58+m54_58+m55_58+m56_58+m57_58+m58_58+m59_58+m60_58+m61_58+m62_58+m63_58+m64_58+m65_58+m66_58+m67_58+m68_58+m69_58+m70_58+m71_58+m72_58+m73_58+m74_58+m75_58+m76_58+m77_58+m78_58+m79_58+m80_58+m81_58+m82_58+m83_58+m84_58+m85_58+m86_58+m87_58+m88_58+m89_58+m90_58+m91_58+m92_58+m93_58+m94_58+m95_58+m96_58+m97_58+m98_58+m99_58+m100_58+m101_58+m102_58+m103_58+m104_58+m105_58+m106_58+m107_58+m108_58+m109_58+m110_58+m111_58+m112_58+m113_58+m114_58+m115_58+m116_58+m117_58+m118_58+m119_58+m120_58+m121_58+m122_58+m123_58+m124_58+m125_58+m126_58+m127_58+m128_58+m129_58+m130_58+m131_58+m132_58+m133_58+m134_58+m135_58+m136_58+m137_58+m138_58+m139_58+m140_58+m141_58+m142_58+m143_58+m144_58+m145_58+m146_58+m147_58+m148_58+m149_58+m150_58+m151_58+m152_58+m153_58+m154_58+m155_58+m156_58+m157_58+m158_58+m159_58+m160_58+m161_58+m162_58+m163_58+m164_58+m165_58+m166_58+m167_58+m168_58+m169_58+m170_58+m171_58+m172_58+m173_58+m174_58+m175_58+m176_58+m177_58+m178_58+m179_58+m180_58+m181_58+m182_58+m183_58+m184_58+m185_58+m186_58+m187_58+m188_58+m189_58+m190_58+m191_58+m192_58+m193_58+m194_58+m195_58+m196_58+m197_58+m198_58+m199_58+m200_58+m201_58+m202_58+m203_58+m204_58+m205_58+m206_58+m207_58+m208_58+m209_58+m210_58+m211_58+m212_58+m213_58+m214_58+m215_58+m216_58+m217_58+m218_58+m219_58+m220_58+m221_58+m222_58+m223_58+m224_58+m225_58+m226_58+m227_58+m228_58+m229_58+m230_58+m231_58+m232_58+m233_58+m234_58+m235_58+m236_58+m237_58+m238_58+m239_58+m240_58+m241_58+m242_58+m243_58+m244_58+m245_58+m246_58+m247_58+m248_58+m249_58+m250_58+m251_58+m252_58+m253_58+m254_58+m255_58+m256_58+m257_58+m258_58+m259_58+m260_58+m261_58+m262_58+m263_58+b58;
   assign out59 = m1_59+m2_59+m3_59+m4_59+m5_59+m6_59+m7_59+m8_59+m9_59+m10_59+m11_59+m12_59+m13_59+m14_59+m15_59+m16_59+m17_59+m18_59+m19_59+m20_59+m21_59+m22_59+m23_59+m24_59+m25_59+m26_59+m27_59+m28_59+m29_59+m30_59+m31_59+m32_59+m33_59+m34_59+m35_59+m36_59+m37_59+m38_59+m39_59+m40_59+m41_59+m42_59+m43_59+m44_59+m45_59+m46_59+m47_59+m48_59+m49_59+m50_59+m51_59+m52_59+m53_59+m54_59+m55_59+m56_59+m57_59+m58_59+m59_59+m60_59+m61_59+m62_59+m63_59+m64_59+m65_59+m66_59+m67_59+m68_59+m69_59+m70_59+m71_59+m72_59+m73_59+m74_59+m75_59+m76_59+m77_59+m78_59+m79_59+m80_59+m81_59+m82_59+m83_59+m84_59+m85_59+m86_59+m87_59+m88_59+m89_59+m90_59+m91_59+m92_59+m93_59+m94_59+m95_59+m96_59+m97_59+m98_59+m99_59+m100_59+m101_59+m102_59+m103_59+m104_59+m105_59+m106_59+m107_59+m108_59+m109_59+m110_59+m111_59+m112_59+m113_59+m114_59+m115_59+m116_59+m117_59+m118_59+m119_59+m120_59+m121_59+m122_59+m123_59+m124_59+m125_59+m126_59+m127_59+m128_59+m129_59+m130_59+m131_59+m132_59+m133_59+m134_59+m135_59+m136_59+m137_59+m138_59+m139_59+m140_59+m141_59+m142_59+m143_59+m144_59+m145_59+m146_59+m147_59+m148_59+m149_59+m150_59+m151_59+m152_59+m153_59+m154_59+m155_59+m156_59+m157_59+m158_59+m159_59+m160_59+m161_59+m162_59+m163_59+m164_59+m165_59+m166_59+m167_59+m168_59+m169_59+m170_59+m171_59+m172_59+m173_59+m174_59+m175_59+m176_59+m177_59+m178_59+m179_59+m180_59+m181_59+m182_59+m183_59+m184_59+m185_59+m186_59+m187_59+m188_59+m189_59+m190_59+m191_59+m192_59+m193_59+m194_59+m195_59+m196_59+m197_59+m198_59+m199_59+m200_59+m201_59+m202_59+m203_59+m204_59+m205_59+m206_59+m207_59+m208_59+m209_59+m210_59+m211_59+m212_59+m213_59+m214_59+m215_59+m216_59+m217_59+m218_59+m219_59+m220_59+m221_59+m222_59+m223_59+m224_59+m225_59+m226_59+m227_59+m228_59+m229_59+m230_59+m231_59+m232_59+m233_59+m234_59+m235_59+m236_59+m237_59+m238_59+m239_59+m240_59+m241_59+m242_59+m243_59+m244_59+m245_59+m246_59+m247_59+m248_59+m249_59+m250_59+m251_59+m252_59+m253_59+m254_59+m255_59+m256_59+m257_59+m258_59+m259_59+m260_59+m261_59+m262_59+m263_59+b59;
   assign out60 = m1_60+m2_60+m3_60+m4_60+m5_60+m6_60+m7_60+m8_60+m9_60+m10_60+m11_60+m12_60+m13_60+m14_60+m15_60+m16_60+m17_60+m18_60+m19_60+m20_60+m21_60+m22_60+m23_60+m24_60+m25_60+m26_60+m27_60+m28_60+m29_60+m30_60+m31_60+m32_60+m33_60+m34_60+m35_60+m36_60+m37_60+m38_60+m39_60+m40_60+m41_60+m42_60+m43_60+m44_60+m45_60+m46_60+m47_60+m48_60+m49_60+m50_60+m51_60+m52_60+m53_60+m54_60+m55_60+m56_60+m57_60+m58_60+m59_60+m60_60+m61_60+m62_60+m63_60+m64_60+m65_60+m66_60+m67_60+m68_60+m69_60+m70_60+m71_60+m72_60+m73_60+m74_60+m75_60+m76_60+m77_60+m78_60+m79_60+m80_60+m81_60+m82_60+m83_60+m84_60+m85_60+m86_60+m87_60+m88_60+m89_60+m90_60+m91_60+m92_60+m93_60+m94_60+m95_60+m96_60+m97_60+m98_60+m99_60+m100_60+m101_60+m102_60+m103_60+m104_60+m105_60+m106_60+m107_60+m108_60+m109_60+m110_60+m111_60+m112_60+m113_60+m114_60+m115_60+m116_60+m117_60+m118_60+m119_60+m120_60+m121_60+m122_60+m123_60+m124_60+m125_60+m126_60+m127_60+m128_60+m129_60+m130_60+m131_60+m132_60+m133_60+m134_60+m135_60+m136_60+m137_60+m138_60+m139_60+m140_60+m141_60+m142_60+m143_60+m144_60+m145_60+m146_60+m147_60+m148_60+m149_60+m150_60+m151_60+m152_60+m153_60+m154_60+m155_60+m156_60+m157_60+m158_60+m159_60+m160_60+m161_60+m162_60+m163_60+m164_60+m165_60+m166_60+m167_60+m168_60+m169_60+m170_60+m171_60+m172_60+m173_60+m174_60+m175_60+m176_60+m177_60+m178_60+m179_60+m180_60+m181_60+m182_60+m183_60+m184_60+m185_60+m186_60+m187_60+m188_60+m189_60+m190_60+m191_60+m192_60+m193_60+m194_60+m195_60+m196_60+m197_60+m198_60+m199_60+m200_60+m201_60+m202_60+m203_60+m204_60+m205_60+m206_60+m207_60+m208_60+m209_60+m210_60+m211_60+m212_60+m213_60+m214_60+m215_60+m216_60+m217_60+m218_60+m219_60+m220_60+m221_60+m222_60+m223_60+m224_60+m225_60+m226_60+m227_60+m228_60+m229_60+m230_60+m231_60+m232_60+m233_60+m234_60+m235_60+m236_60+m237_60+m238_60+m239_60+m240_60+m241_60+m242_60+m243_60+m244_60+m245_60+m246_60+m247_60+m248_60+m249_60+m250_60+m251_60+m252_60+m253_60+m254_60+m255_60+m256_60+m257_60+m258_60+m259_60+m260_60+m261_60+m262_60+m263_60+b60;
   assign out61 = m1_61+m2_61+m3_61+m4_61+m5_61+m6_61+m7_61+m8_61+m9_61+m10_61+m11_61+m12_61+m13_61+m14_61+m15_61+m16_61+m17_61+m18_61+m19_61+m20_61+m21_61+m22_61+m23_61+m24_61+m25_61+m26_61+m27_61+m28_61+m29_61+m30_61+m31_61+m32_61+m33_61+m34_61+m35_61+m36_61+m37_61+m38_61+m39_61+m40_61+m41_61+m42_61+m43_61+m44_61+m45_61+m46_61+m47_61+m48_61+m49_61+m50_61+m51_61+m52_61+m53_61+m54_61+m55_61+m56_61+m57_61+m58_61+m59_61+m60_61+m61_61+m62_61+m63_61+m64_61+m65_61+m66_61+m67_61+m68_61+m69_61+m70_61+m71_61+m72_61+m73_61+m74_61+m75_61+m76_61+m77_61+m78_61+m79_61+m80_61+m81_61+m82_61+m83_61+m84_61+m85_61+m86_61+m87_61+m88_61+m89_61+m90_61+m91_61+m92_61+m93_61+m94_61+m95_61+m96_61+m97_61+m98_61+m99_61+m100_61+m101_61+m102_61+m103_61+m104_61+m105_61+m106_61+m107_61+m108_61+m109_61+m110_61+m111_61+m112_61+m113_61+m114_61+m115_61+m116_61+m117_61+m118_61+m119_61+m120_61+m121_61+m122_61+m123_61+m124_61+m125_61+m126_61+m127_61+m128_61+m129_61+m130_61+m131_61+m132_61+m133_61+m134_61+m135_61+m136_61+m137_61+m138_61+m139_61+m140_61+m141_61+m142_61+m143_61+m144_61+m145_61+m146_61+m147_61+m148_61+m149_61+m150_61+m151_61+m152_61+m153_61+m154_61+m155_61+m156_61+m157_61+m158_61+m159_61+m160_61+m161_61+m162_61+m163_61+m164_61+m165_61+m166_61+m167_61+m168_61+m169_61+m170_61+m171_61+m172_61+m173_61+m174_61+m175_61+m176_61+m177_61+m178_61+m179_61+m180_61+m181_61+m182_61+m183_61+m184_61+m185_61+m186_61+m187_61+m188_61+m189_61+m190_61+m191_61+m192_61+m193_61+m194_61+m195_61+m196_61+m197_61+m198_61+m199_61+m200_61+m201_61+m202_61+m203_61+m204_61+m205_61+m206_61+m207_61+m208_61+m209_61+m210_61+m211_61+m212_61+m213_61+m214_61+m215_61+m216_61+m217_61+m218_61+m219_61+m220_61+m221_61+m222_61+m223_61+m224_61+m225_61+m226_61+m227_61+m228_61+m229_61+m230_61+m231_61+m232_61+m233_61+m234_61+m235_61+m236_61+m237_61+m238_61+m239_61+m240_61+m241_61+m242_61+m243_61+m244_61+m245_61+m246_61+m247_61+m248_61+m249_61+m250_61+m251_61+m252_61+m253_61+m254_61+m255_61+m256_61+m257_61+m258_61+m259_61+m260_61+m261_61+m262_61+m263_61+b61;
   assign out62 = m1_62+m2_62+m3_62+m4_62+m5_62+m6_62+m7_62+m8_62+m9_62+m10_62+m11_62+m12_62+m13_62+m14_62+m15_62+m16_62+m17_62+m18_62+m19_62+m20_62+m21_62+m22_62+m23_62+m24_62+m25_62+m26_62+m27_62+m28_62+m29_62+m30_62+m31_62+m32_62+m33_62+m34_62+m35_62+m36_62+m37_62+m38_62+m39_62+m40_62+m41_62+m42_62+m43_62+m44_62+m45_62+m46_62+m47_62+m48_62+m49_62+m50_62+m51_62+m52_62+m53_62+m54_62+m55_62+m56_62+m57_62+m58_62+m59_62+m60_62+m61_62+m62_62+m63_62+m64_62+m65_62+m66_62+m67_62+m68_62+m69_62+m70_62+m71_62+m72_62+m73_62+m74_62+m75_62+m76_62+m77_62+m78_62+m79_62+m80_62+m81_62+m82_62+m83_62+m84_62+m85_62+m86_62+m87_62+m88_62+m89_62+m90_62+m91_62+m92_62+m93_62+m94_62+m95_62+m96_62+m97_62+m98_62+m99_62+m100_62+m101_62+m102_62+m103_62+m104_62+m105_62+m106_62+m107_62+m108_62+m109_62+m110_62+m111_62+m112_62+m113_62+m114_62+m115_62+m116_62+m117_62+m118_62+m119_62+m120_62+m121_62+m122_62+m123_62+m124_62+m125_62+m126_62+m127_62+m128_62+m129_62+m130_62+m131_62+m132_62+m133_62+m134_62+m135_62+m136_62+m137_62+m138_62+m139_62+m140_62+m141_62+m142_62+m143_62+m144_62+m145_62+m146_62+m147_62+m148_62+m149_62+m150_62+m151_62+m152_62+m153_62+m154_62+m155_62+m156_62+m157_62+m158_62+m159_62+m160_62+m161_62+m162_62+m163_62+m164_62+m165_62+m166_62+m167_62+m168_62+m169_62+m170_62+m171_62+m172_62+m173_62+m174_62+m175_62+m176_62+m177_62+m178_62+m179_62+m180_62+m181_62+m182_62+m183_62+m184_62+m185_62+m186_62+m187_62+m188_62+m189_62+m190_62+m191_62+m192_62+m193_62+m194_62+m195_62+m196_62+m197_62+m198_62+m199_62+m200_62+m201_62+m202_62+m203_62+m204_62+m205_62+m206_62+m207_62+m208_62+m209_62+m210_62+m211_62+m212_62+m213_62+m214_62+m215_62+m216_62+m217_62+m218_62+m219_62+m220_62+m221_62+m222_62+m223_62+m224_62+m225_62+m226_62+m227_62+m228_62+m229_62+m230_62+m231_62+m232_62+m233_62+m234_62+m235_62+m236_62+m237_62+m238_62+m239_62+m240_62+m241_62+m242_62+m243_62+m244_62+m245_62+m246_62+m247_62+m248_62+m249_62+m250_62+m251_62+m252_62+m253_62+m254_62+m255_62+m256_62+m257_62+m258_62+m259_62+m260_62+m261_62+m262_62+m263_62+b62;
   assign out63 = m1_63+m2_63+m3_63+m4_63+m5_63+m6_63+m7_63+m8_63+m9_63+m10_63+m11_63+m12_63+m13_63+m14_63+m15_63+m16_63+m17_63+m18_63+m19_63+m20_63+m21_63+m22_63+m23_63+m24_63+m25_63+m26_63+m27_63+m28_63+m29_63+m30_63+m31_63+m32_63+m33_63+m34_63+m35_63+m36_63+m37_63+m38_63+m39_63+m40_63+m41_63+m42_63+m43_63+m44_63+m45_63+m46_63+m47_63+m48_63+m49_63+m50_63+m51_63+m52_63+m53_63+m54_63+m55_63+m56_63+m57_63+m58_63+m59_63+m60_63+m61_63+m62_63+m63_63+m64_63+m65_63+m66_63+m67_63+m68_63+m69_63+m70_63+m71_63+m72_63+m73_63+m74_63+m75_63+m76_63+m77_63+m78_63+m79_63+m80_63+m81_63+m82_63+m83_63+m84_63+m85_63+m86_63+m87_63+m88_63+m89_63+m90_63+m91_63+m92_63+m93_63+m94_63+m95_63+m96_63+m97_63+m98_63+m99_63+m100_63+m101_63+m102_63+m103_63+m104_63+m105_63+m106_63+m107_63+m108_63+m109_63+m110_63+m111_63+m112_63+m113_63+m114_63+m115_63+m116_63+m117_63+m118_63+m119_63+m120_63+m121_63+m122_63+m123_63+m124_63+m125_63+m126_63+m127_63+m128_63+m129_63+m130_63+m131_63+m132_63+m133_63+m134_63+m135_63+m136_63+m137_63+m138_63+m139_63+m140_63+m141_63+m142_63+m143_63+m144_63+m145_63+m146_63+m147_63+m148_63+m149_63+m150_63+m151_63+m152_63+m153_63+m154_63+m155_63+m156_63+m157_63+m158_63+m159_63+m160_63+m161_63+m162_63+m163_63+m164_63+m165_63+m166_63+m167_63+m168_63+m169_63+m170_63+m171_63+m172_63+m173_63+m174_63+m175_63+m176_63+m177_63+m178_63+m179_63+m180_63+m181_63+m182_63+m183_63+m184_63+m185_63+m186_63+m187_63+m188_63+m189_63+m190_63+m191_63+m192_63+m193_63+m194_63+m195_63+m196_63+m197_63+m198_63+m199_63+m200_63+m201_63+m202_63+m203_63+m204_63+m205_63+m206_63+m207_63+m208_63+m209_63+m210_63+m211_63+m212_63+m213_63+m214_63+m215_63+m216_63+m217_63+m218_63+m219_63+m220_63+m221_63+m222_63+m223_63+m224_63+m225_63+m226_63+m227_63+m228_63+m229_63+m230_63+m231_63+m232_63+m233_63+m234_63+m235_63+m236_63+m237_63+m238_63+m239_63+m240_63+m241_63+m242_63+m243_63+m244_63+m245_63+m246_63+m247_63+m248_63+m249_63+m250_63+m251_63+m252_63+m253_63+m254_63+m255_63+m256_63+m257_63+m258_63+m259_63+m260_63+m261_63+m262_63+m263_63+b63;
   assign out64 = m1_64+m2_64+m3_64+m4_64+m5_64+m6_64+m7_64+m8_64+m9_64+m10_64+m11_64+m12_64+m13_64+m14_64+m15_64+m16_64+m17_64+m18_64+m19_64+m20_64+m21_64+m22_64+m23_64+m24_64+m25_64+m26_64+m27_64+m28_64+m29_64+m30_64+m31_64+m32_64+m33_64+m34_64+m35_64+m36_64+m37_64+m38_64+m39_64+m40_64+m41_64+m42_64+m43_64+m44_64+m45_64+m46_64+m47_64+m48_64+m49_64+m50_64+m51_64+m52_64+m53_64+m54_64+m55_64+m56_64+m57_64+m58_64+m59_64+m60_64+m61_64+m62_64+m63_64+m64_64+m65_64+m66_64+m67_64+m68_64+m69_64+m70_64+m71_64+m72_64+m73_64+m74_64+m75_64+m76_64+m77_64+m78_64+m79_64+m80_64+m81_64+m82_64+m83_64+m84_64+m85_64+m86_64+m87_64+m88_64+m89_64+m90_64+m91_64+m92_64+m93_64+m94_64+m95_64+m96_64+m97_64+m98_64+m99_64+m100_64+m101_64+m102_64+m103_64+m104_64+m105_64+m106_64+m107_64+m108_64+m109_64+m110_64+m111_64+m112_64+m113_64+m114_64+m115_64+m116_64+m117_64+m118_64+m119_64+m120_64+m121_64+m122_64+m123_64+m124_64+m125_64+m126_64+m127_64+m128_64+m129_64+m130_64+m131_64+m132_64+m133_64+m134_64+m135_64+m136_64+m137_64+m138_64+m139_64+m140_64+m141_64+m142_64+m143_64+m144_64+m145_64+m146_64+m147_64+m148_64+m149_64+m150_64+m151_64+m152_64+m153_64+m154_64+m155_64+m156_64+m157_64+m158_64+m159_64+m160_64+m161_64+m162_64+m163_64+m164_64+m165_64+m166_64+m167_64+m168_64+m169_64+m170_64+m171_64+m172_64+m173_64+m174_64+m175_64+m176_64+m177_64+m178_64+m179_64+m180_64+m181_64+m182_64+m183_64+m184_64+m185_64+m186_64+m187_64+m188_64+m189_64+m190_64+m191_64+m192_64+m193_64+m194_64+m195_64+m196_64+m197_64+m198_64+m199_64+m200_64+m201_64+m202_64+m203_64+m204_64+m205_64+m206_64+m207_64+m208_64+m209_64+m210_64+m211_64+m212_64+m213_64+m214_64+m215_64+m216_64+m217_64+m218_64+m219_64+m220_64+m221_64+m222_64+m223_64+m224_64+m225_64+m226_64+m227_64+m228_64+m229_64+m230_64+m231_64+m232_64+m233_64+m234_64+m235_64+m236_64+m237_64+m238_64+m239_64+m240_64+m241_64+m242_64+m243_64+m244_64+m245_64+m246_64+m247_64+m248_64+m249_64+m250_64+m251_64+m252_64+m253_64+m254_64+m255_64+m256_64+m257_64+m258_64+m259_64+m260_64+m261_64+m262_64+m263_64+b64;
   assign out65 = m1_65+m2_65+m3_65+m4_65+m5_65+m6_65+m7_65+m8_65+m9_65+m10_65+m11_65+m12_65+m13_65+m14_65+m15_65+m16_65+m17_65+m18_65+m19_65+m20_65+m21_65+m22_65+m23_65+m24_65+m25_65+m26_65+m27_65+m28_65+m29_65+m30_65+m31_65+m32_65+m33_65+m34_65+m35_65+m36_65+m37_65+m38_65+m39_65+m40_65+m41_65+m42_65+m43_65+m44_65+m45_65+m46_65+m47_65+m48_65+m49_65+m50_65+m51_65+m52_65+m53_65+m54_65+m55_65+m56_65+m57_65+m58_65+m59_65+m60_65+m61_65+m62_65+m63_65+m64_65+m65_65+m66_65+m67_65+m68_65+m69_65+m70_65+m71_65+m72_65+m73_65+m74_65+m75_65+m76_65+m77_65+m78_65+m79_65+m80_65+m81_65+m82_65+m83_65+m84_65+m85_65+m86_65+m87_65+m88_65+m89_65+m90_65+m91_65+m92_65+m93_65+m94_65+m95_65+m96_65+m97_65+m98_65+m99_65+m100_65+m101_65+m102_65+m103_65+m104_65+m105_65+m106_65+m107_65+m108_65+m109_65+m110_65+m111_65+m112_65+m113_65+m114_65+m115_65+m116_65+m117_65+m118_65+m119_65+m120_65+m121_65+m122_65+m123_65+m124_65+m125_65+m126_65+m127_65+m128_65+m129_65+m130_65+m131_65+m132_65+m133_65+m134_65+m135_65+m136_65+m137_65+m138_65+m139_65+m140_65+m141_65+m142_65+m143_65+m144_65+m145_65+m146_65+m147_65+m148_65+m149_65+m150_65+m151_65+m152_65+m153_65+m154_65+m155_65+m156_65+m157_65+m158_65+m159_65+m160_65+m161_65+m162_65+m163_65+m164_65+m165_65+m166_65+m167_65+m168_65+m169_65+m170_65+m171_65+m172_65+m173_65+m174_65+m175_65+m176_65+m177_65+m178_65+m179_65+m180_65+m181_65+m182_65+m183_65+m184_65+m185_65+m186_65+m187_65+m188_65+m189_65+m190_65+m191_65+m192_65+m193_65+m194_65+m195_65+m196_65+m197_65+m198_65+m199_65+m200_65+m201_65+m202_65+m203_65+m204_65+m205_65+m206_65+m207_65+m208_65+m209_65+m210_65+m211_65+m212_65+m213_65+m214_65+m215_65+m216_65+m217_65+m218_65+m219_65+m220_65+m221_65+m222_65+m223_65+m224_65+m225_65+m226_65+m227_65+m228_65+m229_65+m230_65+m231_65+m232_65+m233_65+m234_65+m235_65+m236_65+m237_65+m238_65+m239_65+m240_65+m241_65+m242_65+m243_65+m244_65+m245_65+m246_65+m247_65+m248_65+m249_65+m250_65+m251_65+m252_65+m253_65+m254_65+m255_65+m256_65+m257_65+m258_65+m259_65+m260_65+m261_65+m262_65+m263_65+b65;
   assign out66 = m1_66+m2_66+m3_66+m4_66+m5_66+m6_66+m7_66+m8_66+m9_66+m10_66+m11_66+m12_66+m13_66+m14_66+m15_66+m16_66+m17_66+m18_66+m19_66+m20_66+m21_66+m22_66+m23_66+m24_66+m25_66+m26_66+m27_66+m28_66+m29_66+m30_66+m31_66+m32_66+m33_66+m34_66+m35_66+m36_66+m37_66+m38_66+m39_66+m40_66+m41_66+m42_66+m43_66+m44_66+m45_66+m46_66+m47_66+m48_66+m49_66+m50_66+m51_66+m52_66+m53_66+m54_66+m55_66+m56_66+m57_66+m58_66+m59_66+m60_66+m61_66+m62_66+m63_66+m64_66+m65_66+m66_66+m67_66+m68_66+m69_66+m70_66+m71_66+m72_66+m73_66+m74_66+m75_66+m76_66+m77_66+m78_66+m79_66+m80_66+m81_66+m82_66+m83_66+m84_66+m85_66+m86_66+m87_66+m88_66+m89_66+m90_66+m91_66+m92_66+m93_66+m94_66+m95_66+m96_66+m97_66+m98_66+m99_66+m100_66+m101_66+m102_66+m103_66+m104_66+m105_66+m106_66+m107_66+m108_66+m109_66+m110_66+m111_66+m112_66+m113_66+m114_66+m115_66+m116_66+m117_66+m118_66+m119_66+m120_66+m121_66+m122_66+m123_66+m124_66+m125_66+m126_66+m127_66+m128_66+m129_66+m130_66+m131_66+m132_66+m133_66+m134_66+m135_66+m136_66+m137_66+m138_66+m139_66+m140_66+m141_66+m142_66+m143_66+m144_66+m145_66+m146_66+m147_66+m148_66+m149_66+m150_66+m151_66+m152_66+m153_66+m154_66+m155_66+m156_66+m157_66+m158_66+m159_66+m160_66+m161_66+m162_66+m163_66+m164_66+m165_66+m166_66+m167_66+m168_66+m169_66+m170_66+m171_66+m172_66+m173_66+m174_66+m175_66+m176_66+m177_66+m178_66+m179_66+m180_66+m181_66+m182_66+m183_66+m184_66+m185_66+m186_66+m187_66+m188_66+m189_66+m190_66+m191_66+m192_66+m193_66+m194_66+m195_66+m196_66+m197_66+m198_66+m199_66+m200_66+m201_66+m202_66+m203_66+m204_66+m205_66+m206_66+m207_66+m208_66+m209_66+m210_66+m211_66+m212_66+m213_66+m214_66+m215_66+m216_66+m217_66+m218_66+m219_66+m220_66+m221_66+m222_66+m223_66+m224_66+m225_66+m226_66+m227_66+m228_66+m229_66+m230_66+m231_66+m232_66+m233_66+m234_66+m235_66+m236_66+m237_66+m238_66+m239_66+m240_66+m241_66+m242_66+m243_66+m244_66+m245_66+m246_66+m247_66+m248_66+m249_66+m250_66+m251_66+m252_66+m253_66+m254_66+m255_66+m256_66+m257_66+m258_66+m259_66+m260_66+m261_66+m262_66+m263_66+b66;
   assign out67 = m1_67+m2_67+m3_67+m4_67+m5_67+m6_67+m7_67+m8_67+m9_67+m10_67+m11_67+m12_67+m13_67+m14_67+m15_67+m16_67+m17_67+m18_67+m19_67+m20_67+m21_67+m22_67+m23_67+m24_67+m25_67+m26_67+m27_67+m28_67+m29_67+m30_67+m31_67+m32_67+m33_67+m34_67+m35_67+m36_67+m37_67+m38_67+m39_67+m40_67+m41_67+m42_67+m43_67+m44_67+m45_67+m46_67+m47_67+m48_67+m49_67+m50_67+m51_67+m52_67+m53_67+m54_67+m55_67+m56_67+m57_67+m58_67+m59_67+m60_67+m61_67+m62_67+m63_67+m64_67+m65_67+m66_67+m67_67+m68_67+m69_67+m70_67+m71_67+m72_67+m73_67+m74_67+m75_67+m76_67+m77_67+m78_67+m79_67+m80_67+m81_67+m82_67+m83_67+m84_67+m85_67+m86_67+m87_67+m88_67+m89_67+m90_67+m91_67+m92_67+m93_67+m94_67+m95_67+m96_67+m97_67+m98_67+m99_67+m100_67+m101_67+m102_67+m103_67+m104_67+m105_67+m106_67+m107_67+m108_67+m109_67+m110_67+m111_67+m112_67+m113_67+m114_67+m115_67+m116_67+m117_67+m118_67+m119_67+m120_67+m121_67+m122_67+m123_67+m124_67+m125_67+m126_67+m127_67+m128_67+m129_67+m130_67+m131_67+m132_67+m133_67+m134_67+m135_67+m136_67+m137_67+m138_67+m139_67+m140_67+m141_67+m142_67+m143_67+m144_67+m145_67+m146_67+m147_67+m148_67+m149_67+m150_67+m151_67+m152_67+m153_67+m154_67+m155_67+m156_67+m157_67+m158_67+m159_67+m160_67+m161_67+m162_67+m163_67+m164_67+m165_67+m166_67+m167_67+m168_67+m169_67+m170_67+m171_67+m172_67+m173_67+m174_67+m175_67+m176_67+m177_67+m178_67+m179_67+m180_67+m181_67+m182_67+m183_67+m184_67+m185_67+m186_67+m187_67+m188_67+m189_67+m190_67+m191_67+m192_67+m193_67+m194_67+m195_67+m196_67+m197_67+m198_67+m199_67+m200_67+m201_67+m202_67+m203_67+m204_67+m205_67+m206_67+m207_67+m208_67+m209_67+m210_67+m211_67+m212_67+m213_67+m214_67+m215_67+m216_67+m217_67+m218_67+m219_67+m220_67+m221_67+m222_67+m223_67+m224_67+m225_67+m226_67+m227_67+m228_67+m229_67+m230_67+m231_67+m232_67+m233_67+m234_67+m235_67+m236_67+m237_67+m238_67+m239_67+m240_67+m241_67+m242_67+m243_67+m244_67+m245_67+m246_67+m247_67+m248_67+m249_67+m250_67+m251_67+m252_67+m253_67+m254_67+m255_67+m256_67+m257_67+m258_67+m259_67+m260_67+m261_67+m262_67+m263_67+b67;
   assign out68 = m1_68+m2_68+m3_68+m4_68+m5_68+m6_68+m7_68+m8_68+m9_68+m10_68+m11_68+m12_68+m13_68+m14_68+m15_68+m16_68+m17_68+m18_68+m19_68+m20_68+m21_68+m22_68+m23_68+m24_68+m25_68+m26_68+m27_68+m28_68+m29_68+m30_68+m31_68+m32_68+m33_68+m34_68+m35_68+m36_68+m37_68+m38_68+m39_68+m40_68+m41_68+m42_68+m43_68+m44_68+m45_68+m46_68+m47_68+m48_68+m49_68+m50_68+m51_68+m52_68+m53_68+m54_68+m55_68+m56_68+m57_68+m58_68+m59_68+m60_68+m61_68+m62_68+m63_68+m64_68+m65_68+m66_68+m67_68+m68_68+m69_68+m70_68+m71_68+m72_68+m73_68+m74_68+m75_68+m76_68+m77_68+m78_68+m79_68+m80_68+m81_68+m82_68+m83_68+m84_68+m85_68+m86_68+m87_68+m88_68+m89_68+m90_68+m91_68+m92_68+m93_68+m94_68+m95_68+m96_68+m97_68+m98_68+m99_68+m100_68+m101_68+m102_68+m103_68+m104_68+m105_68+m106_68+m107_68+m108_68+m109_68+m110_68+m111_68+m112_68+m113_68+m114_68+m115_68+m116_68+m117_68+m118_68+m119_68+m120_68+m121_68+m122_68+m123_68+m124_68+m125_68+m126_68+m127_68+m128_68+m129_68+m130_68+m131_68+m132_68+m133_68+m134_68+m135_68+m136_68+m137_68+m138_68+m139_68+m140_68+m141_68+m142_68+m143_68+m144_68+m145_68+m146_68+m147_68+m148_68+m149_68+m150_68+m151_68+m152_68+m153_68+m154_68+m155_68+m156_68+m157_68+m158_68+m159_68+m160_68+m161_68+m162_68+m163_68+m164_68+m165_68+m166_68+m167_68+m168_68+m169_68+m170_68+m171_68+m172_68+m173_68+m174_68+m175_68+m176_68+m177_68+m178_68+m179_68+m180_68+m181_68+m182_68+m183_68+m184_68+m185_68+m186_68+m187_68+m188_68+m189_68+m190_68+m191_68+m192_68+m193_68+m194_68+m195_68+m196_68+m197_68+m198_68+m199_68+m200_68+m201_68+m202_68+m203_68+m204_68+m205_68+m206_68+m207_68+m208_68+m209_68+m210_68+m211_68+m212_68+m213_68+m214_68+m215_68+m216_68+m217_68+m218_68+m219_68+m220_68+m221_68+m222_68+m223_68+m224_68+m225_68+m226_68+m227_68+m228_68+m229_68+m230_68+m231_68+m232_68+m233_68+m234_68+m235_68+m236_68+m237_68+m238_68+m239_68+m240_68+m241_68+m242_68+m243_68+m244_68+m245_68+m246_68+m247_68+m248_68+m249_68+m250_68+m251_68+m252_68+m253_68+m254_68+m255_68+m256_68+m257_68+m258_68+m259_68+m260_68+m261_68+m262_68+m263_68+b68;
   assign out69 = m1_69+m2_69+m3_69+m4_69+m5_69+m6_69+m7_69+m8_69+m9_69+m10_69+m11_69+m12_69+m13_69+m14_69+m15_69+m16_69+m17_69+m18_69+m19_69+m20_69+m21_69+m22_69+m23_69+m24_69+m25_69+m26_69+m27_69+m28_69+m29_69+m30_69+m31_69+m32_69+m33_69+m34_69+m35_69+m36_69+m37_69+m38_69+m39_69+m40_69+m41_69+m42_69+m43_69+m44_69+m45_69+m46_69+m47_69+m48_69+m49_69+m50_69+m51_69+m52_69+m53_69+m54_69+m55_69+m56_69+m57_69+m58_69+m59_69+m60_69+m61_69+m62_69+m63_69+m64_69+m65_69+m66_69+m67_69+m68_69+m69_69+m70_69+m71_69+m72_69+m73_69+m74_69+m75_69+m76_69+m77_69+m78_69+m79_69+m80_69+m81_69+m82_69+m83_69+m84_69+m85_69+m86_69+m87_69+m88_69+m89_69+m90_69+m91_69+m92_69+m93_69+m94_69+m95_69+m96_69+m97_69+m98_69+m99_69+m100_69+m101_69+m102_69+m103_69+m104_69+m105_69+m106_69+m107_69+m108_69+m109_69+m110_69+m111_69+m112_69+m113_69+m114_69+m115_69+m116_69+m117_69+m118_69+m119_69+m120_69+m121_69+m122_69+m123_69+m124_69+m125_69+m126_69+m127_69+m128_69+m129_69+m130_69+m131_69+m132_69+m133_69+m134_69+m135_69+m136_69+m137_69+m138_69+m139_69+m140_69+m141_69+m142_69+m143_69+m144_69+m145_69+m146_69+m147_69+m148_69+m149_69+m150_69+m151_69+m152_69+m153_69+m154_69+m155_69+m156_69+m157_69+m158_69+m159_69+m160_69+m161_69+m162_69+m163_69+m164_69+m165_69+m166_69+m167_69+m168_69+m169_69+m170_69+m171_69+m172_69+m173_69+m174_69+m175_69+m176_69+m177_69+m178_69+m179_69+m180_69+m181_69+m182_69+m183_69+m184_69+m185_69+m186_69+m187_69+m188_69+m189_69+m190_69+m191_69+m192_69+m193_69+m194_69+m195_69+m196_69+m197_69+m198_69+m199_69+m200_69+m201_69+m202_69+m203_69+m204_69+m205_69+m206_69+m207_69+m208_69+m209_69+m210_69+m211_69+m212_69+m213_69+m214_69+m215_69+m216_69+m217_69+m218_69+m219_69+m220_69+m221_69+m222_69+m223_69+m224_69+m225_69+m226_69+m227_69+m228_69+m229_69+m230_69+m231_69+m232_69+m233_69+m234_69+m235_69+m236_69+m237_69+m238_69+m239_69+m240_69+m241_69+m242_69+m243_69+m244_69+m245_69+m246_69+m247_69+m248_69+m249_69+m250_69+m251_69+m252_69+m253_69+m254_69+m255_69+m256_69+m257_69+m258_69+m259_69+m260_69+m261_69+m262_69+m263_69+b69;
   assign out70 = m1_70+m2_70+m3_70+m4_70+m5_70+m6_70+m7_70+m8_70+m9_70+m10_70+m11_70+m12_70+m13_70+m14_70+m15_70+m16_70+m17_70+m18_70+m19_70+m20_70+m21_70+m22_70+m23_70+m24_70+m25_70+m26_70+m27_70+m28_70+m29_70+m30_70+m31_70+m32_70+m33_70+m34_70+m35_70+m36_70+m37_70+m38_70+m39_70+m40_70+m41_70+m42_70+m43_70+m44_70+m45_70+m46_70+m47_70+m48_70+m49_70+m50_70+m51_70+m52_70+m53_70+m54_70+m55_70+m56_70+m57_70+m58_70+m59_70+m60_70+m61_70+m62_70+m63_70+m64_70+m65_70+m66_70+m67_70+m68_70+m69_70+m70_70+m71_70+m72_70+m73_70+m74_70+m75_70+m76_70+m77_70+m78_70+m79_70+m80_70+m81_70+m82_70+m83_70+m84_70+m85_70+m86_70+m87_70+m88_70+m89_70+m90_70+m91_70+m92_70+m93_70+m94_70+m95_70+m96_70+m97_70+m98_70+m99_70+m100_70+m101_70+m102_70+m103_70+m104_70+m105_70+m106_70+m107_70+m108_70+m109_70+m110_70+m111_70+m112_70+m113_70+m114_70+m115_70+m116_70+m117_70+m118_70+m119_70+m120_70+m121_70+m122_70+m123_70+m124_70+m125_70+m126_70+m127_70+m128_70+m129_70+m130_70+m131_70+m132_70+m133_70+m134_70+m135_70+m136_70+m137_70+m138_70+m139_70+m140_70+m141_70+m142_70+m143_70+m144_70+m145_70+m146_70+m147_70+m148_70+m149_70+m150_70+m151_70+m152_70+m153_70+m154_70+m155_70+m156_70+m157_70+m158_70+m159_70+m160_70+m161_70+m162_70+m163_70+m164_70+m165_70+m166_70+m167_70+m168_70+m169_70+m170_70+m171_70+m172_70+m173_70+m174_70+m175_70+m176_70+m177_70+m178_70+m179_70+m180_70+m181_70+m182_70+m183_70+m184_70+m185_70+m186_70+m187_70+m188_70+m189_70+m190_70+m191_70+m192_70+m193_70+m194_70+m195_70+m196_70+m197_70+m198_70+m199_70+m200_70+m201_70+m202_70+m203_70+m204_70+m205_70+m206_70+m207_70+m208_70+m209_70+m210_70+m211_70+m212_70+m213_70+m214_70+m215_70+m216_70+m217_70+m218_70+m219_70+m220_70+m221_70+m222_70+m223_70+m224_70+m225_70+m226_70+m227_70+m228_70+m229_70+m230_70+m231_70+m232_70+m233_70+m234_70+m235_70+m236_70+m237_70+m238_70+m239_70+m240_70+m241_70+m242_70+m243_70+m244_70+m245_70+m246_70+m247_70+m248_70+m249_70+m250_70+m251_70+m252_70+m253_70+m254_70+m255_70+m256_70+m257_70+m258_70+m259_70+m260_70+m261_70+m262_70+m263_70+b70;
   assign out71 = m1_71+m2_71+m3_71+m4_71+m5_71+m6_71+m7_71+m8_71+m9_71+m10_71+m11_71+m12_71+m13_71+m14_71+m15_71+m16_71+m17_71+m18_71+m19_71+m20_71+m21_71+m22_71+m23_71+m24_71+m25_71+m26_71+m27_71+m28_71+m29_71+m30_71+m31_71+m32_71+m33_71+m34_71+m35_71+m36_71+m37_71+m38_71+m39_71+m40_71+m41_71+m42_71+m43_71+m44_71+m45_71+m46_71+m47_71+m48_71+m49_71+m50_71+m51_71+m52_71+m53_71+m54_71+m55_71+m56_71+m57_71+m58_71+m59_71+m60_71+m61_71+m62_71+m63_71+m64_71+m65_71+m66_71+m67_71+m68_71+m69_71+m70_71+m71_71+m72_71+m73_71+m74_71+m75_71+m76_71+m77_71+m78_71+m79_71+m80_71+m81_71+m82_71+m83_71+m84_71+m85_71+m86_71+m87_71+m88_71+m89_71+m90_71+m91_71+m92_71+m93_71+m94_71+m95_71+m96_71+m97_71+m98_71+m99_71+m100_71+m101_71+m102_71+m103_71+m104_71+m105_71+m106_71+m107_71+m108_71+m109_71+m110_71+m111_71+m112_71+m113_71+m114_71+m115_71+m116_71+m117_71+m118_71+m119_71+m120_71+m121_71+m122_71+m123_71+m124_71+m125_71+m126_71+m127_71+m128_71+m129_71+m130_71+m131_71+m132_71+m133_71+m134_71+m135_71+m136_71+m137_71+m138_71+m139_71+m140_71+m141_71+m142_71+m143_71+m144_71+m145_71+m146_71+m147_71+m148_71+m149_71+m150_71+m151_71+m152_71+m153_71+m154_71+m155_71+m156_71+m157_71+m158_71+m159_71+m160_71+m161_71+m162_71+m163_71+m164_71+m165_71+m166_71+m167_71+m168_71+m169_71+m170_71+m171_71+m172_71+m173_71+m174_71+m175_71+m176_71+m177_71+m178_71+m179_71+m180_71+m181_71+m182_71+m183_71+m184_71+m185_71+m186_71+m187_71+m188_71+m189_71+m190_71+m191_71+m192_71+m193_71+m194_71+m195_71+m196_71+m197_71+m198_71+m199_71+m200_71+m201_71+m202_71+m203_71+m204_71+m205_71+m206_71+m207_71+m208_71+m209_71+m210_71+m211_71+m212_71+m213_71+m214_71+m215_71+m216_71+m217_71+m218_71+m219_71+m220_71+m221_71+m222_71+m223_71+m224_71+m225_71+m226_71+m227_71+m228_71+m229_71+m230_71+m231_71+m232_71+m233_71+m234_71+m235_71+m236_71+m237_71+m238_71+m239_71+m240_71+m241_71+m242_71+m243_71+m244_71+m245_71+m246_71+m247_71+m248_71+m249_71+m250_71+m251_71+m252_71+m253_71+m254_71+m255_71+m256_71+m257_71+m258_71+m259_71+m260_71+m261_71+m262_71+m263_71+b71;
   assign out72 = m1_72+m2_72+m3_72+m4_72+m5_72+m6_72+m7_72+m8_72+m9_72+m10_72+m11_72+m12_72+m13_72+m14_72+m15_72+m16_72+m17_72+m18_72+m19_72+m20_72+m21_72+m22_72+m23_72+m24_72+m25_72+m26_72+m27_72+m28_72+m29_72+m30_72+m31_72+m32_72+m33_72+m34_72+m35_72+m36_72+m37_72+m38_72+m39_72+m40_72+m41_72+m42_72+m43_72+m44_72+m45_72+m46_72+m47_72+m48_72+m49_72+m50_72+m51_72+m52_72+m53_72+m54_72+m55_72+m56_72+m57_72+m58_72+m59_72+m60_72+m61_72+m62_72+m63_72+m64_72+m65_72+m66_72+m67_72+m68_72+m69_72+m70_72+m71_72+m72_72+m73_72+m74_72+m75_72+m76_72+m77_72+m78_72+m79_72+m80_72+m81_72+m82_72+m83_72+m84_72+m85_72+m86_72+m87_72+m88_72+m89_72+m90_72+m91_72+m92_72+m93_72+m94_72+m95_72+m96_72+m97_72+m98_72+m99_72+m100_72+m101_72+m102_72+m103_72+m104_72+m105_72+m106_72+m107_72+m108_72+m109_72+m110_72+m111_72+m112_72+m113_72+m114_72+m115_72+m116_72+m117_72+m118_72+m119_72+m120_72+m121_72+m122_72+m123_72+m124_72+m125_72+m126_72+m127_72+m128_72+m129_72+m130_72+m131_72+m132_72+m133_72+m134_72+m135_72+m136_72+m137_72+m138_72+m139_72+m140_72+m141_72+m142_72+m143_72+m144_72+m145_72+m146_72+m147_72+m148_72+m149_72+m150_72+m151_72+m152_72+m153_72+m154_72+m155_72+m156_72+m157_72+m158_72+m159_72+m160_72+m161_72+m162_72+m163_72+m164_72+m165_72+m166_72+m167_72+m168_72+m169_72+m170_72+m171_72+m172_72+m173_72+m174_72+m175_72+m176_72+m177_72+m178_72+m179_72+m180_72+m181_72+m182_72+m183_72+m184_72+m185_72+m186_72+m187_72+m188_72+m189_72+m190_72+m191_72+m192_72+m193_72+m194_72+m195_72+m196_72+m197_72+m198_72+m199_72+m200_72+m201_72+m202_72+m203_72+m204_72+m205_72+m206_72+m207_72+m208_72+m209_72+m210_72+m211_72+m212_72+m213_72+m214_72+m215_72+m216_72+m217_72+m218_72+m219_72+m220_72+m221_72+m222_72+m223_72+m224_72+m225_72+m226_72+m227_72+m228_72+m229_72+m230_72+m231_72+m232_72+m233_72+m234_72+m235_72+m236_72+m237_72+m238_72+m239_72+m240_72+m241_72+m242_72+m243_72+m244_72+m245_72+m246_72+m247_72+m248_72+m249_72+m250_72+m251_72+m252_72+m253_72+m254_72+m255_72+m256_72+m257_72+m258_72+m259_72+m260_72+m261_72+m262_72+m263_72+b72;
   assign out73 = m1_73+m2_73+m3_73+m4_73+m5_73+m6_73+m7_73+m8_73+m9_73+m10_73+m11_73+m12_73+m13_73+m14_73+m15_73+m16_73+m17_73+m18_73+m19_73+m20_73+m21_73+m22_73+m23_73+m24_73+m25_73+m26_73+m27_73+m28_73+m29_73+m30_73+m31_73+m32_73+m33_73+m34_73+m35_73+m36_73+m37_73+m38_73+m39_73+m40_73+m41_73+m42_73+m43_73+m44_73+m45_73+m46_73+m47_73+m48_73+m49_73+m50_73+m51_73+m52_73+m53_73+m54_73+m55_73+m56_73+m57_73+m58_73+m59_73+m60_73+m61_73+m62_73+m63_73+m64_73+m65_73+m66_73+m67_73+m68_73+m69_73+m70_73+m71_73+m72_73+m73_73+m74_73+m75_73+m76_73+m77_73+m78_73+m79_73+m80_73+m81_73+m82_73+m83_73+m84_73+m85_73+m86_73+m87_73+m88_73+m89_73+m90_73+m91_73+m92_73+m93_73+m94_73+m95_73+m96_73+m97_73+m98_73+m99_73+m100_73+m101_73+m102_73+m103_73+m104_73+m105_73+m106_73+m107_73+m108_73+m109_73+m110_73+m111_73+m112_73+m113_73+m114_73+m115_73+m116_73+m117_73+m118_73+m119_73+m120_73+m121_73+m122_73+m123_73+m124_73+m125_73+m126_73+m127_73+m128_73+m129_73+m130_73+m131_73+m132_73+m133_73+m134_73+m135_73+m136_73+m137_73+m138_73+m139_73+m140_73+m141_73+m142_73+m143_73+m144_73+m145_73+m146_73+m147_73+m148_73+m149_73+m150_73+m151_73+m152_73+m153_73+m154_73+m155_73+m156_73+m157_73+m158_73+m159_73+m160_73+m161_73+m162_73+m163_73+m164_73+m165_73+m166_73+m167_73+m168_73+m169_73+m170_73+m171_73+m172_73+m173_73+m174_73+m175_73+m176_73+m177_73+m178_73+m179_73+m180_73+m181_73+m182_73+m183_73+m184_73+m185_73+m186_73+m187_73+m188_73+m189_73+m190_73+m191_73+m192_73+m193_73+m194_73+m195_73+m196_73+m197_73+m198_73+m199_73+m200_73+m201_73+m202_73+m203_73+m204_73+m205_73+m206_73+m207_73+m208_73+m209_73+m210_73+m211_73+m212_73+m213_73+m214_73+m215_73+m216_73+m217_73+m218_73+m219_73+m220_73+m221_73+m222_73+m223_73+m224_73+m225_73+m226_73+m227_73+m228_73+m229_73+m230_73+m231_73+m232_73+m233_73+m234_73+m235_73+m236_73+m237_73+m238_73+m239_73+m240_73+m241_73+m242_73+m243_73+m244_73+m245_73+m246_73+m247_73+m248_73+m249_73+m250_73+m251_73+m252_73+m253_73+m254_73+m255_73+m256_73+m257_73+m258_73+m259_73+m260_73+m261_73+m262_73+m263_73+b73;
   assign out74 = m1_74+m2_74+m3_74+m4_74+m5_74+m6_74+m7_74+m8_74+m9_74+m10_74+m11_74+m12_74+m13_74+m14_74+m15_74+m16_74+m17_74+m18_74+m19_74+m20_74+m21_74+m22_74+m23_74+m24_74+m25_74+m26_74+m27_74+m28_74+m29_74+m30_74+m31_74+m32_74+m33_74+m34_74+m35_74+m36_74+m37_74+m38_74+m39_74+m40_74+m41_74+m42_74+m43_74+m44_74+m45_74+m46_74+m47_74+m48_74+m49_74+m50_74+m51_74+m52_74+m53_74+m54_74+m55_74+m56_74+m57_74+m58_74+m59_74+m60_74+m61_74+m62_74+m63_74+m64_74+m65_74+m66_74+m67_74+m68_74+m69_74+m70_74+m71_74+m72_74+m73_74+m74_74+m75_74+m76_74+m77_74+m78_74+m79_74+m80_74+m81_74+m82_74+m83_74+m84_74+m85_74+m86_74+m87_74+m88_74+m89_74+m90_74+m91_74+m92_74+m93_74+m94_74+m95_74+m96_74+m97_74+m98_74+m99_74+m100_74+m101_74+m102_74+m103_74+m104_74+m105_74+m106_74+m107_74+m108_74+m109_74+m110_74+m111_74+m112_74+m113_74+m114_74+m115_74+m116_74+m117_74+m118_74+m119_74+m120_74+m121_74+m122_74+m123_74+m124_74+m125_74+m126_74+m127_74+m128_74+m129_74+m130_74+m131_74+m132_74+m133_74+m134_74+m135_74+m136_74+m137_74+m138_74+m139_74+m140_74+m141_74+m142_74+m143_74+m144_74+m145_74+m146_74+m147_74+m148_74+m149_74+m150_74+m151_74+m152_74+m153_74+m154_74+m155_74+m156_74+m157_74+m158_74+m159_74+m160_74+m161_74+m162_74+m163_74+m164_74+m165_74+m166_74+m167_74+m168_74+m169_74+m170_74+m171_74+m172_74+m173_74+m174_74+m175_74+m176_74+m177_74+m178_74+m179_74+m180_74+m181_74+m182_74+m183_74+m184_74+m185_74+m186_74+m187_74+m188_74+m189_74+m190_74+m191_74+m192_74+m193_74+m194_74+m195_74+m196_74+m197_74+m198_74+m199_74+m200_74+m201_74+m202_74+m203_74+m204_74+m205_74+m206_74+m207_74+m208_74+m209_74+m210_74+m211_74+m212_74+m213_74+m214_74+m215_74+m216_74+m217_74+m218_74+m219_74+m220_74+m221_74+m222_74+m223_74+m224_74+m225_74+m226_74+m227_74+m228_74+m229_74+m230_74+m231_74+m232_74+m233_74+m234_74+m235_74+m236_74+m237_74+m238_74+m239_74+m240_74+m241_74+m242_74+m243_74+m244_74+m245_74+m246_74+m247_74+m248_74+m249_74+m250_74+m251_74+m252_74+m253_74+m254_74+m255_74+m256_74+m257_74+m258_74+m259_74+m260_74+m261_74+m262_74+m263_74+b74;
   assign out75 = m1_75+m2_75+m3_75+m4_75+m5_75+m6_75+m7_75+m8_75+m9_75+m10_75+m11_75+m12_75+m13_75+m14_75+m15_75+m16_75+m17_75+m18_75+m19_75+m20_75+m21_75+m22_75+m23_75+m24_75+m25_75+m26_75+m27_75+m28_75+m29_75+m30_75+m31_75+m32_75+m33_75+m34_75+m35_75+m36_75+m37_75+m38_75+m39_75+m40_75+m41_75+m42_75+m43_75+m44_75+m45_75+m46_75+m47_75+m48_75+m49_75+m50_75+m51_75+m52_75+m53_75+m54_75+m55_75+m56_75+m57_75+m58_75+m59_75+m60_75+m61_75+m62_75+m63_75+m64_75+m65_75+m66_75+m67_75+m68_75+m69_75+m70_75+m71_75+m72_75+m73_75+m74_75+m75_75+m76_75+m77_75+m78_75+m79_75+m80_75+m81_75+m82_75+m83_75+m84_75+m85_75+m86_75+m87_75+m88_75+m89_75+m90_75+m91_75+m92_75+m93_75+m94_75+m95_75+m96_75+m97_75+m98_75+m99_75+m100_75+m101_75+m102_75+m103_75+m104_75+m105_75+m106_75+m107_75+m108_75+m109_75+m110_75+m111_75+m112_75+m113_75+m114_75+m115_75+m116_75+m117_75+m118_75+m119_75+m120_75+m121_75+m122_75+m123_75+m124_75+m125_75+m126_75+m127_75+m128_75+m129_75+m130_75+m131_75+m132_75+m133_75+m134_75+m135_75+m136_75+m137_75+m138_75+m139_75+m140_75+m141_75+m142_75+m143_75+m144_75+m145_75+m146_75+m147_75+m148_75+m149_75+m150_75+m151_75+m152_75+m153_75+m154_75+m155_75+m156_75+m157_75+m158_75+m159_75+m160_75+m161_75+m162_75+m163_75+m164_75+m165_75+m166_75+m167_75+m168_75+m169_75+m170_75+m171_75+m172_75+m173_75+m174_75+m175_75+m176_75+m177_75+m178_75+m179_75+m180_75+m181_75+m182_75+m183_75+m184_75+m185_75+m186_75+m187_75+m188_75+m189_75+m190_75+m191_75+m192_75+m193_75+m194_75+m195_75+m196_75+m197_75+m198_75+m199_75+m200_75+m201_75+m202_75+m203_75+m204_75+m205_75+m206_75+m207_75+m208_75+m209_75+m210_75+m211_75+m212_75+m213_75+m214_75+m215_75+m216_75+m217_75+m218_75+m219_75+m220_75+m221_75+m222_75+m223_75+m224_75+m225_75+m226_75+m227_75+m228_75+m229_75+m230_75+m231_75+m232_75+m233_75+m234_75+m235_75+m236_75+m237_75+m238_75+m239_75+m240_75+m241_75+m242_75+m243_75+m244_75+m245_75+m246_75+m247_75+m248_75+m249_75+m250_75+m251_75+m252_75+m253_75+m254_75+m255_75+m256_75+m257_75+m258_75+m259_75+m260_75+m261_75+m262_75+m263_75+b75;
   assign out76 = m1_76+m2_76+m3_76+m4_76+m5_76+m6_76+m7_76+m8_76+m9_76+m10_76+m11_76+m12_76+m13_76+m14_76+m15_76+m16_76+m17_76+m18_76+m19_76+m20_76+m21_76+m22_76+m23_76+m24_76+m25_76+m26_76+m27_76+m28_76+m29_76+m30_76+m31_76+m32_76+m33_76+m34_76+m35_76+m36_76+m37_76+m38_76+m39_76+m40_76+m41_76+m42_76+m43_76+m44_76+m45_76+m46_76+m47_76+m48_76+m49_76+m50_76+m51_76+m52_76+m53_76+m54_76+m55_76+m56_76+m57_76+m58_76+m59_76+m60_76+m61_76+m62_76+m63_76+m64_76+m65_76+m66_76+m67_76+m68_76+m69_76+m70_76+m71_76+m72_76+m73_76+m74_76+m75_76+m76_76+m77_76+m78_76+m79_76+m80_76+m81_76+m82_76+m83_76+m84_76+m85_76+m86_76+m87_76+m88_76+m89_76+m90_76+m91_76+m92_76+m93_76+m94_76+m95_76+m96_76+m97_76+m98_76+m99_76+m100_76+m101_76+m102_76+m103_76+m104_76+m105_76+m106_76+m107_76+m108_76+m109_76+m110_76+m111_76+m112_76+m113_76+m114_76+m115_76+m116_76+m117_76+m118_76+m119_76+m120_76+m121_76+m122_76+m123_76+m124_76+m125_76+m126_76+m127_76+m128_76+m129_76+m130_76+m131_76+m132_76+m133_76+m134_76+m135_76+m136_76+m137_76+m138_76+m139_76+m140_76+m141_76+m142_76+m143_76+m144_76+m145_76+m146_76+m147_76+m148_76+m149_76+m150_76+m151_76+m152_76+m153_76+m154_76+m155_76+m156_76+m157_76+m158_76+m159_76+m160_76+m161_76+m162_76+m163_76+m164_76+m165_76+m166_76+m167_76+m168_76+m169_76+m170_76+m171_76+m172_76+m173_76+m174_76+m175_76+m176_76+m177_76+m178_76+m179_76+m180_76+m181_76+m182_76+m183_76+m184_76+m185_76+m186_76+m187_76+m188_76+m189_76+m190_76+m191_76+m192_76+m193_76+m194_76+m195_76+m196_76+m197_76+m198_76+m199_76+m200_76+m201_76+m202_76+m203_76+m204_76+m205_76+m206_76+m207_76+m208_76+m209_76+m210_76+m211_76+m212_76+m213_76+m214_76+m215_76+m216_76+m217_76+m218_76+m219_76+m220_76+m221_76+m222_76+m223_76+m224_76+m225_76+m226_76+m227_76+m228_76+m229_76+m230_76+m231_76+m232_76+m233_76+m234_76+m235_76+m236_76+m237_76+m238_76+m239_76+m240_76+m241_76+m242_76+m243_76+m244_76+m245_76+m246_76+m247_76+m248_76+m249_76+m250_76+m251_76+m252_76+m253_76+m254_76+m255_76+m256_76+m257_76+m258_76+m259_76+m260_76+m261_76+m262_76+m263_76+b76;
   assign out77 = m1_77+m2_77+m3_77+m4_77+m5_77+m6_77+m7_77+m8_77+m9_77+m10_77+m11_77+m12_77+m13_77+m14_77+m15_77+m16_77+m17_77+m18_77+m19_77+m20_77+m21_77+m22_77+m23_77+m24_77+m25_77+m26_77+m27_77+m28_77+m29_77+m30_77+m31_77+m32_77+m33_77+m34_77+m35_77+m36_77+m37_77+m38_77+m39_77+m40_77+m41_77+m42_77+m43_77+m44_77+m45_77+m46_77+m47_77+m48_77+m49_77+m50_77+m51_77+m52_77+m53_77+m54_77+m55_77+m56_77+m57_77+m58_77+m59_77+m60_77+m61_77+m62_77+m63_77+m64_77+m65_77+m66_77+m67_77+m68_77+m69_77+m70_77+m71_77+m72_77+m73_77+m74_77+m75_77+m76_77+m77_77+m78_77+m79_77+m80_77+m81_77+m82_77+m83_77+m84_77+m85_77+m86_77+m87_77+m88_77+m89_77+m90_77+m91_77+m92_77+m93_77+m94_77+m95_77+m96_77+m97_77+m98_77+m99_77+m100_77+m101_77+m102_77+m103_77+m104_77+m105_77+m106_77+m107_77+m108_77+m109_77+m110_77+m111_77+m112_77+m113_77+m114_77+m115_77+m116_77+m117_77+m118_77+m119_77+m120_77+m121_77+m122_77+m123_77+m124_77+m125_77+m126_77+m127_77+m128_77+m129_77+m130_77+m131_77+m132_77+m133_77+m134_77+m135_77+m136_77+m137_77+m138_77+m139_77+m140_77+m141_77+m142_77+m143_77+m144_77+m145_77+m146_77+m147_77+m148_77+m149_77+m150_77+m151_77+m152_77+m153_77+m154_77+m155_77+m156_77+m157_77+m158_77+m159_77+m160_77+m161_77+m162_77+m163_77+m164_77+m165_77+m166_77+m167_77+m168_77+m169_77+m170_77+m171_77+m172_77+m173_77+m174_77+m175_77+m176_77+m177_77+m178_77+m179_77+m180_77+m181_77+m182_77+m183_77+m184_77+m185_77+m186_77+m187_77+m188_77+m189_77+m190_77+m191_77+m192_77+m193_77+m194_77+m195_77+m196_77+m197_77+m198_77+m199_77+m200_77+m201_77+m202_77+m203_77+m204_77+m205_77+m206_77+m207_77+m208_77+m209_77+m210_77+m211_77+m212_77+m213_77+m214_77+m215_77+m216_77+m217_77+m218_77+m219_77+m220_77+m221_77+m222_77+m223_77+m224_77+m225_77+m226_77+m227_77+m228_77+m229_77+m230_77+m231_77+m232_77+m233_77+m234_77+m235_77+m236_77+m237_77+m238_77+m239_77+m240_77+m241_77+m242_77+m243_77+m244_77+m245_77+m246_77+m247_77+m248_77+m249_77+m250_77+m251_77+m252_77+m253_77+m254_77+m255_77+m256_77+m257_77+m258_77+m259_77+m260_77+m261_77+m262_77+m263_77+b77;
   assign out78 = m1_78+m2_78+m3_78+m4_78+m5_78+m6_78+m7_78+m8_78+m9_78+m10_78+m11_78+m12_78+m13_78+m14_78+m15_78+m16_78+m17_78+m18_78+m19_78+m20_78+m21_78+m22_78+m23_78+m24_78+m25_78+m26_78+m27_78+m28_78+m29_78+m30_78+m31_78+m32_78+m33_78+m34_78+m35_78+m36_78+m37_78+m38_78+m39_78+m40_78+m41_78+m42_78+m43_78+m44_78+m45_78+m46_78+m47_78+m48_78+m49_78+m50_78+m51_78+m52_78+m53_78+m54_78+m55_78+m56_78+m57_78+m58_78+m59_78+m60_78+m61_78+m62_78+m63_78+m64_78+m65_78+m66_78+m67_78+m68_78+m69_78+m70_78+m71_78+m72_78+m73_78+m74_78+m75_78+m76_78+m77_78+m78_78+m79_78+m80_78+m81_78+m82_78+m83_78+m84_78+m85_78+m86_78+m87_78+m88_78+m89_78+m90_78+m91_78+m92_78+m93_78+m94_78+m95_78+m96_78+m97_78+m98_78+m99_78+m100_78+m101_78+m102_78+m103_78+m104_78+m105_78+m106_78+m107_78+m108_78+m109_78+m110_78+m111_78+m112_78+m113_78+m114_78+m115_78+m116_78+m117_78+m118_78+m119_78+m120_78+m121_78+m122_78+m123_78+m124_78+m125_78+m126_78+m127_78+m128_78+m129_78+m130_78+m131_78+m132_78+m133_78+m134_78+m135_78+m136_78+m137_78+m138_78+m139_78+m140_78+m141_78+m142_78+m143_78+m144_78+m145_78+m146_78+m147_78+m148_78+m149_78+m150_78+m151_78+m152_78+m153_78+m154_78+m155_78+m156_78+m157_78+m158_78+m159_78+m160_78+m161_78+m162_78+m163_78+m164_78+m165_78+m166_78+m167_78+m168_78+m169_78+m170_78+m171_78+m172_78+m173_78+m174_78+m175_78+m176_78+m177_78+m178_78+m179_78+m180_78+m181_78+m182_78+m183_78+m184_78+m185_78+m186_78+m187_78+m188_78+m189_78+m190_78+m191_78+m192_78+m193_78+m194_78+m195_78+m196_78+m197_78+m198_78+m199_78+m200_78+m201_78+m202_78+m203_78+m204_78+m205_78+m206_78+m207_78+m208_78+m209_78+m210_78+m211_78+m212_78+m213_78+m214_78+m215_78+m216_78+m217_78+m218_78+m219_78+m220_78+m221_78+m222_78+m223_78+m224_78+m225_78+m226_78+m227_78+m228_78+m229_78+m230_78+m231_78+m232_78+m233_78+m234_78+m235_78+m236_78+m237_78+m238_78+m239_78+m240_78+m241_78+m242_78+m243_78+m244_78+m245_78+m246_78+m247_78+m248_78+m249_78+m250_78+m251_78+m252_78+m253_78+m254_78+m255_78+m256_78+m257_78+m258_78+m259_78+m260_78+m261_78+m262_78+m263_78+b78;
   assign out79 = m1_79+m2_79+m3_79+m4_79+m5_79+m6_79+m7_79+m8_79+m9_79+m10_79+m11_79+m12_79+m13_79+m14_79+m15_79+m16_79+m17_79+m18_79+m19_79+m20_79+m21_79+m22_79+m23_79+m24_79+m25_79+m26_79+m27_79+m28_79+m29_79+m30_79+m31_79+m32_79+m33_79+m34_79+m35_79+m36_79+m37_79+m38_79+m39_79+m40_79+m41_79+m42_79+m43_79+m44_79+m45_79+m46_79+m47_79+m48_79+m49_79+m50_79+m51_79+m52_79+m53_79+m54_79+m55_79+m56_79+m57_79+m58_79+m59_79+m60_79+m61_79+m62_79+m63_79+m64_79+m65_79+m66_79+m67_79+m68_79+m69_79+m70_79+m71_79+m72_79+m73_79+m74_79+m75_79+m76_79+m77_79+m78_79+m79_79+m80_79+m81_79+m82_79+m83_79+m84_79+m85_79+m86_79+m87_79+m88_79+m89_79+m90_79+m91_79+m92_79+m93_79+m94_79+m95_79+m96_79+m97_79+m98_79+m99_79+m100_79+m101_79+m102_79+m103_79+m104_79+m105_79+m106_79+m107_79+m108_79+m109_79+m110_79+m111_79+m112_79+m113_79+m114_79+m115_79+m116_79+m117_79+m118_79+m119_79+m120_79+m121_79+m122_79+m123_79+m124_79+m125_79+m126_79+m127_79+m128_79+m129_79+m130_79+m131_79+m132_79+m133_79+m134_79+m135_79+m136_79+m137_79+m138_79+m139_79+m140_79+m141_79+m142_79+m143_79+m144_79+m145_79+m146_79+m147_79+m148_79+m149_79+m150_79+m151_79+m152_79+m153_79+m154_79+m155_79+m156_79+m157_79+m158_79+m159_79+m160_79+m161_79+m162_79+m163_79+m164_79+m165_79+m166_79+m167_79+m168_79+m169_79+m170_79+m171_79+m172_79+m173_79+m174_79+m175_79+m176_79+m177_79+m178_79+m179_79+m180_79+m181_79+m182_79+m183_79+m184_79+m185_79+m186_79+m187_79+m188_79+m189_79+m190_79+m191_79+m192_79+m193_79+m194_79+m195_79+m196_79+m197_79+m198_79+m199_79+m200_79+m201_79+m202_79+m203_79+m204_79+m205_79+m206_79+m207_79+m208_79+m209_79+m210_79+m211_79+m212_79+m213_79+m214_79+m215_79+m216_79+m217_79+m218_79+m219_79+m220_79+m221_79+m222_79+m223_79+m224_79+m225_79+m226_79+m227_79+m228_79+m229_79+m230_79+m231_79+m232_79+m233_79+m234_79+m235_79+m236_79+m237_79+m238_79+m239_79+m240_79+m241_79+m242_79+m243_79+m244_79+m245_79+m246_79+m247_79+m248_79+m249_79+m250_79+m251_79+m252_79+m253_79+m254_79+m255_79+m256_79+m257_79+m258_79+m259_79+m260_79+m261_79+m262_79+m263_79+b79;
   assign out80 = m1_80+m2_80+m3_80+m4_80+m5_80+m6_80+m7_80+m8_80+m9_80+m10_80+m11_80+m12_80+m13_80+m14_80+m15_80+m16_80+m17_80+m18_80+m19_80+m20_80+m21_80+m22_80+m23_80+m24_80+m25_80+m26_80+m27_80+m28_80+m29_80+m30_80+m31_80+m32_80+m33_80+m34_80+m35_80+m36_80+m37_80+m38_80+m39_80+m40_80+m41_80+m42_80+m43_80+m44_80+m45_80+m46_80+m47_80+m48_80+m49_80+m50_80+m51_80+m52_80+m53_80+m54_80+m55_80+m56_80+m57_80+m58_80+m59_80+m60_80+m61_80+m62_80+m63_80+m64_80+m65_80+m66_80+m67_80+m68_80+m69_80+m70_80+m71_80+m72_80+m73_80+m74_80+m75_80+m76_80+m77_80+m78_80+m79_80+m80_80+m81_80+m82_80+m83_80+m84_80+m85_80+m86_80+m87_80+m88_80+m89_80+m90_80+m91_80+m92_80+m93_80+m94_80+m95_80+m96_80+m97_80+m98_80+m99_80+m100_80+m101_80+m102_80+m103_80+m104_80+m105_80+m106_80+m107_80+m108_80+m109_80+m110_80+m111_80+m112_80+m113_80+m114_80+m115_80+m116_80+m117_80+m118_80+m119_80+m120_80+m121_80+m122_80+m123_80+m124_80+m125_80+m126_80+m127_80+m128_80+m129_80+m130_80+m131_80+m132_80+m133_80+m134_80+m135_80+m136_80+m137_80+m138_80+m139_80+m140_80+m141_80+m142_80+m143_80+m144_80+m145_80+m146_80+m147_80+m148_80+m149_80+m150_80+m151_80+m152_80+m153_80+m154_80+m155_80+m156_80+m157_80+m158_80+m159_80+m160_80+m161_80+m162_80+m163_80+m164_80+m165_80+m166_80+m167_80+m168_80+m169_80+m170_80+m171_80+m172_80+m173_80+m174_80+m175_80+m176_80+m177_80+m178_80+m179_80+m180_80+m181_80+m182_80+m183_80+m184_80+m185_80+m186_80+m187_80+m188_80+m189_80+m190_80+m191_80+m192_80+m193_80+m194_80+m195_80+m196_80+m197_80+m198_80+m199_80+m200_80+m201_80+m202_80+m203_80+m204_80+m205_80+m206_80+m207_80+m208_80+m209_80+m210_80+m211_80+m212_80+m213_80+m214_80+m215_80+m216_80+m217_80+m218_80+m219_80+m220_80+m221_80+m222_80+m223_80+m224_80+m225_80+m226_80+m227_80+m228_80+m229_80+m230_80+m231_80+m232_80+m233_80+m234_80+m235_80+m236_80+m237_80+m238_80+m239_80+m240_80+m241_80+m242_80+m243_80+m244_80+m245_80+m246_80+m247_80+m248_80+m249_80+m250_80+m251_80+m252_80+m253_80+m254_80+m255_80+m256_80+m257_80+m258_80+m259_80+m260_80+m261_80+m262_80+m263_80+b80;
   assign out81 = m1_81+m2_81+m3_81+m4_81+m5_81+m6_81+m7_81+m8_81+m9_81+m10_81+m11_81+m12_81+m13_81+m14_81+m15_81+m16_81+m17_81+m18_81+m19_81+m20_81+m21_81+m22_81+m23_81+m24_81+m25_81+m26_81+m27_81+m28_81+m29_81+m30_81+m31_81+m32_81+m33_81+m34_81+m35_81+m36_81+m37_81+m38_81+m39_81+m40_81+m41_81+m42_81+m43_81+m44_81+m45_81+m46_81+m47_81+m48_81+m49_81+m50_81+m51_81+m52_81+m53_81+m54_81+m55_81+m56_81+m57_81+m58_81+m59_81+m60_81+m61_81+m62_81+m63_81+m64_81+m65_81+m66_81+m67_81+m68_81+m69_81+m70_81+m71_81+m72_81+m73_81+m74_81+m75_81+m76_81+m77_81+m78_81+m79_81+m80_81+m81_81+m82_81+m83_81+m84_81+m85_81+m86_81+m87_81+m88_81+m89_81+m90_81+m91_81+m92_81+m93_81+m94_81+m95_81+m96_81+m97_81+m98_81+m99_81+m100_81+m101_81+m102_81+m103_81+m104_81+m105_81+m106_81+m107_81+m108_81+m109_81+m110_81+m111_81+m112_81+m113_81+m114_81+m115_81+m116_81+m117_81+m118_81+m119_81+m120_81+m121_81+m122_81+m123_81+m124_81+m125_81+m126_81+m127_81+m128_81+m129_81+m130_81+m131_81+m132_81+m133_81+m134_81+m135_81+m136_81+m137_81+m138_81+m139_81+m140_81+m141_81+m142_81+m143_81+m144_81+m145_81+m146_81+m147_81+m148_81+m149_81+m150_81+m151_81+m152_81+m153_81+m154_81+m155_81+m156_81+m157_81+m158_81+m159_81+m160_81+m161_81+m162_81+m163_81+m164_81+m165_81+m166_81+m167_81+m168_81+m169_81+m170_81+m171_81+m172_81+m173_81+m174_81+m175_81+m176_81+m177_81+m178_81+m179_81+m180_81+m181_81+m182_81+m183_81+m184_81+m185_81+m186_81+m187_81+m188_81+m189_81+m190_81+m191_81+m192_81+m193_81+m194_81+m195_81+m196_81+m197_81+m198_81+m199_81+m200_81+m201_81+m202_81+m203_81+m204_81+m205_81+m206_81+m207_81+m208_81+m209_81+m210_81+m211_81+m212_81+m213_81+m214_81+m215_81+m216_81+m217_81+m218_81+m219_81+m220_81+m221_81+m222_81+m223_81+m224_81+m225_81+m226_81+m227_81+m228_81+m229_81+m230_81+m231_81+m232_81+m233_81+m234_81+m235_81+m236_81+m237_81+m238_81+m239_81+m240_81+m241_81+m242_81+m243_81+m244_81+m245_81+m246_81+m247_81+m248_81+m249_81+m250_81+m251_81+m252_81+m253_81+m254_81+m255_81+m256_81+m257_81+m258_81+m259_81+m260_81+m261_81+m262_81+m263_81+b81;
   assign out82 = m1_82+m2_82+m3_82+m4_82+m5_82+m6_82+m7_82+m8_82+m9_82+m10_82+m11_82+m12_82+m13_82+m14_82+m15_82+m16_82+m17_82+m18_82+m19_82+m20_82+m21_82+m22_82+m23_82+m24_82+m25_82+m26_82+m27_82+m28_82+m29_82+m30_82+m31_82+m32_82+m33_82+m34_82+m35_82+m36_82+m37_82+m38_82+m39_82+m40_82+m41_82+m42_82+m43_82+m44_82+m45_82+m46_82+m47_82+m48_82+m49_82+m50_82+m51_82+m52_82+m53_82+m54_82+m55_82+m56_82+m57_82+m58_82+m59_82+m60_82+m61_82+m62_82+m63_82+m64_82+m65_82+m66_82+m67_82+m68_82+m69_82+m70_82+m71_82+m72_82+m73_82+m74_82+m75_82+m76_82+m77_82+m78_82+m79_82+m80_82+m81_82+m82_82+m83_82+m84_82+m85_82+m86_82+m87_82+m88_82+m89_82+m90_82+m91_82+m92_82+m93_82+m94_82+m95_82+m96_82+m97_82+m98_82+m99_82+m100_82+m101_82+m102_82+m103_82+m104_82+m105_82+m106_82+m107_82+m108_82+m109_82+m110_82+m111_82+m112_82+m113_82+m114_82+m115_82+m116_82+m117_82+m118_82+m119_82+m120_82+m121_82+m122_82+m123_82+m124_82+m125_82+m126_82+m127_82+m128_82+m129_82+m130_82+m131_82+m132_82+m133_82+m134_82+m135_82+m136_82+m137_82+m138_82+m139_82+m140_82+m141_82+m142_82+m143_82+m144_82+m145_82+m146_82+m147_82+m148_82+m149_82+m150_82+m151_82+m152_82+m153_82+m154_82+m155_82+m156_82+m157_82+m158_82+m159_82+m160_82+m161_82+m162_82+m163_82+m164_82+m165_82+m166_82+m167_82+m168_82+m169_82+m170_82+m171_82+m172_82+m173_82+m174_82+m175_82+m176_82+m177_82+m178_82+m179_82+m180_82+m181_82+m182_82+m183_82+m184_82+m185_82+m186_82+m187_82+m188_82+m189_82+m190_82+m191_82+m192_82+m193_82+m194_82+m195_82+m196_82+m197_82+m198_82+m199_82+m200_82+m201_82+m202_82+m203_82+m204_82+m205_82+m206_82+m207_82+m208_82+m209_82+m210_82+m211_82+m212_82+m213_82+m214_82+m215_82+m216_82+m217_82+m218_82+m219_82+m220_82+m221_82+m222_82+m223_82+m224_82+m225_82+m226_82+m227_82+m228_82+m229_82+m230_82+m231_82+m232_82+m233_82+m234_82+m235_82+m236_82+m237_82+m238_82+m239_82+m240_82+m241_82+m242_82+m243_82+m244_82+m245_82+m246_82+m247_82+m248_82+m249_82+m250_82+m251_82+m252_82+m253_82+m254_82+m255_82+m256_82+m257_82+m258_82+m259_82+m260_82+m261_82+m262_82+m263_82+b82;
   assign out83 = m1_83+m2_83+m3_83+m4_83+m5_83+m6_83+m7_83+m8_83+m9_83+m10_83+m11_83+m12_83+m13_83+m14_83+m15_83+m16_83+m17_83+m18_83+m19_83+m20_83+m21_83+m22_83+m23_83+m24_83+m25_83+m26_83+m27_83+m28_83+m29_83+m30_83+m31_83+m32_83+m33_83+m34_83+m35_83+m36_83+m37_83+m38_83+m39_83+m40_83+m41_83+m42_83+m43_83+m44_83+m45_83+m46_83+m47_83+m48_83+m49_83+m50_83+m51_83+m52_83+m53_83+m54_83+m55_83+m56_83+m57_83+m58_83+m59_83+m60_83+m61_83+m62_83+m63_83+m64_83+m65_83+m66_83+m67_83+m68_83+m69_83+m70_83+m71_83+m72_83+m73_83+m74_83+m75_83+m76_83+m77_83+m78_83+m79_83+m80_83+m81_83+m82_83+m83_83+m84_83+m85_83+m86_83+m87_83+m88_83+m89_83+m90_83+m91_83+m92_83+m93_83+m94_83+m95_83+m96_83+m97_83+m98_83+m99_83+m100_83+m101_83+m102_83+m103_83+m104_83+m105_83+m106_83+m107_83+m108_83+m109_83+m110_83+m111_83+m112_83+m113_83+m114_83+m115_83+m116_83+m117_83+m118_83+m119_83+m120_83+m121_83+m122_83+m123_83+m124_83+m125_83+m126_83+m127_83+m128_83+m129_83+m130_83+m131_83+m132_83+m133_83+m134_83+m135_83+m136_83+m137_83+m138_83+m139_83+m140_83+m141_83+m142_83+m143_83+m144_83+m145_83+m146_83+m147_83+m148_83+m149_83+m150_83+m151_83+m152_83+m153_83+m154_83+m155_83+m156_83+m157_83+m158_83+m159_83+m160_83+m161_83+m162_83+m163_83+m164_83+m165_83+m166_83+m167_83+m168_83+m169_83+m170_83+m171_83+m172_83+m173_83+m174_83+m175_83+m176_83+m177_83+m178_83+m179_83+m180_83+m181_83+m182_83+m183_83+m184_83+m185_83+m186_83+m187_83+m188_83+m189_83+m190_83+m191_83+m192_83+m193_83+m194_83+m195_83+m196_83+m197_83+m198_83+m199_83+m200_83+m201_83+m202_83+m203_83+m204_83+m205_83+m206_83+m207_83+m208_83+m209_83+m210_83+m211_83+m212_83+m213_83+m214_83+m215_83+m216_83+m217_83+m218_83+m219_83+m220_83+m221_83+m222_83+m223_83+m224_83+m225_83+m226_83+m227_83+m228_83+m229_83+m230_83+m231_83+m232_83+m233_83+m234_83+m235_83+m236_83+m237_83+m238_83+m239_83+m240_83+m241_83+m242_83+m243_83+m244_83+m245_83+m246_83+m247_83+m248_83+m249_83+m250_83+m251_83+m252_83+m253_83+m254_83+m255_83+m256_83+m257_83+m258_83+m259_83+m260_83+m261_83+m262_83+m263_83+b83;
   assign out84 = m1_84+m2_84+m3_84+m4_84+m5_84+m6_84+m7_84+m8_84+m9_84+m10_84+m11_84+m12_84+m13_84+m14_84+m15_84+m16_84+m17_84+m18_84+m19_84+m20_84+m21_84+m22_84+m23_84+m24_84+m25_84+m26_84+m27_84+m28_84+m29_84+m30_84+m31_84+m32_84+m33_84+m34_84+m35_84+m36_84+m37_84+m38_84+m39_84+m40_84+m41_84+m42_84+m43_84+m44_84+m45_84+m46_84+m47_84+m48_84+m49_84+m50_84+m51_84+m52_84+m53_84+m54_84+m55_84+m56_84+m57_84+m58_84+m59_84+m60_84+m61_84+m62_84+m63_84+m64_84+m65_84+m66_84+m67_84+m68_84+m69_84+m70_84+m71_84+m72_84+m73_84+m74_84+m75_84+m76_84+m77_84+m78_84+m79_84+m80_84+m81_84+m82_84+m83_84+m84_84+m85_84+m86_84+m87_84+m88_84+m89_84+m90_84+m91_84+m92_84+m93_84+m94_84+m95_84+m96_84+m97_84+m98_84+m99_84+m100_84+m101_84+m102_84+m103_84+m104_84+m105_84+m106_84+m107_84+m108_84+m109_84+m110_84+m111_84+m112_84+m113_84+m114_84+m115_84+m116_84+m117_84+m118_84+m119_84+m120_84+m121_84+m122_84+m123_84+m124_84+m125_84+m126_84+m127_84+m128_84+m129_84+m130_84+m131_84+m132_84+m133_84+m134_84+m135_84+m136_84+m137_84+m138_84+m139_84+m140_84+m141_84+m142_84+m143_84+m144_84+m145_84+m146_84+m147_84+m148_84+m149_84+m150_84+m151_84+m152_84+m153_84+m154_84+m155_84+m156_84+m157_84+m158_84+m159_84+m160_84+m161_84+m162_84+m163_84+m164_84+m165_84+m166_84+m167_84+m168_84+m169_84+m170_84+m171_84+m172_84+m173_84+m174_84+m175_84+m176_84+m177_84+m178_84+m179_84+m180_84+m181_84+m182_84+m183_84+m184_84+m185_84+m186_84+m187_84+m188_84+m189_84+m190_84+m191_84+m192_84+m193_84+m194_84+m195_84+m196_84+m197_84+m198_84+m199_84+m200_84+m201_84+m202_84+m203_84+m204_84+m205_84+m206_84+m207_84+m208_84+m209_84+m210_84+m211_84+m212_84+m213_84+m214_84+m215_84+m216_84+m217_84+m218_84+m219_84+m220_84+m221_84+m222_84+m223_84+m224_84+m225_84+m226_84+m227_84+m228_84+m229_84+m230_84+m231_84+m232_84+m233_84+m234_84+m235_84+m236_84+m237_84+m238_84+m239_84+m240_84+m241_84+m242_84+m243_84+m244_84+m245_84+m246_84+m247_84+m248_84+m249_84+m250_84+m251_84+m252_84+m253_84+m254_84+m255_84+m256_84+m257_84+m258_84+m259_84+m260_84+m261_84+m262_84+m263_84+b84;
   assign out85 = m1_85+m2_85+m3_85+m4_85+m5_85+m6_85+m7_85+m8_85+m9_85+m10_85+m11_85+m12_85+m13_85+m14_85+m15_85+m16_85+m17_85+m18_85+m19_85+m20_85+m21_85+m22_85+m23_85+m24_85+m25_85+m26_85+m27_85+m28_85+m29_85+m30_85+m31_85+m32_85+m33_85+m34_85+m35_85+m36_85+m37_85+m38_85+m39_85+m40_85+m41_85+m42_85+m43_85+m44_85+m45_85+m46_85+m47_85+m48_85+m49_85+m50_85+m51_85+m52_85+m53_85+m54_85+m55_85+m56_85+m57_85+m58_85+m59_85+m60_85+m61_85+m62_85+m63_85+m64_85+m65_85+m66_85+m67_85+m68_85+m69_85+m70_85+m71_85+m72_85+m73_85+m74_85+m75_85+m76_85+m77_85+m78_85+m79_85+m80_85+m81_85+m82_85+m83_85+m84_85+m85_85+m86_85+m87_85+m88_85+m89_85+m90_85+m91_85+m92_85+m93_85+m94_85+m95_85+m96_85+m97_85+m98_85+m99_85+m100_85+m101_85+m102_85+m103_85+m104_85+m105_85+m106_85+m107_85+m108_85+m109_85+m110_85+m111_85+m112_85+m113_85+m114_85+m115_85+m116_85+m117_85+m118_85+m119_85+m120_85+m121_85+m122_85+m123_85+m124_85+m125_85+m126_85+m127_85+m128_85+m129_85+m130_85+m131_85+m132_85+m133_85+m134_85+m135_85+m136_85+m137_85+m138_85+m139_85+m140_85+m141_85+m142_85+m143_85+m144_85+m145_85+m146_85+m147_85+m148_85+m149_85+m150_85+m151_85+m152_85+m153_85+m154_85+m155_85+m156_85+m157_85+m158_85+m159_85+m160_85+m161_85+m162_85+m163_85+m164_85+m165_85+m166_85+m167_85+m168_85+m169_85+m170_85+m171_85+m172_85+m173_85+m174_85+m175_85+m176_85+m177_85+m178_85+m179_85+m180_85+m181_85+m182_85+m183_85+m184_85+m185_85+m186_85+m187_85+m188_85+m189_85+m190_85+m191_85+m192_85+m193_85+m194_85+m195_85+m196_85+m197_85+m198_85+m199_85+m200_85+m201_85+m202_85+m203_85+m204_85+m205_85+m206_85+m207_85+m208_85+m209_85+m210_85+m211_85+m212_85+m213_85+m214_85+m215_85+m216_85+m217_85+m218_85+m219_85+m220_85+m221_85+m222_85+m223_85+m224_85+m225_85+m226_85+m227_85+m228_85+m229_85+m230_85+m231_85+m232_85+m233_85+m234_85+m235_85+m236_85+m237_85+m238_85+m239_85+m240_85+m241_85+m242_85+m243_85+m244_85+m245_85+m246_85+m247_85+m248_85+m249_85+m250_85+m251_85+m252_85+m253_85+m254_85+m255_85+m256_85+m257_85+m258_85+m259_85+m260_85+m261_85+m262_85+m263_85+b85;
   assign out86 = m1_86+m2_86+m3_86+m4_86+m5_86+m6_86+m7_86+m8_86+m9_86+m10_86+m11_86+m12_86+m13_86+m14_86+m15_86+m16_86+m17_86+m18_86+m19_86+m20_86+m21_86+m22_86+m23_86+m24_86+m25_86+m26_86+m27_86+m28_86+m29_86+m30_86+m31_86+m32_86+m33_86+m34_86+m35_86+m36_86+m37_86+m38_86+m39_86+m40_86+m41_86+m42_86+m43_86+m44_86+m45_86+m46_86+m47_86+m48_86+m49_86+m50_86+m51_86+m52_86+m53_86+m54_86+m55_86+m56_86+m57_86+m58_86+m59_86+m60_86+m61_86+m62_86+m63_86+m64_86+m65_86+m66_86+m67_86+m68_86+m69_86+m70_86+m71_86+m72_86+m73_86+m74_86+m75_86+m76_86+m77_86+m78_86+m79_86+m80_86+m81_86+m82_86+m83_86+m84_86+m85_86+m86_86+m87_86+m88_86+m89_86+m90_86+m91_86+m92_86+m93_86+m94_86+m95_86+m96_86+m97_86+m98_86+m99_86+m100_86+m101_86+m102_86+m103_86+m104_86+m105_86+m106_86+m107_86+m108_86+m109_86+m110_86+m111_86+m112_86+m113_86+m114_86+m115_86+m116_86+m117_86+m118_86+m119_86+m120_86+m121_86+m122_86+m123_86+m124_86+m125_86+m126_86+m127_86+m128_86+m129_86+m130_86+m131_86+m132_86+m133_86+m134_86+m135_86+m136_86+m137_86+m138_86+m139_86+m140_86+m141_86+m142_86+m143_86+m144_86+m145_86+m146_86+m147_86+m148_86+m149_86+m150_86+m151_86+m152_86+m153_86+m154_86+m155_86+m156_86+m157_86+m158_86+m159_86+m160_86+m161_86+m162_86+m163_86+m164_86+m165_86+m166_86+m167_86+m168_86+m169_86+m170_86+m171_86+m172_86+m173_86+m174_86+m175_86+m176_86+m177_86+m178_86+m179_86+m180_86+m181_86+m182_86+m183_86+m184_86+m185_86+m186_86+m187_86+m188_86+m189_86+m190_86+m191_86+m192_86+m193_86+m194_86+m195_86+m196_86+m197_86+m198_86+m199_86+m200_86+m201_86+m202_86+m203_86+m204_86+m205_86+m206_86+m207_86+m208_86+m209_86+m210_86+m211_86+m212_86+m213_86+m214_86+m215_86+m216_86+m217_86+m218_86+m219_86+m220_86+m221_86+m222_86+m223_86+m224_86+m225_86+m226_86+m227_86+m228_86+m229_86+m230_86+m231_86+m232_86+m233_86+m234_86+m235_86+m236_86+m237_86+m238_86+m239_86+m240_86+m241_86+m242_86+m243_86+m244_86+m245_86+m246_86+m247_86+m248_86+m249_86+m250_86+m251_86+m252_86+m253_86+m254_86+m255_86+m256_86+m257_86+m258_86+m259_86+m260_86+m261_86+m262_86+m263_86+b86;
   assign out87 = m1_87+m2_87+m3_87+m4_87+m5_87+m6_87+m7_87+m8_87+m9_87+m10_87+m11_87+m12_87+m13_87+m14_87+m15_87+m16_87+m17_87+m18_87+m19_87+m20_87+m21_87+m22_87+m23_87+m24_87+m25_87+m26_87+m27_87+m28_87+m29_87+m30_87+m31_87+m32_87+m33_87+m34_87+m35_87+m36_87+m37_87+m38_87+m39_87+m40_87+m41_87+m42_87+m43_87+m44_87+m45_87+m46_87+m47_87+m48_87+m49_87+m50_87+m51_87+m52_87+m53_87+m54_87+m55_87+m56_87+m57_87+m58_87+m59_87+m60_87+m61_87+m62_87+m63_87+m64_87+m65_87+m66_87+m67_87+m68_87+m69_87+m70_87+m71_87+m72_87+m73_87+m74_87+m75_87+m76_87+m77_87+m78_87+m79_87+m80_87+m81_87+m82_87+m83_87+m84_87+m85_87+m86_87+m87_87+m88_87+m89_87+m90_87+m91_87+m92_87+m93_87+m94_87+m95_87+m96_87+m97_87+m98_87+m99_87+m100_87+m101_87+m102_87+m103_87+m104_87+m105_87+m106_87+m107_87+m108_87+m109_87+m110_87+m111_87+m112_87+m113_87+m114_87+m115_87+m116_87+m117_87+m118_87+m119_87+m120_87+m121_87+m122_87+m123_87+m124_87+m125_87+m126_87+m127_87+m128_87+m129_87+m130_87+m131_87+m132_87+m133_87+m134_87+m135_87+m136_87+m137_87+m138_87+m139_87+m140_87+m141_87+m142_87+m143_87+m144_87+m145_87+m146_87+m147_87+m148_87+m149_87+m150_87+m151_87+m152_87+m153_87+m154_87+m155_87+m156_87+m157_87+m158_87+m159_87+m160_87+m161_87+m162_87+m163_87+m164_87+m165_87+m166_87+m167_87+m168_87+m169_87+m170_87+m171_87+m172_87+m173_87+m174_87+m175_87+m176_87+m177_87+m178_87+m179_87+m180_87+m181_87+m182_87+m183_87+m184_87+m185_87+m186_87+m187_87+m188_87+m189_87+m190_87+m191_87+m192_87+m193_87+m194_87+m195_87+m196_87+m197_87+m198_87+m199_87+m200_87+m201_87+m202_87+m203_87+m204_87+m205_87+m206_87+m207_87+m208_87+m209_87+m210_87+m211_87+m212_87+m213_87+m214_87+m215_87+m216_87+m217_87+m218_87+m219_87+m220_87+m221_87+m222_87+m223_87+m224_87+m225_87+m226_87+m227_87+m228_87+m229_87+m230_87+m231_87+m232_87+m233_87+m234_87+m235_87+m236_87+m237_87+m238_87+m239_87+m240_87+m241_87+m242_87+m243_87+m244_87+m245_87+m246_87+m247_87+m248_87+m249_87+m250_87+m251_87+m252_87+m253_87+m254_87+m255_87+m256_87+m257_87+m258_87+m259_87+m260_87+m261_87+m262_87+m263_87+b87;
   assign out88 = m1_88+m2_88+m3_88+m4_88+m5_88+m6_88+m7_88+m8_88+m9_88+m10_88+m11_88+m12_88+m13_88+m14_88+m15_88+m16_88+m17_88+m18_88+m19_88+m20_88+m21_88+m22_88+m23_88+m24_88+m25_88+m26_88+m27_88+m28_88+m29_88+m30_88+m31_88+m32_88+m33_88+m34_88+m35_88+m36_88+m37_88+m38_88+m39_88+m40_88+m41_88+m42_88+m43_88+m44_88+m45_88+m46_88+m47_88+m48_88+m49_88+m50_88+m51_88+m52_88+m53_88+m54_88+m55_88+m56_88+m57_88+m58_88+m59_88+m60_88+m61_88+m62_88+m63_88+m64_88+m65_88+m66_88+m67_88+m68_88+m69_88+m70_88+m71_88+m72_88+m73_88+m74_88+m75_88+m76_88+m77_88+m78_88+m79_88+m80_88+m81_88+m82_88+m83_88+m84_88+m85_88+m86_88+m87_88+m88_88+m89_88+m90_88+m91_88+m92_88+m93_88+m94_88+m95_88+m96_88+m97_88+m98_88+m99_88+m100_88+m101_88+m102_88+m103_88+m104_88+m105_88+m106_88+m107_88+m108_88+m109_88+m110_88+m111_88+m112_88+m113_88+m114_88+m115_88+m116_88+m117_88+m118_88+m119_88+m120_88+m121_88+m122_88+m123_88+m124_88+m125_88+m126_88+m127_88+m128_88+m129_88+m130_88+m131_88+m132_88+m133_88+m134_88+m135_88+m136_88+m137_88+m138_88+m139_88+m140_88+m141_88+m142_88+m143_88+m144_88+m145_88+m146_88+m147_88+m148_88+m149_88+m150_88+m151_88+m152_88+m153_88+m154_88+m155_88+m156_88+m157_88+m158_88+m159_88+m160_88+m161_88+m162_88+m163_88+m164_88+m165_88+m166_88+m167_88+m168_88+m169_88+m170_88+m171_88+m172_88+m173_88+m174_88+m175_88+m176_88+m177_88+m178_88+m179_88+m180_88+m181_88+m182_88+m183_88+m184_88+m185_88+m186_88+m187_88+m188_88+m189_88+m190_88+m191_88+m192_88+m193_88+m194_88+m195_88+m196_88+m197_88+m198_88+m199_88+m200_88+m201_88+m202_88+m203_88+m204_88+m205_88+m206_88+m207_88+m208_88+m209_88+m210_88+m211_88+m212_88+m213_88+m214_88+m215_88+m216_88+m217_88+m218_88+m219_88+m220_88+m221_88+m222_88+m223_88+m224_88+m225_88+m226_88+m227_88+m228_88+m229_88+m230_88+m231_88+m232_88+m233_88+m234_88+m235_88+m236_88+m237_88+m238_88+m239_88+m240_88+m241_88+m242_88+m243_88+m244_88+m245_88+m246_88+m247_88+m248_88+m249_88+m250_88+m251_88+m252_88+m253_88+m254_88+m255_88+m256_88+m257_88+m258_88+m259_88+m260_88+m261_88+m262_88+m263_88+b88;
   assign out89 = m1_89+m2_89+m3_89+m4_89+m5_89+m6_89+m7_89+m8_89+m9_89+m10_89+m11_89+m12_89+m13_89+m14_89+m15_89+m16_89+m17_89+m18_89+m19_89+m20_89+m21_89+m22_89+m23_89+m24_89+m25_89+m26_89+m27_89+m28_89+m29_89+m30_89+m31_89+m32_89+m33_89+m34_89+m35_89+m36_89+m37_89+m38_89+m39_89+m40_89+m41_89+m42_89+m43_89+m44_89+m45_89+m46_89+m47_89+m48_89+m49_89+m50_89+m51_89+m52_89+m53_89+m54_89+m55_89+m56_89+m57_89+m58_89+m59_89+m60_89+m61_89+m62_89+m63_89+m64_89+m65_89+m66_89+m67_89+m68_89+m69_89+m70_89+m71_89+m72_89+m73_89+m74_89+m75_89+m76_89+m77_89+m78_89+m79_89+m80_89+m81_89+m82_89+m83_89+m84_89+m85_89+m86_89+m87_89+m88_89+m89_89+m90_89+m91_89+m92_89+m93_89+m94_89+m95_89+m96_89+m97_89+m98_89+m99_89+m100_89+m101_89+m102_89+m103_89+m104_89+m105_89+m106_89+m107_89+m108_89+m109_89+m110_89+m111_89+m112_89+m113_89+m114_89+m115_89+m116_89+m117_89+m118_89+m119_89+m120_89+m121_89+m122_89+m123_89+m124_89+m125_89+m126_89+m127_89+m128_89+m129_89+m130_89+m131_89+m132_89+m133_89+m134_89+m135_89+m136_89+m137_89+m138_89+m139_89+m140_89+m141_89+m142_89+m143_89+m144_89+m145_89+m146_89+m147_89+m148_89+m149_89+m150_89+m151_89+m152_89+m153_89+m154_89+m155_89+m156_89+m157_89+m158_89+m159_89+m160_89+m161_89+m162_89+m163_89+m164_89+m165_89+m166_89+m167_89+m168_89+m169_89+m170_89+m171_89+m172_89+m173_89+m174_89+m175_89+m176_89+m177_89+m178_89+m179_89+m180_89+m181_89+m182_89+m183_89+m184_89+m185_89+m186_89+m187_89+m188_89+m189_89+m190_89+m191_89+m192_89+m193_89+m194_89+m195_89+m196_89+m197_89+m198_89+m199_89+m200_89+m201_89+m202_89+m203_89+m204_89+m205_89+m206_89+m207_89+m208_89+m209_89+m210_89+m211_89+m212_89+m213_89+m214_89+m215_89+m216_89+m217_89+m218_89+m219_89+m220_89+m221_89+m222_89+m223_89+m224_89+m225_89+m226_89+m227_89+m228_89+m229_89+m230_89+m231_89+m232_89+m233_89+m234_89+m235_89+m236_89+m237_89+m238_89+m239_89+m240_89+m241_89+m242_89+m243_89+m244_89+m245_89+m246_89+m247_89+m248_89+m249_89+m250_89+m251_89+m252_89+m253_89+m254_89+m255_89+m256_89+m257_89+m258_89+m259_89+m260_89+m261_89+m262_89+m263_89+b89;
   assign out90 = m1_90+m2_90+m3_90+m4_90+m5_90+m6_90+m7_90+m8_90+m9_90+m10_90+m11_90+m12_90+m13_90+m14_90+m15_90+m16_90+m17_90+m18_90+m19_90+m20_90+m21_90+m22_90+m23_90+m24_90+m25_90+m26_90+m27_90+m28_90+m29_90+m30_90+m31_90+m32_90+m33_90+m34_90+m35_90+m36_90+m37_90+m38_90+m39_90+m40_90+m41_90+m42_90+m43_90+m44_90+m45_90+m46_90+m47_90+m48_90+m49_90+m50_90+m51_90+m52_90+m53_90+m54_90+m55_90+m56_90+m57_90+m58_90+m59_90+m60_90+m61_90+m62_90+m63_90+m64_90+m65_90+m66_90+m67_90+m68_90+m69_90+m70_90+m71_90+m72_90+m73_90+m74_90+m75_90+m76_90+m77_90+m78_90+m79_90+m80_90+m81_90+m82_90+m83_90+m84_90+m85_90+m86_90+m87_90+m88_90+m89_90+m90_90+m91_90+m92_90+m93_90+m94_90+m95_90+m96_90+m97_90+m98_90+m99_90+m100_90+m101_90+m102_90+m103_90+m104_90+m105_90+m106_90+m107_90+m108_90+m109_90+m110_90+m111_90+m112_90+m113_90+m114_90+m115_90+m116_90+m117_90+m118_90+m119_90+m120_90+m121_90+m122_90+m123_90+m124_90+m125_90+m126_90+m127_90+m128_90+m129_90+m130_90+m131_90+m132_90+m133_90+m134_90+m135_90+m136_90+m137_90+m138_90+m139_90+m140_90+m141_90+m142_90+m143_90+m144_90+m145_90+m146_90+m147_90+m148_90+m149_90+m150_90+m151_90+m152_90+m153_90+m154_90+m155_90+m156_90+m157_90+m158_90+m159_90+m160_90+m161_90+m162_90+m163_90+m164_90+m165_90+m166_90+m167_90+m168_90+m169_90+m170_90+m171_90+m172_90+m173_90+m174_90+m175_90+m176_90+m177_90+m178_90+m179_90+m180_90+m181_90+m182_90+m183_90+m184_90+m185_90+m186_90+m187_90+m188_90+m189_90+m190_90+m191_90+m192_90+m193_90+m194_90+m195_90+m196_90+m197_90+m198_90+m199_90+m200_90+m201_90+m202_90+m203_90+m204_90+m205_90+m206_90+m207_90+m208_90+m209_90+m210_90+m211_90+m212_90+m213_90+m214_90+m215_90+m216_90+m217_90+m218_90+m219_90+m220_90+m221_90+m222_90+m223_90+m224_90+m225_90+m226_90+m227_90+m228_90+m229_90+m230_90+m231_90+m232_90+m233_90+m234_90+m235_90+m236_90+m237_90+m238_90+m239_90+m240_90+m241_90+m242_90+m243_90+m244_90+m245_90+m246_90+m247_90+m248_90+m249_90+m250_90+m251_90+m252_90+m253_90+m254_90+m255_90+m256_90+m257_90+m258_90+m259_90+m260_90+m261_90+m262_90+m263_90+b90;
   assign out91 = m1_91+m2_91+m3_91+m4_91+m5_91+m6_91+m7_91+m8_91+m9_91+m10_91+m11_91+m12_91+m13_91+m14_91+m15_91+m16_91+m17_91+m18_91+m19_91+m20_91+m21_91+m22_91+m23_91+m24_91+m25_91+m26_91+m27_91+m28_91+m29_91+m30_91+m31_91+m32_91+m33_91+m34_91+m35_91+m36_91+m37_91+m38_91+m39_91+m40_91+m41_91+m42_91+m43_91+m44_91+m45_91+m46_91+m47_91+m48_91+m49_91+m50_91+m51_91+m52_91+m53_91+m54_91+m55_91+m56_91+m57_91+m58_91+m59_91+m60_91+m61_91+m62_91+m63_91+m64_91+m65_91+m66_91+m67_91+m68_91+m69_91+m70_91+m71_91+m72_91+m73_91+m74_91+m75_91+m76_91+m77_91+m78_91+m79_91+m80_91+m81_91+m82_91+m83_91+m84_91+m85_91+m86_91+m87_91+m88_91+m89_91+m90_91+m91_91+m92_91+m93_91+m94_91+m95_91+m96_91+m97_91+m98_91+m99_91+m100_91+m101_91+m102_91+m103_91+m104_91+m105_91+m106_91+m107_91+m108_91+m109_91+m110_91+m111_91+m112_91+m113_91+m114_91+m115_91+m116_91+m117_91+m118_91+m119_91+m120_91+m121_91+m122_91+m123_91+m124_91+m125_91+m126_91+m127_91+m128_91+m129_91+m130_91+m131_91+m132_91+m133_91+m134_91+m135_91+m136_91+m137_91+m138_91+m139_91+m140_91+m141_91+m142_91+m143_91+m144_91+m145_91+m146_91+m147_91+m148_91+m149_91+m150_91+m151_91+m152_91+m153_91+m154_91+m155_91+m156_91+m157_91+m158_91+m159_91+m160_91+m161_91+m162_91+m163_91+m164_91+m165_91+m166_91+m167_91+m168_91+m169_91+m170_91+m171_91+m172_91+m173_91+m174_91+m175_91+m176_91+m177_91+m178_91+m179_91+m180_91+m181_91+m182_91+m183_91+m184_91+m185_91+m186_91+m187_91+m188_91+m189_91+m190_91+m191_91+m192_91+m193_91+m194_91+m195_91+m196_91+m197_91+m198_91+m199_91+m200_91+m201_91+m202_91+m203_91+m204_91+m205_91+m206_91+m207_91+m208_91+m209_91+m210_91+m211_91+m212_91+m213_91+m214_91+m215_91+m216_91+m217_91+m218_91+m219_91+m220_91+m221_91+m222_91+m223_91+m224_91+m225_91+m226_91+m227_91+m228_91+m229_91+m230_91+m231_91+m232_91+m233_91+m234_91+m235_91+m236_91+m237_91+m238_91+m239_91+m240_91+m241_91+m242_91+m243_91+m244_91+m245_91+m246_91+m247_91+m248_91+m249_91+m250_91+m251_91+m252_91+m253_91+m254_91+m255_91+m256_91+m257_91+m258_91+m259_91+m260_91+m261_91+m262_91+m263_91+b91;
   assign out92 = m1_92+m2_92+m3_92+m4_92+m5_92+m6_92+m7_92+m8_92+m9_92+m10_92+m11_92+m12_92+m13_92+m14_92+m15_92+m16_92+m17_92+m18_92+m19_92+m20_92+m21_92+m22_92+m23_92+m24_92+m25_92+m26_92+m27_92+m28_92+m29_92+m30_92+m31_92+m32_92+m33_92+m34_92+m35_92+m36_92+m37_92+m38_92+m39_92+m40_92+m41_92+m42_92+m43_92+m44_92+m45_92+m46_92+m47_92+m48_92+m49_92+m50_92+m51_92+m52_92+m53_92+m54_92+m55_92+m56_92+m57_92+m58_92+m59_92+m60_92+m61_92+m62_92+m63_92+m64_92+m65_92+m66_92+m67_92+m68_92+m69_92+m70_92+m71_92+m72_92+m73_92+m74_92+m75_92+m76_92+m77_92+m78_92+m79_92+m80_92+m81_92+m82_92+m83_92+m84_92+m85_92+m86_92+m87_92+m88_92+m89_92+m90_92+m91_92+m92_92+m93_92+m94_92+m95_92+m96_92+m97_92+m98_92+m99_92+m100_92+m101_92+m102_92+m103_92+m104_92+m105_92+m106_92+m107_92+m108_92+m109_92+m110_92+m111_92+m112_92+m113_92+m114_92+m115_92+m116_92+m117_92+m118_92+m119_92+m120_92+m121_92+m122_92+m123_92+m124_92+m125_92+m126_92+m127_92+m128_92+m129_92+m130_92+m131_92+m132_92+m133_92+m134_92+m135_92+m136_92+m137_92+m138_92+m139_92+m140_92+m141_92+m142_92+m143_92+m144_92+m145_92+m146_92+m147_92+m148_92+m149_92+m150_92+m151_92+m152_92+m153_92+m154_92+m155_92+m156_92+m157_92+m158_92+m159_92+m160_92+m161_92+m162_92+m163_92+m164_92+m165_92+m166_92+m167_92+m168_92+m169_92+m170_92+m171_92+m172_92+m173_92+m174_92+m175_92+m176_92+m177_92+m178_92+m179_92+m180_92+m181_92+m182_92+m183_92+m184_92+m185_92+m186_92+m187_92+m188_92+m189_92+m190_92+m191_92+m192_92+m193_92+m194_92+m195_92+m196_92+m197_92+m198_92+m199_92+m200_92+m201_92+m202_92+m203_92+m204_92+m205_92+m206_92+m207_92+m208_92+m209_92+m210_92+m211_92+m212_92+m213_92+m214_92+m215_92+m216_92+m217_92+m218_92+m219_92+m220_92+m221_92+m222_92+m223_92+m224_92+m225_92+m226_92+m227_92+m228_92+m229_92+m230_92+m231_92+m232_92+m233_92+m234_92+m235_92+m236_92+m237_92+m238_92+m239_92+m240_92+m241_92+m242_92+m243_92+m244_92+m245_92+m246_92+m247_92+m248_92+m249_92+m250_92+m251_92+m252_92+m253_92+m254_92+m255_92+m256_92+m257_92+m258_92+m259_92+m260_92+m261_92+m262_92+m263_92+b92;
   assign out93 = m1_93+m2_93+m3_93+m4_93+m5_93+m6_93+m7_93+m8_93+m9_93+m10_93+m11_93+m12_93+m13_93+m14_93+m15_93+m16_93+m17_93+m18_93+m19_93+m20_93+m21_93+m22_93+m23_93+m24_93+m25_93+m26_93+m27_93+m28_93+m29_93+m30_93+m31_93+m32_93+m33_93+m34_93+m35_93+m36_93+m37_93+m38_93+m39_93+m40_93+m41_93+m42_93+m43_93+m44_93+m45_93+m46_93+m47_93+m48_93+m49_93+m50_93+m51_93+m52_93+m53_93+m54_93+m55_93+m56_93+m57_93+m58_93+m59_93+m60_93+m61_93+m62_93+m63_93+m64_93+m65_93+m66_93+m67_93+m68_93+m69_93+m70_93+m71_93+m72_93+m73_93+m74_93+m75_93+m76_93+m77_93+m78_93+m79_93+m80_93+m81_93+m82_93+m83_93+m84_93+m85_93+m86_93+m87_93+m88_93+m89_93+m90_93+m91_93+m92_93+m93_93+m94_93+m95_93+m96_93+m97_93+m98_93+m99_93+m100_93+m101_93+m102_93+m103_93+m104_93+m105_93+m106_93+m107_93+m108_93+m109_93+m110_93+m111_93+m112_93+m113_93+m114_93+m115_93+m116_93+m117_93+m118_93+m119_93+m120_93+m121_93+m122_93+m123_93+m124_93+m125_93+m126_93+m127_93+m128_93+m129_93+m130_93+m131_93+m132_93+m133_93+m134_93+m135_93+m136_93+m137_93+m138_93+m139_93+m140_93+m141_93+m142_93+m143_93+m144_93+m145_93+m146_93+m147_93+m148_93+m149_93+m150_93+m151_93+m152_93+m153_93+m154_93+m155_93+m156_93+m157_93+m158_93+m159_93+m160_93+m161_93+m162_93+m163_93+m164_93+m165_93+m166_93+m167_93+m168_93+m169_93+m170_93+m171_93+m172_93+m173_93+m174_93+m175_93+m176_93+m177_93+m178_93+m179_93+m180_93+m181_93+m182_93+m183_93+m184_93+m185_93+m186_93+m187_93+m188_93+m189_93+m190_93+m191_93+m192_93+m193_93+m194_93+m195_93+m196_93+m197_93+m198_93+m199_93+m200_93+m201_93+m202_93+m203_93+m204_93+m205_93+m206_93+m207_93+m208_93+m209_93+m210_93+m211_93+m212_93+m213_93+m214_93+m215_93+m216_93+m217_93+m218_93+m219_93+m220_93+m221_93+m222_93+m223_93+m224_93+m225_93+m226_93+m227_93+m228_93+m229_93+m230_93+m231_93+m232_93+m233_93+m234_93+m235_93+m236_93+m237_93+m238_93+m239_93+m240_93+m241_93+m242_93+m243_93+m244_93+m245_93+m246_93+m247_93+m248_93+m249_93+m250_93+m251_93+m252_93+m253_93+m254_93+m255_93+m256_93+m257_93+m258_93+m259_93+m260_93+m261_93+m262_93+m263_93+b93;
   assign out94 = m1_94+m2_94+m3_94+m4_94+m5_94+m6_94+m7_94+m8_94+m9_94+m10_94+m11_94+m12_94+m13_94+m14_94+m15_94+m16_94+m17_94+m18_94+m19_94+m20_94+m21_94+m22_94+m23_94+m24_94+m25_94+m26_94+m27_94+m28_94+m29_94+m30_94+m31_94+m32_94+m33_94+m34_94+m35_94+m36_94+m37_94+m38_94+m39_94+m40_94+m41_94+m42_94+m43_94+m44_94+m45_94+m46_94+m47_94+m48_94+m49_94+m50_94+m51_94+m52_94+m53_94+m54_94+m55_94+m56_94+m57_94+m58_94+m59_94+m60_94+m61_94+m62_94+m63_94+m64_94+m65_94+m66_94+m67_94+m68_94+m69_94+m70_94+m71_94+m72_94+m73_94+m74_94+m75_94+m76_94+m77_94+m78_94+m79_94+m80_94+m81_94+m82_94+m83_94+m84_94+m85_94+m86_94+m87_94+m88_94+m89_94+m90_94+m91_94+m92_94+m93_94+m94_94+m95_94+m96_94+m97_94+m98_94+m99_94+m100_94+m101_94+m102_94+m103_94+m104_94+m105_94+m106_94+m107_94+m108_94+m109_94+m110_94+m111_94+m112_94+m113_94+m114_94+m115_94+m116_94+m117_94+m118_94+m119_94+m120_94+m121_94+m122_94+m123_94+m124_94+m125_94+m126_94+m127_94+m128_94+m129_94+m130_94+m131_94+m132_94+m133_94+m134_94+m135_94+m136_94+m137_94+m138_94+m139_94+m140_94+m141_94+m142_94+m143_94+m144_94+m145_94+m146_94+m147_94+m148_94+m149_94+m150_94+m151_94+m152_94+m153_94+m154_94+m155_94+m156_94+m157_94+m158_94+m159_94+m160_94+m161_94+m162_94+m163_94+m164_94+m165_94+m166_94+m167_94+m168_94+m169_94+m170_94+m171_94+m172_94+m173_94+m174_94+m175_94+m176_94+m177_94+m178_94+m179_94+m180_94+m181_94+m182_94+m183_94+m184_94+m185_94+m186_94+m187_94+m188_94+m189_94+m190_94+m191_94+m192_94+m193_94+m194_94+m195_94+m196_94+m197_94+m198_94+m199_94+m200_94+m201_94+m202_94+m203_94+m204_94+m205_94+m206_94+m207_94+m208_94+m209_94+m210_94+m211_94+m212_94+m213_94+m214_94+m215_94+m216_94+m217_94+m218_94+m219_94+m220_94+m221_94+m222_94+m223_94+m224_94+m225_94+m226_94+m227_94+m228_94+m229_94+m230_94+m231_94+m232_94+m233_94+m234_94+m235_94+m236_94+m237_94+m238_94+m239_94+m240_94+m241_94+m242_94+m243_94+m244_94+m245_94+m246_94+m247_94+m248_94+m249_94+m250_94+m251_94+m252_94+m253_94+m254_94+m255_94+m256_94+m257_94+m258_94+m259_94+m260_94+m261_94+m262_94+m263_94+b94;
   assign out95 = m1_95+m2_95+m3_95+m4_95+m5_95+m6_95+m7_95+m8_95+m9_95+m10_95+m11_95+m12_95+m13_95+m14_95+m15_95+m16_95+m17_95+m18_95+m19_95+m20_95+m21_95+m22_95+m23_95+m24_95+m25_95+m26_95+m27_95+m28_95+m29_95+m30_95+m31_95+m32_95+m33_95+m34_95+m35_95+m36_95+m37_95+m38_95+m39_95+m40_95+m41_95+m42_95+m43_95+m44_95+m45_95+m46_95+m47_95+m48_95+m49_95+m50_95+m51_95+m52_95+m53_95+m54_95+m55_95+m56_95+m57_95+m58_95+m59_95+m60_95+m61_95+m62_95+m63_95+m64_95+m65_95+m66_95+m67_95+m68_95+m69_95+m70_95+m71_95+m72_95+m73_95+m74_95+m75_95+m76_95+m77_95+m78_95+m79_95+m80_95+m81_95+m82_95+m83_95+m84_95+m85_95+m86_95+m87_95+m88_95+m89_95+m90_95+m91_95+m92_95+m93_95+m94_95+m95_95+m96_95+m97_95+m98_95+m99_95+m100_95+m101_95+m102_95+m103_95+m104_95+m105_95+m106_95+m107_95+m108_95+m109_95+m110_95+m111_95+m112_95+m113_95+m114_95+m115_95+m116_95+m117_95+m118_95+m119_95+m120_95+m121_95+m122_95+m123_95+m124_95+m125_95+m126_95+m127_95+m128_95+m129_95+m130_95+m131_95+m132_95+m133_95+m134_95+m135_95+m136_95+m137_95+m138_95+m139_95+m140_95+m141_95+m142_95+m143_95+m144_95+m145_95+m146_95+m147_95+m148_95+m149_95+m150_95+m151_95+m152_95+m153_95+m154_95+m155_95+m156_95+m157_95+m158_95+m159_95+m160_95+m161_95+m162_95+m163_95+m164_95+m165_95+m166_95+m167_95+m168_95+m169_95+m170_95+m171_95+m172_95+m173_95+m174_95+m175_95+m176_95+m177_95+m178_95+m179_95+m180_95+m181_95+m182_95+m183_95+m184_95+m185_95+m186_95+m187_95+m188_95+m189_95+m190_95+m191_95+m192_95+m193_95+m194_95+m195_95+m196_95+m197_95+m198_95+m199_95+m200_95+m201_95+m202_95+m203_95+m204_95+m205_95+m206_95+m207_95+m208_95+m209_95+m210_95+m211_95+m212_95+m213_95+m214_95+m215_95+m216_95+m217_95+m218_95+m219_95+m220_95+m221_95+m222_95+m223_95+m224_95+m225_95+m226_95+m227_95+m228_95+m229_95+m230_95+m231_95+m232_95+m233_95+m234_95+m235_95+m236_95+m237_95+m238_95+m239_95+m240_95+m241_95+m242_95+m243_95+m244_95+m245_95+m246_95+m247_95+m248_95+m249_95+m250_95+m251_95+m252_95+m253_95+m254_95+m255_95+m256_95+m257_95+m258_95+m259_95+m260_95+m261_95+m262_95+m263_95+b95;
   assign out96 = m1_96+m2_96+m3_96+m4_96+m5_96+m6_96+m7_96+m8_96+m9_96+m10_96+m11_96+m12_96+m13_96+m14_96+m15_96+m16_96+m17_96+m18_96+m19_96+m20_96+m21_96+m22_96+m23_96+m24_96+m25_96+m26_96+m27_96+m28_96+m29_96+m30_96+m31_96+m32_96+m33_96+m34_96+m35_96+m36_96+m37_96+m38_96+m39_96+m40_96+m41_96+m42_96+m43_96+m44_96+m45_96+m46_96+m47_96+m48_96+m49_96+m50_96+m51_96+m52_96+m53_96+m54_96+m55_96+m56_96+m57_96+m58_96+m59_96+m60_96+m61_96+m62_96+m63_96+m64_96+m65_96+m66_96+m67_96+m68_96+m69_96+m70_96+m71_96+m72_96+m73_96+m74_96+m75_96+m76_96+m77_96+m78_96+m79_96+m80_96+m81_96+m82_96+m83_96+m84_96+m85_96+m86_96+m87_96+m88_96+m89_96+m90_96+m91_96+m92_96+m93_96+m94_96+m95_96+m96_96+m97_96+m98_96+m99_96+m100_96+m101_96+m102_96+m103_96+m104_96+m105_96+m106_96+m107_96+m108_96+m109_96+m110_96+m111_96+m112_96+m113_96+m114_96+m115_96+m116_96+m117_96+m118_96+m119_96+m120_96+m121_96+m122_96+m123_96+m124_96+m125_96+m126_96+m127_96+m128_96+m129_96+m130_96+m131_96+m132_96+m133_96+m134_96+m135_96+m136_96+m137_96+m138_96+m139_96+m140_96+m141_96+m142_96+m143_96+m144_96+m145_96+m146_96+m147_96+m148_96+m149_96+m150_96+m151_96+m152_96+m153_96+m154_96+m155_96+m156_96+m157_96+m158_96+m159_96+m160_96+m161_96+m162_96+m163_96+m164_96+m165_96+m166_96+m167_96+m168_96+m169_96+m170_96+m171_96+m172_96+m173_96+m174_96+m175_96+m176_96+m177_96+m178_96+m179_96+m180_96+m181_96+m182_96+m183_96+m184_96+m185_96+m186_96+m187_96+m188_96+m189_96+m190_96+m191_96+m192_96+m193_96+m194_96+m195_96+m196_96+m197_96+m198_96+m199_96+m200_96+m201_96+m202_96+m203_96+m204_96+m205_96+m206_96+m207_96+m208_96+m209_96+m210_96+m211_96+m212_96+m213_96+m214_96+m215_96+m216_96+m217_96+m218_96+m219_96+m220_96+m221_96+m222_96+m223_96+m224_96+m225_96+m226_96+m227_96+m228_96+m229_96+m230_96+m231_96+m232_96+m233_96+m234_96+m235_96+m236_96+m237_96+m238_96+m239_96+m240_96+m241_96+m242_96+m243_96+m244_96+m245_96+m246_96+m247_96+m248_96+m249_96+m250_96+m251_96+m252_96+m253_96+m254_96+m255_96+m256_96+m257_96+m258_96+m259_96+m260_96+m261_96+m262_96+m263_96+b96;
   assign out97 = m1_97+m2_97+m3_97+m4_97+m5_97+m6_97+m7_97+m8_97+m9_97+m10_97+m11_97+m12_97+m13_97+m14_97+m15_97+m16_97+m17_97+m18_97+m19_97+m20_97+m21_97+m22_97+m23_97+m24_97+m25_97+m26_97+m27_97+m28_97+m29_97+m30_97+m31_97+m32_97+m33_97+m34_97+m35_97+m36_97+m37_97+m38_97+m39_97+m40_97+m41_97+m42_97+m43_97+m44_97+m45_97+m46_97+m47_97+m48_97+m49_97+m50_97+m51_97+m52_97+m53_97+m54_97+m55_97+m56_97+m57_97+m58_97+m59_97+m60_97+m61_97+m62_97+m63_97+m64_97+m65_97+m66_97+m67_97+m68_97+m69_97+m70_97+m71_97+m72_97+m73_97+m74_97+m75_97+m76_97+m77_97+m78_97+m79_97+m80_97+m81_97+m82_97+m83_97+m84_97+m85_97+m86_97+m87_97+m88_97+m89_97+m90_97+m91_97+m92_97+m93_97+m94_97+m95_97+m96_97+m97_97+m98_97+m99_97+m100_97+m101_97+m102_97+m103_97+m104_97+m105_97+m106_97+m107_97+m108_97+m109_97+m110_97+m111_97+m112_97+m113_97+m114_97+m115_97+m116_97+m117_97+m118_97+m119_97+m120_97+m121_97+m122_97+m123_97+m124_97+m125_97+m126_97+m127_97+m128_97+m129_97+m130_97+m131_97+m132_97+m133_97+m134_97+m135_97+m136_97+m137_97+m138_97+m139_97+m140_97+m141_97+m142_97+m143_97+m144_97+m145_97+m146_97+m147_97+m148_97+m149_97+m150_97+m151_97+m152_97+m153_97+m154_97+m155_97+m156_97+m157_97+m158_97+m159_97+m160_97+m161_97+m162_97+m163_97+m164_97+m165_97+m166_97+m167_97+m168_97+m169_97+m170_97+m171_97+m172_97+m173_97+m174_97+m175_97+m176_97+m177_97+m178_97+m179_97+m180_97+m181_97+m182_97+m183_97+m184_97+m185_97+m186_97+m187_97+m188_97+m189_97+m190_97+m191_97+m192_97+m193_97+m194_97+m195_97+m196_97+m197_97+m198_97+m199_97+m200_97+m201_97+m202_97+m203_97+m204_97+m205_97+m206_97+m207_97+m208_97+m209_97+m210_97+m211_97+m212_97+m213_97+m214_97+m215_97+m216_97+m217_97+m218_97+m219_97+m220_97+m221_97+m222_97+m223_97+m224_97+m225_97+m226_97+m227_97+m228_97+m229_97+m230_97+m231_97+m232_97+m233_97+m234_97+m235_97+m236_97+m237_97+m238_97+m239_97+m240_97+m241_97+m242_97+m243_97+m244_97+m245_97+m246_97+m247_97+m248_97+m249_97+m250_97+m251_97+m252_97+m253_97+m254_97+m255_97+m256_97+m257_97+m258_97+m259_97+m260_97+m261_97+m262_97+m263_97+b97;
   assign out98 = m1_98+m2_98+m3_98+m4_98+m5_98+m6_98+m7_98+m8_98+m9_98+m10_98+m11_98+m12_98+m13_98+m14_98+m15_98+m16_98+m17_98+m18_98+m19_98+m20_98+m21_98+m22_98+m23_98+m24_98+m25_98+m26_98+m27_98+m28_98+m29_98+m30_98+m31_98+m32_98+m33_98+m34_98+m35_98+m36_98+m37_98+m38_98+m39_98+m40_98+m41_98+m42_98+m43_98+m44_98+m45_98+m46_98+m47_98+m48_98+m49_98+m50_98+m51_98+m52_98+m53_98+m54_98+m55_98+m56_98+m57_98+m58_98+m59_98+m60_98+m61_98+m62_98+m63_98+m64_98+m65_98+m66_98+m67_98+m68_98+m69_98+m70_98+m71_98+m72_98+m73_98+m74_98+m75_98+m76_98+m77_98+m78_98+m79_98+m80_98+m81_98+m82_98+m83_98+m84_98+m85_98+m86_98+m87_98+m88_98+m89_98+m90_98+m91_98+m92_98+m93_98+m94_98+m95_98+m96_98+m97_98+m98_98+m99_98+m100_98+m101_98+m102_98+m103_98+m104_98+m105_98+m106_98+m107_98+m108_98+m109_98+m110_98+m111_98+m112_98+m113_98+m114_98+m115_98+m116_98+m117_98+m118_98+m119_98+m120_98+m121_98+m122_98+m123_98+m124_98+m125_98+m126_98+m127_98+m128_98+m129_98+m130_98+m131_98+m132_98+m133_98+m134_98+m135_98+m136_98+m137_98+m138_98+m139_98+m140_98+m141_98+m142_98+m143_98+m144_98+m145_98+m146_98+m147_98+m148_98+m149_98+m150_98+m151_98+m152_98+m153_98+m154_98+m155_98+m156_98+m157_98+m158_98+m159_98+m160_98+m161_98+m162_98+m163_98+m164_98+m165_98+m166_98+m167_98+m168_98+m169_98+m170_98+m171_98+m172_98+m173_98+m174_98+m175_98+m176_98+m177_98+m178_98+m179_98+m180_98+m181_98+m182_98+m183_98+m184_98+m185_98+m186_98+m187_98+m188_98+m189_98+m190_98+m191_98+m192_98+m193_98+m194_98+m195_98+m196_98+m197_98+m198_98+m199_98+m200_98+m201_98+m202_98+m203_98+m204_98+m205_98+m206_98+m207_98+m208_98+m209_98+m210_98+m211_98+m212_98+m213_98+m214_98+m215_98+m216_98+m217_98+m218_98+m219_98+m220_98+m221_98+m222_98+m223_98+m224_98+m225_98+m226_98+m227_98+m228_98+m229_98+m230_98+m231_98+m232_98+m233_98+m234_98+m235_98+m236_98+m237_98+m238_98+m239_98+m240_98+m241_98+m242_98+m243_98+m244_98+m245_98+m246_98+m247_98+m248_98+m249_98+m250_98+m251_98+m252_98+m253_98+m254_98+m255_98+m256_98+m257_98+m258_98+m259_98+m260_98+m261_98+m262_98+m263_98+b98;
   assign out99 = m1_99+m2_99+m3_99+m4_99+m5_99+m6_99+m7_99+m8_99+m9_99+m10_99+m11_99+m12_99+m13_99+m14_99+m15_99+m16_99+m17_99+m18_99+m19_99+m20_99+m21_99+m22_99+m23_99+m24_99+m25_99+m26_99+m27_99+m28_99+m29_99+m30_99+m31_99+m32_99+m33_99+m34_99+m35_99+m36_99+m37_99+m38_99+m39_99+m40_99+m41_99+m42_99+m43_99+m44_99+m45_99+m46_99+m47_99+m48_99+m49_99+m50_99+m51_99+m52_99+m53_99+m54_99+m55_99+m56_99+m57_99+m58_99+m59_99+m60_99+m61_99+m62_99+m63_99+m64_99+m65_99+m66_99+m67_99+m68_99+m69_99+m70_99+m71_99+m72_99+m73_99+m74_99+m75_99+m76_99+m77_99+m78_99+m79_99+m80_99+m81_99+m82_99+m83_99+m84_99+m85_99+m86_99+m87_99+m88_99+m89_99+m90_99+m91_99+m92_99+m93_99+m94_99+m95_99+m96_99+m97_99+m98_99+m99_99+m100_99+m101_99+m102_99+m103_99+m104_99+m105_99+m106_99+m107_99+m108_99+m109_99+m110_99+m111_99+m112_99+m113_99+m114_99+m115_99+m116_99+m117_99+m118_99+m119_99+m120_99+m121_99+m122_99+m123_99+m124_99+m125_99+m126_99+m127_99+m128_99+m129_99+m130_99+m131_99+m132_99+m133_99+m134_99+m135_99+m136_99+m137_99+m138_99+m139_99+m140_99+m141_99+m142_99+m143_99+m144_99+m145_99+m146_99+m147_99+m148_99+m149_99+m150_99+m151_99+m152_99+m153_99+m154_99+m155_99+m156_99+m157_99+m158_99+m159_99+m160_99+m161_99+m162_99+m163_99+m164_99+m165_99+m166_99+m167_99+m168_99+m169_99+m170_99+m171_99+m172_99+m173_99+m174_99+m175_99+m176_99+m177_99+m178_99+m179_99+m180_99+m181_99+m182_99+m183_99+m184_99+m185_99+m186_99+m187_99+m188_99+m189_99+m190_99+m191_99+m192_99+m193_99+m194_99+m195_99+m196_99+m197_99+m198_99+m199_99+m200_99+m201_99+m202_99+m203_99+m204_99+m205_99+m206_99+m207_99+m208_99+m209_99+m210_99+m211_99+m212_99+m213_99+m214_99+m215_99+m216_99+m217_99+m218_99+m219_99+m220_99+m221_99+m222_99+m223_99+m224_99+m225_99+m226_99+m227_99+m228_99+m229_99+m230_99+m231_99+m232_99+m233_99+m234_99+m235_99+m236_99+m237_99+m238_99+m239_99+m240_99+m241_99+m242_99+m243_99+m244_99+m245_99+m246_99+m247_99+m248_99+m249_99+m250_99+m251_99+m252_99+m253_99+m254_99+m255_99+m256_99+m257_99+m258_99+m259_99+m260_99+m261_99+m262_99+m263_99+b99;
   assign out100 = m1_100+m2_100+m3_100+m4_100+m5_100+m6_100+m7_100+m8_100+m9_100+m10_100+m11_100+m12_100+m13_100+m14_100+m15_100+m16_100+m17_100+m18_100+m19_100+m20_100+m21_100+m22_100+m23_100+m24_100+m25_100+m26_100+m27_100+m28_100+m29_100+m30_100+m31_100+m32_100+m33_100+m34_100+m35_100+m36_100+m37_100+m38_100+m39_100+m40_100+m41_100+m42_100+m43_100+m44_100+m45_100+m46_100+m47_100+m48_100+m49_100+m50_100+m51_100+m52_100+m53_100+m54_100+m55_100+m56_100+m57_100+m58_100+m59_100+m60_100+m61_100+m62_100+m63_100+m64_100+m65_100+m66_100+m67_100+m68_100+m69_100+m70_100+m71_100+m72_100+m73_100+m74_100+m75_100+m76_100+m77_100+m78_100+m79_100+m80_100+m81_100+m82_100+m83_100+m84_100+m85_100+m86_100+m87_100+m88_100+m89_100+m90_100+m91_100+m92_100+m93_100+m94_100+m95_100+m96_100+m97_100+m98_100+m99_100+m100_100+m101_100+m102_100+m103_100+m104_100+m105_100+m106_100+m107_100+m108_100+m109_100+m110_100+m111_100+m112_100+m113_100+m114_100+m115_100+m116_100+m117_100+m118_100+m119_100+m120_100+m121_100+m122_100+m123_100+m124_100+m125_100+m126_100+m127_100+m128_100+m129_100+m130_100+m131_100+m132_100+m133_100+m134_100+m135_100+m136_100+m137_100+m138_100+m139_100+m140_100+m141_100+m142_100+m143_100+m144_100+m145_100+m146_100+m147_100+m148_100+m149_100+m150_100+m151_100+m152_100+m153_100+m154_100+m155_100+m156_100+m157_100+m158_100+m159_100+m160_100+m161_100+m162_100+m163_100+m164_100+m165_100+m166_100+m167_100+m168_100+m169_100+m170_100+m171_100+m172_100+m173_100+m174_100+m175_100+m176_100+m177_100+m178_100+m179_100+m180_100+m181_100+m182_100+m183_100+m184_100+m185_100+m186_100+m187_100+m188_100+m189_100+m190_100+m191_100+m192_100+m193_100+m194_100+m195_100+m196_100+m197_100+m198_100+m199_100+m200_100+m201_100+m202_100+m203_100+m204_100+m205_100+m206_100+m207_100+m208_100+m209_100+m210_100+m211_100+m212_100+m213_100+m214_100+m215_100+m216_100+m217_100+m218_100+m219_100+m220_100+m221_100+m222_100+m223_100+m224_100+m225_100+m226_100+m227_100+m228_100+m229_100+m230_100+m231_100+m232_100+m233_100+m234_100+m235_100+m236_100+m237_100+m238_100+m239_100+m240_100+m241_100+m242_100+m243_100+m244_100+m245_100+m246_100+m247_100+m248_100+m249_100+m250_100+m251_100+m252_100+m253_100+m254_100+m255_100+m256_100+m257_100+m258_100+m259_100+m260_100+m261_100+m262_100+m263_100+b100;
endmodule