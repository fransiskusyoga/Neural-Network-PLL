module test_layer_1(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27);
   input signed [5:0] in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80;
   output signed [6:0] out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27;
   wire signed [5:0] neg1,neg2,neg3,neg4,neg5,neg6,neg7,neg8,neg9,neg10,neg11,neg12,neg13,neg14,neg15,neg16,neg17,neg18,neg19,neg20,neg21,neg22,neg23,neg24,neg25,neg26,neg27,neg28,neg29,neg30,neg31,neg32,neg33,neg34,neg35,neg36,neg37,neg38,neg39,neg40,neg41,neg42,neg43,neg44,neg45,neg46,neg47,neg48,neg49,neg50,neg51,neg52,neg53,neg54,neg55,neg56,neg57,neg58,neg59,neg60,neg61,neg62,neg63,neg64,neg65,neg66,neg67,neg68,neg69,neg70,neg71,neg72,neg73,neg74,neg75,neg76,neg77,neg78,neg79,neg80;

   //Bias value
   wire signed [6:0] b1 = $signed(7'h0);
   wire signed [6:0] b2 = $signed(7'h1);
   wire signed [6:0] b3 = $signed(7'h1);
   wire signed [6:0] b4 = $signed(7'h0);
   wire signed [6:0] b5 = $signed(7'h1);
   wire signed [6:0] b6 = $signed(7'h1);
   wire signed [6:0] b7 = $signed(7'h1);
   wire signed [6:0] b8 = $signed(7'h0);
   wire signed [6:0] b9 = $signed(7'h1);
   wire signed [6:0] b10 = $signed(7'h0);
   wire signed [6:0] b11 = $signed(7'h1);
   wire signed [6:0] b12 = $signed(7'h1);
   wire signed [6:0] b13 = $signed(7'h2);
   wire signed [6:0] b14 = $signed(7'h1);
   wire signed [6:0] b15 = $signed(7'h0);
   wire signed [6:0] b16 = $signed(7'h0);
   wire signed [6:0] b17 = $signed(7'h0);
   wire signed [6:0] b18 = $signed(7'h0);
   wire signed [6:0] b19 = $signed(7'h3);
   wire signed [6:0] b20 = $signed(7'h0);
   wire signed [6:0] b21 = $signed(7'h1);
   wire signed [6:0] b22 = $signed(7'h1);
   wire signed [6:0] b23 = $signed(7'h0);
   wire signed [6:0] b24 = $signed(7'h1);
   wire signed [6:0] b25 = $signed(7'h0);
   wire signed [6:0] b26 = $signed(7'h0);
   wire signed [6:0] b27 = $signed(7'h1);

   //Negation modules
   negate #(6) N1(in1,neg1);
   negate #(6) N2(in2,neg2);
   negate #(6) N3(in3,neg3);
   negate #(6) N4(in4,neg4);
   negate #(6) N5(in5,neg5);
   negate #(6) N6(in6,neg6);
   negate #(6) N7(in7,neg7);
   negate #(6) N8(in8,neg8);
   negate #(6) N9(in9,neg9);
   negate #(6) N10(in10,neg10);
   negate #(6) N11(in11,neg11);
   negate #(6) N12(in12,neg12);
   negate #(6) N13(in13,neg13);
   negate #(6) N14(in14,neg14);
   negate #(6) N15(in15,neg15);
   negate #(6) N16(in16,neg16);
   negate #(6) N17(in17,neg17);
   negate #(6) N18(in18,neg18);
   negate #(6) N19(in19,neg19);
   negate #(6) N20(in20,neg20);
   negate #(6) N21(in21,neg21);
   negate #(6) N22(in22,neg22);
   negate #(6) N23(in23,neg23);
   negate #(6) N24(in24,neg24);
   negate #(6) N25(in25,neg25);
   negate #(6) N26(in26,neg26);
   negate #(6) N27(in27,neg27);
   negate #(6) N28(in28,neg28);
   negate #(6) N29(in29,neg29);
   negate #(6) N30(in30,neg30);
   negate #(6) N31(in31,neg31);
   negate #(6) N32(in32,neg32);
   negate #(6) N33(in33,neg33);
   negate #(6) N34(in34,neg34);
   negate #(6) N35(in35,neg35);
   negate #(6) N36(in36,neg36);
   negate #(6) N37(in37,neg37);
   negate #(6) N38(in38,neg38);
   negate #(6) N39(in39,neg39);
   negate #(6) N40(in40,neg40);
   negate #(6) N41(in41,neg41);
   negate #(6) N42(in42,neg42);
   negate #(6) N43(in43,neg43);
   negate #(6) N44(in44,neg44);
   negate #(6) N45(in45,neg45);
   negate #(6) N46(in46,neg46);
   negate #(6) N47(in47,neg47);
   negate #(6) N48(in48,neg48);
   negate #(6) N49(in49,neg49);
   negate #(6) N50(in50,neg50);
   negate #(6) N51(in51,neg51);
   negate #(6) N52(in52,neg52);
   negate #(6) N53(in53,neg53);
   negate #(6) N54(in54,neg54);
   negate #(6) N55(in55,neg55);
   negate #(6) N56(in56,neg56);
   negate #(6) N57(in57,neg57);
   negate #(6) N58(in58,neg58);
   negate #(6) N59(in59,neg59);
   negate #(6) N60(in60,neg60);
   negate #(6) N61(in61,neg61);
   negate #(6) N62(in62,neg62);
   negate #(6) N63(in63,neg63);
   negate #(6) N64(in64,neg64);
   negate #(6) N65(in65,neg65);
   negate #(6) N66(in66,neg66);
   negate #(6) N67(in67,neg67);
   negate #(6) N68(in68,neg68);
   negate #(6) N69(in69,neg69);
   negate #(6) N70(in70,neg70);
   negate #(6) N71(in71,neg71);
   negate #(6) N72(in72,neg72);
   negate #(6) N73(in73,neg73);
   negate #(6) N74(in74,neg74);
   negate #(6) N75(in75,neg75);
   negate #(6) N76(in76,neg76);
   negate #(6) N77(in77,neg77);
   negate #(6) N78(in78,neg78);
   negate #(6) N79(in79,neg79);
   negate #(6) N80(in80,neg80);

   // m1_1 = W*in
   wire signed [6:0] m1_1;
   assign m1_1 =7'b0;

   // m1_2 = W*in
   wire signed [6:0] m1_2;
   assign m1_2 =7'b0;

   // m1_3 = W*in
   wire signed [6:0] m1_3;
   assign m1_3 =7'b0;

   // m1_4 = W*in
   wire signed [6:0] m1_4;
   assign m1_4 =7'b0;

   // m1_5 = W*in
   wire signed [6:0] m1_5;
   assign m1_5 =7'b0;

   // m1_6 = W*in
   wire signed [6:0] m1_6;
   assign m1_6 =7'b0;

   // m1_7 = W*in
   wire signed [6:0] m1_7;
   assign m1_7 =7'b0;

   // m1_8 = W*in
   wire signed [6:0] m1_8;
   assign m1_8 =7'b0;

   // m1_9 = W*in
   wire signed [6:0] m1_9;
   assign m1_9 =7'b0;

   // m1_10 = W*in
   wire signed [6:0] m1_10;
   assign m1_10 =7'b0;

   // m1_11 = W*in
   wire signed [6:0] m1_11;
   assign m1_11 =7'b0;

   // m1_12 = W*in
   wire signed [6:0] m1_12;
   assign m1_12 =7'b0;

   // m1_13 = W*in
   wire signed [6:0] m1_13;
   assign m1_13 =7'b0;

   // m1_14 = W*in
   wire signed [6:0] m1_14;
   assign m1_14 =7'b0;

   // m1_15 = W*in
   wire signed [6:0] m1_15;
   assign m1_15 =7'b0;

   // m1_16 = W*in
   wire signed [6:0] m1_16;
   assign m1_16 =7'b0;

   // m1_17 = W*in
   wire signed [6:0] m1_17;
   assign m1_17 =7'b0;

   // m1_18 = W*in
   wire signed [6:0] m1_18;
   assign m1_18 ={ {2{in1[5]}} , in1[5:1] };

   // m1_19 = W*in
   wire signed [6:0] m1_19;
   assign m1_19 =7'b0;

   // m1_20 = W*in
   wire signed [6:0] m1_20;
   assign m1_20 =7'b0;

   // m1_21 = W*in
   wire signed [6:0] m1_21;
   assign m1_21 =7'b0;

   // m1_22 = W*in
   wire signed [6:0] m1_22;
   assign m1_22 =7'b0;

   // m1_23 = W*in
   wire signed [6:0] m1_23;
   assign m1_23 =7'b0;

   // m1_24 = W*in
   wire signed [6:0] m1_24;
   assign m1_24 =7'b0;

   // m1_25 = W*in
   wire signed [6:0] m1_25;
   assign m1_25 =7'b0;

   // m1_26 = W*in
   wire signed [6:0] m1_26;
   assign m1_26 =7'b0;

   // m1_27 = W*in
   wire signed [6:0] m1_27;
   assign m1_27 =7'b0;

   // m2_1 = W*in
   wire signed [6:0] m2_1;
   assign m2_1 =7'b0;

   // m2_2 = W*in
   wire signed [6:0] m2_2;
   assign m2_2 =7'b0;

   // m2_3 = W*in
   wire signed [6:0] m2_3;
   assign m2_3 =7'b0;

   // m2_4 = W*in
   wire signed [6:0] m2_4;
   assign m2_4 ={ {2{in2[5]}} , in2[5:1] };

   // m2_5 = W*in
   wire signed [6:0] m2_5;
   assign m2_5 =7'b0;

   // m2_6 = W*in
   wire signed [6:0] m2_6;
   assign m2_6 =7'b0;

   // m2_7 = W*in
   wire signed [6:0] m2_7;
   assign m2_7 =7'b0;

   // m2_8 = W*in
   wire signed [6:0] m2_8;
   assign m2_8 =7'b0;

   // m2_9 = W*in
   wire signed [6:0] m2_9;
   assign m2_9 =7'b0;

   // m2_10 = W*in
   wire signed [6:0] m2_10;
   assign m2_10 =7'b0;

   // m2_11 = W*in
   wire signed [6:0] m2_11;
   assign m2_11 =7'b0;

   // m2_12 = W*in
   wire signed [6:0] m2_12;
   assign m2_12 =7'b0;

   // m2_13 = W*in
   wire signed [6:0] m2_13;
   assign m2_13 =7'b0;

   // m2_14 = W*in
   wire signed [6:0] m2_14;
   assign m2_14 =7'b0;

   // m2_15 = W*in
   wire signed [6:0] m2_15;
   assign m2_15 =7'b0;

   // m2_16 = W*in
   wire signed [6:0] m2_16;
   assign m2_16 =7'b0;

   // m2_17 = W*in
   wire signed [6:0] m2_17;
   assign m2_17 =7'b0;

   // m2_18 = W*in
   wire signed [6:0] m2_18;
   assign m2_18 =7'b0;

   // m2_19 = W*in
   wire signed [6:0] m2_19;
   assign m2_19 =7'b0;

   // m2_20 = W*in
   wire signed [6:0] m2_20;
   assign m2_20 =7'b0;

   // m2_21 = W*in
   wire signed [6:0] m2_21;
   assign m2_21 =7'b0;

   // m2_22 = W*in
   wire signed [6:0] m2_22;
   assign m2_22 =7'b0;

   // m2_23 = W*in
   wire signed [6:0] m2_23;
   assign m2_23 =7'b0;

   // m2_24 = W*in
   wire signed [6:0] m2_24;
   assign m2_24 =7'b0;

   // m2_25 = W*in
   wire signed [6:0] m2_25;
   assign m2_25 =7'b0;

   // m2_26 = W*in
   wire signed [6:0] m2_26;
   assign m2_26 =7'b0;

   // m2_27 = W*in
   wire signed [6:0] m2_27;
   assign m2_27 =7'b0;

   // m3_1 = W*in
   wire signed [6:0] m3_1;
   assign m3_1 =7'b0;

   // m3_2 = W*in
   wire signed [6:0] m3_2;
   assign m3_2 =7'b0;

   // m3_3 = W*in
   wire signed [6:0] m3_3;
   assign m3_3 =7'b0;

   // m3_4 = W*in
   wire signed [6:0] m3_4;
   assign m3_4 =7'b0;

   // m3_5 = W*in
   wire signed [6:0] m3_5;
   assign m3_5 =7'b0;

   // m3_6 = W*in
   wire signed [6:0] m3_6;
   assign m3_6 =7'b0;

   // m3_7 = W*in
   wire signed [6:0] m3_7;
   assign m3_7 ={ {2{in3[5]}} , in3[5:1] };

   // m3_8 = W*in
   wire signed [6:0] m3_8;
   assign m3_8 =7'b0;

   // m3_9 = W*in
   wire signed [6:0] m3_9;
   assign m3_9 =7'b0;

   // m3_10 = W*in
   wire signed [6:0] m3_10;
   assign m3_10 =7'b0;

   // m3_11 = W*in
   wire signed [6:0] m3_11;
   assign m3_11 =7'b0;

   // m3_12 = W*in
   wire signed [6:0] m3_12;
   assign m3_12 =7'b0;

   // m3_13 = W*in
   wire signed [6:0] m3_13;
   assign m3_13 =7'b0;

   // m3_14 = W*in
   wire signed [6:0] m3_14;
   assign m3_14 =7'b0;

   // m3_15 = W*in
   wire signed [6:0] m3_15;
   assign m3_15 =7'b0;

   // m3_16 = W*in
   wire signed [6:0] m3_16;
   assign m3_16 =7'b0;

   // m3_17 = W*in
   wire signed [6:0] m3_17;
   assign m3_17 =7'b0;

   // m3_18 = W*in
   wire signed [6:0] m3_18;
   assign m3_18 =7'b0;

   // m3_19 = W*in
   wire signed [6:0] m3_19;
   assign m3_19 =7'b0;

   // m3_20 = W*in
   wire signed [6:0] m3_20;
   assign m3_20 =7'b0;

   // m3_21 = W*in
   wire signed [6:0] m3_21;
   assign m3_21 =7'b0;

   // m3_22 = W*in
   wire signed [6:0] m3_22;
   assign m3_22 =7'b0;

   // m3_23 = W*in
   wire signed [6:0] m3_23;
   assign m3_23 =7'b0;

   // m3_24 = W*in
   wire signed [6:0] m3_24;
   assign m3_24 =7'b0;

   // m3_25 = W*in
   wire signed [6:0] m3_25;
   assign m3_25 =7'b0;

   // m3_26 = W*in
   wire signed [6:0] m3_26;
   assign m3_26 =7'b0;

   // m3_27 = W*in
   wire signed [6:0] m3_27;
   assign m3_27 ={ {1{in3[5]}} , in3[5:0] };

   // m4_1 = W*in
   wire signed [6:0] m4_1;
   assign m4_1 =7'b0;

   // m4_2 = W*in
   wire signed [6:0] m4_2;
   assign m4_2 =7'b0;

   // m4_3 = W*in
   wire signed [6:0] m4_3;
   assign m4_3 =7'b0;

   // m4_4 = W*in
   wire signed [6:0] m4_4;
   assign m4_4 =7'b0;

   // m4_5 = W*in
   wire signed [6:0] m4_5;
   assign m4_5 =7'b0;

   // m4_6 = W*in
   wire signed [6:0] m4_6;
   assign m4_6 =7'b0;

   // m4_7 = W*in
   wire signed [6:0] m4_7;
   assign m4_7 =7'b0;

   // m4_8 = W*in
   wire signed [6:0] m4_8;
   assign m4_8 =7'b0;

   // m4_9 = W*in
   wire signed [6:0] m4_9;
   assign m4_9 =7'b0;

   // m4_10 = W*in
   wire signed [6:0] m4_10;
   assign m4_10 =7'b0;

   // m4_11 = W*in
   wire signed [6:0] m4_11;
   assign m4_11 =7'b0;

   // m4_12 = W*in
   wire signed [6:0] m4_12;
   assign m4_12 =7'b0;

   // m4_13 = W*in
   wire signed [6:0] m4_13;
   assign m4_13 =7'b0;

   // m4_14 = W*in
   wire signed [6:0] m4_14;
   assign m4_14 =7'b0;

   // m4_15 = W*in
   wire signed [6:0] m4_15;
   assign m4_15 =7'b0;

   // m4_16 = W*in
   wire signed [6:0] m4_16;
   assign m4_16 ={ {1{in4[5]}} , in4[5:0] };

   // m4_17 = W*in
   wire signed [6:0] m4_17;
   assign m4_17 =7'b0;

   // m4_18 = W*in
   wire signed [6:0] m4_18;
   assign m4_18 =7'b0;

   // m4_19 = W*in
   wire signed [6:0] m4_19;
   assign m4_19 =7'b0;

   // m4_20 = W*in
   wire signed [6:0] m4_20;
   assign m4_20 =7'b0;

   // m4_21 = W*in
   wire signed [6:0] m4_21;
   assign m4_21 =7'b0;

   // m4_22 = W*in
   wire signed [6:0] m4_22;
   assign m4_22 =7'b0;

   // m4_23 = W*in
   wire signed [6:0] m4_23;
   assign m4_23 =7'b0;

   // m4_24 = W*in
   wire signed [6:0] m4_24;
   assign m4_24 =7'b0;

   // m4_25 = W*in
   wire signed [6:0] m4_25;
   assign m4_25 =7'b0;

   // m4_26 = W*in
   wire signed [6:0] m4_26;
   assign m4_26 =7'b0;

   // m4_27 = W*in
   wire signed [6:0] m4_27;
   assign m4_27 =7'b0;

   // m5_1 = W*in
   wire signed [6:0] m5_1;
   assign m5_1 =7'b0;

   // m5_2 = W*in
   wire signed [6:0] m5_2;
   assign m5_2 =7'b0;

   // m5_3 = W*in
   wire signed [6:0] m5_3;
   assign m5_3 =7'b0;

   // m5_4 = W*in
   wire signed [6:0] m5_4;
   assign m5_4 =7'b0;

   // m5_5 = W*in
   wire signed [6:0] m5_5;
   assign m5_5 =7'b0;

   // m5_6 = W*in
   wire signed [6:0] m5_6;
   assign m5_6 =7'b0;

   // m5_7 = W*in
   wire signed [6:0] m5_7;
   assign m5_7 =7'b0;

   // m5_8 = W*in
   wire signed [6:0] m5_8;
   assign m5_8 =7'b0;

   // m5_9 = W*in
   wire signed [6:0] m5_9;
   assign m5_9 =7'b0;

   // m5_10 = W*in
   wire signed [6:0] m5_10;
   assign m5_10 =7'b0;

   // m5_11 = W*in
   wire signed [6:0] m5_11;
   assign m5_11 =7'b0;

   // m5_12 = W*in
   wire signed [6:0] m5_12;
   assign m5_12 =7'b0;

   // m5_13 = W*in
   wire signed [6:0] m5_13;
   assign m5_13 =7'b0;

   // m5_14 = W*in
   wire signed [6:0] m5_14;
   assign m5_14 =7'b0;

   // m5_15 = W*in
   wire signed [6:0] m5_15;
   assign m5_15 =7'b0;

   // m5_16 = W*in
   wire signed [6:0] m5_16;
   assign m5_16 =7'b0;

   // m5_17 = W*in
   wire signed [6:0] m5_17;
   assign m5_17 =7'b0;

   // m5_18 = W*in
   wire signed [6:0] m5_18;
   assign m5_18 =7'b0;

   // m5_19 = W*in
   wire signed [6:0] m5_19;
   assign m5_19 =7'b0;

   // m5_20 = W*in
   wire signed [6:0] m5_20;
   assign m5_20 =7'b0;

   // m5_21 = W*in
   wire signed [6:0] m5_21;
   wire signed [7:0] tm5_21;
   assign tm5_21[0:0] = in5[0:0];
   assign tm5_21[7:1] = { {1{in5[5]}} , in5[5:0] } + { {2{in5[5]}} , in5[5:1] };
   assign m5_21 ={ {1{tm5_21[7]}} , tm5_21[7:2] };

   // m5_22 = W*in
   wire signed [6:0] m5_22;
   assign m5_22 =7'b0;

   // m5_23 = W*in
   wire signed [6:0] m5_23;
   assign m5_23 =7'b0;

   // m5_24 = W*in
   wire signed [6:0] m5_24;
   assign m5_24 =7'b0;

   // m5_25 = W*in
   wire signed [6:0] m5_25;
   assign m5_25 =7'b0;

   // m5_26 = W*in
   wire signed [6:0] m5_26;
   assign m5_26 =7'b0;

   // m5_27 = W*in
   wire signed [6:0] m5_27;
   assign m5_27 =7'b0;

   // m6_1 = W*in
   wire signed [6:0] m6_1;
   assign m6_1 =7'b0;

   // m6_2 = W*in
   wire signed [6:0] m6_2;
   assign m6_2 =7'b0;

   // m6_3 = W*in
   wire signed [6:0] m6_3;
   assign m6_3 =7'b0;

   // m6_4 = W*in
   wire signed [6:0] m6_4;
   assign m6_4 =7'b0;

   // m6_5 = W*in
   wire signed [6:0] m6_5;
   assign m6_5 =7'b0;

   // m6_6 = W*in
   wire signed [6:0] m6_6;
   assign m6_6 =7'b0;

   // m6_7 = W*in
   wire signed [6:0] m6_7;
   assign m6_7 =7'b0;

   // m6_8 = W*in
   wire signed [6:0] m6_8;
   assign m6_8 =7'b0;

   // m6_9 = W*in
   wire signed [6:0] m6_9;
   assign m6_9 =7'b0;

   // m6_10 = W*in
   wire signed [6:0] m6_10;
   assign m6_10 =7'b0;

   // m6_11 = W*in
   wire signed [6:0] m6_11;
   assign m6_11 =7'b0;

   // m6_12 = W*in
   wire signed [6:0] m6_12;
   assign m6_12 ={ {2{neg6[5]}} , neg6[5:1] };

   // m6_13 = W*in
   wire signed [6:0] m6_13;
   assign m6_13 =7'b0;

   // m6_14 = W*in
   wire signed [6:0] m6_14;
   assign m6_14 =7'b0;

   // m6_15 = W*in
   wire signed [6:0] m6_15;
   assign m6_15 =7'b0;

   // m6_16 = W*in
   wire signed [6:0] m6_16;
   assign m6_16 =7'b0;

   // m6_17 = W*in
   wire signed [6:0] m6_17;
   assign m6_17 =7'b0;

   // m6_18 = W*in
   wire signed [6:0] m6_18;
   assign m6_18 =7'b0;

   // m6_19 = W*in
   wire signed [6:0] m6_19;
   assign m6_19 =7'b0;

   // m6_20 = W*in
   wire signed [6:0] m6_20;
   assign m6_20 =7'b0;

   // m6_21 = W*in
   wire signed [6:0] m6_21;
   assign m6_21 =7'b0;

   // m6_22 = W*in
   wire signed [6:0] m6_22;
   assign m6_22 =7'b0;

   // m6_23 = W*in
   wire signed [6:0] m6_23;
   assign m6_23 =7'b0;

   // m6_24 = W*in
   wire signed [6:0] m6_24;
   assign m6_24 =7'b0;

   // m6_25 = W*in
   wire signed [6:0] m6_25;
   assign m6_25 =7'b0;

   // m6_26 = W*in
   wire signed [6:0] m6_26;
   assign m6_26 =7'b0;

   // m6_27 = W*in
   wire signed [6:0] m6_27;
   assign m6_27 =7'b0;

   // m7_1 = W*in
   wire signed [6:0] m7_1;
   assign m7_1 =7'b0;

   // m7_2 = W*in
   wire signed [6:0] m7_2;
   assign m7_2 =7'b0;

   // m7_3 = W*in
   wire signed [6:0] m7_3;
   assign m7_3 =7'b0;

   // m7_4 = W*in
   wire signed [6:0] m7_4;
   assign m7_4 =7'b0;

   // m7_5 = W*in
   wire signed [6:0] m7_5;
   assign m7_5 =7'b0;

   // m7_6 = W*in
   wire signed [6:0] m7_6;
   assign m7_6 =7'b0;

   // m7_7 = W*in
   wire signed [6:0] m7_7;
   assign m7_7 =7'b0;

   // m7_8 = W*in
   wire signed [6:0] m7_8;
   assign m7_8 =7'b0;

   // m7_9 = W*in
   wire signed [6:0] m7_9;
   assign m7_9 =7'b0;

   // m7_10 = W*in
   wire signed [6:0] m7_10;
   assign m7_10 =7'b0;

   // m7_11 = W*in
   wire signed [6:0] m7_11;
   assign m7_11 =7'b0;

   // m7_12 = W*in
   wire signed [6:0] m7_12;
   assign m7_12 =7'b0;

   // m7_13 = W*in
   wire signed [6:0] m7_13;
   assign m7_13 =7'b0;

   // m7_14 = W*in
   wire signed [6:0] m7_14;
   assign m7_14 =7'b0;

   // m7_15 = W*in
   wire signed [6:0] m7_15;
   assign m7_15 =7'b0;

   // m7_16 = W*in
   wire signed [6:0] m7_16;
   assign m7_16 =7'b0;

   // m7_17 = W*in
   wire signed [6:0] m7_17;
   assign m7_17 =7'b0;

   // m7_18 = W*in
   wire signed [6:0] m7_18;
   assign m7_18 =7'b0;

   // m7_19 = W*in
   wire signed [6:0] m7_19;
   assign m7_19 =7'b0;

   // m7_20 = W*in
   wire signed [6:0] m7_20;
   assign m7_20 =7'b0;

   // m7_21 = W*in
   wire signed [6:0] m7_21;
   assign m7_21 ={ {2{in7[5]}} , in7[5:1] };

   // m7_22 = W*in
   wire signed [6:0] m7_22;
   assign m7_22 ={ {2{in7[5]}} , in7[5:1] };

   // m7_23 = W*in
   wire signed [6:0] m7_23;
   assign m7_23 =7'b0;

   // m7_24 = W*in
   wire signed [6:0] m7_24;
   assign m7_24 =7'b0;

   // m7_25 = W*in
   wire signed [6:0] m7_25;
   assign m7_25 =7'b0;

   // m7_26 = W*in
   wire signed [6:0] m7_26;
   assign m7_26 =7'b0;

   // m7_27 = W*in
   wire signed [6:0] m7_27;
   assign m7_27 =7'b0;

   // m8_1 = W*in
   wire signed [6:0] m8_1;
   assign m8_1 =7'b0;

   // m8_2 = W*in
   wire signed [6:0] m8_2;
   assign m8_2 ={ {2{in8[5]}} , in8[5:1] };

   // m8_3 = W*in
   wire signed [6:0] m8_3;
   assign m8_3 =7'b0;

   // m8_4 = W*in
   wire signed [6:0] m8_4;
   assign m8_4 =7'b0;

   // m8_5 = W*in
   wire signed [6:0] m8_5;
   assign m8_5 =7'b0;

   // m8_6 = W*in
   wire signed [6:0] m8_6;
   assign m8_6 =7'b0;

   // m8_7 = W*in
   wire signed [6:0] m8_7;
   assign m8_7 =7'b0;

   // m8_8 = W*in
   wire signed [6:0] m8_8;
   assign m8_8 =7'b0;

   // m8_9 = W*in
   wire signed [6:0] m8_9;
   assign m8_9 =7'b0;

   // m8_10 = W*in
   wire signed [6:0] m8_10;
   assign m8_10 =7'b0;

   // m8_11 = W*in
   wire signed [6:0] m8_11;
   assign m8_11 =7'b0;

   // m8_12 = W*in
   wire signed [6:0] m8_12;
   assign m8_12 =7'b0;

   // m8_13 = W*in
   wire signed [6:0] m8_13;
   assign m8_13 =7'b0;

   // m8_14 = W*in
   wire signed [6:0] m8_14;
   assign m8_14 =7'b0;

   // m8_15 = W*in
   wire signed [6:0] m8_15;
   assign m8_15 =7'b0;

   // m8_16 = W*in
   wire signed [6:0] m8_16;
   assign m8_16 =7'b0;

   // m8_17 = W*in
   wire signed [6:0] m8_17;
   assign m8_17 =7'b0;

   // m8_18 = W*in
   wire signed [6:0] m8_18;
   assign m8_18 =7'b0;

   // m8_19 = W*in
   wire signed [6:0] m8_19;
   assign m8_19 =7'b0;

   // m8_20 = W*in
   wire signed [6:0] m8_20;
   assign m8_20 =7'b0;

   // m8_21 = W*in
   wire signed [6:0] m8_21;
   assign m8_21 =7'b0;

   // m8_22 = W*in
   wire signed [6:0] m8_22;
   assign m8_22 =7'b0;

   // m8_23 = W*in
   wire signed [6:0] m8_23;
   assign m8_23 =7'b0;

   // m8_24 = W*in
   wire signed [6:0] m8_24;
   assign m8_24 =7'b0;

   // m8_25 = W*in
   wire signed [6:0] m8_25;
   assign m8_25 =7'b0;

   // m8_26 = W*in
   wire signed [6:0] m8_26;
   assign m8_26 =7'b0;

   // m8_27 = W*in
   wire signed [6:0] m8_27;
   assign m8_27 =7'b0;

   // m9_1 = W*in
   wire signed [6:0] m9_1;
   assign m9_1 =7'b0;

   // m9_2 = W*in
   wire signed [6:0] m9_2;
   assign m9_2 =7'b0;

   // m9_3 = W*in
   wire signed [6:0] m9_3;
   assign m9_3 =7'b0;

   // m9_4 = W*in
   wire signed [6:0] m9_4;
   assign m9_4 =7'b0;

   // m9_5 = W*in
   wire signed [6:0] m9_5;
   assign m9_5 =7'b0;

   // m9_6 = W*in
   wire signed [6:0] m9_6;
   assign m9_6 =7'b0;

   // m9_7 = W*in
   wire signed [6:0] m9_7;
   assign m9_7 =7'b0;

   // m9_8 = W*in
   wire signed [6:0] m9_8;
   assign m9_8 =7'b0;

   // m9_9 = W*in
   wire signed [6:0] m9_9;
   assign m9_9 =7'b0;

   // m9_10 = W*in
   wire signed [6:0] m9_10;
   assign m9_10 =7'b0;

   // m9_11 = W*in
   wire signed [6:0] m9_11;
   assign m9_11 =7'b0;

   // m9_12 = W*in
   wire signed [6:0] m9_12;
   assign m9_12 ={ {1{in9[5]}} , in9[5:0] };

   // m9_13 = W*in
   wire signed [6:0] m9_13;
   assign m9_13 =7'b0;

   // m9_14 = W*in
   wire signed [6:0] m9_14;
   assign m9_14 =7'b0;

   // m9_15 = W*in
   wire signed [6:0] m9_15;
   assign m9_15 =7'b0;

   // m9_16 = W*in
   wire signed [6:0] m9_16;
   assign m9_16 =7'b0;

   // m9_17 = W*in
   wire signed [6:0] m9_17;
   assign m9_17 =7'b0;

   // m9_18 = W*in
   wire signed [6:0] m9_18;
   assign m9_18 =7'b0;

   // m9_19 = W*in
   wire signed [6:0] m9_19;
   assign m9_19 =7'b0;

   // m9_20 = W*in
   wire signed [6:0] m9_20;
   assign m9_20 =7'b0;

   // m9_21 = W*in
   wire signed [6:0] m9_21;
   assign m9_21 =7'b0;

   // m9_22 = W*in
   wire signed [6:0] m9_22;
   assign m9_22 =7'b0;

   // m9_23 = W*in
   wire signed [6:0] m9_23;
   assign m9_23 =7'b0;

   // m9_24 = W*in
   wire signed [6:0] m9_24;
   assign m9_24 =7'b0;

   // m9_25 = W*in
   wire signed [6:0] m9_25;
   assign m9_25 =7'b0;

   // m9_26 = W*in
   wire signed [6:0] m9_26;
   assign m9_26 =7'b0;

   // m9_27 = W*in
   wire signed [6:0] m9_27;
   assign m9_27 =7'b0;

   // m10_1 = W*in
   wire signed [6:0] m10_1;
   assign m10_1 =7'b0;

   // m10_2 = W*in
   wire signed [6:0] m10_2;
   assign m10_2 =7'b0;

   // m10_3 = W*in
   wire signed [6:0] m10_3;
   assign m10_3 =7'b0;

   // m10_4 = W*in
   wire signed [6:0] m10_4;
   assign m10_4 =7'b0;

   // m10_5 = W*in
   wire signed [6:0] m10_5;
   assign m10_5 =7'b0;

   // m10_6 = W*in
   wire signed [6:0] m10_6;
   assign m10_6 =7'b0;

   // m10_7 = W*in
   wire signed [6:0] m10_7;
   assign m10_7 =7'b0;

   // m10_8 = W*in
   wire signed [6:0] m10_8;
   assign m10_8 =7'b0;

   // m10_9 = W*in
   wire signed [6:0] m10_9;
   assign m10_9 =7'b0;

   // m10_10 = W*in
   wire signed [6:0] m10_10;
   assign m10_10 =7'b0;

   // m10_11 = W*in
   wire signed [6:0] m10_11;
   assign m10_11 =7'b0;

   // m10_12 = W*in
   wire signed [6:0] m10_12;
   assign m10_12 =7'b0;

   // m10_13 = W*in
   wire signed [6:0] m10_13;
   assign m10_13 =7'b0;

   // m10_14 = W*in
   wire signed [6:0] m10_14;
   assign m10_14 =7'b0;

   // m10_15 = W*in
   wire signed [6:0] m10_15;
   assign m10_15 =7'b0;

   // m10_16 = W*in
   wire signed [6:0] m10_16;
   wire signed [7:0] tm10_16;
   assign tm10_16[0:0] = in10[0:0];
   assign tm10_16[7:1] = { {1{in10[5]}} , in10[5:0] } + { {2{in10[5]}} , in10[5:1] };
   assign m10_16 ={ {1{tm10_16[7]}} , tm10_16[7:2] };

   // m10_17 = W*in
   wire signed [6:0] m10_17;
   assign m10_17 =7'b0;

   // m10_18 = W*in
   wire signed [6:0] m10_18;
   assign m10_18 =7'b0;

   // m10_19 = W*in
   wire signed [6:0] m10_19;
   assign m10_19 =7'b0;

   // m10_20 = W*in
   wire signed [6:0] m10_20;
   assign m10_20 =7'b0;

   // m10_21 = W*in
   wire signed [6:0] m10_21;
   assign m10_21 =7'b0;

   // m10_22 = W*in
   wire signed [6:0] m10_22;
   assign m10_22 =7'b0;

   // m10_23 = W*in
   wire signed [6:0] m10_23;
   assign m10_23 =7'b0;

   // m10_24 = W*in
   wire signed [6:0] m10_24;
   assign m10_24 =7'b0;

   // m10_25 = W*in
   wire signed [6:0] m10_25;
   assign m10_25 =7'b0;

   // m10_26 = W*in
   wire signed [6:0] m10_26;
   assign m10_26 =7'b0;

   // m10_27 = W*in
   wire signed [6:0] m10_27;
   assign m10_27 =7'b0;

   // m11_1 = W*in
   wire signed [6:0] m11_1;
   assign m11_1 ={ {2{in11[5]}} , in11[5:1] };

   // m11_2 = W*in
   wire signed [6:0] m11_2;
   assign m11_2 =7'b0;

   // m11_3 = W*in
   wire signed [6:0] m11_3;
   assign m11_3 =7'b0;

   // m11_4 = W*in
   wire signed [6:0] m11_4;
   assign m11_4 =7'b0;

   // m11_5 = W*in
   wire signed [6:0] m11_5;
   assign m11_5 =7'b0;

   // m11_6 = W*in
   wire signed [6:0] m11_6;
   assign m11_6 =7'b0;

   // m11_7 = W*in
   wire signed [6:0] m11_7;
   assign m11_7 =7'b0;

   // m11_8 = W*in
   wire signed [6:0] m11_8;
   assign m11_8 =7'b0;

   // m11_9 = W*in
   wire signed [6:0] m11_9;
   assign m11_9 =7'b0;

   // m11_10 = W*in
   wire signed [6:0] m11_10;
   assign m11_10 =7'b0;

   // m11_11 = W*in
   wire signed [6:0] m11_11;
   assign m11_11 =7'b0;

   // m11_12 = W*in
   wire signed [6:0] m11_12;
   assign m11_12 =7'b0;

   // m11_13 = W*in
   wire signed [6:0] m11_13;
   assign m11_13 =7'b0;

   // m11_14 = W*in
   wire signed [6:0] m11_14;
   assign m11_14 =7'b0;

   // m11_15 = W*in
   wire signed [6:0] m11_15;
   assign m11_15 ={ {2{in11[5]}} , in11[5:1] };

   // m11_16 = W*in
   wire signed [6:0] m11_16;
   assign m11_16 =7'b0;

   // m11_17 = W*in
   wire signed [6:0] m11_17;
   assign m11_17 =7'b0;

   // m11_18 = W*in
   wire signed [6:0] m11_18;
   assign m11_18 =7'b0;

   // m11_19 = W*in
   wire signed [6:0] m11_19;
   assign m11_19 =7'b0;

   // m11_20 = W*in
   wire signed [6:0] m11_20;
   assign m11_20 =7'b0;

   // m11_21 = W*in
   wire signed [6:0] m11_21;
   assign m11_21 =7'b0;

   // m11_22 = W*in
   wire signed [6:0] m11_22;
   assign m11_22 =7'b0;

   // m11_23 = W*in
   wire signed [6:0] m11_23;
   assign m11_23 =7'b0;

   // m11_24 = W*in
   wire signed [6:0] m11_24;
   assign m11_24 =7'b0;

   // m11_25 = W*in
   wire signed [6:0] m11_25;
   assign m11_25 =7'b0;

   // m11_26 = W*in
   wire signed [6:0] m11_26;
   assign m11_26 =7'b0;

   // m11_27 = W*in
   wire signed [6:0] m11_27;
   assign m11_27 =7'b0;

   // m12_1 = W*in
   wire signed [6:0] m12_1;
   assign m12_1 =7'b0;

   // m12_2 = W*in
   wire signed [6:0] m12_2;
   assign m12_2 =7'b0;

   // m12_3 = W*in
   wire signed [6:0] m12_3;
   assign m12_3 =7'b0;

   // m12_4 = W*in
   wire signed [6:0] m12_4;
   assign m12_4 =7'b0;

   // m12_5 = W*in
   wire signed [6:0] m12_5;
   assign m12_5 =7'b0;

   // m12_6 = W*in
   wire signed [6:0] m12_6;
   assign m12_6 =7'b0;

   // m12_7 = W*in
   wire signed [6:0] m12_7;
   assign m12_7 =7'b0;

   // m12_8 = W*in
   wire signed [6:0] m12_8;
   assign m12_8 =7'b0;

   // m12_9 = W*in
   wire signed [6:0] m12_9;
   wire signed [7:0] tm12_9;
   assign tm12_9[0:0] = in12[0:0];
   assign tm12_9[7:1] = { {1{in12[5]}} , in12[5:0] } + { {2{in12[5]}} , in12[5:1] };
   assign m12_9 ={ {1{tm12_9[7]}} , tm12_9[7:2] };

   // m12_10 = W*in
   wire signed [6:0] m12_10;
   assign m12_10 =7'b0;

   // m12_11 = W*in
   wire signed [6:0] m12_11;
   assign m12_11 =7'b0;

   // m12_12 = W*in
   wire signed [6:0] m12_12;
   assign m12_12 =7'b0;

   // m12_13 = W*in
   wire signed [6:0] m12_13;
   assign m12_13 =7'b0;

   // m12_14 = W*in
   wire signed [6:0] m12_14;
   assign m12_14 =7'b0;

   // m12_15 = W*in
   wire signed [6:0] m12_15;
   assign m12_15 =7'b0;

   // m12_16 = W*in
   wire signed [6:0] m12_16;
   assign m12_16 =7'b0;

   // m12_17 = W*in
   wire signed [6:0] m12_17;
   assign m12_17 =7'b0;

   // m12_18 = W*in
   wire signed [6:0] m12_18;
   assign m12_18 =7'b0;

   // m12_19 = W*in
   wire signed [6:0] m12_19;
   assign m12_19 =7'b0;

   // m12_20 = W*in
   wire signed [6:0] m12_20;
   assign m12_20 =7'b0;

   // m12_21 = W*in
   wire signed [6:0] m12_21;
   assign m12_21 ={ {2{in12[5]}} , in12[5:1] };

   // m12_22 = W*in
   wire signed [6:0] m12_22;
   assign m12_22 =7'b0;

   // m12_23 = W*in
   wire signed [6:0] m12_23;
   assign m12_23 =7'b0;

   // m12_24 = W*in
   wire signed [6:0] m12_24;
   assign m12_24 =7'b0;

   // m12_25 = W*in
   wire signed [6:0] m12_25;
   assign m12_25 =7'b0;

   // m12_26 = W*in
   wire signed [6:0] m12_26;
   assign m12_26 =7'b0;

   // m12_27 = W*in
   wire signed [6:0] m12_27;
   assign m12_27 =7'b0;

   // m13_1 = W*in
   wire signed [6:0] m13_1;
   assign m13_1 =7'b0;

   // m13_2 = W*in
   wire signed [6:0] m13_2;
   assign m13_2 =7'b0;

   // m13_3 = W*in
   wire signed [6:0] m13_3;
   assign m13_3 =7'b0;

   // m13_4 = W*in
   wire signed [6:0] m13_4;
   assign m13_4 =7'b0;

   // m13_5 = W*in
   wire signed [6:0] m13_5;
   assign m13_5 =7'b0;

   // m13_6 = W*in
   wire signed [6:0] m13_6;
   assign m13_6 =7'b0;

   // m13_7 = W*in
   wire signed [6:0] m13_7;
   assign m13_7 =7'b0;

   // m13_8 = W*in
   wire signed [6:0] m13_8;
   assign m13_8 =7'b0;

   // m13_9 = W*in
   wire signed [6:0] m13_9;
   assign m13_9 =7'b0;

   // m13_10 = W*in
   wire signed [6:0] m13_10;
   assign m13_10 =7'b0;

   // m13_11 = W*in
   wire signed [6:0] m13_11;
   assign m13_11 =7'b0;

   // m13_12 = W*in
   wire signed [6:0] m13_12;
   assign m13_12 =7'b0;

   // m13_13 = W*in
   wire signed [6:0] m13_13;
   assign m13_13 =7'b0;

   // m13_14 = W*in
   wire signed [6:0] m13_14;
   assign m13_14 =7'b0;

   // m13_15 = W*in
   wire signed [6:0] m13_15;
   assign m13_15 =7'b0;

   // m13_16 = W*in
   wire signed [6:0] m13_16;
   assign m13_16 =7'b0;

   // m13_17 = W*in
   wire signed [6:0] m13_17;
   assign m13_17 =7'b0;

   // m13_18 = W*in
   wire signed [6:0] m13_18;
   assign m13_18 =7'b0;

   // m13_19 = W*in
   wire signed [6:0] m13_19;
   assign m13_19 =7'b0;

   // m13_20 = W*in
   wire signed [6:0] m13_20;
   assign m13_20 =7'b0;

   // m13_21 = W*in
   wire signed [6:0] m13_21;
   assign m13_21 =7'b0;

   // m13_22 = W*in
   wire signed [6:0] m13_22;
   assign m13_22 =7'b0;

   // m13_23 = W*in
   wire signed [6:0] m13_23;
   assign m13_23 =7'b0;

   // m13_24 = W*in
   wire signed [6:0] m13_24;
   assign m13_24 ={ {2{in13[5]}} , in13[5:1] };

   // m13_25 = W*in
   wire signed [6:0] m13_25;
   assign m13_25 =7'b0;

   // m13_26 = W*in
   wire signed [6:0] m13_26;
   assign m13_26 =7'b0;

   // m13_27 = W*in
   wire signed [6:0] m13_27;
   assign m13_27 =7'b0;

   // m14_1 = W*in
   wire signed [6:0] m14_1;
   assign m14_1 =7'b0;

   // m14_2 = W*in
   wire signed [6:0] m14_2;
   assign m14_2 =7'b0;

   // m14_3 = W*in
   wire signed [6:0] m14_3;
   assign m14_3 =7'b0;

   // m14_4 = W*in
   wire signed [6:0] m14_4;
   assign m14_4 =7'b0;

   // m14_5 = W*in
   wire signed [6:0] m14_5;
   assign m14_5 =7'b0;

   // m14_6 = W*in
   wire signed [6:0] m14_6;
   assign m14_6 =7'b0;

   // m14_7 = W*in
   wire signed [6:0] m14_7;
   assign m14_7 =7'b0;

   // m14_8 = W*in
   wire signed [6:0] m14_8;
   assign m14_8 =7'b0;

   // m14_9 = W*in
   wire signed [6:0] m14_9;
   assign m14_9 =7'b0;

   // m14_10 = W*in
   wire signed [6:0] m14_10;
   assign m14_10 =7'b0;

   // m14_11 = W*in
   wire signed [6:0] m14_11;
   assign m14_11 =7'b0;

   // m14_12 = W*in
   wire signed [6:0] m14_12;
   assign m14_12 =7'b0;

   // m14_13 = W*in
   wire signed [6:0] m14_13;
   assign m14_13 =7'b0;

   // m14_14 = W*in
   wire signed [6:0] m14_14;
   assign m14_14 =7'b0;

   // m14_15 = W*in
   wire signed [6:0] m14_15;
   assign m14_15 =7'b0;

   // m14_16 = W*in
   wire signed [6:0] m14_16;
   assign m14_16 =7'b0;

   // m14_17 = W*in
   wire signed [6:0] m14_17;
   assign m14_17 =7'b0;

   // m14_18 = W*in
   wire signed [6:0] m14_18;
   assign m14_18 =7'b0;

   // m14_19 = W*in
   wire signed [6:0] m14_19;
   assign m14_19 ={ {2{neg14[5]}} , neg14[5:1] };

   // m14_20 = W*in
   wire signed [6:0] m14_20;
   assign m14_20 =7'b0;

   // m14_21 = W*in
   wire signed [6:0] m14_21;
   assign m14_21 =7'b0;

   // m14_22 = W*in
   wire signed [6:0] m14_22;
   assign m14_22 =7'b0;

   // m14_23 = W*in
   wire signed [6:0] m14_23;
   assign m14_23 ={ {2{in14[5]}} , in14[5:1] };

   // m14_24 = W*in
   wire signed [6:0] m14_24;
   assign m14_24 =7'b0;

   // m14_25 = W*in
   wire signed [6:0] m14_25;
   assign m14_25 =7'b0;

   // m14_26 = W*in
   wire signed [6:0] m14_26;
   assign m14_26 =7'b0;

   // m14_27 = W*in
   wire signed [6:0] m14_27;
   assign m14_27 =7'b0;

   // m15_1 = W*in
   wire signed [6:0] m15_1;
   assign m15_1 =7'b0;

   // m15_2 = W*in
   wire signed [6:0] m15_2;
   assign m15_2 =7'b0;

   // m15_3 = W*in
   wire signed [6:0] m15_3;
   assign m15_3 =7'b0;

   // m15_4 = W*in
   wire signed [6:0] m15_4;
   assign m15_4 =7'b0;

   // m15_5 = W*in
   wire signed [6:0] m15_5;
   assign m15_5 =7'b0;

   // m15_6 = W*in
   wire signed [6:0] m15_6;
   assign m15_6 =7'b0;

   // m15_7 = W*in
   wire signed [6:0] m15_7;
   assign m15_7 =7'b0;

   // m15_8 = W*in
   wire signed [6:0] m15_8;
   assign m15_8 =7'b0;

   // m15_9 = W*in
   wire signed [6:0] m15_9;
   assign m15_9 =7'b0;

   // m15_10 = W*in
   wire signed [6:0] m15_10;
   assign m15_10 =7'b0;

   // m15_11 = W*in
   wire signed [6:0] m15_11;
   assign m15_11 =7'b0;

   // m15_12 = W*in
   wire signed [6:0] m15_12;
   assign m15_12 =7'b0;

   // m15_13 = W*in
   wire signed [6:0] m15_13;
   assign m15_13 ={ {2{in15[5]}} , in15[5:1] };

   // m15_14 = W*in
   wire signed [6:0] m15_14;
   assign m15_14 =7'b0;

   // m15_15 = W*in
   wire signed [6:0] m15_15;
   assign m15_15 =7'b0;

   // m15_16 = W*in
   wire signed [6:0] m15_16;
   assign m15_16 =7'b0;

   // m15_17 = W*in
   wire signed [6:0] m15_17;
   assign m15_17 =7'b0;

   // m15_18 = W*in
   wire signed [6:0] m15_18;
   assign m15_18 =7'b0;

   // m15_19 = W*in
   wire signed [6:0] m15_19;
   assign m15_19 =7'b0;

   // m15_20 = W*in
   wire signed [6:0] m15_20;
   assign m15_20 =7'b0;

   // m15_21 = W*in
   wire signed [6:0] m15_21;
   assign m15_21 =7'b0;

   // m15_22 = W*in
   wire signed [6:0] m15_22;
   assign m15_22 =7'b0;

   // m15_23 = W*in
   wire signed [6:0] m15_23;
   assign m15_23 =7'b0;

   // m15_24 = W*in
   wire signed [6:0] m15_24;
   assign m15_24 =7'b0;

   // m15_25 = W*in
   wire signed [6:0] m15_25;
   assign m15_25 =7'b0;

   // m15_26 = W*in
   wire signed [6:0] m15_26;
   assign m15_26 =7'b0;

   // m15_27 = W*in
   wire signed [6:0] m15_27;
   assign m15_27 =7'b0;

   // m16_1 = W*in
   wire signed [6:0] m16_1;
   assign m16_1 =7'b0;

   // m16_2 = W*in
   wire signed [6:0] m16_2;
   assign m16_2 =7'b0;

   // m16_3 = W*in
   wire signed [6:0] m16_3;
   assign m16_3 =7'b0;

   // m16_4 = W*in
   wire signed [6:0] m16_4;
   assign m16_4 =7'b0;

   // m16_5 = W*in
   wire signed [6:0] m16_5;
   assign m16_5 =7'b0;

   // m16_6 = W*in
   wire signed [6:0] m16_6;
   assign m16_6 =7'b0;

   // m16_7 = W*in
   wire signed [6:0] m16_7;
   assign m16_7 =7'b0;

   // m16_8 = W*in
   wire signed [6:0] m16_8;
   assign m16_8 =7'b0;

   // m16_9 = W*in
   wire signed [6:0] m16_9;
   assign m16_9 ={ {2{in16[5]}} , in16[5:1] };

   // m16_10 = W*in
   wire signed [6:0] m16_10;
   assign m16_10 =7'b0;

   // m16_11 = W*in
   wire signed [6:0] m16_11;
   assign m16_11 =7'b0;

   // m16_12 = W*in
   wire signed [6:0] m16_12;
   assign m16_12 =7'b0;

   // m16_13 = W*in
   wire signed [6:0] m16_13;
   assign m16_13 =7'b0;

   // m16_14 = W*in
   wire signed [6:0] m16_14;
   assign m16_14 =7'b0;

   // m16_15 = W*in
   wire signed [6:0] m16_15;
   assign m16_15 =7'b0;

   // m16_16 = W*in
   wire signed [6:0] m16_16;
   assign m16_16 =7'b0;

   // m16_17 = W*in
   wire signed [6:0] m16_17;
   assign m16_17 =7'b0;

   // m16_18 = W*in
   wire signed [6:0] m16_18;
   assign m16_18 =7'b0;

   // m16_19 = W*in
   wire signed [6:0] m16_19;
   assign m16_19 =7'b0;

   // m16_20 = W*in
   wire signed [6:0] m16_20;
   assign m16_20 =7'b0;

   // m16_21 = W*in
   wire signed [6:0] m16_21;
   assign m16_21 =7'b0;

   // m16_22 = W*in
   wire signed [6:0] m16_22;
   assign m16_22 =7'b0;

   // m16_23 = W*in
   wire signed [6:0] m16_23;
   assign m16_23 =7'b0;

   // m16_24 = W*in
   wire signed [6:0] m16_24;
   assign m16_24 =7'b0;

   // m16_25 = W*in
   wire signed [6:0] m16_25;
   assign m16_25 =7'b0;

   // m16_26 = W*in
   wire signed [6:0] m16_26;
   assign m16_26 =7'b0;

   // m16_27 = W*in
   wire signed [6:0] m16_27;
   assign m16_27 =7'b0;

   // m17_1 = W*in
   wire signed [6:0] m17_1;
   assign m17_1 =7'b0;

   // m17_2 = W*in
   wire signed [6:0] m17_2;
   assign m17_2 =7'b0;

   // m17_3 = W*in
   wire signed [6:0] m17_3;
   assign m17_3 =7'b0;

   // m17_4 = W*in
   wire signed [6:0] m17_4;
   assign m17_4 =7'b0;

   // m17_5 = W*in
   wire signed [6:0] m17_5;
   assign m17_5 =7'b0;

   // m17_6 = W*in
   wire signed [6:0] m17_6;
   assign m17_6 =7'b0;

   // m17_7 = W*in
   wire signed [6:0] m17_7;
   assign m17_7 =7'b0;

   // m17_8 = W*in
   wire signed [6:0] m17_8;
   assign m17_8 =7'b0;

   // m17_9 = W*in
   wire signed [6:0] m17_9;
   assign m17_9 =7'b0;

   // m17_10 = W*in
   wire signed [6:0] m17_10;
   assign m17_10 =7'b0;

   // m17_11 = W*in
   wire signed [6:0] m17_11;
   assign m17_11 =7'b0;

   // m17_12 = W*in
   wire signed [6:0] m17_12;
   assign m17_12 =7'b0;

   // m17_13 = W*in
   wire signed [6:0] m17_13;
   assign m17_13 =7'b0;

   // m17_14 = W*in
   wire signed [6:0] m17_14;
   assign m17_14 =7'b0;

   // m17_15 = W*in
   wire signed [6:0] m17_15;
   assign m17_15 =7'b0;

   // m17_16 = W*in
   wire signed [6:0] m17_16;
   assign m17_16 =7'b0;

   // m17_17 = W*in
   wire signed [6:0] m17_17;
   assign m17_17 =7'b0;

   // m17_18 = W*in
   wire signed [6:0] m17_18;
   assign m17_18 =7'b0;

   // m17_19 = W*in
   wire signed [6:0] m17_19;
   assign m17_19 =7'b0;

   // m17_20 = W*in
   wire signed [6:0] m17_20;
   assign m17_20 =7'b0;

   // m17_21 = W*in
   wire signed [6:0] m17_21;
   assign m17_21 =7'b0;

   // m17_22 = W*in
   wire signed [6:0] m17_22;
   assign m17_22 =7'b0;

   // m17_23 = W*in
   wire signed [6:0] m17_23;
   assign m17_23 =7'b0;

   // m17_24 = W*in
   wire signed [6:0] m17_24;
   assign m17_24 =7'b0;

   // m17_25 = W*in
   wire signed [6:0] m17_25;
   assign m17_25 ={ {1{in17[5]}} , in17[5:0] };

   // m17_26 = W*in
   wire signed [6:0] m17_26;
   assign m17_26 =7'b0;

   // m17_27 = W*in
   wire signed [6:0] m17_27;
   assign m17_27 =7'b0;

   // m18_1 = W*in
   wire signed [6:0] m18_1;
   assign m18_1 =7'b0;

   // m18_2 = W*in
   wire signed [6:0] m18_2;
   assign m18_2 =7'b0;

   // m18_3 = W*in
   wire signed [6:0] m18_3;
   assign m18_3 =7'b0;

   // m18_4 = W*in
   wire signed [6:0] m18_4;
   assign m18_4 =7'b0;

   // m18_5 = W*in
   wire signed [6:0] m18_5;
   assign m18_5 =7'b0;

   // m18_6 = W*in
   wire signed [6:0] m18_6;
   assign m18_6 =7'b0;

   // m18_7 = W*in
   wire signed [6:0] m18_7;
   assign m18_7 =7'b0;

   // m18_8 = W*in
   wire signed [6:0] m18_8;
   assign m18_8 =7'b0;

   // m18_9 = W*in
   wire signed [6:0] m18_9;
   assign m18_9 =7'b0;

   // m18_10 = W*in
   wire signed [6:0] m18_10;
   assign m18_10 =7'b0;

   // m18_11 = W*in
   wire signed [6:0] m18_11;
   assign m18_11 =7'b0;

   // m18_12 = W*in
   wire signed [6:0] m18_12;
   assign m18_12 =7'b0;

   // m18_13 = W*in
   wire signed [6:0] m18_13;
   assign m18_13 =7'b0;

   // m18_14 = W*in
   wire signed [6:0] m18_14;
   assign m18_14 =7'b0;

   // m18_15 = W*in
   wire signed [6:0] m18_15;
   assign m18_15 =7'b0;

   // m18_16 = W*in
   wire signed [6:0] m18_16;
   assign m18_16 =7'b0;

   // m18_17 = W*in
   wire signed [6:0] m18_17;
   assign m18_17 =7'b0;

   // m18_18 = W*in
   wire signed [6:0] m18_18;
   assign m18_18 =7'b0;

   // m18_19 = W*in
   wire signed [6:0] m18_19;
   assign m18_19 =7'b0;

   // m18_20 = W*in
   wire signed [6:0] m18_20;
   assign m18_20 =7'b0;

   // m18_21 = W*in
   wire signed [6:0] m18_21;
   assign m18_21 ={ {1{in18[5]}} , in18[5:0] };

   // m18_22 = W*in
   wire signed [6:0] m18_22;
   assign m18_22 =7'b0;

   // m18_23 = W*in
   wire signed [6:0] m18_23;
   assign m18_23 =7'b0;

   // m18_24 = W*in
   wire signed [6:0] m18_24;
   assign m18_24 =7'b0;

   // m18_25 = W*in
   wire signed [6:0] m18_25;
   assign m18_25 =7'b0;

   // m18_26 = W*in
   wire signed [6:0] m18_26;
   assign m18_26 =7'b0;

   // m18_27 = W*in
   wire signed [6:0] m18_27;
   assign m18_27 =7'b0;

   // m19_1 = W*in
   wire signed [6:0] m19_1;
   assign m19_1 =7'b0;

   // m19_2 = W*in
   wire signed [6:0] m19_2;
   assign m19_2 =7'b0;

   // m19_3 = W*in
   wire signed [6:0] m19_3;
   assign m19_3 =7'b0;

   // m19_4 = W*in
   wire signed [6:0] m19_4;
   assign m19_4 =7'b0;

   // m19_5 = W*in
   wire signed [6:0] m19_5;
   assign m19_5 =7'b0;

   // m19_6 = W*in
   wire signed [6:0] m19_6;
   assign m19_6 =7'b0;

   // m19_7 = W*in
   wire signed [6:0] m19_7;
   assign m19_7 =7'b0;

   // m19_8 = W*in
   wire signed [6:0] m19_8;
   assign m19_8 =7'b0;

   // m19_9 = W*in
   wire signed [6:0] m19_9;
   assign m19_9 ={ {2{in19[5]}} , in19[5:1] };

   // m19_10 = W*in
   wire signed [6:0] m19_10;
   assign m19_10 =7'b0;

   // m19_11 = W*in
   wire signed [6:0] m19_11;
   assign m19_11 =7'b0;

   // m19_12 = W*in
   wire signed [6:0] m19_12;
   assign m19_12 =7'b0;

   // m19_13 = W*in
   wire signed [6:0] m19_13;
   assign m19_13 =7'b0;

   // m19_14 = W*in
   wire signed [6:0] m19_14;
   assign m19_14 =7'b0;

   // m19_15 = W*in
   wire signed [6:0] m19_15;
   assign m19_15 =7'b0;

   // m19_16 = W*in
   wire signed [6:0] m19_16;
   assign m19_16 =7'b0;

   // m19_17 = W*in
   wire signed [6:0] m19_17;
   assign m19_17 =7'b0;

   // m19_18 = W*in
   wire signed [6:0] m19_18;
   assign m19_18 =7'b0;

   // m19_19 = W*in
   wire signed [6:0] m19_19;
   assign m19_19 =7'b0;

   // m19_20 = W*in
   wire signed [6:0] m19_20;
   assign m19_20 =7'b0;

   // m19_21 = W*in
   wire signed [6:0] m19_21;
   assign m19_21 =7'b0;

   // m19_22 = W*in
   wire signed [6:0] m19_22;
   assign m19_22 =7'b0;

   // m19_23 = W*in
   wire signed [6:0] m19_23;
   assign m19_23 =7'b0;

   // m19_24 = W*in
   wire signed [6:0] m19_24;
   assign m19_24 =7'b0;

   // m19_25 = W*in
   wire signed [6:0] m19_25;
   assign m19_25 =7'b0;

   // m19_26 = W*in
   wire signed [6:0] m19_26;
   assign m19_26 =7'b0;

   // m19_27 = W*in
   wire signed [6:0] m19_27;
   assign m19_27 =7'b0;

   // m20_1 = W*in
   wire signed [6:0] m20_1;
   assign m20_1 =7'b0;

   // m20_2 = W*in
   wire signed [6:0] m20_2;
   assign m20_2 =7'b0;

   // m20_3 = W*in
   wire signed [6:0] m20_3;
   assign m20_3 =7'b0;

   // m20_4 = W*in
   wire signed [6:0] m20_4;
   assign m20_4 ={ {1{in20[5]}} , in20[5:0] };

   // m20_5 = W*in
   wire signed [6:0] m20_5;
   assign m20_5 =7'b0;

   // m20_6 = W*in
   wire signed [6:0] m20_6;
   assign m20_6 ={ {1{in20[5]}} , in20[5:0] };

   // m20_7 = W*in
   wire signed [6:0] m20_7;
   assign m20_7 =7'b0;

   // m20_8 = W*in
   wire signed [6:0] m20_8;
   assign m20_8 =7'b0;

   // m20_9 = W*in
   wire signed [6:0] m20_9;
   assign m20_9 =7'b0;

   // m20_10 = W*in
   wire signed [6:0] m20_10;
   assign m20_10 =7'b0;

   // m20_11 = W*in
   wire signed [6:0] m20_11;
   assign m20_11 =7'b0;

   // m20_12 = W*in
   wire signed [6:0] m20_12;
   assign m20_12 =7'b0;

   // m20_13 = W*in
   wire signed [6:0] m20_13;
   assign m20_13 =7'b0;

   // m20_14 = W*in
   wire signed [6:0] m20_14;
   assign m20_14 =7'b0;

   // m20_15 = W*in
   wire signed [6:0] m20_15;
   assign m20_15 =7'b0;

   // m20_16 = W*in
   wire signed [6:0] m20_16;
   assign m20_16 =7'b0;

   // m20_17 = W*in
   wire signed [6:0] m20_17;
   assign m20_17 =7'b0;

   // m20_18 = W*in
   wire signed [6:0] m20_18;
   assign m20_18 =7'b0;

   // m20_19 = W*in
   wire signed [6:0] m20_19;
   assign m20_19 =7'b0;

   // m20_20 = W*in
   wire signed [6:0] m20_20;
   assign m20_20 =7'b0;

   // m20_21 = W*in
   wire signed [6:0] m20_21;
   assign m20_21 =7'b0;

   // m20_22 = W*in
   wire signed [6:0] m20_22;
   assign m20_22 =7'b0;

   // m20_23 = W*in
   wire signed [6:0] m20_23;
   assign m20_23 =7'b0;

   // m20_24 = W*in
   wire signed [6:0] m20_24;
   assign m20_24 =7'b0;

   // m20_25 = W*in
   wire signed [6:0] m20_25;
   assign m20_25 =7'b0;

   // m20_26 = W*in
   wire signed [6:0] m20_26;
   assign m20_26 =7'b0;

   // m20_27 = W*in
   wire signed [6:0] m20_27;
   assign m20_27 =7'b0;

   // m21_1 = W*in
   wire signed [6:0] m21_1;
   assign m21_1 =7'b0;

   // m21_2 = W*in
   wire signed [6:0] m21_2;
   assign m21_2 =7'b0;

   // m21_3 = W*in
   wire signed [6:0] m21_3;
   assign m21_3 =7'b0;

   // m21_4 = W*in
   wire signed [6:0] m21_4;
   assign m21_4 =7'b0;

   // m21_5 = W*in
   wire signed [6:0] m21_5;
   assign m21_5 =7'b0;

   // m21_6 = W*in
   wire signed [6:0] m21_6;
   assign m21_6 =7'b0;

   // m21_7 = W*in
   wire signed [6:0] m21_7;
   assign m21_7 =7'b0;

   // m21_8 = W*in
   wire signed [6:0] m21_8;
   assign m21_8 =7'b0;

   // m21_9 = W*in
   wire signed [6:0] m21_9;
   assign m21_9 ={ {1{in21[5]}} , in21[5:0] };

   // m21_10 = W*in
   wire signed [6:0] m21_10;
   assign m21_10 =7'b0;

   // m21_11 = W*in
   wire signed [6:0] m21_11;
   assign m21_11 =7'b0;

   // m21_12 = W*in
   wire signed [6:0] m21_12;
   assign m21_12 =7'b0;

   // m21_13 = W*in
   wire signed [6:0] m21_13;
   assign m21_13 =7'b0;

   // m21_14 = W*in
   wire signed [6:0] m21_14;
   assign m21_14 =7'b0;

   // m21_15 = W*in
   wire signed [6:0] m21_15;
   assign m21_15 =7'b0;

   // m21_16 = W*in
   wire signed [6:0] m21_16;
   assign m21_16 =7'b0;

   // m21_17 = W*in
   wire signed [6:0] m21_17;
   assign m21_17 =7'b0;

   // m21_18 = W*in
   wire signed [6:0] m21_18;
   assign m21_18 =7'b0;

   // m21_19 = W*in
   wire signed [6:0] m21_19;
   assign m21_19 =7'b0;

   // m21_20 = W*in
   wire signed [6:0] m21_20;
   assign m21_20 =7'b0;

   // m21_21 = W*in
   wire signed [6:0] m21_21;
   assign m21_21 =7'b0;

   // m21_22 = W*in
   wire signed [6:0] m21_22;
   assign m21_22 =7'b0;

   // m21_23 = W*in
   wire signed [6:0] m21_23;
   assign m21_23 =7'b0;

   // m21_24 = W*in
   wire signed [6:0] m21_24;
   assign m21_24 =7'b0;

   // m21_25 = W*in
   wire signed [6:0] m21_25;
   assign m21_25 =7'b0;

   // m21_26 = W*in
   wire signed [6:0] m21_26;
   assign m21_26 =7'b0;

   // m21_27 = W*in
   wire signed [6:0] m21_27;
   assign m21_27 =7'b0;

   // m22_1 = W*in
   wire signed [6:0] m22_1;
   assign m22_1 =7'b0;

   // m22_2 = W*in
   wire signed [6:0] m22_2;
   assign m22_2 =7'b0;

   // m22_3 = W*in
   wire signed [6:0] m22_3;
   assign m22_3 =7'b0;

   // m22_4 = W*in
   wire signed [6:0] m22_4;
   assign m22_4 =7'b0;

   // m22_5 = W*in
   wire signed [6:0] m22_5;
   assign m22_5 =7'b0;

   // m22_6 = W*in
   wire signed [6:0] m22_6;
   assign m22_6 =7'b0;

   // m22_7 = W*in
   wire signed [6:0] m22_7;
   assign m22_7 =7'b0;

   // m22_8 = W*in
   wire signed [6:0] m22_8;
   assign m22_8 =7'b0;

   // m22_9 = W*in
   wire signed [6:0] m22_9;
   assign m22_9 =7'b0;

   // m22_10 = W*in
   wire signed [6:0] m22_10;
   assign m22_10 =7'b0;

   // m22_11 = W*in
   wire signed [6:0] m22_11;
   assign m22_11 =7'b0;

   // m22_12 = W*in
   wire signed [6:0] m22_12;
   assign m22_12 =7'b0;

   // m22_13 = W*in
   wire signed [6:0] m22_13;
   assign m22_13 =7'b0;

   // m22_14 = W*in
   wire signed [6:0] m22_14;
   assign m22_14 =7'b0;

   // m22_15 = W*in
   wire signed [6:0] m22_15;
   assign m22_15 =7'b0;

   // m22_16 = W*in
   wire signed [6:0] m22_16;
   assign m22_16 =7'b0;

   // m22_17 = W*in
   wire signed [6:0] m22_17;
   assign m22_17 ={ {2{in22[5]}} , in22[5:1] };

   // m22_18 = W*in
   wire signed [6:0] m22_18;
   assign m22_18 =7'b0;

   // m22_19 = W*in
   wire signed [6:0] m22_19;
   assign m22_19 =7'b0;

   // m22_20 = W*in
   wire signed [6:0] m22_20;
   assign m22_20 =7'b0;

   // m22_21 = W*in
   wire signed [6:0] m22_21;
   assign m22_21 =7'b0;

   // m22_22 = W*in
   wire signed [6:0] m22_22;
   assign m22_22 =7'b0;

   // m22_23 = W*in
   wire signed [6:0] m22_23;
   assign m22_23 =7'b0;

   // m22_24 = W*in
   wire signed [6:0] m22_24;
   assign m22_24 =7'b0;

   // m22_25 = W*in
   wire signed [6:0] m22_25;
   assign m22_25 =7'b0;

   // m22_26 = W*in
   wire signed [6:0] m22_26;
   assign m22_26 =7'b0;

   // m22_27 = W*in
   wire signed [6:0] m22_27;
   assign m22_27 =7'b0;

   // m23_1 = W*in
   wire signed [6:0] m23_1;
   assign m23_1 =7'b0;

   // m23_2 = W*in
   wire signed [6:0] m23_2;
   assign m23_2 =7'b0;

   // m23_3 = W*in
   wire signed [6:0] m23_3;
   assign m23_3 =7'b0;

   // m23_4 = W*in
   wire signed [6:0] m23_4;
   assign m23_4 =7'b0;

   // m23_5 = W*in
   wire signed [6:0] m23_5;
   assign m23_5 =7'b0;

   // m23_6 = W*in
   wire signed [6:0] m23_6;
   assign m23_6 =7'b0;

   // m23_7 = W*in
   wire signed [6:0] m23_7;
   assign m23_7 =7'b0;

   // m23_8 = W*in
   wire signed [6:0] m23_8;
   assign m23_8 =7'b0;

   // m23_9 = W*in
   wire signed [6:0] m23_9;
   assign m23_9 =7'b0;

   // m23_10 = W*in
   wire signed [6:0] m23_10;
   assign m23_10 =7'b0;

   // m23_11 = W*in
   wire signed [6:0] m23_11;
   assign m23_11 =7'b0;

   // m23_12 = W*in
   wire signed [6:0] m23_12;
   assign m23_12 =7'b0;

   // m23_13 = W*in
   wire signed [6:0] m23_13;
   wire signed [7:0] tm23_13;
   assign tm23_13[0:0] = in23[0:0];
   assign tm23_13[7:1] = { {1{in23[5]}} , in23[5:0] } + { {2{in23[5]}} , in23[5:1] };
   assign m23_13 ={ {1{tm23_13[7]}} , tm23_13[7:2] };

   // m23_14 = W*in
   wire signed [6:0] m23_14;
   assign m23_14 =7'b0;

   // m23_15 = W*in
   wire signed [6:0] m23_15;
   assign m23_15 =7'b0;

   // m23_16 = W*in
   wire signed [6:0] m23_16;
   assign m23_16 =7'b0;

   // m23_17 = W*in
   wire signed [6:0] m23_17;
   assign m23_17 =7'b0;

   // m23_18 = W*in
   wire signed [6:0] m23_18;
   assign m23_18 =7'b0;

   // m23_19 = W*in
   wire signed [6:0] m23_19;
   assign m23_19 =7'b0;

   // m23_20 = W*in
   wire signed [6:0] m23_20;
   assign m23_20 =7'b0;

   // m23_21 = W*in
   wire signed [6:0] m23_21;
   assign m23_21 =7'b0;

   // m23_22 = W*in
   wire signed [6:0] m23_22;
   assign m23_22 =7'b0;

   // m23_23 = W*in
   wire signed [6:0] m23_23;
   assign m23_23 =7'b0;

   // m23_24 = W*in
   wire signed [6:0] m23_24;
   assign m23_24 =7'b0;

   // m23_25 = W*in
   wire signed [6:0] m23_25;
   assign m23_25 =7'b0;

   // m23_26 = W*in
   wire signed [6:0] m23_26;
   assign m23_26 =7'b0;

   // m23_27 = W*in
   wire signed [6:0] m23_27;
   assign m23_27 =7'b0;

   // m24_1 = W*in
   wire signed [6:0] m24_1;
   assign m24_1 =7'b0;

   // m24_2 = W*in
   wire signed [6:0] m24_2;
   assign m24_2 =7'b0;

   // m24_3 = W*in
   wire signed [6:0] m24_3;
   assign m24_3 =7'b0;

   // m24_4 = W*in
   wire signed [6:0] m24_4;
   assign m24_4 =7'b0;

   // m24_5 = W*in
   wire signed [6:0] m24_5;
   assign m24_5 =7'b0;

   // m24_6 = W*in
   wire signed [6:0] m24_6;
   assign m24_6 =7'b0;

   // m24_7 = W*in
   wire signed [6:0] m24_7;
   assign m24_7 =7'b0;

   // m24_8 = W*in
   wire signed [6:0] m24_8;
   assign m24_8 =7'b0;

   // m24_9 = W*in
   wire signed [6:0] m24_9;
   assign m24_9 =7'b0;

   // m24_10 = W*in
   wire signed [6:0] m24_10;
   assign m24_10 =7'b0;

   // m24_11 = W*in
   wire signed [6:0] m24_11;
   assign m24_11 =7'b0;

   // m24_12 = W*in
   wire signed [6:0] m24_12;
   assign m24_12 =7'b0;

   // m24_13 = W*in
   wire signed [6:0] m24_13;
   assign m24_13 ={ {1{in24[5]}} , in24[5:0] };

   // m24_14 = W*in
   wire signed [6:0] m24_14;
   assign m24_14 =7'b0;

   // m24_15 = W*in
   wire signed [6:0] m24_15;
   assign m24_15 =7'b0;

   // m24_16 = W*in
   wire signed [6:0] m24_16;
   assign m24_16 =7'b0;

   // m24_17 = W*in
   wire signed [6:0] m24_17;
   assign m24_17 =7'b0;

   // m24_18 = W*in
   wire signed [6:0] m24_18;
   assign m24_18 =7'b0;

   // m24_19 = W*in
   wire signed [6:0] m24_19;
   assign m24_19 =7'b0;

   // m24_20 = W*in
   wire signed [6:0] m24_20;
   assign m24_20 =7'b0;

   // m24_21 = W*in
   wire signed [6:0] m24_21;
   assign m24_21 =7'b0;

   // m24_22 = W*in
   wire signed [6:0] m24_22;
   assign m24_22 ={ {2{in24[5]}} , in24[5:1] };

   // m24_23 = W*in
   wire signed [6:0] m24_23;
   assign m24_23 =7'b0;

   // m24_24 = W*in
   wire signed [6:0] m24_24;
   assign m24_24 =7'b0;

   // m24_25 = W*in
   wire signed [6:0] m24_25;
   assign m24_25 =7'b0;

   // m24_26 = W*in
   wire signed [6:0] m24_26;
   assign m24_26 =7'b0;

   // m24_27 = W*in
   wire signed [6:0] m24_27;
   assign m24_27 =7'b0;

   // m25_1 = W*in
   wire signed [6:0] m25_1;
   assign m25_1 =7'b0;

   // m25_2 = W*in
   wire signed [6:0] m25_2;
   assign m25_2 =7'b0;

   // m25_3 = W*in
   wire signed [6:0] m25_3;
   assign m25_3 ={ {2{neg25[5]}} , neg25[5:1] };

   // m25_4 = W*in
   wire signed [6:0] m25_4;
   assign m25_4 =7'b0;

   // m25_5 = W*in
   wire signed [6:0] m25_5;
   assign m25_5 =7'b0;

   // m25_6 = W*in
   wire signed [6:0] m25_6;
   assign m25_6 =7'b0;

   // m25_7 = W*in
   wire signed [6:0] m25_7;
   assign m25_7 ={ {2{neg25[5]}} , neg25[5:1] };

   // m25_8 = W*in
   wire signed [6:0] m25_8;
   assign m25_8 =7'b0;

   // m25_9 = W*in
   wire signed [6:0] m25_9;
   assign m25_9 =7'b0;

   // m25_10 = W*in
   wire signed [6:0] m25_10;
   assign m25_10 =7'b0;

   // m25_11 = W*in
   wire signed [6:0] m25_11;
   assign m25_11 =7'b0;

   // m25_12 = W*in
   wire signed [6:0] m25_12;
   assign m25_12 =7'b0;

   // m25_13 = W*in
   wire signed [6:0] m25_13;
   assign m25_13 =7'b0;

   // m25_14 = W*in
   wire signed [6:0] m25_14;
   assign m25_14 =7'b0;

   // m25_15 = W*in
   wire signed [6:0] m25_15;
   assign m25_15 =7'b0;

   // m25_16 = W*in
   wire signed [6:0] m25_16;
   assign m25_16 =7'b0;

   // m25_17 = W*in
   wire signed [6:0] m25_17;
   assign m25_17 =7'b0;

   // m25_18 = W*in
   wire signed [6:0] m25_18;
   assign m25_18 =7'b0;

   // m25_19 = W*in
   wire signed [6:0] m25_19;
   assign m25_19 =7'b0;

   // m25_20 = W*in
   wire signed [6:0] m25_20;
   assign m25_20 =7'b0;

   // m25_21 = W*in
   wire signed [6:0] m25_21;
   assign m25_21 =7'b0;

   // m25_22 = W*in
   wire signed [6:0] m25_22;
   assign m25_22 =7'b0;

   // m25_23 = W*in
   wire signed [6:0] m25_23;
   assign m25_23 =7'b0;

   // m25_24 = W*in
   wire signed [6:0] m25_24;
   assign m25_24 =7'b0;

   // m25_25 = W*in
   wire signed [6:0] m25_25;
   assign m25_25 =7'b0;

   // m25_26 = W*in
   wire signed [6:0] m25_26;
   assign m25_26 =7'b0;

   // m25_27 = W*in
   wire signed [6:0] m25_27;
   assign m25_27 =7'b0;

   // m26_1 = W*in
   wire signed [6:0] m26_1;
   assign m26_1 =7'b0;

   // m26_2 = W*in
   wire signed [6:0] m26_2;
   assign m26_2 =7'b0;

   // m26_3 = W*in
   wire signed [6:0] m26_3;
   assign m26_3 =7'b0;

   // m26_4 = W*in
   wire signed [6:0] m26_4;
   assign m26_4 =7'b0;

   // m26_5 = W*in
   wire signed [6:0] m26_5;
   assign m26_5 =7'b0;

   // m26_6 = W*in
   wire signed [6:0] m26_6;
   assign m26_6 =7'b0;

   // m26_7 = W*in
   wire signed [6:0] m26_7;
   assign m26_7 =7'b0;

   // m26_8 = W*in
   wire signed [6:0] m26_8;
   assign m26_8 =7'b0;

   // m26_9 = W*in
   wire signed [6:0] m26_9;
   assign m26_9 =7'b0;

   // m26_10 = W*in
   wire signed [6:0] m26_10;
   assign m26_10 =7'b0;

   // m26_11 = W*in
   wire signed [6:0] m26_11;
   assign m26_11 =7'b0;

   // m26_12 = W*in
   wire signed [6:0] m26_12;
   assign m26_12 =7'b0;

   // m26_13 = W*in
   wire signed [6:0] m26_13;
   assign m26_13 =7'b0;

   // m26_14 = W*in
   wire signed [6:0] m26_14;
   assign m26_14 =7'b0;

   // m26_15 = W*in
   wire signed [6:0] m26_15;
   assign m26_15 ={ {2{in26[5]}} , in26[5:1] };

   // m26_16 = W*in
   wire signed [6:0] m26_16;
   assign m26_16 =7'b0;

   // m26_17 = W*in
   wire signed [6:0] m26_17;
   assign m26_17 =7'b0;

   // m26_18 = W*in
   wire signed [6:0] m26_18;
   assign m26_18 =7'b0;

   // m26_19 = W*in
   wire signed [6:0] m26_19;
   assign m26_19 =7'b0;

   // m26_20 = W*in
   wire signed [6:0] m26_20;
   assign m26_20 =7'b0;

   // m26_21 = W*in
   wire signed [6:0] m26_21;
   assign m26_21 =7'b0;

   // m26_22 = W*in
   wire signed [6:0] m26_22;
   assign m26_22 =7'b0;

   // m26_23 = W*in
   wire signed [6:0] m26_23;
   assign m26_23 =7'b0;

   // m26_24 = W*in
   wire signed [6:0] m26_24;
   assign m26_24 =7'b0;

   // m26_25 = W*in
   wire signed [6:0] m26_25;
   assign m26_25 =7'b0;

   // m26_26 = W*in
   wire signed [6:0] m26_26;
   assign m26_26 =7'b0;

   // m26_27 = W*in
   wire signed [6:0] m26_27;
   assign m26_27 =7'b0;

   // m27_1 = W*in
   wire signed [6:0] m27_1;
   assign m27_1 =7'b0;

   // m27_2 = W*in
   wire signed [6:0] m27_2;
   assign m27_2 ={ {2{in27[5]}} , in27[5:1] };

   // m27_3 = W*in
   wire signed [6:0] m27_3;
   assign m27_3 =7'b0;

   // m27_4 = W*in
   wire signed [6:0] m27_4;
   assign m27_4 =7'b0;

   // m27_5 = W*in
   wire signed [6:0] m27_5;
   assign m27_5 =7'b0;

   // m27_6 = W*in
   wire signed [6:0] m27_6;
   assign m27_6 =7'b0;

   // m27_7 = W*in
   wire signed [6:0] m27_7;
   assign m27_7 =7'b0;

   // m27_8 = W*in
   wire signed [6:0] m27_8;
   assign m27_8 =7'b0;

   // m27_9 = W*in
   wire signed [6:0] m27_9;
   assign m27_9 =7'b0;

   // m27_10 = W*in
   wire signed [6:0] m27_10;
   assign m27_10 =7'b0;

   // m27_11 = W*in
   wire signed [6:0] m27_11;
   assign m27_11 =7'b0;

   // m27_12 = W*in
   wire signed [6:0] m27_12;
   assign m27_12 =7'b0;

   // m27_13 = W*in
   wire signed [6:0] m27_13;
   assign m27_13 =7'b0;

   // m27_14 = W*in
   wire signed [6:0] m27_14;
   assign m27_14 =7'b0;

   // m27_15 = W*in
   wire signed [6:0] m27_15;
   assign m27_15 =7'b0;

   // m27_16 = W*in
   wire signed [6:0] m27_16;
   assign m27_16 =7'b0;

   // m27_17 = W*in
   wire signed [6:0] m27_17;
   assign m27_17 =7'b0;

   // m27_18 = W*in
   wire signed [6:0] m27_18;
   assign m27_18 =7'b0;

   // m27_19 = W*in
   wire signed [6:0] m27_19;
   assign m27_19 =7'b0;

   // m27_20 = W*in
   wire signed [6:0] m27_20;
   assign m27_20 =7'b0;

   // m27_21 = W*in
   wire signed [6:0] m27_21;
   assign m27_21 =7'b0;

   // m27_22 = W*in
   wire signed [6:0] m27_22;
   assign m27_22 =7'b0;

   // m27_23 = W*in
   wire signed [6:0] m27_23;
   assign m27_23 =7'b0;

   // m27_24 = W*in
   wire signed [6:0] m27_24;
   assign m27_24 =7'b0;

   // m27_25 = W*in
   wire signed [6:0] m27_25;
   assign m27_25 ={ {2{in27[5]}} , in27[5:1] };

   // m27_26 = W*in
   wire signed [6:0] m27_26;
   assign m27_26 =7'b0;

   // m27_27 = W*in
   wire signed [6:0] m27_27;
   assign m27_27 =7'b0;

   // m28_1 = W*in
   wire signed [6:0] m28_1;
   assign m28_1 =7'b0;

   // m28_2 = W*in
   wire signed [6:0] m28_2;
   assign m28_2 =7'b0;

   // m28_3 = W*in
   wire signed [6:0] m28_3;
   assign m28_3 =7'b0;

   // m28_4 = W*in
   wire signed [6:0] m28_4;
   assign m28_4 =7'b0;

   // m28_5 = W*in
   wire signed [6:0] m28_5;
   assign m28_5 =7'b0;

   // m28_6 = W*in
   wire signed [6:0] m28_6;
   assign m28_6 =7'b0;

   // m28_7 = W*in
   wire signed [6:0] m28_7;
   assign m28_7 =7'b0;

   // m28_8 = W*in
   wire signed [6:0] m28_8;
   assign m28_8 =7'b0;

   // m28_9 = W*in
   wire signed [6:0] m28_9;
   assign m28_9 =7'b0;

   // m28_10 = W*in
   wire signed [6:0] m28_10;
   assign m28_10 =7'b0;

   // m28_11 = W*in
   wire signed [6:0] m28_11;
   assign m28_11 =7'b0;

   // m28_12 = W*in
   wire signed [6:0] m28_12;
   assign m28_12 =7'b0;

   // m28_13 = W*in
   wire signed [6:0] m28_13;
   assign m28_13 =7'b0;

   // m28_14 = W*in
   wire signed [6:0] m28_14;
   assign m28_14 =7'b0;

   // m28_15 = W*in
   wire signed [6:0] m28_15;
   assign m28_15 =7'b0;

   // m28_16 = W*in
   wire signed [6:0] m28_16;
   assign m28_16 =7'b0;

   // m28_17 = W*in
   wire signed [6:0] m28_17;
   assign m28_17 =7'b0;

   // m28_18 = W*in
   wire signed [6:0] m28_18;
   assign m28_18 =7'b0;

   // m28_19 = W*in
   wire signed [6:0] m28_19;
   assign m28_19 =7'b0;

   // m28_20 = W*in
   wire signed [6:0] m28_20;
   assign m28_20 =7'b0;

   // m28_21 = W*in
   wire signed [6:0] m28_21;
   assign m28_21 ={ {1{in28[5]}} , in28[5:0] };

   // m28_22 = W*in
   wire signed [6:0] m28_22;
   assign m28_22 =7'b0;

   // m28_23 = W*in
   wire signed [6:0] m28_23;
   assign m28_23 =7'b0;

   // m28_24 = W*in
   wire signed [6:0] m28_24;
   assign m28_24 =7'b0;

   // m28_25 = W*in
   wire signed [6:0] m28_25;
   assign m28_25 =7'b0;

   // m28_26 = W*in
   wire signed [6:0] m28_26;
   assign m28_26 =7'b0;

   // m28_27 = W*in
   wire signed [6:0] m28_27;
   assign m28_27 =7'b0;

   // m29_1 = W*in
   wire signed [6:0] m29_1;
   assign m29_1 =7'b0;

   // m29_2 = W*in
   wire signed [6:0] m29_2;
   assign m29_2 =7'b0;

   // m29_3 = W*in
   wire signed [6:0] m29_3;
   assign m29_3 =7'b0;

   // m29_4 = W*in
   wire signed [6:0] m29_4;
   assign m29_4 =7'b0;

   // m29_5 = W*in
   wire signed [6:0] m29_5;
   assign m29_5 =7'b0;

   // m29_6 = W*in
   wire signed [6:0] m29_6;
   assign m29_6 =7'b0;

   // m29_7 = W*in
   wire signed [6:0] m29_7;
   assign m29_7 ={ {1{in29[5]}} , in29[5:0] };

   // m29_8 = W*in
   wire signed [6:0] m29_8;
   assign m29_8 =7'b0;

   // m29_9 = W*in
   wire signed [6:0] m29_9;
   assign m29_9 =7'b0;

   // m29_10 = W*in
   wire signed [6:0] m29_10;
   assign m29_10 =7'b0;

   // m29_11 = W*in
   wire signed [6:0] m29_11;
   assign m29_11 =7'b0;

   // m29_12 = W*in
   wire signed [6:0] m29_12;
   assign m29_12 =7'b0;

   // m29_13 = W*in
   wire signed [6:0] m29_13;
   assign m29_13 =7'b0;

   // m29_14 = W*in
   wire signed [6:0] m29_14;
   assign m29_14 =7'b0;

   // m29_15 = W*in
   wire signed [6:0] m29_15;
   assign m29_15 =7'b0;

   // m29_16 = W*in
   wire signed [6:0] m29_16;
   assign m29_16 =7'b0;

   // m29_17 = W*in
   wire signed [6:0] m29_17;
   assign m29_17 =7'b0;

   // m29_18 = W*in
   wire signed [6:0] m29_18;
   assign m29_18 =7'b0;

   // m29_19 = W*in
   wire signed [6:0] m29_19;
   assign m29_19 =7'b0;

   // m29_20 = W*in
   wire signed [6:0] m29_20;
   assign m29_20 =7'b0;

   // m29_21 = W*in
   wire signed [6:0] m29_21;
   assign m29_21 =7'b0;

   // m29_22 = W*in
   wire signed [6:0] m29_22;
   assign m29_22 =7'b0;

   // m29_23 = W*in
   wire signed [6:0] m29_23;
   assign m29_23 =7'b0;

   // m29_24 = W*in
   wire signed [6:0] m29_24;
   assign m29_24 =7'b0;

   // m29_25 = W*in
   wire signed [6:0] m29_25;
   assign m29_25 =7'b0;

   // m29_26 = W*in
   wire signed [6:0] m29_26;
   assign m29_26 =7'b0;

   // m29_27 = W*in
   wire signed [6:0] m29_27;
   assign m29_27 =7'b0;

   // m30_1 = W*in
   wire signed [6:0] m30_1;
   assign m30_1 =7'b0;

   // m30_2 = W*in
   wire signed [6:0] m30_2;
   assign m30_2 =7'b0;

   // m30_3 = W*in
   wire signed [6:0] m30_3;
   assign m30_3 =7'b0;

   // m30_4 = W*in
   wire signed [6:0] m30_4;
   assign m30_4 =7'b0;

   // m30_5 = W*in
   wire signed [6:0] m30_5;
   assign m30_5 =7'b0;

   // m30_6 = W*in
   wire signed [6:0] m30_6;
   assign m30_6 =7'b0;

   // m30_7 = W*in
   wire signed [6:0] m30_7;
   assign m30_7 =7'b0;

   // m30_8 = W*in
   wire signed [6:0] m30_8;
   assign m30_8 =7'b0;

   // m30_9 = W*in
   wire signed [6:0] m30_9;
   wire signed [7:0] tm30_9;
   assign tm30_9[0:0] = in30[0:0];
   assign tm30_9[7:1] = { {1{in30[5]}} , in30[5:0] } + { {2{in30[5]}} , in30[5:1] };
   assign m30_9 ={ {1{tm30_9[7]}} , tm30_9[7:2] };

   // m30_10 = W*in
   wire signed [6:0] m30_10;
   assign m30_10 =7'b0;

   // m30_11 = W*in
   wire signed [6:0] m30_11;
   assign m30_11 =7'b0;

   // m30_12 = W*in
   wire signed [6:0] m30_12;
   assign m30_12 =7'b0;

   // m30_13 = W*in
   wire signed [6:0] m30_13;
   assign m30_13 =7'b0;

   // m30_14 = W*in
   wire signed [6:0] m30_14;
   assign m30_14 =7'b0;

   // m30_15 = W*in
   wire signed [6:0] m30_15;
   assign m30_15 =7'b0;

   // m30_16 = W*in
   wire signed [6:0] m30_16;
   assign m30_16 =7'b0;

   // m30_17 = W*in
   wire signed [6:0] m30_17;
   assign m30_17 =7'b0;

   // m30_18 = W*in
   wire signed [6:0] m30_18;
   assign m30_18 =7'b0;

   // m30_19 = W*in
   wire signed [6:0] m30_19;
   assign m30_19 =7'b0;

   // m30_20 = W*in
   wire signed [6:0] m30_20;
   assign m30_20 =7'b0;

   // m30_21 = W*in
   wire signed [6:0] m30_21;
   assign m30_21 =7'b0;

   // m30_22 = W*in
   wire signed [6:0] m30_22;
   assign m30_22 =7'b0;

   // m30_23 = W*in
   wire signed [6:0] m30_23;
   assign m30_23 =7'b0;

   // m30_24 = W*in
   wire signed [6:0] m30_24;
   assign m30_24 =7'b0;

   // m30_25 = W*in
   wire signed [6:0] m30_25;
   assign m30_25 =7'b0;

   // m30_26 = W*in
   wire signed [6:0] m30_26;
   assign m30_26 =7'b0;

   // m30_27 = W*in
   wire signed [6:0] m30_27;
   assign m30_27 =7'b0;

   // m31_1 = W*in
   wire signed [6:0] m31_1;
   assign m31_1 =7'b0;

   // m31_2 = W*in
   wire signed [6:0] m31_2;
   assign m31_2 =7'b0;

   // m31_3 = W*in
   wire signed [6:0] m31_3;
   assign m31_3 =7'b0;

   // m31_4 = W*in
   wire signed [6:0] m31_4;
   assign m31_4 =7'b0;

   // m31_5 = W*in
   wire signed [6:0] m31_5;
   assign m31_5 =7'b0;

   // m31_6 = W*in
   wire signed [6:0] m31_6;
   assign m31_6 =7'b0;

   // m31_7 = W*in
   wire signed [6:0] m31_7;
   wire signed [7:0] tm31_7;
   assign tm31_7[0:0] = in31[0:0];
   assign tm31_7[7:1] = { {1{in31[5]}} , in31[5:0] } + { {2{in31[5]}} , in31[5:1] };
   assign m31_7 ={ {1{tm31_7[7]}} , tm31_7[7:2] };

   // m31_8 = W*in
   wire signed [6:0] m31_8;
   assign m31_8 =7'b0;

   // m31_9 = W*in
   wire signed [6:0] m31_9;
   assign m31_9 =7'b0;

   // m31_10 = W*in
   wire signed [6:0] m31_10;
   assign m31_10 =7'b0;

   // m31_11 = W*in
   wire signed [6:0] m31_11;
   assign m31_11 =7'b0;

   // m31_12 = W*in
   wire signed [6:0] m31_12;
   assign m31_12 =7'b0;

   // m31_13 = W*in
   wire signed [6:0] m31_13;
   assign m31_13 =7'b0;

   // m31_14 = W*in
   wire signed [6:0] m31_14;
   assign m31_14 =7'b0;

   // m31_15 = W*in
   wire signed [6:0] m31_15;
   assign m31_15 =7'b0;

   // m31_16 = W*in
   wire signed [6:0] m31_16;
   assign m31_16 =7'b0;

   // m31_17 = W*in
   wire signed [6:0] m31_17;
   assign m31_17 =7'b0;

   // m31_18 = W*in
   wire signed [6:0] m31_18;
   assign m31_18 =7'b0;

   // m31_19 = W*in
   wire signed [6:0] m31_19;
   assign m31_19 =7'b0;

   // m31_20 = W*in
   wire signed [6:0] m31_20;
   assign m31_20 =7'b0;

   // m31_21 = W*in
   wire signed [6:0] m31_21;
   assign m31_21 =7'b0;

   // m31_22 = W*in
   wire signed [6:0] m31_22;
   assign m31_22 =7'b0;

   // m31_23 = W*in
   wire signed [6:0] m31_23;
   assign m31_23 =7'b0;

   // m31_24 = W*in
   wire signed [6:0] m31_24;
   assign m31_24 =7'b0;

   // m31_25 = W*in
   wire signed [6:0] m31_25;
   assign m31_25 =7'b0;

   // m31_26 = W*in
   wire signed [6:0] m31_26;
   assign m31_26 =7'b0;

   // m31_27 = W*in
   wire signed [6:0] m31_27;
   assign m31_27 =7'b0;

   // m32_1 = W*in
   wire signed [6:0] m32_1;
   assign m32_1 =7'b0;

   // m32_2 = W*in
   wire signed [6:0] m32_2;
   assign m32_2 =7'b0;

   // m32_3 = W*in
   wire signed [6:0] m32_3;
   assign m32_3 =7'b0;

   // m32_4 = W*in
   wire signed [6:0] m32_4;
   assign m32_4 =7'b0;

   // m32_5 = W*in
   wire signed [6:0] m32_5;
   assign m32_5 =7'b0;

   // m32_6 = W*in
   wire signed [6:0] m32_6;
   assign m32_6 =7'b0;

   // m32_7 = W*in
   wire signed [6:0] m32_7;
   assign m32_7 =7'b0;

   // m32_8 = W*in
   wire signed [6:0] m32_8;
   assign m32_8 =7'b0;

   // m32_9 = W*in
   wire signed [6:0] m32_9;
   assign m32_9 =7'b0;

   // m32_10 = W*in
   wire signed [6:0] m32_10;
   assign m32_10 =7'b0;

   // m32_11 = W*in
   wire signed [6:0] m32_11;
   assign m32_11 =7'b0;

   // m32_12 = W*in
   wire signed [6:0] m32_12;
   assign m32_12 =7'b0;

   // m32_13 = W*in
   wire signed [6:0] m32_13;
   assign m32_13 =7'b0;

   // m32_14 = W*in
   wire signed [6:0] m32_14;
   assign m32_14 =7'b0;

   // m32_15 = W*in
   wire signed [6:0] m32_15;
   assign m32_15 =7'b0;

   // m32_16 = W*in
   wire signed [6:0] m32_16;
   assign m32_16 =7'b0;

   // m32_17 = W*in
   wire signed [6:0] m32_17;
   assign m32_17 =7'b0;

   // m32_18 = W*in
   wire signed [6:0] m32_18;
   assign m32_18 =7'b0;

   // m32_19 = W*in
   wire signed [6:0] m32_19;
   assign m32_19 =7'b0;

   // m32_20 = W*in
   wire signed [6:0] m32_20;
   assign m32_20 =7'b0;

   // m32_21 = W*in
   wire signed [6:0] m32_21;
   assign m32_21 ={ {2{in32[5]}} , in32[5:1] };

   // m32_22 = W*in
   wire signed [6:0] m32_22;
   assign m32_22 =7'b0;

   // m32_23 = W*in
   wire signed [6:0] m32_23;
   assign m32_23 =7'b0;

   // m32_24 = W*in
   wire signed [6:0] m32_24;
   assign m32_24 =7'b0;

   // m32_25 = W*in
   wire signed [6:0] m32_25;
   assign m32_25 =7'b0;

   // m32_26 = W*in
   wire signed [6:0] m32_26;
   assign m32_26 =7'b0;

   // m32_27 = W*in
   wire signed [6:0] m32_27;
   assign m32_27 =7'b0;

   // m33_1 = W*in
   wire signed [6:0] m33_1;
   assign m33_1 =7'b0;

   // m33_2 = W*in
   wire signed [6:0] m33_2;
   assign m33_2 ={ {2{in33[5]}} , in33[5:1] };

   // m33_3 = W*in
   wire signed [6:0] m33_3;
   assign m33_3 =7'b0;

   // m33_4 = W*in
   wire signed [6:0] m33_4;
   assign m33_4 =7'b0;

   // m33_5 = W*in
   wire signed [6:0] m33_5;
   assign m33_5 =7'b0;

   // m33_6 = W*in
   wire signed [6:0] m33_6;
   assign m33_6 =7'b0;

   // m33_7 = W*in
   wire signed [6:0] m33_7;
   assign m33_7 =7'b0;

   // m33_8 = W*in
   wire signed [6:0] m33_8;
   assign m33_8 =7'b0;

   // m33_9 = W*in
   wire signed [6:0] m33_9;
   assign m33_9 =7'b0;

   // m33_10 = W*in
   wire signed [6:0] m33_10;
   assign m33_10 =7'b0;

   // m33_11 = W*in
   wire signed [6:0] m33_11;
   assign m33_11 =7'b0;

   // m33_12 = W*in
   wire signed [6:0] m33_12;
   assign m33_12 =7'b0;

   // m33_13 = W*in
   wire signed [6:0] m33_13;
   assign m33_13 =7'b0;

   // m33_14 = W*in
   wire signed [6:0] m33_14;
   assign m33_14 =7'b0;

   // m33_15 = W*in
   wire signed [6:0] m33_15;
   assign m33_15 =7'b0;

   // m33_16 = W*in
   wire signed [6:0] m33_16;
   assign m33_16 =7'b0;

   // m33_17 = W*in
   wire signed [6:0] m33_17;
   assign m33_17 =7'b0;

   // m33_18 = W*in
   wire signed [6:0] m33_18;
   assign m33_18 =7'b0;

   // m33_19 = W*in
   wire signed [6:0] m33_19;
   assign m33_19 =7'b0;

   // m33_20 = W*in
   wire signed [6:0] m33_20;
   assign m33_20 =7'b0;

   // m33_21 = W*in
   wire signed [6:0] m33_21;
   assign m33_21 =7'b0;

   // m33_22 = W*in
   wire signed [6:0] m33_22;
   assign m33_22 =7'b0;

   // m33_23 = W*in
   wire signed [6:0] m33_23;
   assign m33_23 =7'b0;

   // m33_24 = W*in
   wire signed [6:0] m33_24;
   assign m33_24 =7'b0;

   // m33_25 = W*in
   wire signed [6:0] m33_25;
   assign m33_25 =7'b0;

   // m33_26 = W*in
   wire signed [6:0] m33_26;
   assign m33_26 =7'b0;

   // m33_27 = W*in
   wire signed [6:0] m33_27;
   assign m33_27 =7'b0;

   // m34_1 = W*in
   wire signed [6:0] m34_1;
   assign m34_1 ={ {2{in34[5]}} , in34[5:1] };

   // m34_2 = W*in
   wire signed [6:0] m34_2;
   assign m34_2 =7'b0;

   // m34_3 = W*in
   wire signed [6:0] m34_3;
   assign m34_3 =7'b0;

   // m34_4 = W*in
   wire signed [6:0] m34_4;
   assign m34_4 =7'b0;

   // m34_5 = W*in
   wire signed [6:0] m34_5;
   assign m34_5 =7'b0;

   // m34_6 = W*in
   wire signed [6:0] m34_6;
   assign m34_6 =7'b0;

   // m34_7 = W*in
   wire signed [6:0] m34_7;
   assign m34_7 =7'b0;

   // m34_8 = W*in
   wire signed [6:0] m34_8;
   assign m34_8 =7'b0;

   // m34_9 = W*in
   wire signed [6:0] m34_9;
   assign m34_9 =7'b0;

   // m34_10 = W*in
   wire signed [6:0] m34_10;
   assign m34_10 =7'b0;

   // m34_11 = W*in
   wire signed [6:0] m34_11;
   assign m34_11 =7'b0;

   // m34_12 = W*in
   wire signed [6:0] m34_12;
   assign m34_12 =7'b0;

   // m34_13 = W*in
   wire signed [6:0] m34_13;
   assign m34_13 =7'b0;

   // m34_14 = W*in
   wire signed [6:0] m34_14;
   assign m34_14 =7'b0;

   // m34_15 = W*in
   wire signed [6:0] m34_15;
   assign m34_15 =7'b0;

   // m34_16 = W*in
   wire signed [6:0] m34_16;
   assign m34_16 =7'b0;

   // m34_17 = W*in
   wire signed [6:0] m34_17;
   assign m34_17 =7'b0;

   // m34_18 = W*in
   wire signed [6:0] m34_18;
   assign m34_18 =7'b0;

   // m34_19 = W*in
   wire signed [6:0] m34_19;
   assign m34_19 =7'b0;

   // m34_20 = W*in
   wire signed [6:0] m34_20;
   assign m34_20 =7'b0;

   // m34_21 = W*in
   wire signed [6:0] m34_21;
   assign m34_21 ={ {1{in34[5]}} , in34[5:0] };

   // m34_22 = W*in
   wire signed [6:0] m34_22;
   assign m34_22 =7'b0;

   // m34_23 = W*in
   wire signed [6:0] m34_23;
   assign m34_23 =7'b0;

   // m34_24 = W*in
   wire signed [6:0] m34_24;
   assign m34_24 ={ {2{neg34[5]}} , neg34[5:1] };

   // m34_25 = W*in
   wire signed [6:0] m34_25;
   assign m34_25 =7'b0;

   // m34_26 = W*in
   wire signed [6:0] m34_26;
   assign m34_26 =7'b0;

   // m34_27 = W*in
   wire signed [6:0] m34_27;
   assign m34_27 =7'b0;

   // m35_1 = W*in
   wire signed [6:0] m35_1;
   assign m35_1 =7'b0;

   // m35_2 = W*in
   wire signed [6:0] m35_2;
   assign m35_2 =7'b0;

   // m35_3 = W*in
   wire signed [6:0] m35_3;
   assign m35_3 =7'b0;

   // m35_4 = W*in
   wire signed [6:0] m35_4;
   assign m35_4 =7'b0;

   // m35_5 = W*in
   wire signed [6:0] m35_5;
   assign m35_5 =7'b0;

   // m35_6 = W*in
   wire signed [6:0] m35_6;
   assign m35_6 =7'b0;

   // m35_7 = W*in
   wire signed [6:0] m35_7;
   assign m35_7 =7'b0;

   // m35_8 = W*in
   wire signed [6:0] m35_8;
   assign m35_8 =7'b0;

   // m35_9 = W*in
   wire signed [6:0] m35_9;
   assign m35_9 =7'b0;

   // m35_10 = W*in
   wire signed [6:0] m35_10;
   assign m35_10 =7'b0;

   // m35_11 = W*in
   wire signed [6:0] m35_11;
   assign m35_11 =7'b0;

   // m35_12 = W*in
   wire signed [6:0] m35_12;
   assign m35_12 =7'b0;

   // m35_13 = W*in
   wire signed [6:0] m35_13;
   assign m35_13 =7'b0;

   // m35_14 = W*in
   wire signed [6:0] m35_14;
   assign m35_14 =7'b0;

   // m35_15 = W*in
   wire signed [6:0] m35_15;
   assign m35_15 ={ {1{in35[5]}} , in35[5:0] };

   // m35_16 = W*in
   wire signed [6:0] m35_16;
   assign m35_16 =7'b0;

   // m35_17 = W*in
   wire signed [6:0] m35_17;
   assign m35_17 =7'b0;

   // m35_18 = W*in
   wire signed [6:0] m35_18;
   assign m35_18 =7'b0;

   // m35_19 = W*in
   wire signed [6:0] m35_19;
   assign m35_19 =7'b0;

   // m35_20 = W*in
   wire signed [6:0] m35_20;
   assign m35_20 =7'b0;

   // m35_21 = W*in
   wire signed [6:0] m35_21;
   assign m35_21 =7'b0;

   // m35_22 = W*in
   wire signed [6:0] m35_22;
   assign m35_22 =7'b0;

   // m35_23 = W*in
   wire signed [6:0] m35_23;
   assign m35_23 =7'b0;

   // m35_24 = W*in
   wire signed [6:0] m35_24;
   assign m35_24 =7'b0;

   // m35_25 = W*in
   wire signed [6:0] m35_25;
   assign m35_25 =7'b0;

   // m35_26 = W*in
   wire signed [6:0] m35_26;
   assign m35_26 =7'b0;

   // m35_27 = W*in
   wire signed [6:0] m35_27;
   assign m35_27 =7'b0;

   // m36_1 = W*in
   wire signed [6:0] m36_1;
   assign m36_1 =7'b0;

   // m36_2 = W*in
   wire signed [6:0] m36_2;
   assign m36_2 =7'b0;

   // m36_3 = W*in
   wire signed [6:0] m36_3;
   assign m36_3 =7'b0;

   // m36_4 = W*in
   wire signed [6:0] m36_4;
   assign m36_4 =7'b0;

   // m36_5 = W*in
   wire signed [6:0] m36_5;
   assign m36_5 =7'b0;

   // m36_6 = W*in
   wire signed [6:0] m36_6;
   assign m36_6 ={ {2{neg36[5]}} , neg36[5:1] };

   // m36_7 = W*in
   wire signed [6:0] m36_7;
   assign m36_7 =7'b0;

   // m36_8 = W*in
   wire signed [6:0] m36_8;
   assign m36_8 =7'b0;

   // m36_9 = W*in
   wire signed [6:0] m36_9;
   assign m36_9 =7'b0;

   // m36_10 = W*in
   wire signed [6:0] m36_10;
   assign m36_10 =7'b0;

   // m36_11 = W*in
   wire signed [6:0] m36_11;
   assign m36_11 =7'b0;

   // m36_12 = W*in
   wire signed [6:0] m36_12;
   assign m36_12 ={ {2{neg36[5]}} , neg36[5:1] };

   // m36_13 = W*in
   wire signed [6:0] m36_13;
   assign m36_13 =7'b0;

   // m36_14 = W*in
   wire signed [6:0] m36_14;
   assign m36_14 =7'b0;

   // m36_15 = W*in
   wire signed [6:0] m36_15;
   assign m36_15 =7'b0;

   // m36_16 = W*in
   wire signed [6:0] m36_16;
   assign m36_16 =7'b0;

   // m36_17 = W*in
   wire signed [6:0] m36_17;
   assign m36_17 =7'b0;

   // m36_18 = W*in
   wire signed [6:0] m36_18;
   assign m36_18 =7'b0;

   // m36_19 = W*in
   wire signed [6:0] m36_19;
   assign m36_19 =7'b0;

   // m36_20 = W*in
   wire signed [6:0] m36_20;
   assign m36_20 =7'b0;

   // m36_21 = W*in
   wire signed [6:0] m36_21;
   assign m36_21 ={ {1{in36[5]}} , in36[5:0] };

   // m36_22 = W*in
   wire signed [6:0] m36_22;
   assign m36_22 =7'b0;

   // m36_23 = W*in
   wire signed [6:0] m36_23;
   assign m36_23 =7'b0;

   // m36_24 = W*in
   wire signed [6:0] m36_24;
   assign m36_24 =7'b0;

   // m36_25 = W*in
   wire signed [6:0] m36_25;
   assign m36_25 =7'b0;

   // m36_26 = W*in
   wire signed [6:0] m36_26;
   assign m36_26 =7'b0;

   // m36_27 = W*in
   wire signed [6:0] m36_27;
   assign m36_27 =7'b0;

   // m37_1 = W*in
   wire signed [6:0] m37_1;
   assign m37_1 =7'b0;

   // m37_2 = W*in
   wire signed [6:0] m37_2;
   assign m37_2 =7'b0;

   // m37_3 = W*in
   wire signed [6:0] m37_3;
   assign m37_3 =7'b0;

   // m37_4 = W*in
   wire signed [6:0] m37_4;
   assign m37_4 =7'b0;

   // m37_5 = W*in
   wire signed [6:0] m37_5;
   assign m37_5 =7'b0;

   // m37_6 = W*in
   wire signed [6:0] m37_6;
   assign m37_6 =7'b0;

   // m37_7 = W*in
   wire signed [6:0] m37_7;
   assign m37_7 =7'b0;

   // m37_8 = W*in
   wire signed [6:0] m37_8;
   assign m37_8 =7'b0;

   // m37_9 = W*in
   wire signed [6:0] m37_9;
   assign m37_9 =7'b0;

   // m37_10 = W*in
   wire signed [6:0] m37_10;
   assign m37_10 =7'b0;

   // m37_11 = W*in
   wire signed [6:0] m37_11;
   assign m37_11 =7'b0;

   // m37_12 = W*in
   wire signed [6:0] m37_12;
   assign m37_12 =7'b0;

   // m37_13 = W*in
   wire signed [6:0] m37_13;
   assign m37_13 =7'b0;

   // m37_14 = W*in
   wire signed [6:0] m37_14;
   assign m37_14 =7'b0;

   // m37_15 = W*in
   wire signed [6:0] m37_15;
   assign m37_15 =7'b0;

   // m37_16 = W*in
   wire signed [6:0] m37_16;
   assign m37_16 =7'b0;

   // m37_17 = W*in
   wire signed [6:0] m37_17;
   assign m37_17 =7'b0;

   // m37_18 = W*in
   wire signed [6:0] m37_18;
   assign m37_18 =7'b0;

   // m37_19 = W*in
   wire signed [6:0] m37_19;
   assign m37_19 =7'b0;

   // m37_20 = W*in
   wire signed [6:0] m37_20;
   assign m37_20 =7'b0;

   // m37_21 = W*in
   wire signed [6:0] m37_21;
   assign m37_21 =7'b0;

   // m37_22 = W*in
   wire signed [6:0] m37_22;
   assign m37_22 =7'b0;

   // m37_23 = W*in
   wire signed [6:0] m37_23;
   assign m37_23 =7'b0;

   // m37_24 = W*in
   wire signed [6:0] m37_24;
   assign m37_24 =7'b0;

   // m37_25 = W*in
   wire signed [6:0] m37_25;
   assign m37_25 =7'b0;

   // m37_26 = W*in
   wire signed [6:0] m37_26;
   assign m37_26 =7'b0;

   // m37_27 = W*in
   wire signed [6:0] m37_27;
   assign m37_27 ={ {2{neg37[5]}} , neg37[5:1] };

   // m38_1 = W*in
   wire signed [6:0] m38_1;
   assign m38_1 =7'b0;

   // m38_2 = W*in
   wire signed [6:0] m38_2;
   assign m38_2 =7'b0;

   // m38_3 = W*in
   wire signed [6:0] m38_3;
   assign m38_3 =7'b0;

   // m38_4 = W*in
   wire signed [6:0] m38_4;
   assign m38_4 =7'b0;

   // m38_5 = W*in
   wire signed [6:0] m38_5;
   assign m38_5 =7'b0;

   // m38_6 = W*in
   wire signed [6:0] m38_6;
   assign m38_6 =7'b0;

   // m38_7 = W*in
   wire signed [6:0] m38_7;
   assign m38_7 =7'b0;

   // m38_8 = W*in
   wire signed [6:0] m38_8;
   assign m38_8 =7'b0;

   // m38_9 = W*in
   wire signed [6:0] m38_9;
   assign m38_9 =7'b0;

   // m38_10 = W*in
   wire signed [6:0] m38_10;
   assign m38_10 =7'b0;

   // m38_11 = W*in
   wire signed [6:0] m38_11;
   assign m38_11 =7'b0;

   // m38_12 = W*in
   wire signed [6:0] m38_12;
   assign m38_12 =7'b0;

   // m38_13 = W*in
   wire signed [6:0] m38_13;
   assign m38_13 =7'b0;

   // m38_14 = W*in
   wire signed [6:0] m38_14;
   assign m38_14 =7'b0;

   // m38_15 = W*in
   wire signed [6:0] m38_15;
   assign m38_15 =7'b0;

   // m38_16 = W*in
   wire signed [6:0] m38_16;
   assign m38_16 =7'b0;

   // m38_17 = W*in
   wire signed [6:0] m38_17;
   assign m38_17 =7'b0;

   // m38_18 = W*in
   wire signed [6:0] m38_18;
   assign m38_18 =7'b0;

   // m38_19 = W*in
   wire signed [6:0] m38_19;
   assign m38_19 ={ {1{in38[5]}} , in38[5:0] };

   // m38_20 = W*in
   wire signed [6:0] m38_20;
   assign m38_20 =7'b0;

   // m38_21 = W*in
   wire signed [6:0] m38_21;
   assign m38_21 =7'b0;

   // m38_22 = W*in
   wire signed [6:0] m38_22;
   assign m38_22 =7'b0;

   // m38_23 = W*in
   wire signed [6:0] m38_23;
   assign m38_23 =7'b0;

   // m38_24 = W*in
   wire signed [6:0] m38_24;
   assign m38_24 =7'b0;

   // m38_25 = W*in
   wire signed [6:0] m38_25;
   assign m38_25 =7'b0;

   // m38_26 = W*in
   wire signed [6:0] m38_26;
   assign m38_26 =7'b0;

   // m38_27 = W*in
   wire signed [6:0] m38_27;
   assign m38_27 =7'b0;

   // m39_1 = W*in
   wire signed [6:0] m39_1;
   assign m39_1 =7'b0;

   // m39_2 = W*in
   wire signed [6:0] m39_2;
   assign m39_2 =7'b0;

   // m39_3 = W*in
   wire signed [6:0] m39_3;
   assign m39_3 ={ {1{in39[5]}} , in39[5:0] };

   // m39_4 = W*in
   wire signed [6:0] m39_4;
   assign m39_4 =7'b0;

   // m39_5 = W*in
   wire signed [6:0] m39_5;
   assign m39_5 =7'b0;

   // m39_6 = W*in
   wire signed [6:0] m39_6;
   assign m39_6 =7'b0;

   // m39_7 = W*in
   wire signed [6:0] m39_7;
   assign m39_7 =7'b0;

   // m39_8 = W*in
   wire signed [6:0] m39_8;
   assign m39_8 =7'b0;

   // m39_9 = W*in
   wire signed [6:0] m39_9;
   assign m39_9 ={ {1{in39[5]}} , in39[5:0] };

   // m39_10 = W*in
   wire signed [6:0] m39_10;
   assign m39_10 =7'b0;

   // m39_11 = W*in
   wire signed [6:0] m39_11;
   assign m39_11 =7'b0;

   // m39_12 = W*in
   wire signed [6:0] m39_12;
   assign m39_12 =7'b0;

   // m39_13 = W*in
   wire signed [6:0] m39_13;
   assign m39_13 =7'b0;

   // m39_14 = W*in
   wire signed [6:0] m39_14;
   assign m39_14 =7'b0;

   // m39_15 = W*in
   wire signed [6:0] m39_15;
   assign m39_15 =7'b0;

   // m39_16 = W*in
   wire signed [6:0] m39_16;
   assign m39_16 =7'b0;

   // m39_17 = W*in
   wire signed [6:0] m39_17;
   assign m39_17 =7'b0;

   // m39_18 = W*in
   wire signed [6:0] m39_18;
   assign m39_18 =7'b0;

   // m39_19 = W*in
   wire signed [6:0] m39_19;
   assign m39_19 =7'b0;

   // m39_20 = W*in
   wire signed [6:0] m39_20;
   assign m39_20 =7'b0;

   // m39_21 = W*in
   wire signed [6:0] m39_21;
   assign m39_21 =7'b0;

   // m39_22 = W*in
   wire signed [6:0] m39_22;
   assign m39_22 =7'b0;

   // m39_23 = W*in
   wire signed [6:0] m39_23;
   assign m39_23 =7'b0;

   // m39_24 = W*in
   wire signed [6:0] m39_24;
   assign m39_24 =7'b0;

   // m39_25 = W*in
   wire signed [6:0] m39_25;
   assign m39_25 =7'b0;

   // m39_26 = W*in
   wire signed [6:0] m39_26;
   assign m39_26 =7'b0;

   // m39_27 = W*in
   wire signed [6:0] m39_27;
   assign m39_27 =7'b0;

   // m40_1 = W*in
   wire signed [6:0] m40_1;
   assign m40_1 ={ {1{in40[5]}} , in40[5:0] };

   // m40_2 = W*in
   wire signed [6:0] m40_2;
   assign m40_2 =7'b0;

   // m40_3 = W*in
   wire signed [6:0] m40_3;
   assign m40_3 =7'b0;

   // m40_4 = W*in
   wire signed [6:0] m40_4;
   assign m40_4 =7'b0;

   // m40_5 = W*in
   wire signed [6:0] m40_5;
   assign m40_5 =7'b0;

   // m40_6 = W*in
   wire signed [6:0] m40_6;
   assign m40_6 =7'b0;

   // m40_7 = W*in
   wire signed [6:0] m40_7;
   assign m40_7 =7'b0;

   // m40_8 = W*in
   wire signed [6:0] m40_8;
   assign m40_8 =7'b0;

   // m40_9 = W*in
   wire signed [6:0] m40_9;
   assign m40_9 =7'b0;

   // m40_10 = W*in
   wire signed [6:0] m40_10;
   assign m40_10 =7'b0;

   // m40_11 = W*in
   wire signed [6:0] m40_11;
   assign m40_11 =7'b0;

   // m40_12 = W*in
   wire signed [6:0] m40_12;
   assign m40_12 =7'b0;

   // m40_13 = W*in
   wire signed [6:0] m40_13;
   assign m40_13 =7'b0;

   // m40_14 = W*in
   wire signed [6:0] m40_14;
   assign m40_14 ={ {2{in40[5]}} , in40[5:1] };

   // m40_15 = W*in
   wire signed [6:0] m40_15;
   assign m40_15 =7'b0;

   // m40_16 = W*in
   wire signed [6:0] m40_16;
   assign m40_16 =7'b0;

   // m40_17 = W*in
   wire signed [6:0] m40_17;
   assign m40_17 =7'b0;

   // m40_18 = W*in
   wire signed [6:0] m40_18;
   assign m40_18 =7'b0;

   // m40_19 = W*in
   wire signed [6:0] m40_19;
   assign m40_19 =7'b0;

   // m40_20 = W*in
   wire signed [6:0] m40_20;
   assign m40_20 =7'b0;

   // m40_21 = W*in
   wire signed [6:0] m40_21;
   assign m40_21 =7'b0;

   // m40_22 = W*in
   wire signed [6:0] m40_22;
   assign m40_22 ={ {2{in40[5]}} , in40[5:1] };

   // m40_23 = W*in
   wire signed [6:0] m40_23;
   assign m40_23 =7'b0;

   // m40_24 = W*in
   wire signed [6:0] m40_24;
   assign m40_24 =7'b0;

   // m40_25 = W*in
   wire signed [6:0] m40_25;
   assign m40_25 =7'b0;

   // m40_26 = W*in
   wire signed [6:0] m40_26;
   assign m40_26 =7'b0;

   // m40_27 = W*in
   wire signed [6:0] m40_27;
   assign m40_27 =7'b0;

   // m41_1 = W*in
   wire signed [6:0] m41_1;
   assign m41_1 =7'b0;

   // m41_2 = W*in
   wire signed [6:0] m41_2;
   assign m41_2 =7'b0;

   // m41_3 = W*in
   wire signed [6:0] m41_3;
   assign m41_3 =7'b0;

   // m41_4 = W*in
   wire signed [6:0] m41_4;
   assign m41_4 =7'b0;

   // m41_5 = W*in
   wire signed [6:0] m41_5;
   assign m41_5 =7'b0;

   // m41_6 = W*in
   wire signed [6:0] m41_6;
   assign m41_6 =7'b0;

   // m41_7 = W*in
   wire signed [6:0] m41_7;
   assign m41_7 =7'b0;

   // m41_8 = W*in
   wire signed [6:0] m41_8;
   assign m41_8 =7'b0;

   // m41_9 = W*in
   wire signed [6:0] m41_9;
   assign m41_9 =7'b0;

   // m41_10 = W*in
   wire signed [6:0] m41_10;
   assign m41_10 =7'b0;

   // m41_11 = W*in
   wire signed [6:0] m41_11;
   assign m41_11 =7'b0;

   // m41_12 = W*in
   wire signed [6:0] m41_12;
   assign m41_12 =7'b0;

   // m41_13 = W*in
   wire signed [6:0] m41_13;
   assign m41_13 =7'b0;

   // m41_14 = W*in
   wire signed [6:0] m41_14;
   assign m41_14 =7'b0;

   // m41_15 = W*in
   wire signed [6:0] m41_15;
   assign m41_15 =7'b0;

   // m41_16 = W*in
   wire signed [6:0] m41_16;
   assign m41_16 =7'b0;

   // m41_17 = W*in
   wire signed [6:0] m41_17;
   assign m41_17 =7'b0;

   // m41_18 = W*in
   wire signed [6:0] m41_18;
   assign m41_18 =7'b0;

   // m41_19 = W*in
   wire signed [6:0] m41_19;
   assign m41_19 =7'b0;

   // m41_20 = W*in
   wire signed [6:0] m41_20;
   assign m41_20 =7'b0;

   // m41_21 = W*in
   wire signed [6:0] m41_21;
   assign m41_21 =7'b0;

   // m41_22 = W*in
   wire signed [6:0] m41_22;
   assign m41_22 ={ {2{in41[5]}} , in41[5:1] };

   // m41_23 = W*in
   wire signed [6:0] m41_23;
   assign m41_23 =7'b0;

   // m41_24 = W*in
   wire signed [6:0] m41_24;
   assign m41_24 =7'b0;

   // m41_25 = W*in
   wire signed [6:0] m41_25;
   assign m41_25 =7'b0;

   // m41_26 = W*in
   wire signed [6:0] m41_26;
   assign m41_26 =7'b0;

   // m41_27 = W*in
   wire signed [6:0] m41_27;
   assign m41_27 =7'b0;

   // m42_1 = W*in
   wire signed [6:0] m42_1;
   assign m42_1 =7'b0;

   // m42_2 = W*in
   wire signed [6:0] m42_2;
   assign m42_2 =7'b0;

   // m42_3 = W*in
   wire signed [6:0] m42_3;
   assign m42_3 =7'b0;

   // m42_4 = W*in
   wire signed [6:0] m42_4;
   assign m42_4 =7'b0;

   // m42_5 = W*in
   wire signed [6:0] m42_5;
   assign m42_5 =7'b0;

   // m42_6 = W*in
   wire signed [6:0] m42_6;
   assign m42_6 =7'b0;

   // m42_7 = W*in
   wire signed [6:0] m42_7;
   assign m42_7 =7'b0;

   // m42_8 = W*in
   wire signed [6:0] m42_8;
   assign m42_8 =7'b0;

   // m42_9 = W*in
   wire signed [6:0] m42_9;
   assign m42_9 =7'b0;

   // m42_10 = W*in
   wire signed [6:0] m42_10;
   assign m42_10 =7'b0;

   // m42_11 = W*in
   wire signed [6:0] m42_11;
   assign m42_11 =7'b0;

   // m42_12 = W*in
   wire signed [6:0] m42_12;
   assign m42_12 =7'b0;

   // m42_13 = W*in
   wire signed [6:0] m42_13;
   assign m42_13 ={ {1{in42[5]}} , in42[5:0] };

   // m42_14 = W*in
   wire signed [6:0] m42_14;
   assign m42_14 =7'b0;

   // m42_15 = W*in
   wire signed [6:0] m42_15;
   assign m42_15 =7'b0;

   // m42_16 = W*in
   wire signed [6:0] m42_16;
   assign m42_16 =7'b0;

   // m42_17 = W*in
   wire signed [6:0] m42_17;
   assign m42_17 =7'b0;

   // m42_18 = W*in
   wire signed [6:0] m42_18;
   assign m42_18 =7'b0;

   // m42_19 = W*in
   wire signed [6:0] m42_19;
   assign m42_19 =7'b0;

   // m42_20 = W*in
   wire signed [6:0] m42_20;
   assign m42_20 =7'b0;

   // m42_21 = W*in
   wire signed [6:0] m42_21;
   assign m42_21 =7'b0;

   // m42_22 = W*in
   wire signed [6:0] m42_22;
   wire signed [7:0] tm42_22;
   assign tm42_22[0:0] = in42[0:0];
   assign tm42_22[7:1] = { {1{in42[5]}} , in42[5:0] } + { {2{in42[5]}} , in42[5:1] };
   assign m42_22 ={ {1{tm42_22[7]}} , tm42_22[7:2] };

   // m42_23 = W*in
   wire signed [6:0] m42_23;
   assign m42_23 =7'b0;

   // m42_24 = W*in
   wire signed [6:0] m42_24;
   assign m42_24 =7'b0;

   // m42_25 = W*in
   wire signed [6:0] m42_25;
   assign m42_25 =7'b0;

   // m42_26 = W*in
   wire signed [6:0] m42_26;
   assign m42_26 =7'b0;

   // m42_27 = W*in
   wire signed [6:0] m42_27;
   assign m42_27 =7'b0;

   // m43_1 = W*in
   wire signed [6:0] m43_1;
   assign m43_1 =7'b0;

   // m43_2 = W*in
   wire signed [6:0] m43_2;
   assign m43_2 =7'b0;

   // m43_3 = W*in
   wire signed [6:0] m43_3;
   assign m43_3 =7'b0;

   // m43_4 = W*in
   wire signed [6:0] m43_4;
   assign m43_4 =7'b0;

   // m43_5 = W*in
   wire signed [6:0] m43_5;
   assign m43_5 =7'b0;

   // m43_6 = W*in
   wire signed [6:0] m43_6;
   assign m43_6 =7'b0;

   // m43_7 = W*in
   wire signed [6:0] m43_7;
   assign m43_7 ={ {1{in43[5]}} , in43[5:0] };

   // m43_8 = W*in
   wire signed [6:0] m43_8;
   assign m43_8 =7'b0;

   // m43_9 = W*in
   wire signed [6:0] m43_9;
   assign m43_9 =7'b0;

   // m43_10 = W*in
   wire signed [6:0] m43_10;
   assign m43_10 =7'b0;

   // m43_11 = W*in
   wire signed [6:0] m43_11;
   assign m43_11 =7'b0;

   // m43_12 = W*in
   wire signed [6:0] m43_12;
   assign m43_12 =7'b0;

   // m43_13 = W*in
   wire signed [6:0] m43_13;
   assign m43_13 =7'b0;

   // m43_14 = W*in
   wire signed [6:0] m43_14;
   assign m43_14 =7'b0;

   // m43_15 = W*in
   wire signed [6:0] m43_15;
   assign m43_15 =7'b0;

   // m43_16 = W*in
   wire signed [6:0] m43_16;
   assign m43_16 =7'b0;

   // m43_17 = W*in
   wire signed [6:0] m43_17;
   assign m43_17 =7'b0;

   // m43_18 = W*in
   wire signed [6:0] m43_18;
   assign m43_18 =7'b0;

   // m43_19 = W*in
   wire signed [6:0] m43_19;
   assign m43_19 =7'b0;

   // m43_20 = W*in
   wire signed [6:0] m43_20;
   assign m43_20 =7'b0;

   // m43_21 = W*in
   wire signed [6:0] m43_21;
   assign m43_21 =7'b0;

   // m43_22 = W*in
   wire signed [6:0] m43_22;
   assign m43_22 =7'b0;

   // m43_23 = W*in
   wire signed [6:0] m43_23;
   assign m43_23 =7'b0;

   // m43_24 = W*in
   wire signed [6:0] m43_24;
   assign m43_24 =7'b0;

   // m43_25 = W*in
   wire signed [6:0] m43_25;
   assign m43_25 =7'b0;

   // m43_26 = W*in
   wire signed [6:0] m43_26;
   assign m43_26 =7'b0;

   // m43_27 = W*in
   wire signed [6:0] m43_27;
   assign m43_27 =7'b0;

   // m44_1 = W*in
   wire signed [6:0] m44_1;
   assign m44_1 =7'b0;

   // m44_2 = W*in
   wire signed [6:0] m44_2;
   assign m44_2 ={ {1{in44[5]}} , in44[5:0] };

   // m44_3 = W*in
   wire signed [6:0] m44_3;
   assign m44_3 =7'b0;

   // m44_4 = W*in
   wire signed [6:0] m44_4;
   assign m44_4 =7'b0;

   // m44_5 = W*in
   wire signed [6:0] m44_5;
   assign m44_5 =7'b0;

   // m44_6 = W*in
   wire signed [6:0] m44_6;
   assign m44_6 =7'b0;

   // m44_7 = W*in
   wire signed [6:0] m44_7;
   assign m44_7 =7'b0;

   // m44_8 = W*in
   wire signed [6:0] m44_8;
   assign m44_8 =7'b0;

   // m44_9 = W*in
   wire signed [6:0] m44_9;
   assign m44_9 =7'b0;

   // m44_10 = W*in
   wire signed [6:0] m44_10;
   assign m44_10 =7'b0;

   // m44_11 = W*in
   wire signed [6:0] m44_11;
   assign m44_11 =7'b0;

   // m44_12 = W*in
   wire signed [6:0] m44_12;
   assign m44_12 =7'b0;

   // m44_13 = W*in
   wire signed [6:0] m44_13;
   assign m44_13 =7'b0;

   // m44_14 = W*in
   wire signed [6:0] m44_14;
   assign m44_14 =7'b0;

   // m44_15 = W*in
   wire signed [6:0] m44_15;
   assign m44_15 =7'b0;

   // m44_16 = W*in
   wire signed [6:0] m44_16;
   assign m44_16 =7'b0;

   // m44_17 = W*in
   wire signed [6:0] m44_17;
   assign m44_17 =7'b0;

   // m44_18 = W*in
   wire signed [6:0] m44_18;
   assign m44_18 =7'b0;

   // m44_19 = W*in
   wire signed [6:0] m44_19;
   assign m44_19 =7'b0;

   // m44_20 = W*in
   wire signed [6:0] m44_20;
   assign m44_20 =7'b0;

   // m44_21 = W*in
   wire signed [6:0] m44_21;
   assign m44_21 =7'b0;

   // m44_22 = W*in
   wire signed [6:0] m44_22;
   assign m44_22 =7'b0;

   // m44_23 = W*in
   wire signed [6:0] m44_23;
   assign m44_23 =7'b0;

   // m44_24 = W*in
   wire signed [6:0] m44_24;
   assign m44_24 =7'b0;

   // m44_25 = W*in
   wire signed [6:0] m44_25;
   assign m44_25 =7'b0;

   // m44_26 = W*in
   wire signed [6:0] m44_26;
   assign m44_26 =7'b0;

   // m44_27 = W*in
   wire signed [6:0] m44_27;
   assign m44_27 =7'b0;

   // m45_1 = W*in
   wire signed [6:0] m45_1;
   assign m45_1 =7'b0;

   // m45_2 = W*in
   wire signed [6:0] m45_2;
   assign m45_2 =7'b0;

   // m45_3 = W*in
   wire signed [6:0] m45_3;
   assign m45_3 =7'b0;

   // m45_4 = W*in
   wire signed [6:0] m45_4;
   assign m45_4 =7'b0;

   // m45_5 = W*in
   wire signed [6:0] m45_5;
   assign m45_5 =7'b0;

   // m45_6 = W*in
   wire signed [6:0] m45_6;
   assign m45_6 =7'b0;

   // m45_7 = W*in
   wire signed [6:0] m45_7;
   assign m45_7 ={ {2{in45[5]}} , in45[5:1] };

   // m45_8 = W*in
   wire signed [6:0] m45_8;
   assign m45_8 =7'b0;

   // m45_9 = W*in
   wire signed [6:0] m45_9;
   assign m45_9 =7'b0;

   // m45_10 = W*in
   wire signed [6:0] m45_10;
   assign m45_10 =7'b0;

   // m45_11 = W*in
   wire signed [6:0] m45_11;
   assign m45_11 =7'b0;

   // m45_12 = W*in
   wire signed [6:0] m45_12;
   assign m45_12 =7'b0;

   // m45_13 = W*in
   wire signed [6:0] m45_13;
   assign m45_13 =7'b0;

   // m45_14 = W*in
   wire signed [6:0] m45_14;
   assign m45_14 =7'b0;

   // m45_15 = W*in
   wire signed [6:0] m45_15;
   assign m45_15 =7'b0;

   // m45_16 = W*in
   wire signed [6:0] m45_16;
   assign m45_16 =7'b0;

   // m45_17 = W*in
   wire signed [6:0] m45_17;
   assign m45_17 =7'b0;

   // m45_18 = W*in
   wire signed [6:0] m45_18;
   assign m45_18 =7'b0;

   // m45_19 = W*in
   wire signed [6:0] m45_19;
   assign m45_19 =7'b0;

   // m45_20 = W*in
   wire signed [6:0] m45_20;
   assign m45_20 =7'b0;

   // m45_21 = W*in
   wire signed [6:0] m45_21;
   assign m45_21 =7'b0;

   // m45_22 = W*in
   wire signed [6:0] m45_22;
   assign m45_22 =7'b0;

   // m45_23 = W*in
   wire signed [6:0] m45_23;
   assign m45_23 =7'b0;

   // m45_24 = W*in
   wire signed [6:0] m45_24;
   assign m45_24 =7'b0;

   // m45_25 = W*in
   wire signed [6:0] m45_25;
   assign m45_25 =7'b0;

   // m45_26 = W*in
   wire signed [6:0] m45_26;
   assign m45_26 =7'b0;

   // m45_27 = W*in
   wire signed [6:0] m45_27;
   assign m45_27 =7'b0;

   // m46_1 = W*in
   wire signed [6:0] m46_1;
   assign m46_1 =7'b0;

   // m46_2 = W*in
   wire signed [6:0] m46_2;
   assign m46_2 =7'b0;

   // m46_3 = W*in
   wire signed [6:0] m46_3;
   assign m46_3 =7'b0;

   // m46_4 = W*in
   wire signed [6:0] m46_4;
   assign m46_4 =7'b0;

   // m46_5 = W*in
   wire signed [6:0] m46_5;
   assign m46_5 =7'b0;

   // m46_6 = W*in
   wire signed [6:0] m46_6;
   assign m46_6 =7'b0;

   // m46_7 = W*in
   wire signed [6:0] m46_7;
   assign m46_7 =7'b0;

   // m46_8 = W*in
   wire signed [6:0] m46_8;
   assign m46_8 =7'b0;

   // m46_9 = W*in
   wire signed [6:0] m46_9;
   assign m46_9 =7'b0;

   // m46_10 = W*in
   wire signed [6:0] m46_10;
   assign m46_10 =7'b0;

   // m46_11 = W*in
   wire signed [6:0] m46_11;
   assign m46_11 =7'b0;

   // m46_12 = W*in
   wire signed [6:0] m46_12;
   assign m46_12 =7'b0;

   // m46_13 = W*in
   wire signed [6:0] m46_13;
   assign m46_13 =7'b0;

   // m46_14 = W*in
   wire signed [6:0] m46_14;
   assign m46_14 =7'b0;

   // m46_15 = W*in
   wire signed [6:0] m46_15;
   assign m46_15 =7'b0;

   // m46_16 = W*in
   wire signed [6:0] m46_16;
   assign m46_16 =7'b0;

   // m46_17 = W*in
   wire signed [6:0] m46_17;
   assign m46_17 =7'b0;

   // m46_18 = W*in
   wire signed [6:0] m46_18;
   assign m46_18 =7'b0;

   // m46_19 = W*in
   wire signed [6:0] m46_19;
   assign m46_19 =7'b0;

   // m46_20 = W*in
   wire signed [6:0] m46_20;
   assign m46_20 =7'b0;

   // m46_21 = W*in
   wire signed [6:0] m46_21;
   assign m46_21 =7'b0;

   // m46_22 = W*in
   wire signed [6:0] m46_22;
   assign m46_22 =7'b0;

   // m46_23 = W*in
   wire signed [6:0] m46_23;
   assign m46_23 ={ {1{in46[5]}} , in46[5:0] };

   // m46_24 = W*in
   wire signed [6:0] m46_24;
   assign m46_24 =7'b0;

   // m46_25 = W*in
   wire signed [6:0] m46_25;
   assign m46_25 =7'b0;

   // m46_26 = W*in
   wire signed [6:0] m46_26;
   assign m46_26 =7'b0;

   // m46_27 = W*in
   wire signed [6:0] m46_27;
   assign m46_27 =7'b0;

   // m47_1 = W*in
   wire signed [6:0] m47_1;
   assign m47_1 =7'b0;

   // m47_2 = W*in
   wire signed [6:0] m47_2;
   assign m47_2 =7'b0;

   // m47_3 = W*in
   wire signed [6:0] m47_3;
   assign m47_3 =7'b0;

   // m47_4 = W*in
   wire signed [6:0] m47_4;
   assign m47_4 =7'b0;

   // m47_5 = W*in
   wire signed [6:0] m47_5;
   assign m47_5 =7'b0;

   // m47_6 = W*in
   wire signed [6:0] m47_6;
   assign m47_6 =7'b0;

   // m47_7 = W*in
   wire signed [6:0] m47_7;
   assign m47_7 =7'b0;

   // m47_8 = W*in
   wire signed [6:0] m47_8;
   assign m47_8 =7'b0;

   // m47_9 = W*in
   wire signed [6:0] m47_9;
   assign m47_9 =7'b0;

   // m47_10 = W*in
   wire signed [6:0] m47_10;
   assign m47_10 =7'b0;

   // m47_11 = W*in
   wire signed [6:0] m47_11;
   assign m47_11 =7'b0;

   // m47_12 = W*in
   wire signed [6:0] m47_12;
   assign m47_12 =7'b0;

   // m47_13 = W*in
   wire signed [6:0] m47_13;
   assign m47_13 =7'b0;

   // m47_14 = W*in
   wire signed [6:0] m47_14;
   assign m47_14 =7'b0;

   // m47_15 = W*in
   wire signed [6:0] m47_15;
   assign m47_15 =7'b0;

   // m47_16 = W*in
   wire signed [6:0] m47_16;
   assign m47_16 =7'b0;

   // m47_17 = W*in
   wire signed [6:0] m47_17;
   assign m47_17 =7'b0;

   // m47_18 = W*in
   wire signed [6:0] m47_18;
   assign m47_18 =7'b0;

   // m47_19 = W*in
   wire signed [6:0] m47_19;
   assign m47_19 =7'b0;

   // m47_20 = W*in
   wire signed [6:0] m47_20;
   assign m47_20 =7'b0;

   // m47_21 = W*in
   wire signed [6:0] m47_21;
   assign m47_21 =7'b0;

   // m47_22 = W*in
   wire signed [6:0] m47_22;
   assign m47_22 =7'b0;

   // m47_23 = W*in
   wire signed [6:0] m47_23;
   assign m47_23 =7'b0;

   // m47_24 = W*in
   wire signed [6:0] m47_24;
   assign m47_24 =7'b0;

   // m47_25 = W*in
   wire signed [6:0] m47_25;
   assign m47_25 ={ {1{in47[5]}} , in47[5:0] };

   // m47_26 = W*in
   wire signed [6:0] m47_26;
   assign m47_26 =7'b0;

   // m47_27 = W*in
   wire signed [6:0] m47_27;
   assign m47_27 =7'b0;

   // m48_1 = W*in
   wire signed [6:0] m48_1;
   assign m48_1 =7'b0;

   // m48_2 = W*in
   wire signed [6:0] m48_2;
   assign m48_2 =7'b0;

   // m48_3 = W*in
   wire signed [6:0] m48_3;
   assign m48_3 =7'b0;

   // m48_4 = W*in
   wire signed [6:0] m48_4;
   assign m48_4 =7'b0;

   // m48_5 = W*in
   wire signed [6:0] m48_5;
   assign m48_5 =7'b0;

   // m48_6 = W*in
   wire signed [6:0] m48_6;
   assign m48_6 =7'b0;

   // m48_7 = W*in
   wire signed [6:0] m48_7;
   assign m48_7 =7'b0;

   // m48_8 = W*in
   wire signed [6:0] m48_8;
   assign m48_8 =7'b0;

   // m48_9 = W*in
   wire signed [6:0] m48_9;
   assign m48_9 =7'b0;

   // m48_10 = W*in
   wire signed [6:0] m48_10;
   assign m48_10 =7'b0;

   // m48_11 = W*in
   wire signed [6:0] m48_11;
   assign m48_11 =7'b0;

   // m48_12 = W*in
   wire signed [6:0] m48_12;
   assign m48_12 =7'b0;

   // m48_13 = W*in
   wire signed [6:0] m48_13;
   assign m48_13 =7'b0;

   // m48_14 = W*in
   wire signed [6:0] m48_14;
   assign m48_14 =7'b0;

   // m48_15 = W*in
   wire signed [6:0] m48_15;
   assign m48_15 =7'b0;

   // m48_16 = W*in
   wire signed [6:0] m48_16;
   assign m48_16 =7'b0;

   // m48_17 = W*in
   wire signed [6:0] m48_17;
   assign m48_17 =7'b0;

   // m48_18 = W*in
   wire signed [6:0] m48_18;
   assign m48_18 =7'b0;

   // m48_19 = W*in
   wire signed [6:0] m48_19;
   assign m48_19 =7'b0;

   // m48_20 = W*in
   wire signed [6:0] m48_20;
   assign m48_20 =7'b0;

   // m48_21 = W*in
   wire signed [6:0] m48_21;
   assign m48_21 ={ {2{in48[5]}} , in48[5:1] };

   // m48_22 = W*in
   wire signed [6:0] m48_22;
   assign m48_22 =7'b0;

   // m48_23 = W*in
   wire signed [6:0] m48_23;
   assign m48_23 =7'b0;

   // m48_24 = W*in
   wire signed [6:0] m48_24;
   assign m48_24 =7'b0;

   // m48_25 = W*in
   wire signed [6:0] m48_25;
   assign m48_25 =7'b0;

   // m48_26 = W*in
   wire signed [6:0] m48_26;
   assign m48_26 =7'b0;

   // m48_27 = W*in
   wire signed [6:0] m48_27;
   assign m48_27 =7'b0;

   // m49_1 = W*in
   wire signed [6:0] m49_1;
   assign m49_1 =7'b0;

   // m49_2 = W*in
   wire signed [6:0] m49_2;
   assign m49_2 =7'b0;

   // m49_3 = W*in
   wire signed [6:0] m49_3;
   assign m49_3 =7'b0;

   // m49_4 = W*in
   wire signed [6:0] m49_4;
   assign m49_4 =7'b0;

   // m49_5 = W*in
   wire signed [6:0] m49_5;
   assign m49_5 =7'b0;

   // m49_6 = W*in
   wire signed [6:0] m49_6;
   assign m49_6 =7'b0;

   // m49_7 = W*in
   wire signed [6:0] m49_7;
   assign m49_7 =7'b0;

   // m49_8 = W*in
   wire signed [6:0] m49_8;
   assign m49_8 =7'b0;

   // m49_9 = W*in
   wire signed [6:0] m49_9;
   assign m49_9 =7'b0;

   // m49_10 = W*in
   wire signed [6:0] m49_10;
   assign m49_10 =7'b0;

   // m49_11 = W*in
   wire signed [6:0] m49_11;
   assign m49_11 =7'b0;

   // m49_12 = W*in
   wire signed [6:0] m49_12;
   assign m49_12 =7'b0;

   // m49_13 = W*in
   wire signed [6:0] m49_13;
   assign m49_13 =7'b0;

   // m49_14 = W*in
   wire signed [6:0] m49_14;
   assign m49_14 =7'b0;

   // m49_15 = W*in
   wire signed [6:0] m49_15;
   assign m49_15 =7'b0;

   // m49_16 = W*in
   wire signed [6:0] m49_16;
   assign m49_16 =7'b0;

   // m49_17 = W*in
   wire signed [6:0] m49_17;
   assign m49_17 =7'b0;

   // m49_18 = W*in
   wire signed [6:0] m49_18;
   assign m49_18 =7'b0;

   // m49_19 = W*in
   wire signed [6:0] m49_19;
   assign m49_19 =7'b0;

   // m49_20 = W*in
   wire signed [6:0] m49_20;
   assign m49_20 ={ {2{in49[5]}} , in49[5:1] };

   // m49_21 = W*in
   wire signed [6:0] m49_21;
   assign m49_21 =7'b0;

   // m49_22 = W*in
   wire signed [6:0] m49_22;
   assign m49_22 =7'b0;

   // m49_23 = W*in
   wire signed [6:0] m49_23;
   assign m49_23 =7'b0;

   // m49_24 = W*in
   wire signed [6:0] m49_24;
   assign m49_24 =7'b0;

   // m49_25 = W*in
   wire signed [6:0] m49_25;
   assign m49_25 =7'b0;

   // m49_26 = W*in
   wire signed [6:0] m49_26;
   assign m49_26 =7'b0;

   // m49_27 = W*in
   wire signed [6:0] m49_27;
   assign m49_27 =7'b0;

   // m50_1 = W*in
   wire signed [6:0] m50_1;
   assign m50_1 =7'b0;

   // m50_2 = W*in
   wire signed [6:0] m50_2;
   assign m50_2 =7'b0;

   // m50_3 = W*in
   wire signed [6:0] m50_3;
   assign m50_3 =7'b0;

   // m50_4 = W*in
   wire signed [6:0] m50_4;
   assign m50_4 =7'b0;

   // m50_5 = W*in
   wire signed [6:0] m50_5;
   assign m50_5 =7'b0;

   // m50_6 = W*in
   wire signed [6:0] m50_6;
   assign m50_6 ={ {2{in50[5]}} , in50[5:1] };

   // m50_7 = W*in
   wire signed [6:0] m50_7;
   assign m50_7 =7'b0;

   // m50_8 = W*in
   wire signed [6:0] m50_8;
   assign m50_8 =7'b0;

   // m50_9 = W*in
   wire signed [6:0] m50_9;
   assign m50_9 =7'b0;

   // m50_10 = W*in
   wire signed [6:0] m50_10;
   assign m50_10 =7'b0;

   // m50_11 = W*in
   wire signed [6:0] m50_11;
   assign m50_11 =7'b0;

   // m50_12 = W*in
   wire signed [6:0] m50_12;
   assign m50_12 =7'b0;

   // m50_13 = W*in
   wire signed [6:0] m50_13;
   assign m50_13 =7'b0;

   // m50_14 = W*in
   wire signed [6:0] m50_14;
   assign m50_14 =7'b0;

   // m50_15 = W*in
   wire signed [6:0] m50_15;
   assign m50_15 =7'b0;

   // m50_16 = W*in
   wire signed [6:0] m50_16;
   assign m50_16 =7'b0;

   // m50_17 = W*in
   wire signed [6:0] m50_17;
   assign m50_17 =7'b0;

   // m50_18 = W*in
   wire signed [6:0] m50_18;
   assign m50_18 =7'b0;

   // m50_19 = W*in
   wire signed [6:0] m50_19;
   assign m50_19 =7'b0;

   // m50_20 = W*in
   wire signed [6:0] m50_20;
   assign m50_20 =7'b0;

   // m50_21 = W*in
   wire signed [6:0] m50_21;
   assign m50_21 =7'b0;

   // m50_22 = W*in
   wire signed [6:0] m50_22;
   assign m50_22 =7'b0;

   // m50_23 = W*in
   wire signed [6:0] m50_23;
   assign m50_23 =7'b0;

   // m50_24 = W*in
   wire signed [6:0] m50_24;
   assign m50_24 =7'b0;

   // m50_25 = W*in
   wire signed [6:0] m50_25;
   assign m50_25 =7'b0;

   // m50_26 = W*in
   wire signed [6:0] m50_26;
   assign m50_26 ={ {2{in50[5]}} , in50[5:1] };

   // m50_27 = W*in
   wire signed [6:0] m50_27;
   assign m50_27 =7'b0;

   // m51_1 = W*in
   wire signed [6:0] m51_1;
   assign m51_1 =7'b0;

   // m51_2 = W*in
   wire signed [6:0] m51_2;
   assign m51_2 ={ {1{in51[5]}} , in51[5:0] };

   // m51_3 = W*in
   wire signed [6:0] m51_3;
   assign m51_3 =7'b0;

   // m51_4 = W*in
   wire signed [6:0] m51_4;
   assign m51_4 =7'b0;

   // m51_5 = W*in
   wire signed [6:0] m51_5;
   assign m51_5 =7'b0;

   // m51_6 = W*in
   wire signed [6:0] m51_6;
   assign m51_6 =7'b0;

   // m51_7 = W*in
   wire signed [6:0] m51_7;
   assign m51_7 =7'b0;

   // m51_8 = W*in
   wire signed [6:0] m51_8;
   assign m51_8 =7'b0;

   // m51_9 = W*in
   wire signed [6:0] m51_9;
   assign m51_9 =7'b0;

   // m51_10 = W*in
   wire signed [6:0] m51_10;
   assign m51_10 =7'b0;

   // m51_11 = W*in
   wire signed [6:0] m51_11;
   assign m51_11 ={ {2{in51[5]}} , in51[5:1] };

   // m51_12 = W*in
   wire signed [6:0] m51_12;
   assign m51_12 =7'b0;

   // m51_13 = W*in
   wire signed [6:0] m51_13;
   assign m51_13 =7'b0;

   // m51_14 = W*in
   wire signed [6:0] m51_14;
   assign m51_14 =7'b0;

   // m51_15 = W*in
   wire signed [6:0] m51_15;
   assign m51_15 =7'b0;

   // m51_16 = W*in
   wire signed [6:0] m51_16;
   assign m51_16 =7'b0;

   // m51_17 = W*in
   wire signed [6:0] m51_17;
   assign m51_17 =7'b0;

   // m51_18 = W*in
   wire signed [6:0] m51_18;
   assign m51_18 =7'b0;

   // m51_19 = W*in
   wire signed [6:0] m51_19;
   assign m51_19 =7'b0;

   // m51_20 = W*in
   wire signed [6:0] m51_20;
   assign m51_20 =7'b0;

   // m51_21 = W*in
   wire signed [6:0] m51_21;
   assign m51_21 =7'b0;

   // m51_22 = W*in
   wire signed [6:0] m51_22;
   assign m51_22 =7'b0;

   // m51_23 = W*in
   wire signed [6:0] m51_23;
   assign m51_23 =7'b0;

   // m51_24 = W*in
   wire signed [6:0] m51_24;
   assign m51_24 =7'b0;

   // m51_25 = W*in
   wire signed [6:0] m51_25;
   assign m51_25 =7'b0;

   // m51_26 = W*in
   wire signed [6:0] m51_26;
   assign m51_26 =7'b0;

   // m51_27 = W*in
   wire signed [6:0] m51_27;
   assign m51_27 =7'b0;

   // m52_1 = W*in
   wire signed [6:0] m52_1;
   assign m52_1 =7'b0;

   // m52_2 = W*in
   wire signed [6:0] m52_2;
   assign m52_2 =7'b0;

   // m52_3 = W*in
   wire signed [6:0] m52_3;
   assign m52_3 =7'b0;

   // m52_4 = W*in
   wire signed [6:0] m52_4;
   assign m52_4 =7'b0;

   // m52_5 = W*in
   wire signed [6:0] m52_5;
   assign m52_5 =7'b0;

   // m52_6 = W*in
   wire signed [6:0] m52_6;
   assign m52_6 =7'b0;

   // m52_7 = W*in
   wire signed [6:0] m52_7;
   assign m52_7 =7'b0;

   // m52_8 = W*in
   wire signed [6:0] m52_8;
   assign m52_8 =7'b0;

   // m52_9 = W*in
   wire signed [6:0] m52_9;
   assign m52_9 =7'b0;

   // m52_10 = W*in
   wire signed [6:0] m52_10;
   assign m52_10 =7'b0;

   // m52_11 = W*in
   wire signed [6:0] m52_11;
   assign m52_11 =7'b0;

   // m52_12 = W*in
   wire signed [6:0] m52_12;
   assign m52_12 =7'b0;

   // m52_13 = W*in
   wire signed [6:0] m52_13;
   assign m52_13 ={ {2{in52[5]}} , in52[5:1] };

   // m52_14 = W*in
   wire signed [6:0] m52_14;
   assign m52_14 =7'b0;

   // m52_15 = W*in
   wire signed [6:0] m52_15;
   assign m52_15 =7'b0;

   // m52_16 = W*in
   wire signed [6:0] m52_16;
   assign m52_16 =7'b0;

   // m52_17 = W*in
   wire signed [6:0] m52_17;
   assign m52_17 =7'b0;

   // m52_18 = W*in
   wire signed [6:0] m52_18;
   assign m52_18 =7'b0;

   // m52_19 = W*in
   wire signed [6:0] m52_19;
   assign m52_19 =7'b0;

   // m52_20 = W*in
   wire signed [6:0] m52_20;
   assign m52_20 =7'b0;

   // m52_21 = W*in
   wire signed [6:0] m52_21;
   assign m52_21 =7'b0;

   // m52_22 = W*in
   wire signed [6:0] m52_22;
   assign m52_22 =7'b0;

   // m52_23 = W*in
   wire signed [6:0] m52_23;
   assign m52_23 =7'b0;

   // m52_24 = W*in
   wire signed [6:0] m52_24;
   assign m52_24 =7'b0;

   // m52_25 = W*in
   wire signed [6:0] m52_25;
   assign m52_25 =7'b0;

   // m52_26 = W*in
   wire signed [6:0] m52_26;
   assign m52_26 =7'b0;

   // m52_27 = W*in
   wire signed [6:0] m52_27;
   assign m52_27 =7'b0;

   // m53_1 = W*in
   wire signed [6:0] m53_1;
   assign m53_1 =7'b0;

   // m53_2 = W*in
   wire signed [6:0] m53_2;
   assign m53_2 =7'b0;

   // m53_3 = W*in
   wire signed [6:0] m53_3;
   assign m53_3 =7'b0;

   // m53_4 = W*in
   wire signed [6:0] m53_4;
   assign m53_4 =7'b0;

   // m53_5 = W*in
   wire signed [6:0] m53_5;
   assign m53_5 =7'b0;

   // m53_6 = W*in
   wire signed [6:0] m53_6;
   assign m53_6 =7'b0;

   // m53_7 = W*in
   wire signed [6:0] m53_7;
   assign m53_7 =7'b0;

   // m53_8 = W*in
   wire signed [6:0] m53_8;
   assign m53_8 =7'b0;

   // m53_9 = W*in
   wire signed [6:0] m53_9;
   assign m53_9 =7'b0;

   // m53_10 = W*in
   wire signed [6:0] m53_10;
   assign m53_10 =7'b0;

   // m53_11 = W*in
   wire signed [6:0] m53_11;
   assign m53_11 =7'b0;

   // m53_12 = W*in
   wire signed [6:0] m53_12;
   assign m53_12 =7'b0;

   // m53_13 = W*in
   wire signed [6:0] m53_13;
   assign m53_13 =7'b0;

   // m53_14 = W*in
   wire signed [6:0] m53_14;
   assign m53_14 =7'b0;

   // m53_15 = W*in
   wire signed [6:0] m53_15;
   assign m53_15 =7'b0;

   // m53_16 = W*in
   wire signed [6:0] m53_16;
   assign m53_16 =7'b0;

   // m53_17 = W*in
   wire signed [6:0] m53_17;
   assign m53_17 =7'b0;

   // m53_18 = W*in
   wire signed [6:0] m53_18;
   assign m53_18 =7'b0;

   // m53_19 = W*in
   wire signed [6:0] m53_19;
   assign m53_19 =7'b0;

   // m53_20 = W*in
   wire signed [6:0] m53_20;
   assign m53_20 =7'b0;

   // m53_21 = W*in
   wire signed [6:0] m53_21;
   assign m53_21 =7'b0;

   // m53_22 = W*in
   wire signed [6:0] m53_22;
   assign m53_22 ={ {1{in53[5]}} , in53[5:0] };

   // m53_23 = W*in
   wire signed [6:0] m53_23;
   assign m53_23 =7'b0;

   // m53_24 = W*in
   wire signed [6:0] m53_24;
   assign m53_24 =7'b0;

   // m53_25 = W*in
   wire signed [6:0] m53_25;
   assign m53_25 =7'b0;

   // m53_26 = W*in
   wire signed [6:0] m53_26;
   assign m53_26 =7'b0;

   // m53_27 = W*in
   wire signed [6:0] m53_27;
   assign m53_27 =7'b0;

   // m54_1 = W*in
   wire signed [6:0] m54_1;
   assign m54_1 =7'b0;

   // m54_2 = W*in
   wire signed [6:0] m54_2;
   assign m54_2 =7'b0;

   // m54_3 = W*in
   wire signed [6:0] m54_3;
   assign m54_3 ={ {1{in54[5]}} , in54[5:0] };

   // m54_4 = W*in
   wire signed [6:0] m54_4;
   assign m54_4 =7'b0;

   // m54_5 = W*in
   wire signed [6:0] m54_5;
   assign m54_5 =7'b0;

   // m54_6 = W*in
   wire signed [6:0] m54_6;
   assign m54_6 =7'b0;

   // m54_7 = W*in
   wire signed [6:0] m54_7;
   assign m54_7 =7'b0;

   // m54_8 = W*in
   wire signed [6:0] m54_8;
   assign m54_8 =7'b0;

   // m54_9 = W*in
   wire signed [6:0] m54_9;
   assign m54_9 =7'b0;

   // m54_10 = W*in
   wire signed [6:0] m54_10;
   assign m54_10 =7'b0;

   // m54_11 = W*in
   wire signed [6:0] m54_11;
   assign m54_11 =7'b0;

   // m54_12 = W*in
   wire signed [6:0] m54_12;
   assign m54_12 =7'b0;

   // m54_13 = W*in
   wire signed [6:0] m54_13;
   assign m54_13 =7'b0;

   // m54_14 = W*in
   wire signed [6:0] m54_14;
   assign m54_14 =7'b0;

   // m54_15 = W*in
   wire signed [6:0] m54_15;
   assign m54_15 =7'b0;

   // m54_16 = W*in
   wire signed [6:0] m54_16;
   assign m54_16 =7'b0;

   // m54_17 = W*in
   wire signed [6:0] m54_17;
   assign m54_17 =7'b0;

   // m54_18 = W*in
   wire signed [6:0] m54_18;
   assign m54_18 =7'b0;

   // m54_19 = W*in
   wire signed [6:0] m54_19;
   assign m54_19 =7'b0;

   // m54_20 = W*in
   wire signed [6:0] m54_20;
   assign m54_20 =7'b0;

   // m54_21 = W*in
   wire signed [6:0] m54_21;
   assign m54_21 =7'b0;

   // m54_22 = W*in
   wire signed [6:0] m54_22;
   assign m54_22 =7'b0;

   // m54_23 = W*in
   wire signed [6:0] m54_23;
   assign m54_23 =7'b0;

   // m54_24 = W*in
   wire signed [6:0] m54_24;
   assign m54_24 =7'b0;

   // m54_25 = W*in
   wire signed [6:0] m54_25;
   assign m54_25 =7'b0;

   // m54_26 = W*in
   wire signed [6:0] m54_26;
   assign m54_26 =7'b0;

   // m54_27 = W*in
   wire signed [6:0] m54_27;
   assign m54_27 =7'b0;

   // m55_1 = W*in
   wire signed [6:0] m55_1;
   assign m55_1 =7'b0;

   // m55_2 = W*in
   wire signed [6:0] m55_2;
   assign m55_2 =7'b0;

   // m55_3 = W*in
   wire signed [6:0] m55_3;
   assign m55_3 =7'b0;

   // m55_4 = W*in
   wire signed [6:0] m55_4;
   assign m55_4 =7'b0;

   // m55_5 = W*in
   wire signed [6:0] m55_5;
   assign m55_5 =7'b0;

   // m55_6 = W*in
   wire signed [6:0] m55_6;
   assign m55_6 =7'b0;

   // m55_7 = W*in
   wire signed [6:0] m55_7;
   assign m55_7 =7'b0;

   // m55_8 = W*in
   wire signed [6:0] m55_8;
   assign m55_8 =7'b0;

   // m55_9 = W*in
   wire signed [6:0] m55_9;
   assign m55_9 =7'b0;

   // m55_10 = W*in
   wire signed [6:0] m55_10;
   assign m55_10 =7'b0;

   // m55_11 = W*in
   wire signed [6:0] m55_11;
   assign m55_11 =7'b0;

   // m55_12 = W*in
   wire signed [6:0] m55_12;
   assign m55_12 =7'b0;

   // m55_13 = W*in
   wire signed [6:0] m55_13;
   assign m55_13 =7'b0;

   // m55_14 = W*in
   wire signed [6:0] m55_14;
   assign m55_14 =7'b0;

   // m55_15 = W*in
   wire signed [6:0] m55_15;
   assign m55_15 =7'b0;

   // m55_16 = W*in
   wire signed [6:0] m55_16;
   assign m55_16 =7'b0;

   // m55_17 = W*in
   wire signed [6:0] m55_17;
   assign m55_17 ={ {2{in55[5]}} , in55[5:1] };

   // m55_18 = W*in
   wire signed [6:0] m55_18;
   assign m55_18 =7'b0;

   // m55_19 = W*in
   wire signed [6:0] m55_19;
   assign m55_19 ={ {1{in55[5]}} , in55[5:0] };

   // m55_20 = W*in
   wire signed [6:0] m55_20;
   assign m55_20 =7'b0;

   // m55_21 = W*in
   wire signed [6:0] m55_21;
   assign m55_21 =7'b0;

   // m55_22 = W*in
   wire signed [6:0] m55_22;
   assign m55_22 =7'b0;

   // m55_23 = W*in
   wire signed [6:0] m55_23;
   assign m55_23 =7'b0;

   // m55_24 = W*in
   wire signed [6:0] m55_24;
   assign m55_24 =7'b0;

   // m55_25 = W*in
   wire signed [6:0] m55_25;
   assign m55_25 =7'b0;

   // m55_26 = W*in
   wire signed [6:0] m55_26;
   assign m55_26 =7'b0;

   // m55_27 = W*in
   wire signed [6:0] m55_27;
   assign m55_27 =7'b0;

   // m56_1 = W*in
   wire signed [6:0] m56_1;
   assign m56_1 =7'b0;

   // m56_2 = W*in
   wire signed [6:0] m56_2;
   assign m56_2 =7'b0;

   // m56_3 = W*in
   wire signed [6:0] m56_3;
   assign m56_3 =7'b0;

   // m56_4 = W*in
   wire signed [6:0] m56_4;
   assign m56_4 =7'b0;

   // m56_5 = W*in
   wire signed [6:0] m56_5;
   assign m56_5 =7'b0;

   // m56_6 = W*in
   wire signed [6:0] m56_6;
   assign m56_6 =7'b0;

   // m56_7 = W*in
   wire signed [6:0] m56_7;
   assign m56_7 =7'b0;

   // m56_8 = W*in
   wire signed [6:0] m56_8;
   assign m56_8 =7'b0;

   // m56_9 = W*in
   wire signed [6:0] m56_9;
   assign m56_9 =7'b0;

   // m56_10 = W*in
   wire signed [6:0] m56_10;
   assign m56_10 =7'b0;

   // m56_11 = W*in
   wire signed [6:0] m56_11;
   assign m56_11 =7'b0;

   // m56_12 = W*in
   wire signed [6:0] m56_12;
   assign m56_12 =7'b0;

   // m56_13 = W*in
   wire signed [6:0] m56_13;
   assign m56_13 =7'b0;

   // m56_14 = W*in
   wire signed [6:0] m56_14;
   assign m56_14 =7'b0;

   // m56_15 = W*in
   wire signed [6:0] m56_15;
   assign m56_15 =7'b0;

   // m56_16 = W*in
   wire signed [6:0] m56_16;
   assign m56_16 =7'b0;

   // m56_17 = W*in
   wire signed [6:0] m56_17;
   assign m56_17 =7'b0;

   // m56_18 = W*in
   wire signed [6:0] m56_18;
   assign m56_18 ={ {1{in56[5]}} , in56[5:0] };

   // m56_19 = W*in
   wire signed [6:0] m56_19;
   assign m56_19 =7'b0;

   // m56_20 = W*in
   wire signed [6:0] m56_20;
   assign m56_20 =7'b0;

   // m56_21 = W*in
   wire signed [6:0] m56_21;
   assign m56_21 =7'b0;

   // m56_22 = W*in
   wire signed [6:0] m56_22;
   assign m56_22 =7'b0;

   // m56_23 = W*in
   wire signed [6:0] m56_23;
   assign m56_23 =7'b0;

   // m56_24 = W*in
   wire signed [6:0] m56_24;
   assign m56_24 =7'b0;

   // m56_25 = W*in
   wire signed [6:0] m56_25;
   assign m56_25 =7'b0;

   // m56_26 = W*in
   wire signed [6:0] m56_26;
   assign m56_26 =7'b0;

   // m56_27 = W*in
   wire signed [6:0] m56_27;
   assign m56_27 =7'b0;

   // m57_1 = W*in
   wire signed [6:0] m57_1;
   assign m57_1 =7'b0;

   // m57_2 = W*in
   wire signed [6:0] m57_2;
   assign m57_2 =7'b0;

   // m57_3 = W*in
   wire signed [6:0] m57_3;
   assign m57_3 =7'b0;

   // m57_4 = W*in
   wire signed [6:0] m57_4;
   assign m57_4 =7'b0;

   // m57_5 = W*in
   wire signed [6:0] m57_5;
   assign m57_5 =7'b0;

   // m57_6 = W*in
   wire signed [6:0] m57_6;
   assign m57_6 =7'b0;

   // m57_7 = W*in
   wire signed [6:0] m57_7;
   assign m57_7 =7'b0;

   // m57_8 = W*in
   wire signed [6:0] m57_8;
   assign m57_8 =7'b0;

   // m57_9 = W*in
   wire signed [6:0] m57_9;
   assign m57_9 =7'b0;

   // m57_10 = W*in
   wire signed [6:0] m57_10;
   assign m57_10 =7'b0;

   // m57_11 = W*in
   wire signed [6:0] m57_11;
   assign m57_11 =7'b0;

   // m57_12 = W*in
   wire signed [6:0] m57_12;
   assign m57_12 =7'b0;

   // m57_13 = W*in
   wire signed [6:0] m57_13;
   wire signed [7:0] tm57_13;
   assign tm57_13[0:0] = in57[0:0];
   assign tm57_13[7:1] = { {1{in57[5]}} , in57[5:0] } + { {2{in57[5]}} , in57[5:1] };
   assign m57_13 ={ {1{tm57_13[7]}} , tm57_13[7:2] };

   // m57_14 = W*in
   wire signed [6:0] m57_14;
   assign m57_14 =7'b0;

   // m57_15 = W*in
   wire signed [6:0] m57_15;
   assign m57_15 =7'b0;

   // m57_16 = W*in
   wire signed [6:0] m57_16;
   assign m57_16 ={ {1{in57[5]}} , in57[5:0] };

   // m57_17 = W*in
   wire signed [6:0] m57_17;
   assign m57_17 =7'b0;

   // m57_18 = W*in
   wire signed [6:0] m57_18;
   assign m57_18 =7'b0;

   // m57_19 = W*in
   wire signed [6:0] m57_19;
   assign m57_19 =7'b0;

   // m57_20 = W*in
   wire signed [6:0] m57_20;
   assign m57_20 =7'b0;

   // m57_21 = W*in
   wire signed [6:0] m57_21;
   assign m57_21 =7'b0;

   // m57_22 = W*in
   wire signed [6:0] m57_22;
   assign m57_22 =7'b0;

   // m57_23 = W*in
   wire signed [6:0] m57_23;
   assign m57_23 =7'b0;

   // m57_24 = W*in
   wire signed [6:0] m57_24;
   assign m57_24 =7'b0;

   // m57_25 = W*in
   wire signed [6:0] m57_25;
   assign m57_25 =7'b0;

   // m57_26 = W*in
   wire signed [6:0] m57_26;
   assign m57_26 =7'b0;

   // m57_27 = W*in
   wire signed [6:0] m57_27;
   assign m57_27 =7'b0;

   // m58_1 = W*in
   wire signed [6:0] m58_1;
   assign m58_1 =7'b0;

   // m58_2 = W*in
   wire signed [6:0] m58_2;
   assign m58_2 =7'b0;

   // m58_3 = W*in
   wire signed [6:0] m58_3;
   assign m58_3 =7'b0;

   // m58_4 = W*in
   wire signed [6:0] m58_4;
   assign m58_4 =7'b0;

   // m58_5 = W*in
   wire signed [6:0] m58_5;
   assign m58_5 =7'b0;

   // m58_6 = W*in
   wire signed [6:0] m58_6;
   assign m58_6 =7'b0;

   // m58_7 = W*in
   wire signed [6:0] m58_7;
   assign m58_7 =7'b0;

   // m58_8 = W*in
   wire signed [6:0] m58_8;
   assign m58_8 =7'b0;

   // m58_9 = W*in
   wire signed [6:0] m58_9;
   assign m58_9 =7'b0;

   // m58_10 = W*in
   wire signed [6:0] m58_10;
   assign m58_10 =7'b0;

   // m58_11 = W*in
   wire signed [6:0] m58_11;
   assign m58_11 =7'b0;

   // m58_12 = W*in
   wire signed [6:0] m58_12;
   assign m58_12 =7'b0;

   // m58_13 = W*in
   wire signed [6:0] m58_13;
   assign m58_13 =7'b0;

   // m58_14 = W*in
   wire signed [6:0] m58_14;
   assign m58_14 =7'b0;

   // m58_15 = W*in
   wire signed [6:0] m58_15;
   assign m58_15 =7'b0;

   // m58_16 = W*in
   wire signed [6:0] m58_16;
   assign m58_16 =7'b0;

   // m58_17 = W*in
   wire signed [6:0] m58_17;
   assign m58_17 =7'b0;

   // m58_18 = W*in
   wire signed [6:0] m58_18;
   assign m58_18 =7'b0;

   // m58_19 = W*in
   wire signed [6:0] m58_19;
   assign m58_19 ={ {2{neg58[5]}} , neg58[5:1] };

   // m58_20 = W*in
   wire signed [6:0] m58_20;
   assign m58_20 =7'b0;

   // m58_21 = W*in
   wire signed [6:0] m58_21;
   assign m58_21 =7'b0;

   // m58_22 = W*in
   wire signed [6:0] m58_22;
   assign m58_22 =7'b0;

   // m58_23 = W*in
   wire signed [6:0] m58_23;
   assign m58_23 =7'b0;

   // m58_24 = W*in
   wire signed [6:0] m58_24;
   assign m58_24 =7'b0;

   // m58_25 = W*in
   wire signed [6:0] m58_25;
   assign m58_25 =7'b0;

   // m58_26 = W*in
   wire signed [6:0] m58_26;
   assign m58_26 =7'b0;

   // m58_27 = W*in
   wire signed [6:0] m58_27;
   assign m58_27 =7'b0;

   // m59_1 = W*in
   wire signed [6:0] m59_1;
   assign m59_1 =7'b0;

   // m59_2 = W*in
   wire signed [6:0] m59_2;
   assign m59_2 =7'b0;

   // m59_3 = W*in
   wire signed [6:0] m59_3;
   assign m59_3 =7'b0;

   // m59_4 = W*in
   wire signed [6:0] m59_4;
   assign m59_4 =7'b0;

   // m59_5 = W*in
   wire signed [6:0] m59_5;
   assign m59_5 ={ {2{in59[5]}} , in59[5:1] };

   // m59_6 = W*in
   wire signed [6:0] m59_6;
   assign m59_6 =7'b0;

   // m59_7 = W*in
   wire signed [6:0] m59_7;
   assign m59_7 =7'b0;

   // m59_8 = W*in
   wire signed [6:0] m59_8;
   assign m59_8 =7'b0;

   // m59_9 = W*in
   wire signed [6:0] m59_9;
   assign m59_9 ={ {2{in59[5]}} , in59[5:1] };

   // m59_10 = W*in
   wire signed [6:0] m59_10;
   assign m59_10 =7'b0;

   // m59_11 = W*in
   wire signed [6:0] m59_11;
   assign m59_11 =7'b0;

   // m59_12 = W*in
   wire signed [6:0] m59_12;
   assign m59_12 =7'b0;

   // m59_13 = W*in
   wire signed [6:0] m59_13;
   assign m59_13 =7'b0;

   // m59_14 = W*in
   wire signed [6:0] m59_14;
   assign m59_14 =7'b0;

   // m59_15 = W*in
   wire signed [6:0] m59_15;
   assign m59_15 =7'b0;

   // m59_16 = W*in
   wire signed [6:0] m59_16;
   assign m59_16 =7'b0;

   // m59_17 = W*in
   wire signed [6:0] m59_17;
   assign m59_17 =7'b0;

   // m59_18 = W*in
   wire signed [6:0] m59_18;
   assign m59_18 =7'b0;

   // m59_19 = W*in
   wire signed [6:0] m59_19;
   assign m59_19 =7'b0;

   // m59_20 = W*in
   wire signed [6:0] m59_20;
   assign m59_20 =7'b0;

   // m59_21 = W*in
   wire signed [6:0] m59_21;
   assign m59_21 =7'b0;

   // m59_22 = W*in
   wire signed [6:0] m59_22;
   assign m59_22 =7'b0;

   // m59_23 = W*in
   wire signed [6:0] m59_23;
   assign m59_23 =7'b0;

   // m59_24 = W*in
   wire signed [6:0] m59_24;
   assign m59_24 =7'b0;

   // m59_25 = W*in
   wire signed [6:0] m59_25;
   assign m59_25 =7'b0;

   // m59_26 = W*in
   wire signed [6:0] m59_26;
   assign m59_26 =7'b0;

   // m59_27 = W*in
   wire signed [6:0] m59_27;
   assign m59_27 =7'b0;

   // m60_1 = W*in
   wire signed [6:0] m60_1;
   assign m60_1 =7'b0;

   // m60_2 = W*in
   wire signed [6:0] m60_2;
   assign m60_2 =7'b0;

   // m60_3 = W*in
   wire signed [6:0] m60_3;
   assign m60_3 =7'b0;

   // m60_4 = W*in
   wire signed [6:0] m60_4;
   assign m60_4 =7'b0;

   // m60_5 = W*in
   wire signed [6:0] m60_5;
   assign m60_5 =7'b0;

   // m60_6 = W*in
   wire signed [6:0] m60_6;
   assign m60_6 =7'b0;

   // m60_7 = W*in
   wire signed [6:0] m60_7;
   assign m60_7 =7'b0;

   // m60_8 = W*in
   wire signed [6:0] m60_8;
   assign m60_8 =7'b0;

   // m60_9 = W*in
   wire signed [6:0] m60_9;
   assign m60_9 ={ {2{in60[5]}} , in60[5:1] };

   // m60_10 = W*in
   wire signed [6:0] m60_10;
   assign m60_10 =7'b0;

   // m60_11 = W*in
   wire signed [6:0] m60_11;
   assign m60_11 =7'b0;

   // m60_12 = W*in
   wire signed [6:0] m60_12;
   assign m60_12 =7'b0;

   // m60_13 = W*in
   wire signed [6:0] m60_13;
   assign m60_13 =7'b0;

   // m60_14 = W*in
   wire signed [6:0] m60_14;
   assign m60_14 =7'b0;

   // m60_15 = W*in
   wire signed [6:0] m60_15;
   assign m60_15 =7'b0;

   // m60_16 = W*in
   wire signed [6:0] m60_16;
   assign m60_16 =7'b0;

   // m60_17 = W*in
   wire signed [6:0] m60_17;
   assign m60_17 =7'b0;

   // m60_18 = W*in
   wire signed [6:0] m60_18;
   assign m60_18 =7'b0;

   // m60_19 = W*in
   wire signed [6:0] m60_19;
   assign m60_19 =7'b0;

   // m60_20 = W*in
   wire signed [6:0] m60_20;
   assign m60_20 =7'b0;

   // m60_21 = W*in
   wire signed [6:0] m60_21;
   assign m60_21 =7'b0;

   // m60_22 = W*in
   wire signed [6:0] m60_22;
   assign m60_22 =7'b0;

   // m60_23 = W*in
   wire signed [6:0] m60_23;
   assign m60_23 =7'b0;

   // m60_24 = W*in
   wire signed [6:0] m60_24;
   assign m60_24 =7'b0;

   // m60_25 = W*in
   wire signed [6:0] m60_25;
   assign m60_25 =7'b0;

   // m60_26 = W*in
   wire signed [6:0] m60_26;
   assign m60_26 ={ {2{in60[5]}} , in60[5:1] };

   // m60_27 = W*in
   wire signed [6:0] m60_27;
   assign m60_27 =7'b0;

   // m61_1 = W*in
   wire signed [6:0] m61_1;
   assign m61_1 =7'b0;

   // m61_2 = W*in
   wire signed [6:0] m61_2;
   assign m61_2 =7'b0;

   // m61_3 = W*in
   wire signed [6:0] m61_3;
   assign m61_3 =7'b0;

   // m61_4 = W*in
   wire signed [6:0] m61_4;
   assign m61_4 =7'b0;

   // m61_5 = W*in
   wire signed [6:0] m61_5;
   assign m61_5 =7'b0;

   // m61_6 = W*in
   wire signed [6:0] m61_6;
   assign m61_6 =7'b0;

   // m61_7 = W*in
   wire signed [6:0] m61_7;
   assign m61_7 =7'b0;

   // m61_8 = W*in
   wire signed [6:0] m61_8;
   assign m61_8 =7'b0;

   // m61_9 = W*in
   wire signed [6:0] m61_9;
   assign m61_9 =7'b0;

   // m61_10 = W*in
   wire signed [6:0] m61_10;
   assign m61_10 =7'b0;

   // m61_11 = W*in
   wire signed [6:0] m61_11;
   assign m61_11 =7'b0;

   // m61_12 = W*in
   wire signed [6:0] m61_12;
   assign m61_12 =7'b0;

   // m61_13 = W*in
   wire signed [6:0] m61_13;
   assign m61_13 ={ {1{in61[5]}} , in61[5:0] };

   // m61_14 = W*in
   wire signed [6:0] m61_14;
   assign m61_14 =7'b0;

   // m61_15 = W*in
   wire signed [6:0] m61_15;
   assign m61_15 =7'b0;

   // m61_16 = W*in
   wire signed [6:0] m61_16;
   assign m61_16 =7'b0;

   // m61_17 = W*in
   wire signed [6:0] m61_17;
   assign m61_17 =7'b0;

   // m61_18 = W*in
   wire signed [6:0] m61_18;
   assign m61_18 =7'b0;

   // m61_19 = W*in
   wire signed [6:0] m61_19;
   assign m61_19 =7'b0;

   // m61_20 = W*in
   wire signed [6:0] m61_20;
   assign m61_20 =7'b0;

   // m61_21 = W*in
   wire signed [6:0] m61_21;
   assign m61_21 ={ {2{in61[5]}} , in61[5:1] };

   // m61_22 = W*in
   wire signed [6:0] m61_22;
   assign m61_22 =7'b0;

   // m61_23 = W*in
   wire signed [6:0] m61_23;
   assign m61_23 =7'b0;

   // m61_24 = W*in
   wire signed [6:0] m61_24;
   assign m61_24 =7'b0;

   // m61_25 = W*in
   wire signed [6:0] m61_25;
   assign m61_25 =7'b0;

   // m61_26 = W*in
   wire signed [6:0] m61_26;
   assign m61_26 =7'b0;

   // m61_27 = W*in
   wire signed [6:0] m61_27;
   assign m61_27 =7'b0;

   // m62_1 = W*in
   wire signed [6:0] m62_1;
   assign m62_1 =7'b0;

   // m62_2 = W*in
   wire signed [6:0] m62_2;
   assign m62_2 =7'b0;

   // m62_3 = W*in
   wire signed [6:0] m62_3;
   assign m62_3 =7'b0;

   // m62_4 = W*in
   wire signed [6:0] m62_4;
   assign m62_4 =7'b0;

   // m62_5 = W*in
   wire signed [6:0] m62_5;
   assign m62_5 =7'b0;

   // m62_6 = W*in
   wire signed [6:0] m62_6;
   assign m62_6 =7'b0;

   // m62_7 = W*in
   wire signed [6:0] m62_7;
   assign m62_7 =7'b0;

   // m62_8 = W*in
   wire signed [6:0] m62_8;
   assign m62_8 =7'b0;

   // m62_9 = W*in
   wire signed [6:0] m62_9;
   assign m62_9 =7'b0;

   // m62_10 = W*in
   wire signed [6:0] m62_10;
   assign m62_10 =7'b0;

   // m62_11 = W*in
   wire signed [6:0] m62_11;
   assign m62_11 =7'b0;

   // m62_12 = W*in
   wire signed [6:0] m62_12;
   assign m62_12 ={ {2{neg62[5]}} , neg62[5:1] };

   // m62_13 = W*in
   wire signed [6:0] m62_13;
   assign m62_13 =7'b0;

   // m62_14 = W*in
   wire signed [6:0] m62_14;
   assign m62_14 =7'b0;

   // m62_15 = W*in
   wire signed [6:0] m62_15;
   assign m62_15 =7'b0;

   // m62_16 = W*in
   wire signed [6:0] m62_16;
   assign m62_16 =7'b0;

   // m62_17 = W*in
   wire signed [6:0] m62_17;
   assign m62_17 =7'b0;

   // m62_18 = W*in
   wire signed [6:0] m62_18;
   assign m62_18 =7'b0;

   // m62_19 = W*in
   wire signed [6:0] m62_19;
   assign m62_19 =7'b0;

   // m62_20 = W*in
   wire signed [6:0] m62_20;
   assign m62_20 =7'b0;

   // m62_21 = W*in
   wire signed [6:0] m62_21;
   assign m62_21 =7'b0;

   // m62_22 = W*in
   wire signed [6:0] m62_22;
   assign m62_22 =7'b0;

   // m62_23 = W*in
   wire signed [6:0] m62_23;
   assign m62_23 =7'b0;

   // m62_24 = W*in
   wire signed [6:0] m62_24;
   assign m62_24 =7'b0;

   // m62_25 = W*in
   wire signed [6:0] m62_25;
   assign m62_25 =7'b0;

   // m62_26 = W*in
   wire signed [6:0] m62_26;
   assign m62_26 =7'b0;

   // m62_27 = W*in
   wire signed [6:0] m62_27;
   assign m62_27 ={ {2{in62[5]}} , in62[5:1] };

   // m63_1 = W*in
   wire signed [6:0] m63_1;
   assign m63_1 =7'b0;

   // m63_2 = W*in
   wire signed [6:0] m63_2;
   assign m63_2 =7'b0;

   // m63_3 = W*in
   wire signed [6:0] m63_3;
   assign m63_3 ={ {2{in63[5]}} , in63[5:1] };

   // m63_4 = W*in
   wire signed [6:0] m63_4;
   assign m63_4 =7'b0;

   // m63_5 = W*in
   wire signed [6:0] m63_5;
   assign m63_5 =7'b0;

   // m63_6 = W*in
   wire signed [6:0] m63_6;
   assign m63_6 =7'b0;

   // m63_7 = W*in
   wire signed [6:0] m63_7;
   assign m63_7 =7'b0;

   // m63_8 = W*in
   wire signed [6:0] m63_8;
   assign m63_8 =7'b0;

   // m63_9 = W*in
   wire signed [6:0] m63_9;
   assign m63_9 =7'b0;

   // m63_10 = W*in
   wire signed [6:0] m63_10;
   assign m63_10 =7'b0;

   // m63_11 = W*in
   wire signed [6:0] m63_11;
   assign m63_11 =7'b0;

   // m63_12 = W*in
   wire signed [6:0] m63_12;
   assign m63_12 =7'b0;

   // m63_13 = W*in
   wire signed [6:0] m63_13;
   assign m63_13 =7'b0;

   // m63_14 = W*in
   wire signed [6:0] m63_14;
   assign m63_14 =7'b0;

   // m63_15 = W*in
   wire signed [6:0] m63_15;
   assign m63_15 =7'b0;

   // m63_16 = W*in
   wire signed [6:0] m63_16;
   assign m63_16 =7'b0;

   // m63_17 = W*in
   wire signed [6:0] m63_17;
   assign m63_17 =7'b0;

   // m63_18 = W*in
   wire signed [6:0] m63_18;
   assign m63_18 ={ {1{in63[5]}} , in63[5:0] };

   // m63_19 = W*in
   wire signed [6:0] m63_19;
   assign m63_19 =7'b0;

   // m63_20 = W*in
   wire signed [6:0] m63_20;
   assign m63_20 =7'b0;

   // m63_21 = W*in
   wire signed [6:0] m63_21;
   assign m63_21 =7'b0;

   // m63_22 = W*in
   wire signed [6:0] m63_22;
   assign m63_22 =7'b0;

   // m63_23 = W*in
   wire signed [6:0] m63_23;
   assign m63_23 =7'b0;

   // m63_24 = W*in
   wire signed [6:0] m63_24;
   assign m63_24 =7'b0;

   // m63_25 = W*in
   wire signed [6:0] m63_25;
   assign m63_25 =7'b0;

   // m63_26 = W*in
   wire signed [6:0] m63_26;
   assign m63_26 =7'b0;

   // m63_27 = W*in
   wire signed [6:0] m63_27;
   assign m63_27 =7'b0;

   // m64_1 = W*in
   wire signed [6:0] m64_1;
   assign m64_1 =7'b0;

   // m64_2 = W*in
   wire signed [6:0] m64_2;
   assign m64_2 =7'b0;

   // m64_3 = W*in
   wire signed [6:0] m64_3;
   assign m64_3 =7'b0;

   // m64_4 = W*in
   wire signed [6:0] m64_4;
   assign m64_4 =7'b0;

   // m64_5 = W*in
   wire signed [6:0] m64_5;
   assign m64_5 =7'b0;

   // m64_6 = W*in
   wire signed [6:0] m64_6;
   assign m64_6 =7'b0;

   // m64_7 = W*in
   wire signed [6:0] m64_7;
   assign m64_7 =7'b0;

   // m64_8 = W*in
   wire signed [6:0] m64_8;
   assign m64_8 =7'b0;

   // m64_9 = W*in
   wire signed [6:0] m64_9;
   assign m64_9 =7'b0;

   // m64_10 = W*in
   wire signed [6:0] m64_10;
   assign m64_10 =7'b0;

   // m64_11 = W*in
   wire signed [6:0] m64_11;
   assign m64_11 =7'b0;

   // m64_12 = W*in
   wire signed [6:0] m64_12;
   assign m64_12 =7'b0;

   // m64_13 = W*in
   wire signed [6:0] m64_13;
   assign m64_13 ={ {2{in64[5]}} , in64[5:1] };

   // m64_14 = W*in
   wire signed [6:0] m64_14;
   assign m64_14 =7'b0;

   // m64_15 = W*in
   wire signed [6:0] m64_15;
   assign m64_15 =7'b0;

   // m64_16 = W*in
   wire signed [6:0] m64_16;
   assign m64_16 =7'b0;

   // m64_17 = W*in
   wire signed [6:0] m64_17;
   assign m64_17 =7'b0;

   // m64_18 = W*in
   wire signed [6:0] m64_18;
   assign m64_18 =7'b0;

   // m64_19 = W*in
   wire signed [6:0] m64_19;
   assign m64_19 =7'b0;

   // m64_20 = W*in
   wire signed [6:0] m64_20;
   assign m64_20 =7'b0;

   // m64_21 = W*in
   wire signed [6:0] m64_21;
   assign m64_21 =7'b0;

   // m64_22 = W*in
   wire signed [6:0] m64_22;
   assign m64_22 =7'b0;

   // m64_23 = W*in
   wire signed [6:0] m64_23;
   assign m64_23 =7'b0;

   // m64_24 = W*in
   wire signed [6:0] m64_24;
   assign m64_24 =7'b0;

   // m64_25 = W*in
   wire signed [6:0] m64_25;
   assign m64_25 =7'b0;

   // m64_26 = W*in
   wire signed [6:0] m64_26;
   assign m64_26 =7'b0;

   // m64_27 = W*in
   wire signed [6:0] m64_27;
   assign m64_27 =7'b0;

   // m65_1 = W*in
   wire signed [6:0] m65_1;
   assign m65_1 =7'b0;

   // m65_2 = W*in
   wire signed [6:0] m65_2;
   assign m65_2 =7'b0;

   // m65_3 = W*in
   wire signed [6:0] m65_3;
   assign m65_3 =7'b0;

   // m65_4 = W*in
   wire signed [6:0] m65_4;
   assign m65_4 =7'b0;

   // m65_5 = W*in
   wire signed [6:0] m65_5;
   assign m65_5 =7'b0;

   // m65_6 = W*in
   wire signed [6:0] m65_6;
   assign m65_6 ={ {2{in65[5]}} , in65[5:1] };

   // m65_7 = W*in
   wire signed [6:0] m65_7;
   assign m65_7 =7'b0;

   // m65_8 = W*in
   wire signed [6:0] m65_8;
   assign m65_8 =7'b0;

   // m65_9 = W*in
   wire signed [6:0] m65_9;
   assign m65_9 =7'b0;

   // m65_10 = W*in
   wire signed [6:0] m65_10;
   assign m65_10 =7'b0;

   // m65_11 = W*in
   wire signed [6:0] m65_11;
   assign m65_11 =7'b0;

   // m65_12 = W*in
   wire signed [6:0] m65_12;
   assign m65_12 =7'b0;

   // m65_13 = W*in
   wire signed [6:0] m65_13;
   assign m65_13 =7'b0;

   // m65_14 = W*in
   wire signed [6:0] m65_14;
   assign m65_14 =7'b0;

   // m65_15 = W*in
   wire signed [6:0] m65_15;
   assign m65_15 =7'b0;

   // m65_16 = W*in
   wire signed [6:0] m65_16;
   assign m65_16 =7'b0;

   // m65_17 = W*in
   wire signed [6:0] m65_17;
   assign m65_17 =7'b0;

   // m65_18 = W*in
   wire signed [6:0] m65_18;
   assign m65_18 =7'b0;

   // m65_19 = W*in
   wire signed [6:0] m65_19;
   assign m65_19 =7'b0;

   // m65_20 = W*in
   wire signed [6:0] m65_20;
   assign m65_20 =7'b0;

   // m65_21 = W*in
   wire signed [6:0] m65_21;
   assign m65_21 =7'b0;

   // m65_22 = W*in
   wire signed [6:0] m65_22;
   assign m65_22 =7'b0;

   // m65_23 = W*in
   wire signed [6:0] m65_23;
   assign m65_23 =7'b0;

   // m65_24 = W*in
   wire signed [6:0] m65_24;
   assign m65_24 =7'b0;

   // m65_25 = W*in
   wire signed [6:0] m65_25;
   assign m65_25 =7'b0;

   // m65_26 = W*in
   wire signed [6:0] m65_26;
   assign m65_26 =7'b0;

   // m65_27 = W*in
   wire signed [6:0] m65_27;
   assign m65_27 =7'b0;

   // m66_1 = W*in
   wire signed [6:0] m66_1;
   assign m66_1 =7'b0;

   // m66_2 = W*in
   wire signed [6:0] m66_2;
   assign m66_2 =7'b0;

   // m66_3 = W*in
   wire signed [6:0] m66_3;
   assign m66_3 =7'b0;

   // m66_4 = W*in
   wire signed [6:0] m66_4;
   assign m66_4 =7'b0;

   // m66_5 = W*in
   wire signed [6:0] m66_5;
   assign m66_5 =7'b0;

   // m66_6 = W*in
   wire signed [6:0] m66_6;
   assign m66_6 =7'b0;

   // m66_7 = W*in
   wire signed [6:0] m66_7;
   assign m66_7 =7'b0;

   // m66_8 = W*in
   wire signed [6:0] m66_8;
   assign m66_8 =7'b0;

   // m66_9 = W*in
   wire signed [6:0] m66_9;
   assign m66_9 =7'b0;

   // m66_10 = W*in
   wire signed [6:0] m66_10;
   assign m66_10 =7'b0;

   // m66_11 = W*in
   wire signed [6:0] m66_11;
   assign m66_11 =7'b0;

   // m66_12 = W*in
   wire signed [6:0] m66_12;
   assign m66_12 =7'b0;

   // m66_13 = W*in
   wire signed [6:0] m66_13;
   assign m66_13 =7'b0;

   // m66_14 = W*in
   wire signed [6:0] m66_14;
   assign m66_14 ={ {2{in66[5]}} , in66[5:1] };

   // m66_15 = W*in
   wire signed [6:0] m66_15;
   assign m66_15 =7'b0;

   // m66_16 = W*in
   wire signed [6:0] m66_16;
   assign m66_16 =7'b0;

   // m66_17 = W*in
   wire signed [6:0] m66_17;
   assign m66_17 ={ {2{in66[5]}} , in66[5:1] };

   // m66_18 = W*in
   wire signed [6:0] m66_18;
   assign m66_18 =7'b0;

   // m66_19 = W*in
   wire signed [6:0] m66_19;
   assign m66_19 =7'b0;

   // m66_20 = W*in
   wire signed [6:0] m66_20;
   assign m66_20 =7'b0;

   // m66_21 = W*in
   wire signed [6:0] m66_21;
   assign m66_21 =7'b0;

   // m66_22 = W*in
   wire signed [6:0] m66_22;
   assign m66_22 =7'b0;

   // m66_23 = W*in
   wire signed [6:0] m66_23;
   assign m66_23 ={ {2{in66[5]}} , in66[5:1] };

   // m66_24 = W*in
   wire signed [6:0] m66_24;
   assign m66_24 =7'b0;

   // m66_25 = W*in
   wire signed [6:0] m66_25;
   assign m66_25 =7'b0;

   // m66_26 = W*in
   wire signed [6:0] m66_26;
   assign m66_26 =7'b0;

   // m66_27 = W*in
   wire signed [6:0] m66_27;
   assign m66_27 =7'b0;

   // m67_1 = W*in
   wire signed [6:0] m67_1;
   assign m67_1 =7'b0;

   // m67_2 = W*in
   wire signed [6:0] m67_2;
   assign m67_2 =7'b0;

   // m67_3 = W*in
   wire signed [6:0] m67_3;
   assign m67_3 =7'b0;

   // m67_4 = W*in
   wire signed [6:0] m67_4;
   assign m67_4 =7'b0;

   // m67_5 = W*in
   wire signed [6:0] m67_5;
   assign m67_5 =7'b0;

   // m67_6 = W*in
   wire signed [6:0] m67_6;
   assign m67_6 =7'b0;

   // m67_7 = W*in
   wire signed [6:0] m67_7;
   assign m67_7 =7'b0;

   // m67_8 = W*in
   wire signed [6:0] m67_8;
   assign m67_8 =7'b0;

   // m67_9 = W*in
   wire signed [6:0] m67_9;
   assign m67_9 =7'b0;

   // m67_10 = W*in
   wire signed [6:0] m67_10;
   assign m67_10 =7'b0;

   // m67_11 = W*in
   wire signed [6:0] m67_11;
   assign m67_11 =7'b0;

   // m67_12 = W*in
   wire signed [6:0] m67_12;
   assign m67_12 =7'b0;

   // m67_13 = W*in
   wire signed [6:0] m67_13;
   assign m67_13 =7'b0;

   // m67_14 = W*in
   wire signed [6:0] m67_14;
   assign m67_14 =7'b0;

   // m67_15 = W*in
   wire signed [6:0] m67_15;
   assign m67_15 =7'b0;

   // m67_16 = W*in
   wire signed [6:0] m67_16;
   assign m67_16 =7'b0;

   // m67_17 = W*in
   wire signed [6:0] m67_17;
   assign m67_17 =7'b0;

   // m67_18 = W*in
   wire signed [6:0] m67_18;
   assign m67_18 =7'b0;

   // m67_19 = W*in
   wire signed [6:0] m67_19;
   assign m67_19 =7'b0;

   // m67_20 = W*in
   wire signed [6:0] m67_20;
   assign m67_20 =7'b0;

   // m67_21 = W*in
   wire signed [6:0] m67_21;
   assign m67_21 ={ {1{in67[5]}} , in67[5:0] };

   // m67_22 = W*in
   wire signed [6:0] m67_22;
   assign m67_22 =7'b0;

   // m67_23 = W*in
   wire signed [6:0] m67_23;
   assign m67_23 =7'b0;

   // m67_24 = W*in
   wire signed [6:0] m67_24;
   assign m67_24 =7'b0;

   // m67_25 = W*in
   wire signed [6:0] m67_25;
   assign m67_25 =7'b0;

   // m67_26 = W*in
   wire signed [6:0] m67_26;
   assign m67_26 =7'b0;

   // m67_27 = W*in
   wire signed [6:0] m67_27;
   assign m67_27 =7'b0;

   // m68_1 = W*in
   wire signed [6:0] m68_1;
   assign m68_1 =7'b0;

   // m68_2 = W*in
   wire signed [6:0] m68_2;
   assign m68_2 =7'b0;

   // m68_3 = W*in
   wire signed [6:0] m68_3;
   assign m68_3 =7'b0;

   // m68_4 = W*in
   wire signed [6:0] m68_4;
   assign m68_4 =7'b0;

   // m68_5 = W*in
   wire signed [6:0] m68_5;
   assign m68_5 =7'b0;

   // m68_6 = W*in
   wire signed [6:0] m68_6;
   assign m68_6 =7'b0;

   // m68_7 = W*in
   wire signed [6:0] m68_7;
   assign m68_7 =7'b0;

   // m68_8 = W*in
   wire signed [6:0] m68_8;
   assign m68_8 ={ {2{in68[5]}} , in68[5:1] };

   // m68_9 = W*in
   wire signed [6:0] m68_9;
   assign m68_9 =7'b0;

   // m68_10 = W*in
   wire signed [6:0] m68_10;
   assign m68_10 ={ {2{in68[5]}} , in68[5:1] };

   // m68_11 = W*in
   wire signed [6:0] m68_11;
   assign m68_11 =7'b0;

   // m68_12 = W*in
   wire signed [6:0] m68_12;
   assign m68_12 =7'b0;

   // m68_13 = W*in
   wire signed [6:0] m68_13;
   assign m68_13 =7'b0;

   // m68_14 = W*in
   wire signed [6:0] m68_14;
   assign m68_14 =7'b0;

   // m68_15 = W*in
   wire signed [6:0] m68_15;
   assign m68_15 =7'b0;

   // m68_16 = W*in
   wire signed [6:0] m68_16;
   assign m68_16 =7'b0;

   // m68_17 = W*in
   wire signed [6:0] m68_17;
   assign m68_17 =7'b0;

   // m68_18 = W*in
   wire signed [6:0] m68_18;
   assign m68_18 =7'b0;

   // m68_19 = W*in
   wire signed [6:0] m68_19;
   assign m68_19 =7'b0;

   // m68_20 = W*in
   wire signed [6:0] m68_20;
   assign m68_20 =7'b0;

   // m68_21 = W*in
   wire signed [6:0] m68_21;
   assign m68_21 =7'b0;

   // m68_22 = W*in
   wire signed [6:0] m68_22;
   assign m68_22 =7'b0;

   // m68_23 = W*in
   wire signed [6:0] m68_23;
   assign m68_23 =7'b0;

   // m68_24 = W*in
   wire signed [6:0] m68_24;
   assign m68_24 =7'b0;

   // m68_25 = W*in
   wire signed [6:0] m68_25;
   assign m68_25 =7'b0;

   // m68_26 = W*in
   wire signed [6:0] m68_26;
   assign m68_26 =7'b0;

   // m68_27 = W*in
   wire signed [6:0] m68_27;
   assign m68_27 =7'b0;

   // m69_1 = W*in
   wire signed [6:0] m69_1;
   assign m69_1 =7'b0;

   // m69_2 = W*in
   wire signed [6:0] m69_2;
   assign m69_2 =7'b0;

   // m69_3 = W*in
   wire signed [6:0] m69_3;
   assign m69_3 =7'b0;

   // m69_4 = W*in
   wire signed [6:0] m69_4;
   assign m69_4 =7'b0;

   // m69_5 = W*in
   wire signed [6:0] m69_5;
   assign m69_5 =7'b0;

   // m69_6 = W*in
   wire signed [6:0] m69_6;
   assign m69_6 =7'b0;

   // m69_7 = W*in
   wire signed [6:0] m69_7;
   assign m69_7 =7'b0;

   // m69_8 = W*in
   wire signed [6:0] m69_8;
   assign m69_8 =7'b0;

   // m69_9 = W*in
   wire signed [6:0] m69_9;
   assign m69_9 =7'b0;

   // m69_10 = W*in
   wire signed [6:0] m69_10;
   assign m69_10 =7'b0;

   // m69_11 = W*in
   wire signed [6:0] m69_11;
   assign m69_11 =7'b0;

   // m69_12 = W*in
   wire signed [6:0] m69_12;
   assign m69_12 =7'b0;

   // m69_13 = W*in
   wire signed [6:0] m69_13;
   assign m69_13 ={ {2{in69[5]}} , in69[5:1] };

   // m69_14 = W*in
   wire signed [6:0] m69_14;
   assign m69_14 =7'b0;

   // m69_15 = W*in
   wire signed [6:0] m69_15;
   assign m69_15 =7'b0;

   // m69_16 = W*in
   wire signed [6:0] m69_16;
   assign m69_16 =7'b0;

   // m69_17 = W*in
   wire signed [6:0] m69_17;
   assign m69_17 =7'b0;

   // m69_18 = W*in
   wire signed [6:0] m69_18;
   assign m69_18 =7'b0;

   // m69_19 = W*in
   wire signed [6:0] m69_19;
   assign m69_19 =7'b0;

   // m69_20 = W*in
   wire signed [6:0] m69_20;
   assign m69_20 =7'b0;

   // m69_21 = W*in
   wire signed [6:0] m69_21;
   assign m69_21 =7'b0;

   // m69_22 = W*in
   wire signed [6:0] m69_22;
   assign m69_22 =7'b0;

   // m69_23 = W*in
   wire signed [6:0] m69_23;
   assign m69_23 =7'b0;

   // m69_24 = W*in
   wire signed [6:0] m69_24;
   assign m69_24 =7'b0;

   // m69_25 = W*in
   wire signed [6:0] m69_25;
   assign m69_25 =7'b0;

   // m69_26 = W*in
   wire signed [6:0] m69_26;
   assign m69_26 =7'b0;

   // m69_27 = W*in
   wire signed [6:0] m69_27;
   assign m69_27 ={ {1{neg69[5]}} , neg69[5:0] };

   // m70_1 = W*in
   wire signed [6:0] m70_1;
   assign m70_1 =7'b0;

   // m70_2 = W*in
   wire signed [6:0] m70_2;
   assign m70_2 ={ {1{neg70[5]}} , neg70[5:0] };

   // m70_3 = W*in
   wire signed [6:0] m70_3;
   assign m70_3 =7'b0;

   // m70_4 = W*in
   wire signed [6:0] m70_4;
   assign m70_4 =7'b0;

   // m70_5 = W*in
   wire signed [6:0] m70_5;
   assign m70_5 =7'b0;

   // m70_6 = W*in
   wire signed [6:0] m70_6;
   assign m70_6 =7'b0;

   // m70_7 = W*in
   wire signed [6:0] m70_7;
   assign m70_7 =7'b0;

   // m70_8 = W*in
   wire signed [6:0] m70_8;
   assign m70_8 =7'b0;

   // m70_9 = W*in
   wire signed [6:0] m70_9;
   assign m70_9 ={ {2{in70[5]}} , in70[5:1] };

   // m70_10 = W*in
   wire signed [6:0] m70_10;
   assign m70_10 =7'b0;

   // m70_11 = W*in
   wire signed [6:0] m70_11;
   assign m70_11 =7'b0;

   // m70_12 = W*in
   wire signed [6:0] m70_12;
   assign m70_12 =7'b0;

   // m70_13 = W*in
   wire signed [6:0] m70_13;
   assign m70_13 =7'b0;

   // m70_14 = W*in
   wire signed [6:0] m70_14;
   assign m70_14 =7'b0;

   // m70_15 = W*in
   wire signed [6:0] m70_15;
   assign m70_15 =7'b0;

   // m70_16 = W*in
   wire signed [6:0] m70_16;
   assign m70_16 =7'b0;

   // m70_17 = W*in
   wire signed [6:0] m70_17;
   assign m70_17 =7'b0;

   // m70_18 = W*in
   wire signed [6:0] m70_18;
   assign m70_18 =7'b0;

   // m70_19 = W*in
   wire signed [6:0] m70_19;
   assign m70_19 =7'b0;

   // m70_20 = W*in
   wire signed [6:0] m70_20;
   assign m70_20 =7'b0;

   // m70_21 = W*in
   wire signed [6:0] m70_21;
   assign m70_21 =7'b0;

   // m70_22 = W*in
   wire signed [6:0] m70_22;
   assign m70_22 =7'b0;

   // m70_23 = W*in
   wire signed [6:0] m70_23;
   assign m70_23 =7'b0;

   // m70_24 = W*in
   wire signed [6:0] m70_24;
   assign m70_24 =7'b0;

   // m70_25 = W*in
   wire signed [6:0] m70_25;
   assign m70_25 =7'b0;

   // m70_26 = W*in
   wire signed [6:0] m70_26;
   assign m70_26 =7'b0;

   // m70_27 = W*in
   wire signed [6:0] m70_27;
   assign m70_27 =7'b0;

   // m71_1 = W*in
   wire signed [6:0] m71_1;
   assign m71_1 =7'b0;

   // m71_2 = W*in
   wire signed [6:0] m71_2;
   assign m71_2 =7'b0;

   // m71_3 = W*in
   wire signed [6:0] m71_3;
   assign m71_3 =7'b0;

   // m71_4 = W*in
   wire signed [6:0] m71_4;
   assign m71_4 =7'b0;

   // m71_5 = W*in
   wire signed [6:0] m71_5;
   assign m71_5 =7'b0;

   // m71_6 = W*in
   wire signed [6:0] m71_6;
   assign m71_6 =7'b0;

   // m71_7 = W*in
   wire signed [6:0] m71_7;
   assign m71_7 =7'b0;

   // m71_8 = W*in
   wire signed [6:0] m71_8;
   assign m71_8 =7'b0;

   // m71_9 = W*in
   wire signed [6:0] m71_9;
   assign m71_9 =7'b0;

   // m71_10 = W*in
   wire signed [6:0] m71_10;
   assign m71_10 =7'b0;

   // m71_11 = W*in
   wire signed [6:0] m71_11;
   assign m71_11 =7'b0;

   // m71_12 = W*in
   wire signed [6:0] m71_12;
   assign m71_12 ={ {2{in71[5]}} , in71[5:1] };

   // m71_13 = W*in
   wire signed [6:0] m71_13;
   assign m71_13 =7'b0;

   // m71_14 = W*in
   wire signed [6:0] m71_14;
   assign m71_14 =7'b0;

   // m71_15 = W*in
   wire signed [6:0] m71_15;
   assign m71_15 =7'b0;

   // m71_16 = W*in
   wire signed [6:0] m71_16;
   assign m71_16 =7'b0;

   // m71_17 = W*in
   wire signed [6:0] m71_17;
   assign m71_17 =7'b0;

   // m71_18 = W*in
   wire signed [6:0] m71_18;
   assign m71_18 =7'b0;

   // m71_19 = W*in
   wire signed [6:0] m71_19;
   assign m71_19 =7'b0;

   // m71_20 = W*in
   wire signed [6:0] m71_20;
   assign m71_20 =7'b0;

   // m71_21 = W*in
   wire signed [6:0] m71_21;
   assign m71_21 =7'b0;

   // m71_22 = W*in
   wire signed [6:0] m71_22;
   assign m71_22 =7'b0;

   // m71_23 = W*in
   wire signed [6:0] m71_23;
   assign m71_23 =7'b0;

   // m71_24 = W*in
   wire signed [6:0] m71_24;
   assign m71_24 =7'b0;

   // m71_25 = W*in
   wire signed [6:0] m71_25;
   assign m71_25 =7'b0;

   // m71_26 = W*in
   wire signed [6:0] m71_26;
   assign m71_26 =7'b0;

   // m71_27 = W*in
   wire signed [6:0] m71_27;
   assign m71_27 =7'b0;

   // m72_1 = W*in
   wire signed [6:0] m72_1;
   assign m72_1 =7'b0;

   // m72_2 = W*in
   wire signed [6:0] m72_2;
   assign m72_2 =7'b0;

   // m72_3 = W*in
   wire signed [6:0] m72_3;
   assign m72_3 =7'b0;

   // m72_4 = W*in
   wire signed [6:0] m72_4;
   assign m72_4 =7'b0;

   // m72_5 = W*in
   wire signed [6:0] m72_5;
   assign m72_5 ={ {2{in72[5]}} , in72[5:1] };

   // m72_6 = W*in
   wire signed [6:0] m72_6;
   assign m72_6 =7'b0;

   // m72_7 = W*in
   wire signed [6:0] m72_7;
   assign m72_7 =7'b0;

   // m72_8 = W*in
   wire signed [6:0] m72_8;
   assign m72_8 =7'b0;

   // m72_9 = W*in
   wire signed [6:0] m72_9;
   assign m72_9 ={ {2{in72[5]}} , in72[5:1] };

   // m72_10 = W*in
   wire signed [6:0] m72_10;
   assign m72_10 =7'b0;

   // m72_11 = W*in
   wire signed [6:0] m72_11;
   assign m72_11 =7'b0;

   // m72_12 = W*in
   wire signed [6:0] m72_12;
   assign m72_12 =7'b0;

   // m72_13 = W*in
   wire signed [6:0] m72_13;
   assign m72_13 =7'b0;

   // m72_14 = W*in
   wire signed [6:0] m72_14;
   assign m72_14 =7'b0;

   // m72_15 = W*in
   wire signed [6:0] m72_15;
   assign m72_15 =7'b0;

   // m72_16 = W*in
   wire signed [6:0] m72_16;
   assign m72_16 =7'b0;

   // m72_17 = W*in
   wire signed [6:0] m72_17;
   assign m72_17 =7'b0;

   // m72_18 = W*in
   wire signed [6:0] m72_18;
   assign m72_18 =7'b0;

   // m72_19 = W*in
   wire signed [6:0] m72_19;
   assign m72_19 =7'b0;

   // m72_20 = W*in
   wire signed [6:0] m72_20;
   assign m72_20 =7'b0;

   // m72_21 = W*in
   wire signed [6:0] m72_21;
   assign m72_21 =7'b0;

   // m72_22 = W*in
   wire signed [6:0] m72_22;
   assign m72_22 =7'b0;

   // m72_23 = W*in
   wire signed [6:0] m72_23;
   assign m72_23 ={ {1{in72[5]}} , in72[5:0] };

   // m72_24 = W*in
   wire signed [6:0] m72_24;
   assign m72_24 =7'b0;

   // m72_25 = W*in
   wire signed [6:0] m72_25;
   assign m72_25 =7'b0;

   // m72_26 = W*in
   wire signed [6:0] m72_26;
   assign m72_26 =7'b0;

   // m72_27 = W*in
   wire signed [6:0] m72_27;
   assign m72_27 =7'b0;

   // m73_1 = W*in
   wire signed [6:0] m73_1;
   wire signed [7:0] tm73_1;
   assign tm73_1[0:0] = in73[0:0];
   assign tm73_1[7:1] = { {1{in73[5]}} , in73[5:0] } + { {2{in73[5]}} , in73[5:1] };
   assign m73_1 ={ {1{tm73_1[7]}} , tm73_1[7:2] };

   // m73_2 = W*in
   wire signed [6:0] m73_2;
   assign m73_2 =7'b0;

   // m73_3 = W*in
   wire signed [6:0] m73_3;
   assign m73_3 =7'b0;

   // m73_4 = W*in
   wire signed [6:0] m73_4;
   assign m73_4 =7'b0;

   // m73_5 = W*in
   wire signed [6:0] m73_5;
   assign m73_5 =7'b0;

   // m73_6 = W*in
   wire signed [6:0] m73_6;
   assign m73_6 =7'b0;

   // m73_7 = W*in
   wire signed [6:0] m73_7;
   assign m73_7 =7'b0;

   // m73_8 = W*in
   wire signed [6:0] m73_8;
   assign m73_8 =7'b0;

   // m73_9 = W*in
   wire signed [6:0] m73_9;
   assign m73_9 =7'b0;

   // m73_10 = W*in
   wire signed [6:0] m73_10;
   assign m73_10 =7'b0;

   // m73_11 = W*in
   wire signed [6:0] m73_11;
   assign m73_11 =7'b0;

   // m73_12 = W*in
   wire signed [6:0] m73_12;
   assign m73_12 =7'b0;

   // m73_13 = W*in
   wire signed [6:0] m73_13;
   assign m73_13 =7'b0;

   // m73_14 = W*in
   wire signed [6:0] m73_14;
   assign m73_14 =7'b0;

   // m73_15 = W*in
   wire signed [6:0] m73_15;
   assign m73_15 =7'b0;

   // m73_16 = W*in
   wire signed [6:0] m73_16;
   assign m73_16 =7'b0;

   // m73_17 = W*in
   wire signed [6:0] m73_17;
   assign m73_17 =7'b0;

   // m73_18 = W*in
   wire signed [6:0] m73_18;
   assign m73_18 =7'b0;

   // m73_19 = W*in
   wire signed [6:0] m73_19;
   assign m73_19 =7'b0;

   // m73_20 = W*in
   wire signed [6:0] m73_20;
   assign m73_20 =7'b0;

   // m73_21 = W*in
   wire signed [6:0] m73_21;
   assign m73_21 =7'b0;

   // m73_22 = W*in
   wire signed [6:0] m73_22;
   assign m73_22 =7'b0;

   // m73_23 = W*in
   wire signed [6:0] m73_23;
   assign m73_23 =7'b0;

   // m73_24 = W*in
   wire signed [6:0] m73_24;
   assign m73_24 =7'b0;

   // m73_25 = W*in
   wire signed [6:0] m73_25;
   assign m73_25 =7'b0;

   // m73_26 = W*in
   wire signed [6:0] m73_26;
   assign m73_26 =7'b0;

   // m73_27 = W*in
   wire signed [6:0] m73_27;
   assign m73_27 =7'b0;

   // m74_1 = W*in
   wire signed [6:0] m74_1;
   assign m74_1 =7'b0;

   // m74_2 = W*in
   wire signed [6:0] m74_2;
   assign m74_2 =7'b0;

   // m74_3 = W*in
   wire signed [6:0] m74_3;
   assign m74_3 =7'b0;

   // m74_4 = W*in
   wire signed [6:0] m74_4;
   assign m74_4 =7'b0;

   // m74_5 = W*in
   wire signed [6:0] m74_5;
   assign m74_5 ={ {2{in74[5]}} , in74[5:1] };

   // m74_6 = W*in
   wire signed [6:0] m74_6;
   assign m74_6 =7'b0;

   // m74_7 = W*in
   wire signed [6:0] m74_7;
   assign m74_7 =7'b0;

   // m74_8 = W*in
   wire signed [6:0] m74_8;
   assign m74_8 =7'b0;

   // m74_9 = W*in
   wire signed [6:0] m74_9;
   assign m74_9 =7'b0;

   // m74_10 = W*in
   wire signed [6:0] m74_10;
   assign m74_10 =7'b0;

   // m74_11 = W*in
   wire signed [6:0] m74_11;
   assign m74_11 =7'b0;

   // m74_12 = W*in
   wire signed [6:0] m74_12;
   assign m74_12 =7'b0;

   // m74_13 = W*in
   wire signed [6:0] m74_13;
   assign m74_13 =7'b0;

   // m74_14 = W*in
   wire signed [6:0] m74_14;
   assign m74_14 =7'b0;

   // m74_15 = W*in
   wire signed [6:0] m74_15;
   assign m74_15 =7'b0;

   // m74_16 = W*in
   wire signed [6:0] m74_16;
   assign m74_16 =7'b0;

   // m74_17 = W*in
   wire signed [6:0] m74_17;
   assign m74_17 =7'b0;

   // m74_18 = W*in
   wire signed [6:0] m74_18;
   assign m74_18 =7'b0;

   // m74_19 = W*in
   wire signed [6:0] m74_19;
   assign m74_19 ={ {2{neg74[5]}} , neg74[5:1] };

   // m74_20 = W*in
   wire signed [6:0] m74_20;
   assign m74_20 =7'b0;

   // m74_21 = W*in
   wire signed [6:0] m74_21;
   assign m74_21 =7'b0;

   // m74_22 = W*in
   wire signed [6:0] m74_22;
   assign m74_22 =7'b0;

   // m74_23 = W*in
   wire signed [6:0] m74_23;
   assign m74_23 =7'b0;

   // m74_24 = W*in
   wire signed [6:0] m74_24;
   assign m74_24 =7'b0;

   // m74_25 = W*in
   wire signed [6:0] m74_25;
   assign m74_25 =7'b0;

   // m74_26 = W*in
   wire signed [6:0] m74_26;
   assign m74_26 ={ {2{in74[5]}} , in74[5:1] };

   // m74_27 = W*in
   wire signed [6:0] m74_27;
   assign m74_27 =7'b0;

   // m75_1 = W*in
   wire signed [6:0] m75_1;
   assign m75_1 =7'b0;

   // m75_2 = W*in
   wire signed [6:0] m75_2;
   assign m75_2 =7'b0;

   // m75_3 = W*in
   wire signed [6:0] m75_3;
   assign m75_3 =7'b0;

   // m75_4 = W*in
   wire signed [6:0] m75_4;
   assign m75_4 =7'b0;

   // m75_5 = W*in
   wire signed [6:0] m75_5;
   assign m75_5 =7'b0;

   // m75_6 = W*in
   wire signed [6:0] m75_6;
   assign m75_6 =7'b0;

   // m75_7 = W*in
   wire signed [6:0] m75_7;
   assign m75_7 =7'b0;

   // m75_8 = W*in
   wire signed [6:0] m75_8;
   assign m75_8 =7'b0;

   // m75_9 = W*in
   wire signed [6:0] m75_9;
   assign m75_9 =7'b0;

   // m75_10 = W*in
   wire signed [6:0] m75_10;
   assign m75_10 =7'b0;

   // m75_11 = W*in
   wire signed [6:0] m75_11;
   assign m75_11 =7'b0;

   // m75_12 = W*in
   wire signed [6:0] m75_12;
   assign m75_12 =7'b0;

   // m75_13 = W*in
   wire signed [6:0] m75_13;
   assign m75_13 =7'b0;

   // m75_14 = W*in
   wire signed [6:0] m75_14;
   assign m75_14 =7'b0;

   // m75_15 = W*in
   wire signed [6:0] m75_15;
   assign m75_15 =7'b0;

   // m75_16 = W*in
   wire signed [6:0] m75_16;
   assign m75_16 =7'b0;

   // m75_17 = W*in
   wire signed [6:0] m75_17;
   assign m75_17 =7'b0;

   // m75_18 = W*in
   wire signed [6:0] m75_18;
   assign m75_18 =7'b0;

   // m75_19 = W*in
   wire signed [6:0] m75_19;
   assign m75_19 =7'b0;

   // m75_20 = W*in
   wire signed [6:0] m75_20;
   assign m75_20 =7'b0;

   // m75_21 = W*in
   wire signed [6:0] m75_21;
   assign m75_21 =7'b0;

   // m75_22 = W*in
   wire signed [6:0] m75_22;
   assign m75_22 =7'b0;

   // m75_23 = W*in
   wire signed [6:0] m75_23;
   assign m75_23 =7'b0;

   // m75_24 = W*in
   wire signed [6:0] m75_24;
   assign m75_24 =7'b0;

   // m75_25 = W*in
   wire signed [6:0] m75_25;
   assign m75_25 ={ {1{in75[5]}} , in75[5:0] };

   // m75_26 = W*in
   wire signed [6:0] m75_26;
   assign m75_26 =7'b0;

   // m75_27 = W*in
   wire signed [6:0] m75_27;
   assign m75_27 =7'b0;

   // m76_1 = W*in
   wire signed [6:0] m76_1;
   assign m76_1 =7'b0;

   // m76_2 = W*in
   wire signed [6:0] m76_2;
   assign m76_2 =7'b0;

   // m76_3 = W*in
   wire signed [6:0] m76_3;
   assign m76_3 =7'b0;

   // m76_4 = W*in
   wire signed [6:0] m76_4;
   assign m76_4 =7'b0;

   // m76_5 = W*in
   wire signed [6:0] m76_5;
   assign m76_5 =7'b0;

   // m76_6 = W*in
   wire signed [6:0] m76_6;
   assign m76_6 =7'b0;

   // m76_7 = W*in
   wire signed [6:0] m76_7;
   assign m76_7 =7'b0;

   // m76_8 = W*in
   wire signed [6:0] m76_8;
   assign m76_8 =7'b0;

   // m76_9 = W*in
   wire signed [6:0] m76_9;
   assign m76_9 =7'b0;

   // m76_10 = W*in
   wire signed [6:0] m76_10;
   assign m76_10 =7'b0;

   // m76_11 = W*in
   wire signed [6:0] m76_11;
   assign m76_11 =7'b0;

   // m76_12 = W*in
   wire signed [6:0] m76_12;
   assign m76_12 =7'b0;

   // m76_13 = W*in
   wire signed [6:0] m76_13;
   assign m76_13 =7'b0;

   // m76_14 = W*in
   wire signed [6:0] m76_14;
   assign m76_14 =7'b0;

   // m76_15 = W*in
   wire signed [6:0] m76_15;
   assign m76_15 =7'b0;

   // m76_16 = W*in
   wire signed [6:0] m76_16;
   assign m76_16 =7'b0;

   // m76_17 = W*in
   wire signed [6:0] m76_17;
   assign m76_17 ={ {2{in76[5]}} , in76[5:1] };

   // m76_18 = W*in
   wire signed [6:0] m76_18;
   assign m76_18 =7'b0;

   // m76_19 = W*in
   wire signed [6:0] m76_19;
   assign m76_19 =7'b0;

   // m76_20 = W*in
   wire signed [6:0] m76_20;
   assign m76_20 =7'b0;

   // m76_21 = W*in
   wire signed [6:0] m76_21;
   assign m76_21 =7'b0;

   // m76_22 = W*in
   wire signed [6:0] m76_22;
   assign m76_22 ={ {2{in76[5]}} , in76[5:1] };

   // m76_23 = W*in
   wire signed [6:0] m76_23;
   assign m76_23 =7'b0;

   // m76_24 = W*in
   wire signed [6:0] m76_24;
   assign m76_24 =7'b0;

   // m76_25 = W*in
   wire signed [6:0] m76_25;
   assign m76_25 =7'b0;

   // m76_26 = W*in
   wire signed [6:0] m76_26;
   assign m76_26 =7'b0;

   // m76_27 = W*in
   wire signed [6:0] m76_27;
   assign m76_27 =7'b0;

   // m77_1 = W*in
   wire signed [6:0] m77_1;
   assign m77_1 =7'b0;

   // m77_2 = W*in
   wire signed [6:0] m77_2;
   assign m77_2 =7'b0;

   // m77_3 = W*in
   wire signed [6:0] m77_3;
   assign m77_3 =7'b0;

   // m77_4 = W*in
   wire signed [6:0] m77_4;
   assign m77_4 =7'b0;

   // m77_5 = W*in
   wire signed [6:0] m77_5;
   assign m77_5 =7'b0;

   // m77_6 = W*in
   wire signed [6:0] m77_6;
   assign m77_6 =7'b0;

   // m77_7 = W*in
   wire signed [6:0] m77_7;
   assign m77_7 =7'b0;

   // m77_8 = W*in
   wire signed [6:0] m77_8;
   assign m77_8 =7'b0;

   // m77_9 = W*in
   wire signed [6:0] m77_9;
   assign m77_9 =7'b0;

   // m77_10 = W*in
   wire signed [6:0] m77_10;
   assign m77_10 =7'b0;

   // m77_11 = W*in
   wire signed [6:0] m77_11;
   assign m77_11 ={ {2{in77[5]}} , in77[5:1] };

   // m77_12 = W*in
   wire signed [6:0] m77_12;
   assign m77_12 ={ {2{in77[5]}} , in77[5:1] };

   // m77_13 = W*in
   wire signed [6:0] m77_13;
   assign m77_13 =7'b0;

   // m77_14 = W*in
   wire signed [6:0] m77_14;
   assign m77_14 =7'b0;

   // m77_15 = W*in
   wire signed [6:0] m77_15;
   assign m77_15 ={ {2{in77[5]}} , in77[5:1] };

   // m77_16 = W*in
   wire signed [6:0] m77_16;
   assign m77_16 =7'b0;

   // m77_17 = W*in
   wire signed [6:0] m77_17;
   assign m77_17 =7'b0;

   // m77_18 = W*in
   wire signed [6:0] m77_18;
   assign m77_18 =7'b0;

   // m77_19 = W*in
   wire signed [6:0] m77_19;
   assign m77_19 =7'b0;

   // m77_20 = W*in
   wire signed [6:0] m77_20;
   assign m77_20 =7'b0;

   // m77_21 = W*in
   wire signed [6:0] m77_21;
   assign m77_21 =7'b0;

   // m77_22 = W*in
   wire signed [6:0] m77_22;
   assign m77_22 =7'b0;

   // m77_23 = W*in
   wire signed [6:0] m77_23;
   assign m77_23 =7'b0;

   // m77_24 = W*in
   wire signed [6:0] m77_24;
   assign m77_24 =7'b0;

   // m77_25 = W*in
   wire signed [6:0] m77_25;
   assign m77_25 =7'b0;

   // m77_26 = W*in
   wire signed [6:0] m77_26;
   assign m77_26 =7'b0;

   // m77_27 = W*in
   wire signed [6:0] m77_27;
   assign m77_27 =7'b0;

   // m78_1 = W*in
   wire signed [6:0] m78_1;
   assign m78_1 =7'b0;

   // m78_2 = W*in
   wire signed [6:0] m78_2;
   assign m78_2 =7'b0;

   // m78_3 = W*in
   wire signed [6:0] m78_3;
   assign m78_3 =7'b0;

   // m78_4 = W*in
   wire signed [6:0] m78_4;
   assign m78_4 =7'b0;

   // m78_5 = W*in
   wire signed [6:0] m78_5;
   assign m78_5 =7'b0;

   // m78_6 = W*in
   wire signed [6:0] m78_6;
   assign m78_6 =7'b0;

   // m78_7 = W*in
   wire signed [6:0] m78_7;
   assign m78_7 ={ {2{neg78[5]}} , neg78[5:1] };

   // m78_8 = W*in
   wire signed [6:0] m78_8;
   assign m78_8 =7'b0;

   // m78_9 = W*in
   wire signed [6:0] m78_9;
   assign m78_9 =7'b0;

   // m78_10 = W*in
   wire signed [6:0] m78_10;
   assign m78_10 =7'b0;

   // m78_11 = W*in
   wire signed [6:0] m78_11;
   assign m78_11 =7'b0;

   // m78_12 = W*in
   wire signed [6:0] m78_12;
   assign m78_12 ={ {2{in78[5]}} , in78[5:1] };

   // m78_13 = W*in
   wire signed [6:0] m78_13;
   assign m78_13 =7'b0;

   // m78_14 = W*in
   wire signed [6:0] m78_14;
   assign m78_14 =7'b0;

   // m78_15 = W*in
   wire signed [6:0] m78_15;
   assign m78_15 =7'b0;

   // m78_16 = W*in
   wire signed [6:0] m78_16;
   assign m78_16 =7'b0;

   // m78_17 = W*in
   wire signed [6:0] m78_17;
   assign m78_17 =7'b0;

   // m78_18 = W*in
   wire signed [6:0] m78_18;
   assign m78_18 =7'b0;

   // m78_19 = W*in
   wire signed [6:0] m78_19;
   assign m78_19 =7'b0;

   // m78_20 = W*in
   wire signed [6:0] m78_20;
   assign m78_20 =7'b0;

   // m78_21 = W*in
   wire signed [6:0] m78_21;
   assign m78_21 =7'b0;

   // m78_22 = W*in
   wire signed [6:0] m78_22;
   assign m78_22 =7'b0;

   // m78_23 = W*in
   wire signed [6:0] m78_23;
   assign m78_23 =7'b0;

   // m78_24 = W*in
   wire signed [6:0] m78_24;
   assign m78_24 =7'b0;

   // m78_25 = W*in
   wire signed [6:0] m78_25;
   assign m78_25 =7'b0;

   // m78_26 = W*in
   wire signed [6:0] m78_26;
   assign m78_26 =7'b0;

   // m78_27 = W*in
   wire signed [6:0] m78_27;
   assign m78_27 =7'b0;

   // m79_1 = W*in
   wire signed [6:0] m79_1;
   assign m79_1 ={ {2{in79[5]}} , in79[5:1] };

   // m79_2 = W*in
   wire signed [6:0] m79_2;
   assign m79_2 =7'b0;

   // m79_3 = W*in
   wire signed [6:0] m79_3;
   assign m79_3 =7'b0;

   // m79_4 = W*in
   wire signed [6:0] m79_4;
   assign m79_4 =7'b0;

   // m79_5 = W*in
   wire signed [6:0] m79_5;
   assign m79_5 =7'b0;

   // m79_6 = W*in
   wire signed [6:0] m79_6;
   assign m79_6 =7'b0;

   // m79_7 = W*in
   wire signed [6:0] m79_7;
   assign m79_7 =7'b0;

   // m79_8 = W*in
   wire signed [6:0] m79_8;
   assign m79_8 =7'b0;

   // m79_9 = W*in
   wire signed [6:0] m79_9;
   assign m79_9 =7'b0;

   // m79_10 = W*in
   wire signed [6:0] m79_10;
   assign m79_10 =7'b0;

   // m79_11 = W*in
   wire signed [6:0] m79_11;
   assign m79_11 =7'b0;

   // m79_12 = W*in
   wire signed [6:0] m79_12;
   assign m79_12 =7'b0;

   // m79_13 = W*in
   wire signed [6:0] m79_13;
   assign m79_13 =7'b0;

   // m79_14 = W*in
   wire signed [6:0] m79_14;
   assign m79_14 =7'b0;

   // m79_15 = W*in
   wire signed [6:0] m79_15;
   assign m79_15 =7'b0;

   // m79_16 = W*in
   wire signed [6:0] m79_16;
   assign m79_16 =7'b0;

   // m79_17 = W*in
   wire signed [6:0] m79_17;
   assign m79_17 =7'b0;

   // m79_18 = W*in
   wire signed [6:0] m79_18;
   assign m79_18 =7'b0;

   // m79_19 = W*in
   wire signed [6:0] m79_19;
   assign m79_19 =7'b0;

   // m79_20 = W*in
   wire signed [6:0] m79_20;
   assign m79_20 =7'b0;

   // m79_21 = W*in
   wire signed [6:0] m79_21;
   assign m79_21 =7'b0;

   // m79_22 = W*in
   wire signed [6:0] m79_22;
   assign m79_22 =7'b0;

   // m79_23 = W*in
   wire signed [6:0] m79_23;
   assign m79_23 =7'b0;

   // m79_24 = W*in
   wire signed [6:0] m79_24;
   assign m79_24 =7'b0;

   // m79_25 = W*in
   wire signed [6:0] m79_25;
   assign m79_25 =7'b0;

   // m79_26 = W*in
   wire signed [6:0] m79_26;
   assign m79_26 =7'b0;

   // m79_27 = W*in
   wire signed [6:0] m79_27;
   assign m79_27 =7'b0;

   // m80_1 = W*in
   wire signed [6:0] m80_1;
   assign m80_1 =7'b0;

   // m80_2 = W*in
   wire signed [6:0] m80_2;
   assign m80_2 =7'b0;

   // m80_3 = W*in
   wire signed [6:0] m80_3;
   assign m80_3 =7'b0;

   // m80_4 = W*in
   wire signed [6:0] m80_4;
   assign m80_4 =7'b0;

   // m80_5 = W*in
   wire signed [6:0] m80_5;
   wire signed [7:0] tm80_5;
   assign tm80_5[0:0] = in80[0:0];
   assign tm80_5[7:1] = { {1{in80[5]}} , in80[5:0] } + { {2{in80[5]}} , in80[5:1] };
   assign m80_5 ={ {1{tm80_5[7]}} , tm80_5[7:2] };

   // m80_6 = W*in
   wire signed [6:0] m80_6;
   assign m80_6 =7'b0;

   // m80_7 = W*in
   wire signed [6:0] m80_7;
   assign m80_7 =7'b0;

   // m80_8 = W*in
   wire signed [6:0] m80_8;
   assign m80_8 =7'b0;

   // m80_9 = W*in
   wire signed [6:0] m80_9;
   assign m80_9 =7'b0;

   // m80_10 = W*in
   wire signed [6:0] m80_10;
   assign m80_10 =7'b0;

   // m80_11 = W*in
   wire signed [6:0] m80_11;
   assign m80_11 =7'b0;

   // m80_12 = W*in
   wire signed [6:0] m80_12;
   assign m80_12 =7'b0;

   // m80_13 = W*in
   wire signed [6:0] m80_13;
   assign m80_13 =7'b0;

   // m80_14 = W*in
   wire signed [6:0] m80_14;
   wire signed [7:0] tm80_14;
   assign tm80_14[0:0] = in80[0:0];
   assign tm80_14[7:1] = { {1{in80[5]}} , in80[5:0] } + { {2{in80[5]}} , in80[5:1] };
   assign m80_14 ={ {1{tm80_14[7]}} , tm80_14[7:2] };

   // m80_15 = W*in
   wire signed [6:0] m80_15;
   assign m80_15 =7'b0;

   // m80_16 = W*in
   wire signed [6:0] m80_16;
   assign m80_16 =7'b0;

   // m80_17 = W*in
   wire signed [6:0] m80_17;
   assign m80_17 ={ {1{in80[5]}} , in80[5:0] };

   // m80_18 = W*in
   wire signed [6:0] m80_18;
   assign m80_18 =7'b0;

   // m80_19 = W*in
   wire signed [6:0] m80_19;
   assign m80_19 =7'b0;

   // m80_20 = W*in
   wire signed [6:0] m80_20;
   assign m80_20 =7'b0;

   // m80_21 = W*in
   wire signed [6:0] m80_21;
   assign m80_21 =7'b0;

   // m80_22 = W*in
   wire signed [6:0] m80_22;
   assign m80_22 =7'b0;

   // m80_23 = W*in
   wire signed [6:0] m80_23;
   assign m80_23 =7'b0;

   // m80_24 = W*in
   wire signed [6:0] m80_24;
   assign m80_24 =7'b0;

   // m80_25 = W*in
   wire signed [6:0] m80_25;
   assign m80_25 =7'b0;

   // m80_26 = W*in
   wire signed [6:0] m80_26;
   assign m80_26 =7'b0;

   // m80_27 = W*in
   wire signed [6:0] m80_27;
   assign m80_27 =7'b0;

   //Perceptron Adders
   assign out1 = m1_1+m2_1+m3_1+m4_1+m5_1+m6_1+m7_1+m8_1+m9_1+m10_1+m11_1+m12_1+m13_1+m14_1+m15_1+m16_1+m17_1+m18_1+m19_1+m20_1+m21_1+m22_1+m23_1+m24_1+m25_1+m26_1+m27_1+m28_1+m29_1+m30_1+m31_1+m32_1+m33_1+m34_1+m35_1+m36_1+m37_1+m38_1+m39_1+m40_1+m41_1+m42_1+m43_1+m44_1+m45_1+m46_1+m47_1+m48_1+m49_1+m50_1+m51_1+m52_1+m53_1+m54_1+m55_1+m56_1+m57_1+m58_1+m59_1+m60_1+m61_1+m62_1+m63_1+m64_1+m65_1+m66_1+m67_1+m68_1+m69_1+m70_1+m71_1+m72_1+m73_1+m74_1+m75_1+m76_1+m77_1+m78_1+m79_1+m80_1+b1;
   assign out2 = m1_2+m2_2+m3_2+m4_2+m5_2+m6_2+m7_2+m8_2+m9_2+m10_2+m11_2+m12_2+m13_2+m14_2+m15_2+m16_2+m17_2+m18_2+m19_2+m20_2+m21_2+m22_2+m23_2+m24_2+m25_2+m26_2+m27_2+m28_2+m29_2+m30_2+m31_2+m32_2+m33_2+m34_2+m35_2+m36_2+m37_2+m38_2+m39_2+m40_2+m41_2+m42_2+m43_2+m44_2+m45_2+m46_2+m47_2+m48_2+m49_2+m50_2+m51_2+m52_2+m53_2+m54_2+m55_2+m56_2+m57_2+m58_2+m59_2+m60_2+m61_2+m62_2+m63_2+m64_2+m65_2+m66_2+m67_2+m68_2+m69_2+m70_2+m71_2+m72_2+m73_2+m74_2+m75_2+m76_2+m77_2+m78_2+m79_2+m80_2+b2;
   assign out3 = m1_3+m2_3+m3_3+m4_3+m5_3+m6_3+m7_3+m8_3+m9_3+m10_3+m11_3+m12_3+m13_3+m14_3+m15_3+m16_3+m17_3+m18_3+m19_3+m20_3+m21_3+m22_3+m23_3+m24_3+m25_3+m26_3+m27_3+m28_3+m29_3+m30_3+m31_3+m32_3+m33_3+m34_3+m35_3+m36_3+m37_3+m38_3+m39_3+m40_3+m41_3+m42_3+m43_3+m44_3+m45_3+m46_3+m47_3+m48_3+m49_3+m50_3+m51_3+m52_3+m53_3+m54_3+m55_3+m56_3+m57_3+m58_3+m59_3+m60_3+m61_3+m62_3+m63_3+m64_3+m65_3+m66_3+m67_3+m68_3+m69_3+m70_3+m71_3+m72_3+m73_3+m74_3+m75_3+m76_3+m77_3+m78_3+m79_3+m80_3+b3;
   assign out4 = m1_4+m2_4+m3_4+m4_4+m5_4+m6_4+m7_4+m8_4+m9_4+m10_4+m11_4+m12_4+m13_4+m14_4+m15_4+m16_4+m17_4+m18_4+m19_4+m20_4+m21_4+m22_4+m23_4+m24_4+m25_4+m26_4+m27_4+m28_4+m29_4+m30_4+m31_4+m32_4+m33_4+m34_4+m35_4+m36_4+m37_4+m38_4+m39_4+m40_4+m41_4+m42_4+m43_4+m44_4+m45_4+m46_4+m47_4+m48_4+m49_4+m50_4+m51_4+m52_4+m53_4+m54_4+m55_4+m56_4+m57_4+m58_4+m59_4+m60_4+m61_4+m62_4+m63_4+m64_4+m65_4+m66_4+m67_4+m68_4+m69_4+m70_4+m71_4+m72_4+m73_4+m74_4+m75_4+m76_4+m77_4+m78_4+m79_4+m80_4+b4;
   assign out5 = m1_5+m2_5+m3_5+m4_5+m5_5+m6_5+m7_5+m8_5+m9_5+m10_5+m11_5+m12_5+m13_5+m14_5+m15_5+m16_5+m17_5+m18_5+m19_5+m20_5+m21_5+m22_5+m23_5+m24_5+m25_5+m26_5+m27_5+m28_5+m29_5+m30_5+m31_5+m32_5+m33_5+m34_5+m35_5+m36_5+m37_5+m38_5+m39_5+m40_5+m41_5+m42_5+m43_5+m44_5+m45_5+m46_5+m47_5+m48_5+m49_5+m50_5+m51_5+m52_5+m53_5+m54_5+m55_5+m56_5+m57_5+m58_5+m59_5+m60_5+m61_5+m62_5+m63_5+m64_5+m65_5+m66_5+m67_5+m68_5+m69_5+m70_5+m71_5+m72_5+m73_5+m74_5+m75_5+m76_5+m77_5+m78_5+m79_5+m80_5+b5;
   assign out6 = m1_6+m2_6+m3_6+m4_6+m5_6+m6_6+m7_6+m8_6+m9_6+m10_6+m11_6+m12_6+m13_6+m14_6+m15_6+m16_6+m17_6+m18_6+m19_6+m20_6+m21_6+m22_6+m23_6+m24_6+m25_6+m26_6+m27_6+m28_6+m29_6+m30_6+m31_6+m32_6+m33_6+m34_6+m35_6+m36_6+m37_6+m38_6+m39_6+m40_6+m41_6+m42_6+m43_6+m44_6+m45_6+m46_6+m47_6+m48_6+m49_6+m50_6+m51_6+m52_6+m53_6+m54_6+m55_6+m56_6+m57_6+m58_6+m59_6+m60_6+m61_6+m62_6+m63_6+m64_6+m65_6+m66_6+m67_6+m68_6+m69_6+m70_6+m71_6+m72_6+m73_6+m74_6+m75_6+m76_6+m77_6+m78_6+m79_6+m80_6+b6;
   assign out7 = m1_7+m2_7+m3_7+m4_7+m5_7+m6_7+m7_7+m8_7+m9_7+m10_7+m11_7+m12_7+m13_7+m14_7+m15_7+m16_7+m17_7+m18_7+m19_7+m20_7+m21_7+m22_7+m23_7+m24_7+m25_7+m26_7+m27_7+m28_7+m29_7+m30_7+m31_7+m32_7+m33_7+m34_7+m35_7+m36_7+m37_7+m38_7+m39_7+m40_7+m41_7+m42_7+m43_7+m44_7+m45_7+m46_7+m47_7+m48_7+m49_7+m50_7+m51_7+m52_7+m53_7+m54_7+m55_7+m56_7+m57_7+m58_7+m59_7+m60_7+m61_7+m62_7+m63_7+m64_7+m65_7+m66_7+m67_7+m68_7+m69_7+m70_7+m71_7+m72_7+m73_7+m74_7+m75_7+m76_7+m77_7+m78_7+m79_7+m80_7+b7;
   assign out8 = m1_8+m2_8+m3_8+m4_8+m5_8+m6_8+m7_8+m8_8+m9_8+m10_8+m11_8+m12_8+m13_8+m14_8+m15_8+m16_8+m17_8+m18_8+m19_8+m20_8+m21_8+m22_8+m23_8+m24_8+m25_8+m26_8+m27_8+m28_8+m29_8+m30_8+m31_8+m32_8+m33_8+m34_8+m35_8+m36_8+m37_8+m38_8+m39_8+m40_8+m41_8+m42_8+m43_8+m44_8+m45_8+m46_8+m47_8+m48_8+m49_8+m50_8+m51_8+m52_8+m53_8+m54_8+m55_8+m56_8+m57_8+m58_8+m59_8+m60_8+m61_8+m62_8+m63_8+m64_8+m65_8+m66_8+m67_8+m68_8+m69_8+m70_8+m71_8+m72_8+m73_8+m74_8+m75_8+m76_8+m77_8+m78_8+m79_8+m80_8+b8;
   assign out9 = m1_9+m2_9+m3_9+m4_9+m5_9+m6_9+m7_9+m8_9+m9_9+m10_9+m11_9+m12_9+m13_9+m14_9+m15_9+m16_9+m17_9+m18_9+m19_9+m20_9+m21_9+m22_9+m23_9+m24_9+m25_9+m26_9+m27_9+m28_9+m29_9+m30_9+m31_9+m32_9+m33_9+m34_9+m35_9+m36_9+m37_9+m38_9+m39_9+m40_9+m41_9+m42_9+m43_9+m44_9+m45_9+m46_9+m47_9+m48_9+m49_9+m50_9+m51_9+m52_9+m53_9+m54_9+m55_9+m56_9+m57_9+m58_9+m59_9+m60_9+m61_9+m62_9+m63_9+m64_9+m65_9+m66_9+m67_9+m68_9+m69_9+m70_9+m71_9+m72_9+m73_9+m74_9+m75_9+m76_9+m77_9+m78_9+m79_9+m80_9+b9;
   assign out10 = m1_10+m2_10+m3_10+m4_10+m5_10+m6_10+m7_10+m8_10+m9_10+m10_10+m11_10+m12_10+m13_10+m14_10+m15_10+m16_10+m17_10+m18_10+m19_10+m20_10+m21_10+m22_10+m23_10+m24_10+m25_10+m26_10+m27_10+m28_10+m29_10+m30_10+m31_10+m32_10+m33_10+m34_10+m35_10+m36_10+m37_10+m38_10+m39_10+m40_10+m41_10+m42_10+m43_10+m44_10+m45_10+m46_10+m47_10+m48_10+m49_10+m50_10+m51_10+m52_10+m53_10+m54_10+m55_10+m56_10+m57_10+m58_10+m59_10+m60_10+m61_10+m62_10+m63_10+m64_10+m65_10+m66_10+m67_10+m68_10+m69_10+m70_10+m71_10+m72_10+m73_10+m74_10+m75_10+m76_10+m77_10+m78_10+m79_10+m80_10+b10;
   assign out11 = m1_11+m2_11+m3_11+m4_11+m5_11+m6_11+m7_11+m8_11+m9_11+m10_11+m11_11+m12_11+m13_11+m14_11+m15_11+m16_11+m17_11+m18_11+m19_11+m20_11+m21_11+m22_11+m23_11+m24_11+m25_11+m26_11+m27_11+m28_11+m29_11+m30_11+m31_11+m32_11+m33_11+m34_11+m35_11+m36_11+m37_11+m38_11+m39_11+m40_11+m41_11+m42_11+m43_11+m44_11+m45_11+m46_11+m47_11+m48_11+m49_11+m50_11+m51_11+m52_11+m53_11+m54_11+m55_11+m56_11+m57_11+m58_11+m59_11+m60_11+m61_11+m62_11+m63_11+m64_11+m65_11+m66_11+m67_11+m68_11+m69_11+m70_11+m71_11+m72_11+m73_11+m74_11+m75_11+m76_11+m77_11+m78_11+m79_11+m80_11+b11;
   assign out12 = m1_12+m2_12+m3_12+m4_12+m5_12+m6_12+m7_12+m8_12+m9_12+m10_12+m11_12+m12_12+m13_12+m14_12+m15_12+m16_12+m17_12+m18_12+m19_12+m20_12+m21_12+m22_12+m23_12+m24_12+m25_12+m26_12+m27_12+m28_12+m29_12+m30_12+m31_12+m32_12+m33_12+m34_12+m35_12+m36_12+m37_12+m38_12+m39_12+m40_12+m41_12+m42_12+m43_12+m44_12+m45_12+m46_12+m47_12+m48_12+m49_12+m50_12+m51_12+m52_12+m53_12+m54_12+m55_12+m56_12+m57_12+m58_12+m59_12+m60_12+m61_12+m62_12+m63_12+m64_12+m65_12+m66_12+m67_12+m68_12+m69_12+m70_12+m71_12+m72_12+m73_12+m74_12+m75_12+m76_12+m77_12+m78_12+m79_12+m80_12+b12;
   assign out13 = m1_13+m2_13+m3_13+m4_13+m5_13+m6_13+m7_13+m8_13+m9_13+m10_13+m11_13+m12_13+m13_13+m14_13+m15_13+m16_13+m17_13+m18_13+m19_13+m20_13+m21_13+m22_13+m23_13+m24_13+m25_13+m26_13+m27_13+m28_13+m29_13+m30_13+m31_13+m32_13+m33_13+m34_13+m35_13+m36_13+m37_13+m38_13+m39_13+m40_13+m41_13+m42_13+m43_13+m44_13+m45_13+m46_13+m47_13+m48_13+m49_13+m50_13+m51_13+m52_13+m53_13+m54_13+m55_13+m56_13+m57_13+m58_13+m59_13+m60_13+m61_13+m62_13+m63_13+m64_13+m65_13+m66_13+m67_13+m68_13+m69_13+m70_13+m71_13+m72_13+m73_13+m74_13+m75_13+m76_13+m77_13+m78_13+m79_13+m80_13+b13;
   assign out14 = m1_14+m2_14+m3_14+m4_14+m5_14+m6_14+m7_14+m8_14+m9_14+m10_14+m11_14+m12_14+m13_14+m14_14+m15_14+m16_14+m17_14+m18_14+m19_14+m20_14+m21_14+m22_14+m23_14+m24_14+m25_14+m26_14+m27_14+m28_14+m29_14+m30_14+m31_14+m32_14+m33_14+m34_14+m35_14+m36_14+m37_14+m38_14+m39_14+m40_14+m41_14+m42_14+m43_14+m44_14+m45_14+m46_14+m47_14+m48_14+m49_14+m50_14+m51_14+m52_14+m53_14+m54_14+m55_14+m56_14+m57_14+m58_14+m59_14+m60_14+m61_14+m62_14+m63_14+m64_14+m65_14+m66_14+m67_14+m68_14+m69_14+m70_14+m71_14+m72_14+m73_14+m74_14+m75_14+m76_14+m77_14+m78_14+m79_14+m80_14+b14;
   assign out15 = m1_15+m2_15+m3_15+m4_15+m5_15+m6_15+m7_15+m8_15+m9_15+m10_15+m11_15+m12_15+m13_15+m14_15+m15_15+m16_15+m17_15+m18_15+m19_15+m20_15+m21_15+m22_15+m23_15+m24_15+m25_15+m26_15+m27_15+m28_15+m29_15+m30_15+m31_15+m32_15+m33_15+m34_15+m35_15+m36_15+m37_15+m38_15+m39_15+m40_15+m41_15+m42_15+m43_15+m44_15+m45_15+m46_15+m47_15+m48_15+m49_15+m50_15+m51_15+m52_15+m53_15+m54_15+m55_15+m56_15+m57_15+m58_15+m59_15+m60_15+m61_15+m62_15+m63_15+m64_15+m65_15+m66_15+m67_15+m68_15+m69_15+m70_15+m71_15+m72_15+m73_15+m74_15+m75_15+m76_15+m77_15+m78_15+m79_15+m80_15+b15;
   assign out16 = m1_16+m2_16+m3_16+m4_16+m5_16+m6_16+m7_16+m8_16+m9_16+m10_16+m11_16+m12_16+m13_16+m14_16+m15_16+m16_16+m17_16+m18_16+m19_16+m20_16+m21_16+m22_16+m23_16+m24_16+m25_16+m26_16+m27_16+m28_16+m29_16+m30_16+m31_16+m32_16+m33_16+m34_16+m35_16+m36_16+m37_16+m38_16+m39_16+m40_16+m41_16+m42_16+m43_16+m44_16+m45_16+m46_16+m47_16+m48_16+m49_16+m50_16+m51_16+m52_16+m53_16+m54_16+m55_16+m56_16+m57_16+m58_16+m59_16+m60_16+m61_16+m62_16+m63_16+m64_16+m65_16+m66_16+m67_16+m68_16+m69_16+m70_16+m71_16+m72_16+m73_16+m74_16+m75_16+m76_16+m77_16+m78_16+m79_16+m80_16+b16;
   assign out17 = m1_17+m2_17+m3_17+m4_17+m5_17+m6_17+m7_17+m8_17+m9_17+m10_17+m11_17+m12_17+m13_17+m14_17+m15_17+m16_17+m17_17+m18_17+m19_17+m20_17+m21_17+m22_17+m23_17+m24_17+m25_17+m26_17+m27_17+m28_17+m29_17+m30_17+m31_17+m32_17+m33_17+m34_17+m35_17+m36_17+m37_17+m38_17+m39_17+m40_17+m41_17+m42_17+m43_17+m44_17+m45_17+m46_17+m47_17+m48_17+m49_17+m50_17+m51_17+m52_17+m53_17+m54_17+m55_17+m56_17+m57_17+m58_17+m59_17+m60_17+m61_17+m62_17+m63_17+m64_17+m65_17+m66_17+m67_17+m68_17+m69_17+m70_17+m71_17+m72_17+m73_17+m74_17+m75_17+m76_17+m77_17+m78_17+m79_17+m80_17+b17;
   assign out18 = m1_18+m2_18+m3_18+m4_18+m5_18+m6_18+m7_18+m8_18+m9_18+m10_18+m11_18+m12_18+m13_18+m14_18+m15_18+m16_18+m17_18+m18_18+m19_18+m20_18+m21_18+m22_18+m23_18+m24_18+m25_18+m26_18+m27_18+m28_18+m29_18+m30_18+m31_18+m32_18+m33_18+m34_18+m35_18+m36_18+m37_18+m38_18+m39_18+m40_18+m41_18+m42_18+m43_18+m44_18+m45_18+m46_18+m47_18+m48_18+m49_18+m50_18+m51_18+m52_18+m53_18+m54_18+m55_18+m56_18+m57_18+m58_18+m59_18+m60_18+m61_18+m62_18+m63_18+m64_18+m65_18+m66_18+m67_18+m68_18+m69_18+m70_18+m71_18+m72_18+m73_18+m74_18+m75_18+m76_18+m77_18+m78_18+m79_18+m80_18+b18;
   assign out19 = m1_19+m2_19+m3_19+m4_19+m5_19+m6_19+m7_19+m8_19+m9_19+m10_19+m11_19+m12_19+m13_19+m14_19+m15_19+m16_19+m17_19+m18_19+m19_19+m20_19+m21_19+m22_19+m23_19+m24_19+m25_19+m26_19+m27_19+m28_19+m29_19+m30_19+m31_19+m32_19+m33_19+m34_19+m35_19+m36_19+m37_19+m38_19+m39_19+m40_19+m41_19+m42_19+m43_19+m44_19+m45_19+m46_19+m47_19+m48_19+m49_19+m50_19+m51_19+m52_19+m53_19+m54_19+m55_19+m56_19+m57_19+m58_19+m59_19+m60_19+m61_19+m62_19+m63_19+m64_19+m65_19+m66_19+m67_19+m68_19+m69_19+m70_19+m71_19+m72_19+m73_19+m74_19+m75_19+m76_19+m77_19+m78_19+m79_19+m80_19+b19;
   assign out20 = m1_20+m2_20+m3_20+m4_20+m5_20+m6_20+m7_20+m8_20+m9_20+m10_20+m11_20+m12_20+m13_20+m14_20+m15_20+m16_20+m17_20+m18_20+m19_20+m20_20+m21_20+m22_20+m23_20+m24_20+m25_20+m26_20+m27_20+m28_20+m29_20+m30_20+m31_20+m32_20+m33_20+m34_20+m35_20+m36_20+m37_20+m38_20+m39_20+m40_20+m41_20+m42_20+m43_20+m44_20+m45_20+m46_20+m47_20+m48_20+m49_20+m50_20+m51_20+m52_20+m53_20+m54_20+m55_20+m56_20+m57_20+m58_20+m59_20+m60_20+m61_20+m62_20+m63_20+m64_20+m65_20+m66_20+m67_20+m68_20+m69_20+m70_20+m71_20+m72_20+m73_20+m74_20+m75_20+m76_20+m77_20+m78_20+m79_20+m80_20+b20;
   assign out21 = m1_21+m2_21+m3_21+m4_21+m5_21+m6_21+m7_21+m8_21+m9_21+m10_21+m11_21+m12_21+m13_21+m14_21+m15_21+m16_21+m17_21+m18_21+m19_21+m20_21+m21_21+m22_21+m23_21+m24_21+m25_21+m26_21+m27_21+m28_21+m29_21+m30_21+m31_21+m32_21+m33_21+m34_21+m35_21+m36_21+m37_21+m38_21+m39_21+m40_21+m41_21+m42_21+m43_21+m44_21+m45_21+m46_21+m47_21+m48_21+m49_21+m50_21+m51_21+m52_21+m53_21+m54_21+m55_21+m56_21+m57_21+m58_21+m59_21+m60_21+m61_21+m62_21+m63_21+m64_21+m65_21+m66_21+m67_21+m68_21+m69_21+m70_21+m71_21+m72_21+m73_21+m74_21+m75_21+m76_21+m77_21+m78_21+m79_21+m80_21+b21;
   assign out22 = m1_22+m2_22+m3_22+m4_22+m5_22+m6_22+m7_22+m8_22+m9_22+m10_22+m11_22+m12_22+m13_22+m14_22+m15_22+m16_22+m17_22+m18_22+m19_22+m20_22+m21_22+m22_22+m23_22+m24_22+m25_22+m26_22+m27_22+m28_22+m29_22+m30_22+m31_22+m32_22+m33_22+m34_22+m35_22+m36_22+m37_22+m38_22+m39_22+m40_22+m41_22+m42_22+m43_22+m44_22+m45_22+m46_22+m47_22+m48_22+m49_22+m50_22+m51_22+m52_22+m53_22+m54_22+m55_22+m56_22+m57_22+m58_22+m59_22+m60_22+m61_22+m62_22+m63_22+m64_22+m65_22+m66_22+m67_22+m68_22+m69_22+m70_22+m71_22+m72_22+m73_22+m74_22+m75_22+m76_22+m77_22+m78_22+m79_22+m80_22+b22;
   assign out23 = m1_23+m2_23+m3_23+m4_23+m5_23+m6_23+m7_23+m8_23+m9_23+m10_23+m11_23+m12_23+m13_23+m14_23+m15_23+m16_23+m17_23+m18_23+m19_23+m20_23+m21_23+m22_23+m23_23+m24_23+m25_23+m26_23+m27_23+m28_23+m29_23+m30_23+m31_23+m32_23+m33_23+m34_23+m35_23+m36_23+m37_23+m38_23+m39_23+m40_23+m41_23+m42_23+m43_23+m44_23+m45_23+m46_23+m47_23+m48_23+m49_23+m50_23+m51_23+m52_23+m53_23+m54_23+m55_23+m56_23+m57_23+m58_23+m59_23+m60_23+m61_23+m62_23+m63_23+m64_23+m65_23+m66_23+m67_23+m68_23+m69_23+m70_23+m71_23+m72_23+m73_23+m74_23+m75_23+m76_23+m77_23+m78_23+m79_23+m80_23+b23;
   assign out24 = m1_24+m2_24+m3_24+m4_24+m5_24+m6_24+m7_24+m8_24+m9_24+m10_24+m11_24+m12_24+m13_24+m14_24+m15_24+m16_24+m17_24+m18_24+m19_24+m20_24+m21_24+m22_24+m23_24+m24_24+m25_24+m26_24+m27_24+m28_24+m29_24+m30_24+m31_24+m32_24+m33_24+m34_24+m35_24+m36_24+m37_24+m38_24+m39_24+m40_24+m41_24+m42_24+m43_24+m44_24+m45_24+m46_24+m47_24+m48_24+m49_24+m50_24+m51_24+m52_24+m53_24+m54_24+m55_24+m56_24+m57_24+m58_24+m59_24+m60_24+m61_24+m62_24+m63_24+m64_24+m65_24+m66_24+m67_24+m68_24+m69_24+m70_24+m71_24+m72_24+m73_24+m74_24+m75_24+m76_24+m77_24+m78_24+m79_24+m80_24+b24;
   assign out25 = m1_25+m2_25+m3_25+m4_25+m5_25+m6_25+m7_25+m8_25+m9_25+m10_25+m11_25+m12_25+m13_25+m14_25+m15_25+m16_25+m17_25+m18_25+m19_25+m20_25+m21_25+m22_25+m23_25+m24_25+m25_25+m26_25+m27_25+m28_25+m29_25+m30_25+m31_25+m32_25+m33_25+m34_25+m35_25+m36_25+m37_25+m38_25+m39_25+m40_25+m41_25+m42_25+m43_25+m44_25+m45_25+m46_25+m47_25+m48_25+m49_25+m50_25+m51_25+m52_25+m53_25+m54_25+m55_25+m56_25+m57_25+m58_25+m59_25+m60_25+m61_25+m62_25+m63_25+m64_25+m65_25+m66_25+m67_25+m68_25+m69_25+m70_25+m71_25+m72_25+m73_25+m74_25+m75_25+m76_25+m77_25+m78_25+m79_25+m80_25+b25;
   assign out26 = m1_26+m2_26+m3_26+m4_26+m5_26+m6_26+m7_26+m8_26+m9_26+m10_26+m11_26+m12_26+m13_26+m14_26+m15_26+m16_26+m17_26+m18_26+m19_26+m20_26+m21_26+m22_26+m23_26+m24_26+m25_26+m26_26+m27_26+m28_26+m29_26+m30_26+m31_26+m32_26+m33_26+m34_26+m35_26+m36_26+m37_26+m38_26+m39_26+m40_26+m41_26+m42_26+m43_26+m44_26+m45_26+m46_26+m47_26+m48_26+m49_26+m50_26+m51_26+m52_26+m53_26+m54_26+m55_26+m56_26+m57_26+m58_26+m59_26+m60_26+m61_26+m62_26+m63_26+m64_26+m65_26+m66_26+m67_26+m68_26+m69_26+m70_26+m71_26+m72_26+m73_26+m74_26+m75_26+m76_26+m77_26+m78_26+m79_26+m80_26+b26;
   assign out27 = m1_27+m2_27+m3_27+m4_27+m5_27+m6_27+m7_27+m8_27+m9_27+m10_27+m11_27+m12_27+m13_27+m14_27+m15_27+m16_27+m17_27+m18_27+m19_27+m20_27+m21_27+m22_27+m23_27+m24_27+m25_27+m26_27+m27_27+m28_27+m29_27+m30_27+m31_27+m32_27+m33_27+m34_27+m35_27+m36_27+m37_27+m38_27+m39_27+m40_27+m41_27+m42_27+m43_27+m44_27+m45_27+m46_27+m47_27+m48_27+m49_27+m50_27+m51_27+m52_27+m53_27+m54_27+m55_27+m56_27+m57_27+m58_27+m59_27+m60_27+m61_27+m62_27+m63_27+m64_27+m65_27+m66_27+m67_27+m68_27+m69_27+m70_27+m71_27+m72_27+m73_27+m74_27+m75_27+m76_27+m77_27+m78_27+m79_27+m80_27+b27;
endmodule